
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_SPEEDY_Top is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_SPEEDY_Top;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Rounds7_0 is

   port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : out
         std_logic_vector (191 downto 0));

end SPEEDY_Rounds7_0;

architecture SYN_Behavioral of SPEEDY_Rounds7_0 is

   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n19, 
      n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n39
      , n40, n41, n42, n43, n44, n46, n48, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n63, n64, n66, n69, n71, n72, n73, n75, n76, n77, n79
      , n80, n81, n82, n84, n85, n87, n88, n89, n91, n92, n96, n97, n100, n101,
      n104, n105, n106, n107, n109, n111, n112, n113, n114, n117, n118, n119, 
      n120, n121, n122, n123, n125, n127, n128, n130, n132, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n153, n155, n156, n157, n159, n161, n162, n163, n165, n167, n168, 
      n169, n170, n171, n172, n174, n175, n178, n179, n180, n181, n182, n183, 
      n184, n186, n187, n188, n189, n190, n191, n192, n193, n195, n196, n197, 
      n198, n199, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n215, n216, n217, n219, n220, n221, n223, n224, n225, 
      n226, n227, n229, n231, n232, n233, n235, n237, n238, n240, n241, n242, 
      n243, n244, n245, n248, n249, n250, n251, n252, n253, n255, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n283, n284, 
      n285, n287, n292, n293, n294, n295, n296, n297, n300, n301, n303, n306, 
      n307, n308, n320, n321, n323, n324, n325, n326, n329, n333, n336, n337, 
      n339, n341, n342, n349, n351, n355, n359, n363, n365, n370, n371, n373, 
      n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
      n386, n387, n388, n389, n390, n391, n393, n394, n395, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n412, n413, 
      n414, n415, n416, n417, n418, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n449, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n468, 
      n469, n470, n471, n473, n474, n475, n476, n477, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n538, n539, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n577, n578, n579, n580, n581, n582, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n612, n613, n614, n615, n616, n617, n618, n619, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n678, n679, n680, n681, n683, n686, n688, n689, n690, n691, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n705, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n717, n719, 
      n720, n721, n722, n724, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n753, n754, n755, n756, n757, n758, n760, 
      n761, n762, n763, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
      n786, n787, n788, n790, n792, n794, n795, n796, n797, n798, n799, n800, 
      n801, n802, n803, n804, n805, n806, n807, n808, n810, n811, n812, n813, 
      n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, 
      n826, n827, n828, n829, n830, n831, n832, n834, n835, n836, n837, n839, 
      n840, n841, n842, n843, n844, n846, n847, n848, n850, n851, n852, n853, 
      n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, 
      n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, 
      n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, 
      n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, 
      n903, n905, n906, n907, n908, n909, n910, n912, n913, n914, n916, n917, 
      n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, 
      n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
      n942, n943, n944, n945, n946, n947, n948, n949, n951, n952, n953, n954, 
      n956, n957, n958, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n977, n980, n981, n983, n984, 
      n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n996, n997, 
      n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008
      , n1009, n1010, n1011, n1012, n1013, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1028, n1029, n1030, 
      n1032, n1033, n1034, n1035, n1037, n1040, n1041, n1042, n1043, n1044, 
      n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
      n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1073, n1075, n1076, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1094, n1095, n1096, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1137, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1169, n1170, n1171, n1172, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1196, n1198, n1199, n1200, n1201, 
      n1202, n1203, n1204, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1223, 
      n1224, n1225, n1226, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1306, n1307, 
      n1308, n1309, n1310, n1311, n1312, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1326, n1327, n1328, n1329, 
      n1330, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1342, n1344, n1345, n1346, n1348, n1349, n1350, n1351, n1352, n1353, 
      n1354, n1355, n1356, n1357, n1358, n1359, n1361, n1362, n1363, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387, 
      n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1410, n1411, n1412, n1413, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1433, 
      n1434, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1487, n1489, n1490, 
      n1491, n1493, n1494, n1495, n1496, n1497, n1498, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1521, n1522, n1523, 
      n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, 
      n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, 
      n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, 
      n1554, n1555, n1556, n1558, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1574, n1575, n1576, n1577, 
      n1580, n1581, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, 
      n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, 
      n1602, n1603, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, 
      n1614, n1615, n1616, n1617, n1619, n1620, n1621, n1622, n1623, n1624, 
      n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1634, n1635, 
      n1637, n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, 
      n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
      n1668, n1669, n1670, n1671, n1673, n1674, n1675, n1676, n1679, n1681, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1690, n1691, n1692, n1693, 
      n1694, n1695, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
      n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
      n1715, n1716, n1717, n1718, n1720, n1721, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1755, n1756, n1757, 
      n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1807, n1808, n1809, n1810, 
      n1811, n1812, n1813, n1814, n1816, n1817, n1818, n1819, n1820, n1821, 
      n1822, n1823, n1824, n1825, n1826, n1828, n1829, n1830, n1831, n1832, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1844, n1845, n1846, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
      n1855, n1856, n1857, n1858, n1859, n1861, n1862, n1863, n1864, n1865, 
      n1868, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1883, n1884, n1885, n1886, n1887, n1888, n1890, n1891, 
      n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, 
      n1902, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1933, 
      n1934, n1938, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, 
      n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, 
      n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
      n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2078, n2079, 
      n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
      n2090, n2091, n2092, n2093, n2094, n2096, n2097, n2098, n2099, n2101, 
      n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2127, n2128, n2129, n2130, n2131, n2132, n2133, 
      n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
      n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, 
      n2154, n2155, n2157, n2158, n2159, n2160, n2161, n2162, n2164, n2165, 
      n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, 
      n2176, n2177, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2196, n2199, 
      n2200, n2201, n2202, n2203, n2205, n2206, n2207, n2208, n2209, n2210, 
      n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2234, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2246, n2247, n2248, n2250, n2251, n2255, n2256, n2257, 
      n2258, n2259, n2260, n2261, n2262, n2263, n2265, n2266, n2267, n2268, 
      n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2278, n2281, 
      n2282, n2283, n2285, n2286, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2299, n2300, n2301, n2302, n2303, n2304, 
      n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, 
      n2315, n2316, n2317, n2318, n2319, n2320, n2323, n2324, n2325, n2326, 
      n2327, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
      n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, 
      n2348, n2349, n2350, n2351, n2352, n2353, n2355, n2357, n2358, n2359, 
      n2360, n2361, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2371, 
      n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, 
      n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, 
      n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, 
      n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, 
      n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2437, n2438, n2439, n2440, n2441, n2442, n2444, 
      n2445, n2446, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, 
      n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, 
      n2466, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2480, n2481, n2482, n2483, n2484, n2485, n2487, n2488, n2489, 
      n2490, n2491, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
      n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, 
      n2511, n2514, n2516, n2518, n2519, n2520, n2521, n2522, n2523, n2524, 
      n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, 
      n2538, n2539, n2541, n2542, n2544, n2545, n2546, n2547, n2549, n2551, 
      n2552, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2589, n2590, n2591, n2592, n2593, 
      n2594, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2617, 
      n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
      n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
      n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, 
      n2648, n2649, n2650, n2651, n2652, n2653, n2655, n2656, n2657, n2658, 
      n2659, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2675, n2676, n2677, n2678, n2680, n2681, n2682, n2683, 
      n2684, n2685, n2687, n2688, n2689, n2690, n2691, n2692, n2694, n2695, 
      n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2704, n2705, n2707, 
      n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
      n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
      n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, 
      n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, 
      n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, 
      n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
      n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2870, 
      n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
      n2882, n2883, n2884, n2885, n2887, n2888, n2889, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2911, n2912, n2913, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2934, n2935, n2937, n2938, n2939, 
      n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
      n2950, n2951, n2952, n2954, n2956, n2957, n2958, n2959, n2960, n2961, 
      n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2999, n3001, n3002, n3003, n3004, n3005, 
      n3006, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, 
      n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, 
      n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3097, n3099, n3100, 
      n3101, n3103, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3121, n3123, n3124, 
      n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3134, n3135, 
      n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, 
      n3146, n3147, n3148, n3149, n3150, n3151, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3174, n3175, n3176, n3177, 
      n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3196, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3210, 
      n3211, n3212, n3213, n3214, n3216, n3217, n3218, n3219, n3220, n3221, 
      n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3254, 
      n3255, n3256, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3266, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3279, n3280, 
      n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, 
      n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, 
      n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, 
      n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, 
      n3321, n3322, n3323, n3325, n3326, n3328, n3329, n3330, n3331, n3332, 
      n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, 
      n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
      n3354, n3356, n3357, n3359, n3360, n3361, n3362, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3382, n3383, n3384, n3385, n3386, n3387, n3390, n3391, 
      n3392, n3393, n3395, n3396, n3397, n3400, n3401, n3402, n3403, n3405, 
      n3406, n3407, n3408, n3409, n3410, n3411, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, 
      n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, 
      n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, 
      n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, 
      n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3473, n3474, n3475, n3477, n3478, n3479, n3480, 
      n3481, n3482, n3483, n3484, n3486, n3487, n3488, n3489, n3490, n3491, 
      n3492, n3493, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3523, n3524, 
      n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, 
      n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, 
      n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, 
      n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, 
      n3565, n3566, n3567, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
      n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3592, n3593, n3594, n3595, n3596, n3597, 
      n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3629, 
      n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, 
      n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, 
      n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, 
      n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, 
      n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, 
      n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, 
      n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, 
      n3701, n3702, n3703, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, 
      n3745, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, 
      n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, 
      n3766, n3768, n3770, n3771, n3773, n3774, n3775, n3776, n3777, n3778, 
      n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, 
      n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, 
      n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, 
      n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, 
      n3819, n3820, n3821, n3823, n3824, n3825, n3826, n3827, n3828, n3829, 
      n3830, n3831, n3832, n3833, n3834, n3836, n3837, n3838, n3839, n3840, 
      n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, 
      n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, 
      n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, 
      n3871, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, 
      n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, 
      n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, 
      n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, 
      n3912, n3913, n3914, n3915, n3917, n3918, n3919, n3921, n3922, n3923, 
      n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, 
      n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, 
      n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, 
      n3954, n3955, n3956, n3957, n3958, n3960, n3961, n3962, n3963, n3964, 
      n3965, n3966, n3967, n3968, n3969, n3971, n3972, n3973, n3974, n3975, 
      n3976, n3977, n3978, n3979, n3980, n3981, n3983, n3984, n3985, n3986, 
      n3987, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, 
      n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, 
      n4008, n4009, n4010, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
      n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, 
      n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, 
      n4060, n4061, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, 
      n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, 
      n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, 
      n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4099, n4100, n4101, 
      n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, 
      n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, 
      n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4132, 
      n4133, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, 
      n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, 
      n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, 
      n4165, n4166, n4167, n4168, n4169, n4171, n4172, n4173, n4174, n4175, 
      n4176, n4177, n4178, n4179, n4180, n4181, n4184, n4185, n4186, n4188, 
      n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4197, n4198, n4199, 
      n4200, n4201, n4202, n4203, n4206, n4209, n4210, n4211, n4212, n4213, 
      n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, 
      n4224, n4225, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
      n4235, n4236, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, 
      n4246, n4247, n4248, n4250, n4251, n4252, n4253, n4254, n4255, n4256, 
      n4258, n4259, n4260, n4261, n4263, n4264, n4265, n4266, n4267, n4268, 
      n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, 
      n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, 
      n4290, n4291, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, 
      n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, 
      n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, 
      n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, 
      n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, 
      n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, 
      n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, 
      n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, 
      n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, 
      n4382, n4383, n4384, n4385, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4409, n4410, n4411, n4412, n4413, n4414, 
      n4415, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, 
      n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, 
      n4436, n4438, n4439, n4440, n4441, n4442, n4443, n4446, n4447, n4448, 
      n4449, n4450, n4451, n4452, n4453, n4455, n4456, n4457, n4458, n4459, 
      n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, 
      n4470, n4472, n4473, n4474, n4476, n4477, n4478, n4479, n4480, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4519, n4520, n4521, n4522, n4523, n4524, 
      n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4535, 
      n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4545, n4546, 
      n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, 
      n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, 
      n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, 
      n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, 
      n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, 
      n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, 
      n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, 
      n4617, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, 
      n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4638, n4639, 
      n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, 
      n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, 
      n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4669, n4670, 
      n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, 
      n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, 
      n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, 
      n4701, n4702, n4703, n4705, n4706, n4707, n4708, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4741, n4744, n4745, n4746, 
      n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, 
      n4757, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, 
      n4768, n4769, n4770, n4772, n4773, n4774, n4776, n4777, n4778, n4779, 
      n4780, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4819, n4820, n4821, n4822, n4823, n4824, 
      n4825, n4826, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, 
      n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, 
      n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, 
      n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, 
      n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, 
      n4876, n4877, n4878, n4880, n4881, n4882, n4883, n4884, n4885, n4886, 
      n4887, n4888, n4889, n4891, n4892, n4893, n4894, n4895, n4896, n4897, 
      n4900, n4901, n4902, n4903, n4904, n4905, n4907, n4908, n4909, n4910, 
      n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4921, 
      n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, 
      n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, 
      n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4950, n4951, n4953, 
      n4954, n4955, n4956, n4957, n4959, n4960, n4961, n4962, n4963, n4965, 
      n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, 
      n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4984, n4985, n4986, 
      n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, 
      n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, 
      n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, 
      n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5028, 
      n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, 
      n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, 
      n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, 
      n5059, n5060, n5061, n5062, n5063, n5064, n5066, n5067, n5068, n5069, 
      n5070, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, 
      n5081, n5082, n5083, n5084, n5086, n5087, n5088, n5089, n5090, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5109, n5112, n5113, n5114, n5115, 
      n5116, n5117, n5118, n5120, n5121, n5122, n5123, n5124, n5125, n5126, 
      n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5136, n5137, 
      n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5146, n5147, n5148, 
      n5149, n5150, n5151, n5154, n5155, n5157, n5158, n5159, n5160, n5161, 
      n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, 
      n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, 
      n5182, n5184, n5185, n5186, n5188, n5189, n5190, n5191, n5192, n5193, 
      n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5203, n5204, 
      n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, 
      n5215, n5216, n5217, n5218, n5219, n5221, n5222, n5223, n5224, n5225, 
      n5226, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, 
      n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, 
      n5248, n5250, n5251, n5252, n5253, n5255, n5256, n5257, n5258, n5259, 
      n5260, n5261, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5272, 
      n5273, n5274, n5275, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5287, n5288, n5289, n5291, n5292, n5293, n5294, n5295, 
      n5297, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, 
      n5308, n5309, n5310, n5312, n5313, n5314, n5315, n5316, n5317, n5318, 
      n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, 
      n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
      n5341, n5342, n5343, n5344, n5346, n5347, n5348, n5349, n5350, n5351, 
      n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, 
      n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, 
      n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5381, n5382, 
      n5383, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, 
      n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5424, n5425, n5426, 
      n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, 
      n5437, n5439, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, 
      n5449, n5450, n5451, n5452, n5453, n5454, n5456, n5457, n5458, n5459, 
      n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
      n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, 
      n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, 
      n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, 
      n5500, n5501, n5502, n5504, n5505, n5507, n5508, n5509, n5510, n5511, 
      n5512, n5513, n5514, n5515, n5517, n5518, n5519, n5520, n5521, n5522, 
      n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, 
      n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, 
      n5543, n5544, n5545, n5546, n5547, n5548, n5550, n5551, n5552, n5553, 
      n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, 
      n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, 
      n5574, n5575, n5576, n5577, n5578, n5579, n5581, n5582, n5584, n5585, 
      n5586, n5587, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, 
      n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, 
      n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, 
      n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, 
      n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, 
      n5637, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, 
      n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, 
      n5659, n5660, n5661, n5663, n5664, n5665, n5666, n5667, n5668, n5669, 
      n5670, n5671, n5672, n5673, n5674, n5676, n5677, n5678, n5679, n5680, 
      n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, 
      n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, 
      n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5709, n5710, n5712, 
      n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, 
      n5723, n5724, n5725, n5726, n5728, n5729, n5730, n5731, n5732, n5733, 
      n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, 
      n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, 
      n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5763, n5764, n5767, 
      n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, 
      n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5788, 
      n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, 
      n5799, n5801, n5802, n5803, n5804, n5805, n5807, n5808, n5809, n5810, 
      n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, 
      n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5830, n5831, n5832, 
      n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, 
      n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, 
      n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5862, n5863, n5865, 
      n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5877, 
      n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, 
      n5888, n5889, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, 
      n5899, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, 
      n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, 
      n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, 
      n5930, n5931, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, 
      n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, 
      n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, 
      n5961, n5962, n5963, n5964, n5966, n5967, n5968, n5969, n5970, n5971, 
      n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, 
      n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5992, n5993, n5994, n5995, n5996, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, 
      n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, 
      n6025, n6026, n6027, n6028, n6029, n6030, n6032, n6033, n6034, n6035, 
      n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, 
      n6046, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, 
      n6057, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, 
      n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
      n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, 
      n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6097, n6098, 
      n6099, n6100, n6101, n6103, n6104, n6105, n6106, n6107, n6108, n6109, 
      n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, 
      n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6128, n6130, n6132, 
      n6133, n6134, n6135, n6136, n6137, n6139, n6140, n6141, n6142, n6143, 
      n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, 
      n6154, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, 
      n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, 
      n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, 
      n6185, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, 
      n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, 
      n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6215, n6216, n6217, 
      n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, 
      n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, 
      n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, 
      n6248, n6249, n6250, n6252, n6253, n6254, n6255, n6256, n6257, n6259, 
      n6260, n6261, n6262, n6264, n6265, n6266, n6267, n6268, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6304, n6305, n6306, n6307, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6332, n6333, n6335, 
      n6336, n6337, n6338, n6341, n6342, n6343, n6344, n6345, n6346, n6347, 
      n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, 
      n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, 
      n6368, n6369, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, 
      n6379, n6380, n6381, n6382, n6384, n6385, n6386, n6387, n6388, n6389, 
      n6390, n6391, n6392, n6393, n6394, n6396, n6397, n6398, n6399, n6400, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6429, n6430, n6431, n6432, 
      n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, 
      n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, 
      n6453, n6454, n6455, n6456, n6457, n6458, n6461, n6462, n6464, n6465, 
      n6466, n6467, n6468, n6469, n6472, n6474, n6476, n6477, n6478, n6479, 
      n6480, n6481, n6482, n6483, n6484, n6485, n6487, n6488, n6489, n6490, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6500, n6501, n6502, 
      n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, 
      n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, 
      n6524, n6526, n6527, n6528, n6530, n6531, n6532, n6533, n6534, n6535, 
      n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6545, n6546, 
      n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, 
      n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, 
      n6567, n6568, n6569, n6571, n6572, n6573, n6574, n6575, n6576, n6577, 
      n6578, n6579, n6580, n6581, n6582, n6584, n6585, n6586, n6587, n6588, 
      n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6599, n6600, 
      n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, 
      n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, 
      n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6631, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6642, n6643, n6644, 
      n6645, n6646, n6647, n6649, n6650, n6651, n6652, n6653, n6654, n6655, 
      n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, 
      n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, 
      n6677, n6678, n6679, n6680, n6681, n6683, n6685, n6686, n6687, n6688, 
      n6689, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, 
      n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, 
      n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, 
      n6721, n6722, n6723, n6724, n6725, n6727, n6728, n6729, n6730, n6731, 
      n6733, n6734, n6735, n6736, n6737, n6738, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6777, n6778, n6779, n6780, n6782, n6783, n6785, n6786, 
      n6787, n6788, n6789, n6790, n6793, n6794, n6795, n6796, n6797, n6798, 
      n6799, n6800, n6801, n6802, n6803, n6804, n6806, n6807, n6808, n6809, 
      n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, 
      n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, 
      n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, 
      n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, 
      n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, 
      n6860, n6861, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, 
      n6871, n6872, n6873, n6874, n6875, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, 
      n6892, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, 
      n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, 
      n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
      n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
      n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
      n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, 
      n6954, n6955, n6956, n6957, n6958, n6960, n6961, n6962, n6963, n6964, 
      n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, 
      n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, 
      n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, 
      n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, 
      n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7013, n7014, n7015, 
      n7016, n7017, n7018, n7020, n7021, n7022, n7023, n7024, n7025, n7026, 
      n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, 
      n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, 
      n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, 
      n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, 
      n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, 
      n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, 
      n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, 
      n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, 
      n7107, n7108, n7109, n7110, n7112, n7113, n7114, n7115, n7116, n7117, 
      n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, 
      n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, 
      n7138, n7139, n7140, n7141, n7142, n7143, n7145, n7146, n7147, n7148, 
      n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, 
      n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, 
      n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, 
      n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, 
      n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, 
      n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, 
      n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, 
      n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, 
      n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, 
      n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, 
      n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, 
      n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, 
      n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, 
      n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, 
      n7289, n7290, n7291, n7292, n7293, n7294, n7296, n7297, n7298, n7299, 
      n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, 
      n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, 
      n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, 
      n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, 
      n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, 
      n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7360, 
      n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, 
      n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, 
      n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, 
      n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, 
      n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, 
      n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7419, n7420, n7421, 
      n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, 
      n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, 
      n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7451, n7452, n7454, 
      n7456, n7457, n7458, n7459, n7460, n7461, n7463, n7464, n7465, n7466, 
      n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, 
      n7477, n7478, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, 
      n7488, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, 
      n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, 
      n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, 
      n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7528, n7529, 
      n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, 
      n7540, n7541, n7542, n7544, n7545, n7546, n7547, n7548, n7549, n7550, 
      n7551, n7552, n7553, n7554, n7555, n7556, n7558, n7559, n7560, n7561, 
      n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, 
      n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, 
      n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, 
      n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, 
      n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, 
      n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, 
      n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7630, n7631, n7632, 
      n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, 
      n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, 
      n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, 
      n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, 
      n7775, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, 
      n7786, n7787, n7788, n7789, n7790, n7792, n7793, n7794, n7795, n7796, 
      n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, 
      n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, 
      n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, 
      n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, 
      n7837, n7838, n7839, n7840, n7842, n7843, n7844, n7845, n7846, n7847, 
      n7848, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, 
      n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, 
      n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, 
      n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, 
      n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, 
      n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, 
      n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, 
      n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, 
      n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, 
      n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, 
      n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, 
      n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7970, 
      n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, 
      n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, 
      n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, 
      n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, 
      n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, 
      n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, 
      n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8094, 
      n8097, n8098, n8099, n8100, n8101, n8102, n8104, n8105, n8106, n8107, 
      n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, 
      n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, 
      n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, 
      n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, 
      n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, 
      n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, 
      n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, 
      n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, 
      n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, 
      n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, 
      n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, 
      n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, 
      n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, 
      n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, 
      n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, 
      n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, 
      n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, 
      n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, 
      n8288, n8289, n8290, n8291, n8292, n8293, n8296, n8297, n8298, n8299, 
      n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, 
      n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, 
      n8320, n8321, n8322, n8323, n8326, n8327, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8350, n8351, n8352, n8353, n8354, 
      n8355, n8356, n8357, n8359, n8360, n8361, n8362, n8364, n8365, n8366, 
      n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, 
      n8377, n8378, n8379, n8381, n8382, n8383, n8384, n8385, n8386, n8387, 
      n8388, n8389, n8390, n8391, n8392, n8393, n8395, n8396, n8397, n8398, 
      n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, 
      n8409, n8410, n8411, n8413, n8414, n8415, n8416, n8417, n8418, n8419, 
      n8420, n8421, n8422, n8423, n8424, n8426, n8427, n8428, n8430, n8431, 
      n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, 
      n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, 
      n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, 
      n8462, n8463, n8464, n8465, n8467, n8468, n8469, n8470, n8471, n8472, 
      n8473, n8474, n8475, n8476, n8477, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8523, n8524, 
      n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, 
      n8535, n8536, n8537, n8538, n8540, n8542, n8543, n8544, n8545, n8546, 
      n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, 
      n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, 
      n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, 
      n8577, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, 
      n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, 
      n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, 
      n8608, n8609, n8610, n8611, n8613, n8614, n8615, n8616, n8617, n8618, 
      n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, 
      n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, 
      n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, 
      n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, 
      n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, 
      n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, 
      n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, 
      n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, 
      n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, 
      n8709, n8710, n8711, n8712, n8713, n8715, n8716, n8717, n8718, n8719, 
      n8720, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, 
      n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, 
      n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, 
      n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, 
      n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, 
      n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8779, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
      n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, 
      n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
      n8814, n8815, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, 
      n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, 
      n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, 
      n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, 
      n8855, n8856, n8857, n8859, n8860, n8861, n8862, n8863, n8864, n8865, 
      n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, 
      n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, 
      n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, 
      n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, 
      n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, 
      n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
      n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, 
      n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, 
      n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, 
      n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
      n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
      n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, 
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9044, n9045, n9046, 
      n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, 
      n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, 
      n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, 
      n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, 
      n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, 
      n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, 
      n9107, n9108, n9109, n9111, n9112, n9113, n9114, n9115, n9116, n9117, 
      n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, 
      n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, 
      n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, 
      n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, 
      n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, 
      n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, 
      n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
      n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
      n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, 
      n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, 
      n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, 
      n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, 
      n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, 
      n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9256, n9257, n9258, 
      n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, 
      n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, 
      n9279, n9280, n9281, n9282, n9283, n9285, n9286, n9287, n9288, n9289, 
      n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, 
      n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, 
      n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, 
      n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, 
      n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, 
      n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, 
      n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, 
      n9360, n9361, n9362, n9363, n9364, n9365, n9368, n9369, n9370, n9372, 
      n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, 
      n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, 
      n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, 
      n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9412, n9413, 
      n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, 
      n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, 
      n9434, n9435, n9436, n9437, n9438, n9440, n9441, n9442, n9443, n9444, 
      n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, 
      n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, 
      n9465, n9466, n9467, n9469, n9470, n9471, n9472, n9473, n9474, n9475, 
      n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, 
      n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, 
      n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, 
      n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, 
      n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, 
      n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9535, n9536, 
      n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, 
      n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, 
      n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, 
      n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, 
      n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, 
      n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, 
      n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, 
      n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, 
      n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, 
      n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, 
      n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, 
      n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, 
      n9657, n9658, n9659, n9660, n9661, n9663, n9664, n9665, n9666, n9667, 
      n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, 
      n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, 
      n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, 
      n9698, n9699, n9700, n9701, n9702, n9703, n9705, n9706, n9707, n9708, 
      n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, 
      n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, 
      n9729, n9730, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, 
      n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, 
      n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, 
      n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, 
      n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, 
      n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, 
      n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, 
      n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, 
      n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, 
      n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, 
      n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, 
      n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, 
      n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, 
      n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, 
      n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, 
      n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, 
      n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, 
      n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, 
      n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, 
      n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, 
      n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, 
      n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, 
      n9950, n9951, n9952, n9954, n9955, n9956, n9957, n9958, n9959, n9960, 
      n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, 
      n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, 
      n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, 
      n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, 
      n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, 
      n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, 
      n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, 
      n10028, n10029, n10030, n10031, n10033, n10034, n10035, n10036, n10037, 
      n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, 
      n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, 
      n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, 
      n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, 
      n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, 
      n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10092, 
      n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, 
      n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, 
      n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, 
      n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, 
      n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, 
      n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, 
      n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, 
      n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, 
      n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, 
      n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, 
      n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, 
      n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, 
      n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, 
      n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, 
      n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, 
      n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, 
      n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, 
      n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, 
      n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, 
      n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, 
      n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10282, 
      n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, 
      n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, 
      n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, 
      n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, 
      n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, 
      n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, 
      n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, 
      n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, 
      n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, 
      n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, 
      n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, 
      n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, 
      n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, 
      n10400, n10401, n10402, n10403, n10406, n10407, n10408, n10409, n10411, 
      n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, 
      n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, 
      n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, 
      n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, 
      n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, 
      n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, 
      n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, 
      n10475, n10476, n10477, n10478, n10479, n10480, n10482, n10484, n10485, 
      n10486, n10487, n10488, n10489, n10490, n10492, n10494, n10495, n10496, 
      n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, 
      n10506, n10507, n10508, n10509, n10511, n10512, n10515, n10516, n10517, 
      n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, 
      n10527, n10528, n10530, n10531, n10532, n10533, n10534, n10535, n10536, 
      n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, 
      n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, 
      n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10563, n10564, 
      n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, 
      n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, 
      n10583, n10584, n10585, n10586, n10587, n10589, n10590, n10591, n10592, 
      n10593, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, 
      n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10611, n10612, 
      n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, 
      n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, 
      n10633, n10634, n10635, n10637, n10638, n10639, n10640, n10641, n10642, 
      n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, 
      n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, 
      n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, 
      n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, 
      n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, 
      n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, 
      n10697, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, 
      n10707, n10708, n10710, n10711, n10712, n10713, n10714, n10715, n10716, 
      n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, 
      n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, 
      n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10744, 
      n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, 
      n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, 
      n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, 
      n10772, n10773, n10775, n10776, n10777, n10778, n10779, n10780, n10781, 
      n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, 
      n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, 
      n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, 
      n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, 
      n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, 
      n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, 
      n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, 
      n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, 
      n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, 
      n10863, n10864, n10865, n10867, n10868, n10869, n10870, n10871, n10872, 
      n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, 
      n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, 
      n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, 
      n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, 
      n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, 
      n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, 
      n10928, n10929, n10930, n10931, n10932, n10933, n10935, n10936, n10937, 
      n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, 
      n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, 
      n10956, n10957, n10958, n10959, n10961, n10962, n10963, n10964, n10965, 
      n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, 
      n10976, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, 
      n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, 
      n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, 
      n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, 
      n11013, n11014, n11015, n11016, n11018, n11019, n11020, n11021, n11022, 
      n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, 
      n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, 
      n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, 
      n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, 
      n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, 
      n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, 
      n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, 
      n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, 
      n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, 
      n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, 
      n11114, n11115, n11116, n11118, n11119, n11120, n11121, n11122, n11123, 
      n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, 
      n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11142, 
      n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, 
      n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, 
      n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, 
      n11170, n11171, n11172, n11174, n11175, n11176, n11178, n11179, n11180, 
      n11181, n11183, n11184, n11185, n11186, n11187, n11188, n11190, n11191, 
      n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, 
      n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, 
      n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, 
      n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, 
      n11228, n11229, n11231, n11232, n11233, n11234, n11235, n11236, n11237, 
      n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, 
      n11248, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, 
      n11258, n11259, n11260, n11261, n11262, n11264, n11265, n11266, n11267, 
      n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, 
      n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, 
      n11287, n11288, n11289, n11290, n11291, n11292, n11294, n11295, n11296, 
      n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, 
      n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, 
      n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, 
      n11324, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
      n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, 
      n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, 
      n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, 
      n11361, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, 
      n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, 
      n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, 
      n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, 
      n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, 
      n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, 
      n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, 
      n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, 
      n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, 
      n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, 
      n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, 
      n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, 
      n11470, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, 
      n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, 
      n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, 
      n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, 
      n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, 
      n11517, n11518, n11520, n11521, n11522, n11523, n11524, n11525, n11526, 
      n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, 
      n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, 
      n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, 
      n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, 
      n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, 
      n11572, n11573, n11574, n11575, n11577, n11578, n11579, n11580, n11581, 
      n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, 
      n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, 
      n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, 
      n11609, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, 
      n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, 
      n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, 
      n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, 
      n11647, n11648, n11650, n11652, n11653, n11654, n11655, n11656, n11657, 
      n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, 
      n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, 
      n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, 
      n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, 
      n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, 
      n11703, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, 
      n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, 
      n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, 
      n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, 
      n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, 
      n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, 
      n11758, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, 
      n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, 
      n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, 
      n11786, n11787, n11789, n11790, n11791, n11792, n11793, n11794, n11795, 
      n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, 
      n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, 
      n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, 
      n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11831, n11832, 
      n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11841, n11843, 
      n11844, n11845, n11846, n11848, n11849, n11850, n11851, n11852, n11853, 
      n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, 
      n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, 
      n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, 
      n11882, n11883, n11884, n11886, n11887, n11888, n11889, n11890, n11891, 
      n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, 
      n11901, n11902, n11903, n11904, n11905, n11907, n11908, n11909, n11911, 
      n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, 
      n11921, n11922, n11924, n11925, n11926, n11927, n11928, n11929, n11930, 
      n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, 
      n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, 
      n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, 
      n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, 
      n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, 
      n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, 
      n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, 
      n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, 
      n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, 
      n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, 
      n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, 
      n12031, n12032, n12033, n12034, n12035, n12037, n12039, n12040, n12041, 
      n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, 
      n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12060, 
      n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, 
      n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, 
      n12079, n12080, n12081, n12083, n12085, n12086, n12087, n12088, n12089, 
      n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, 
      n12099, n12100, n12101, n12102, n12103, n12104, n12106, n12107, n12109, 
      n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, 
      n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, 
      n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, 
      n12137, n12138, n12139, n12140, n12142, n12143, n12144, n12145, n12146, 
      n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, 
      n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, 
      n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, 
      n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, 
      n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, 
      n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, 
      n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, 
      n12211, n12212, n12213, n12214, n12215, n12216, n12218, n12219, n12220, 
      n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, 
      n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, 
      n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, 
      n12248, n12249, n12250, n12251, n12252, n12253, n12255, n12256, n12257, 
      n12258, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, 
      n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, 
      n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, 
      n12286, n12287, n12288, n12289, n12290, n12291, n12293, n12294, n12295, 
      n12296, n12297, n12298, n12299, n12300, n12302, n12303, n12304, n12305, 
      n12306, n12307, n12308, n12309, n12310, n12312, n12313, n12314, n12315, 
      n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, 
      n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, 
      n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12343, 
      n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, 
      n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, 
      n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, 
      n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, 
      n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, 
      n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, 
      n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, 
      n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, 
      n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, 
      n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, 
      n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, 
      n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, 
      n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, 
      n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, 
      n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, 
      n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, 
      n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, 
      n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, 
      n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, 
      n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, 
      n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, 
      n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12542, n12543, 
      n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, 
      n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, 
      n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, 
      n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, 
      n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, 
      n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, 
      n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, 
      n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, 
      n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, 
      n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, 
      n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, 
      n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, 
      n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, 
      n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, 
      n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, 
      n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, 
      n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, 
      n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, 
      n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, 
      n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, 
      n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, 
      n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, 
      n12742, n12743, n12744, n12746, n12747, n12748, n12749, n12750, n12751, 
      n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12760, n12761, 
      n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, 
      n12771, n12772, n12773, n12775, n12776, n12777, n12778, n12779, n12780, 
      n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, 
      n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, 
      n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, 
      n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, 
      n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, 
      n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, 
      n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, 
      n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, 
      n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, 
      n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, 
      n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, 
      n12880, n12881, n12882, n12883, n12884, n12885, n12887, n12888, n12889, 
      n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, 
      n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12907, n12908, 
      n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, 
      n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, 
      n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, 
      n12936, n12938, n12939, n12940, n12941, n12943, n12944, n12945, n12946, 
      n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, 
      n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, 
      n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, 
      n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, 
      n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, 
      n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, 
      n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, 
      n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, 
      n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, 
      n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, 
      n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, 
      n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, 
      n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, 
      n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, 
      n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, 
      n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, 
      n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, 
      n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, 
      n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, 
      n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, 
      n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, 
      n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, 
      n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, 
      n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, 
      n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, 
      n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, 
      n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, 
      n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, 
      n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, 
      n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, 
      n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, 
      n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, 
      n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, 
      n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, 
      n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, 
      n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, 
      n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, 
      n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, 
      n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, 
      n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, 
      n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, 
      n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, 
      n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, 
      n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, 
      n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, 
      n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, 
      n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, 
      n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, 
      n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, 
      n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, 
      n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, 
      n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, 
      n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, 
      n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, 
      n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, 
      n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, 
      n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, 
      n13460, n13461, n13462, n13464, n13465, n13466, n13467, n13468, n13469, 
      n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, 
      n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, 
      n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, 
      n13497, n13498, n13499, n13501, n13502, n13503, n13504, n13505, n13506, 
      n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, 
      n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, 
      n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, 
      n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, 
      n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, 
      n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, 
      n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, 
      n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, 
      n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, 
      n13589, n13590, n13592, n13593, n13594, n13595, n13596, n13597, n13598, 
      n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, 
      n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, 
      n13617, n13618, n13620, n13621, n13624, n13625, n13626, n13627, n13628, 
      n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, 
      n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, 
      n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, 
      n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, 
      n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, 
      n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, 
      n13683, n13684, n13685, n13686, n13687, n13688, n13692, n13693, n13694, 
      n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, 
      n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, 
      n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13722, 
      n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13732, 
      n13733, n13734, n13735, n13736, n13739, n13740, n13741, n13742, n13743, 
      n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, 
      n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, 
      n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, 
      n13771, n13772, n13773, n13774, n13775, n13776, n13778, n13779, n13781, 
      n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, 
      n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, 
      n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, 
      n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, 
      n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, 
      n13827, n13828, n13829, n13830, n13831, n13832, n13834, n13835, n13836, 
      n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, 
      n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13854, n13855, 
      n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, 
      n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, 
      n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, 
      n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, 
      n13892, n13893, n13894, n13898, n13900, n13901, n13902, n13903, n13904, 
      n13905, n13906, n13907, n13908, n13909, n13910, n13912, n13913, n13914, 
      n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, 
      n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, 
      n13933, n13934, n13935, n13936, n13938, n13939, n13940, n13941, n13943, 
      n13944, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, 
      n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, 
      n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, 
      n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, 
      n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, 
      n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, 
      n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, 
      n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, 
      n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, 
      n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, 
      n14035, n14036, n14037, n14038, n14039, n14041, n14042, n14043, n14044, 
      n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, 
      n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14063, 
      n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, 
      n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, 
      n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, 
      n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, 
      n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, 
      n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, 
      n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, 
      n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, 
      n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, 
      n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, 
      n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, 
      n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, 
      n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14181, 
      n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, 
      n14191, n14192, n14193, n14194, n14195, n14197, n14198, n14199, n14200, 
      n14202, n14203, n14204, n14206, n14207, n14208, n14209, n14210, n14211, 
      n14212, n14213, n14214, n14215, n14216, n14217, n14219, n14220, n14221, 
      n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, 
      n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, 
      n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, 
      n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, 
      n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, 
      n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, 
      n14276, n14277, n14278, n14281, n14282, n14283, n14284, n14285, n14286, 
      n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, 
      n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, 
      n14305, n14306, n14309, n14310, n14311, n14312, n14313, n14314, n14315, 
      n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, 
      n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, 
      n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, 
      n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, 
      n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, 
      n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, 
      n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, 
      n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, 
      n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14397, n14398, 
      n14399, n14400, n14401, n14402, n14403, n14405, n14406, n14407, n14408, 
      n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, 
      n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, 
      n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, 
      n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, 
      n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14455, 
      n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, 
      n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, 
      n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, 
      n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, 
      n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14500, n14501, 
      n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14511, 
      n14512, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, 
      n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, 
      n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, 
      n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, 
      n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, 
      n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, 
      n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, 
      n14576, n14577, n14578, n14580, n14581, n14582, n14583, n14584, n14585, 
      n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, 
      n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, 
      n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, 
      n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14621, n14622, 
      n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, 
      n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, 
      n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, 
      n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, 
      n14659, n14660, n14662, n14663, n14664, n14665, n14666, n14667, n14668, 
      n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, 
      n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, 
      n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, 
      n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, 
      n14706, n14707, n14709, n14710, n14711, n14712, n14713, n14714, n14715, 
      n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, 
      n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, 
      n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, 
      n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, 
      n14753, n14754, n14756, n14757, n14758, n14759, n14760, n14761, n14762, 
      n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, 
      n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, 
      n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, 
      n14790, n14791, n14792, n14793, n14794, n14796, n14797, n14798, n14799, 
      n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, 
      n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, 
      n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, 
      n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, 
      n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, 
      n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, 
      n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, 
      n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, 
      n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, 
      n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, 
      n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, 
      n14899, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, 
      n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, 
      n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14927, 
      n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, 
      n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, 
      n14946, n14947, n14948, n14949, n14951, n14952, n14953, n14954, n14955, 
      n14956, n14957, n14958, n14960, n14961, n14962, n14963, n14964, n14966, 
      n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, 
      n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, 
      n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, 
      n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, 
      n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, 
      n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, 
      n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, 
      n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, 
      n15040, n15041, n15042, n15043, n15044, n15046, n15047, n15051, n15052, 
      n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, 
      n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, 
      n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, 
      n15080, n15081, n15082, n15083, n15084, n15085, n15087, n15088, n15089, 
      n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, 
      n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, 
      n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, 
      n15117, n15118, n15119, n15120, n15123, n15124, n15125, n15126, n15127, 
      n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, 
      n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, 
      n15146, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, 
      n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15164, n15165, 
      n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, 
      n15175, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, 
      n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, 
      n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, 
      n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15212, 
      n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, 
      n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, 
      n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, 
      n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, 
      n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, 
      n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, 
      n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, 
      n15276, n15277, n15278, n15279, n15280, n15281, n15284, n15285, n15286, 
      n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, 
      n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, 
      n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, 
      n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, 
      n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, 
      n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, 
      n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, 
      n15350, n15351, n15352, n15353, n15354, n15355, n15357, n15358, n15359, 
      n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, 
      n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, 
      n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, 
      n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, 
      n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, 
      n15405, n15406, n15407, n15409, n15410, n15411, n15412, n15413, n15414, 
      n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, 
      n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, 
      n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, 
      n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, 
      n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, 
      n15460, n15461, n15462, n15463, n15464, n15466, n15467, n15468, n15469, 
      n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, 
      n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, 
      n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, 
      n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, 
      n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, 
      n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, 
      n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, 
      n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, 
      n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, 
      n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, 
      n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, 
      n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, 
      n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, 
      n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, 
      n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, 
      n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, 
      n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, 
      n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, 
      n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, 
      n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, 
      n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, 
      n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, 
      n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, 
      n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, 
      n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, 
      n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, 
      n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, 
      n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, 
      n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, 
      n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, 
      n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, 
      n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, 
      n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, 
      n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, 
      n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, 
      n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, 
      n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, 
      n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, 
      n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, 
      n15822, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, 
      n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, 
      n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, 
      n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, 
      n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, 
      n15868, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, 
      n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, 
      n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, 
      n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, 
      n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, 
      n15914, n15915, n15916, n15917, n15918, n15920, n15922, n15923, n15924, 
      n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, 
      n15934, n15935, n15936, n15938, n15939, n15940, n15941, n15942, n15943, 
      n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, 
      n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, 
      n15962, n15963, n15965, n15966, n15967, n15968, n15969, n15970, n15971, 
      n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, 
      n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, 
      n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, 
      n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, 
      n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, 
      n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16026, 
      n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, 
      n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, 
      n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, 
      n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, 
      n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, 
      n16072, n16073, n16074, n16076, n16077, n16078, n16079, n16080, n16081, 
      n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, 
      n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, 
      n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, 
      n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, 
      n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, 
      n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, 
      n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, 
      n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16154, 
      n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, 
      n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, 
      n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, 
      n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, 
      n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, 
      n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, 
      n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, 
      n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, 
      n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, 
      n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, 
      n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, 
      n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, 
      n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, 
      n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, 
      n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, 
      n16290, n16291, n16293, n16294, n16295, n16296, n16297, n16298, n16299, 
      n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, 
      n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, 
      n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, 
      n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, 
      n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, 
      n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, 
      n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, 
      n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, 
      n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, 
      n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, 
      n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, 
      n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, 
      n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, 
      n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, 
      n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, 
      n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, 
      n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, 
      n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, 
      n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, 
      n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, 
      n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, 
      n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, 
      n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, 
      n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, 
      n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, 
      n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, 
      n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, 
      n16543, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, 
      n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, 
      n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, 
      n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, 
      n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, 
      n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, 
      n16598, n16599, n16601, n16602, n16603, n16604, n16605, n16606, n16607, 
      n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, 
      n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, 
      n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, 
      n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, 
      n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, 
      n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, 
      n16662, n16663, n16664, n16665, n16667, n16668, n16669, n16670, n16671, 
      n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, 
      n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, 
      n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, 
      n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, 
      n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, 
      n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, 
      n16727, n16728, n16729, n16730, n16732, n16733, n16734, n16735, n16736, 
      n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, 
      n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, 
      n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, 
      n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, 
      n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, 
      n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, 
      n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, 
      n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16809, n16810, 
      n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, 
      n16820, n16821, n16822, n16823, n16824, n16825, n16828, n16829, n16830, 
      n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16839, n16840, 
      n16841, n16842, n16843, n16844, n16845, n16846, n16848, n16849, n16850, 
      n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, 
      n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, 
      n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, 
      n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, 
      n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, 
      n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, 
      n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, 
      n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, 
      n16925, n16926, n16927, n16928, n16929, n16930, n16932, n16933, n16934, 
      n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, 
      n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, 
      n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, 
      n16962, n16964, n16965, n16966, n16968, n16969, n16970, n16971, n16972, 
      n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, 
      n16982, n16983, n16985, n16986, n16987, n16988, n16990, n16991, n16992, 
      n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, 
      n17002, n17003, n17004, n17005, n17006, n17008, n17009, n17010, n17011, 
      n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, 
      n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17029, n17030, 
      n17031, n17033, n17035, n17036, n17037, n17038, n17039, n17040, n17041, 
      n17042, n17043, n17044, n17045, n17046, n17047, n17049, n17051, n17052, 
      n17053, n17054, n17055, n17057, n17058, n17059, n17060, n17061, n17062, 
      n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, 
      n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, 
      n17081, n17082, n17083, n17084, n17085, n17087, n17088, n17089, n17090, 
      n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17101, 
      n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, 
      n17111, n17112, n17113, n17116, n17117, n17118, n17119, n17120, n17121, 
      n17122, n17123, n17124, n17125, n17126, n17128, n17129, n17130, n17131, 
      n17132, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, 
      n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, 
      n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, 
      n17161, n17162, n17164, n17165, n17166, n17167, n17169, n17170, n17171, 
      n17172, n17173, n17175, n17176, n17177, n17178, n17179, n17180, n17181, 
      n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, 
      n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, 
      n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, 
      n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, 
      n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, 
      n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, 
      n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, 
      n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, 
      n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, 
      n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, 
      n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, 
      n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, 
      n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, 
      n17301, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, 
      n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, 
      n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17329, n17330, 
      n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, 
      n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, 
      n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, 
      n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, 
      n17368, n17369, n17370, n17371, n17372, n17374, n17375, n17376, n17377, 
      n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, 
      n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, 
      n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, 
      n17406, n17407, n17408, n17410, n17411, n17412, n17413, n17414, n17415, 
      n17416, n17417, n17418, n17419, n17421, n17422, n17423, n17424, n17425, 
      n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, 
      n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, 
      n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, 
      n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, 
      n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, 
      n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, 
      n17480, n17481, n17482, n17484, n17485, n17486, n17487, n17488, n17489, 
      n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, 
      n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, 
      n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, 
      n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17526, 
      n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, 
      n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, 
      n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, 
      n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, 
      n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, 
      n17572, n17573, n17574, n17575, n17577, n17578, n17579, n17580, n17581, 
      n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, 
      n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, 
      n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, 
      n17610, n17611, n17613, n17614, n17615, n17616, n17617, n17618, n17619, 
      n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, 
      n17629, n17630, n17631, n17632, n17635, n17636, n17637, n17638, n17639, 
      n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, 
      n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, 
      n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, 
      n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, 
      n17680, n17681, n17682, n17683, n17684, n17686, n17687, n17688, n17689, 
      n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17699, 
      n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, 
      n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, 
      n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, 
      n17727, n17728, n17729, n17730, n17731, n17732, n17734, n17735, n17736, 
      n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, 
      n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, 
      n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, 
      n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, 
      n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, 
      n17782, n17783, n17785, n17788, n17789, n17792, n17793, n17794, n17795, 
      n17796, n17797, n17798, n17799, n17801, n17802, n17803, n17804, n17808, 
      n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, 
      n17818, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, 
      n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, 
      n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, 
      n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, 
      n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, 
      n17864, n17865, n17866, n17868, n17869, n17870, n17871, n17872, n17873, 
      n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, 
      n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, 
      n17892, n17893, n17895, n17896, n17897, n17898, n17899, n17900, n17902, 
      n17903, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, 
      n17913, n17915, n17916, n17917, n17918, n17919, n17920, n17922, n17923, 
      n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, 
      n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, 
      n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, 
      n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, 
      n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, 
      n17969, n17970, n17972, n17973, n17974, n17975, n17976, n17977, n17978, 
      n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, 
      n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, 
      n17997, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, 
      n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18015, n18016, 
      n18017, n18018, n18019, n18020, n18022, n18023, n18024, n18025, n18027, 
      n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, 
      n18037, n18038, n18039, n18040, n18042, n18043, n18044, n18045, n18046, 
      n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, 
      n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, 
      n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, 
      n18074, n18075, n18076, n18078, n18079, n18080, n18081, n18082, n18083, 
      n18084, n18085, n18086, n18087, n18088, n18090, n18091, n18092, n18093, 
      n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18103, 
      n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, 
      n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, 
      n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, 
      n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, 
      n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, 
      n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, 
      n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, 
      n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, 
      n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, 
      n18187, n18188, n18189, n18190, n18191, n18193, n18194, n18195, n18196, 
      n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, 
      n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, 
      n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, 
      n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, 
      n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, 
      n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, 
      n18251, n18252, n18253, n18254, n18256, n18257, n18258, n18259, n18260, 
      n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, 
      n18270, n18271, n18273, n18274, n18275, n18276, n18277, n18278, n18279, 
      n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18289, 
      n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, 
      n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, 
      n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, 
      n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, 
      n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, 
      n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, 
      n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, 
      n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, 
      n18363, n18364, n18365, n18366, n18367, n18369, n18370, n18371, n18372, 
      n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, 
      n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, 
      n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, 
      n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, 
      n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, 
      n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, 
      n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, 
      n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, 
      n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, 
      n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, 
      n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, 
      n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, 
      n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, 
      n18490, n18491, n18492, n18493, n18495, n18496, n18497, n18498, n18499, 
      n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, 
      n18509, n18510, n18511, n18512, n18513, n18514, n18516, n18517, n18518, 
      n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, 
      n18528, n18529, n18530, n18534, n18535, n18536, n18537, n18538, n18539, 
      n18540, n18541, n18543, n18544, n18545, n18546, n18547, n18548, n18549, 
      n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, 
      n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, 
      n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18576, n18577, 
      n18578, n18579, n18581, n18582, n18583, n18584, n18585, n18586, n18587, 
      n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, 
      n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, 
      n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, 
      n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, 
      n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, 
      n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, 
      n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, 
      n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18660, 
      n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, 
      n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, 
      n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, 
      n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, 
      n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, 
      n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, 
      n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, 
      n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, 
      n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, 
      n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, 
      n18751, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, 
      n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, 
      n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, 
      n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, 
      n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, 
      n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, 
      n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, 
      n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, 
      n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18833, 
      n18834, n18835, n18836, n18837, n18838, n18840, n18841, n18842, n18843, 
      n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, 
      n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, 
      n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, 
      n18871, n18872, n18873, n18875, n18876, n18877, n18878, n18879, n18880, 
      n18881, n18882, n18884, n18885, n18886, n18887, n18888, n18889, n18890, 
      n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, 
      n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, 
      n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, 
      n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, 
      n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, 
      n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, 
      n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, 
      n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, 
      n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, 
      n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, 
      n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, 
      n18990, n18991, n18992, n18994, n18995, n18996, n18997, n18998, n18999, 
      n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, 
      n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, 
      n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, 
      n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, 
      n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, 
      n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19054, 
      n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, 
      n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, 
      n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, 
      n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, 
      n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, 
      n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, 
      n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, 
      n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, 
      n19127, n19128, n19130, n19131, n19132, n19133, n19134, n19135, n19136, 
      n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, 
      n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, 
      n19155, n19156, n19157, n19158, n19160, n19161, n19162, n19163, n19164, 
      n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, 
      n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, 
      n19183, n19184, n19185, n19187, n19188, n19191, n19192, n19193, n19194, 
      n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, 
      n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19212, n19213, 
      n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, 
      n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, 
      n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, 
      n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, 
      n19250, n19251, n19252, n19254, n19256, n19257, n19258, n19259, n19261, 
      n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, 
      n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, 
      n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, 
      n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, 
      n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, 
      n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, 
      n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, 
      n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, 
      n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, 
      n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, 
      n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19361, 
      n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, 
      n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, 
      n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, 
      n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, 
      n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, 
      n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, 
      n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, 
      n19425, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, 
      n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, 
      n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, 
      n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, 
      n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, 
      n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, 
      n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, 
      n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, 
      n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, 
      n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, 
      n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, 
      n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, 
      n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, 
      n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, 
      n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, 
      n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, 
      n19570, n19571, n19572, n19573, n19574, n19575, n19577, n19578, n19579, 
      n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, 
      n19589, n19590, n19591, n19592, n19593, n19595, n19596, n19597, n19598, 
      n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, 
      n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, 
      n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, 
      n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, 
      n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, 
      n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, 
      n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, 
      n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, 
      n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, 
      n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19690, 
      n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, 
      n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, 
      n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, 
      n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, 
      n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, 
      n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, 
      n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, 
      n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, 
      n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, 
      n19772, n19773, n19774, n19775, n19777, n19778, n19779, n19780, n19781, 
      n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, 
      n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, 
      n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, 
      n19809, n19810, n19811, n19813, n19814, n19815, n19816, n19817, n19818, 
      n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, 
      n19828, n19829, n19830, n19832, n19833, n19834, n19836, n19837, n19838, 
      n19839, n19841, n19842, n19843, n19844, n19846, n19848, n19849, n19850, 
      n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, 
      n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, 
      n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, 
      n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, 
      n19887, n19888, n19889, n19890, n19891, n19893, n19894, n19895, n19896, 
      n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19906, 
      n19907, n19908, n19909, n19911, n19912, n19914, n19915, n19916, n19917, 
      n19918, n19919, n19920, n19921, n19923, n19924, n19925, n19926, n19927, 
      n19928, n19930, n19931, n19935, n19936, n19937, n19938, n19939, n19940, 
      n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, 
      n19950, n19951, n19952, n19953, n19955, n19956, n19957, n19958, n19959, 
      n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, 
      n19969, n19970, n19972, n19973, n19974, n19975, n19976, n19977, n19978, 
      n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19987, n19988, 
      n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, 
      n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, 
      n20007, n20008, n20010, n20011, n20012, n20013, n20014, n20015, n20016, 
      n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, 
      n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20035, 
      n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, 
      n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, 
      n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, 
      n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, 
      n20072, n20073, n20074, n20075, n20077, n20078, n20079, n20081, n20082, 
      n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, 
      n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, 
      n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, 
      n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, 
      n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, 
      n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20136, n20137, 
      n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, 
      n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20155, n20156, 
      n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, 
      n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, 
      n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, 
      n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, 
      n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, 
      n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, 
      n20211, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20221, 
      n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, 
      n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, 
      n20240, n20241, n20242, n20243, n20244, n20246, n20247, n20248, n20249, 
      n20250, n20251, n20252, n20254, n20255, n20256, n20257, n20258, n20259, 
      n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20268, n20269, 
      n20270, n20271, n20272, n20273, n20275, n20276, n20277, n20278, n20279, 
      n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, 
      n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, 
      n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, 
      n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, 
      n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, 
      n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, 
      n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20342, n20343, 
      n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, 
      n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, 
      n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, 
      n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20379, n20380, 
      n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, 
      n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, 
      n20400, n20401, n20402, n20404, n20405, n20406, n20407, n20408, n20409, 
      n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, 
      n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, 
      n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, 
      n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, 
      n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, 
      n20455, n20456, n20457, n20458, n20459, n20460, n20462, n20463, n20464, 
      n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, 
      n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, 
      n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, 
      n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, 
      n20501, n20502, n20503, n20504, n20506, n20507, n20508, n20509, n20510, 
      n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20520, 
      n20521, n20522, n20523, n20524, n20526, n20527, n20528, n20529, n20530, 
      n20531, n20532, n20533, n20534, n20535, n20537, n20539, n20541, n20542, 
      n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, 
      n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, 
      n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20570, 
      n20571, n20572, n20573, n20574, n20575, n20577, n20578, n20579, n20580, 
      n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, 
      n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, 
      n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, 
      n20609, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, 
      n20619, n20620, n20621, n20622, n20623, n20625, n20626, n20627, n20628, 
      n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, 
      n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, 
      n20647, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, 
      n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, 
      n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, 
      n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, 
      n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, 
      n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, 
      n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, 
      n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, 
      n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, 
      n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, 
      n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, 
      n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, 
      n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, 
      n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, 
      n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, 
      n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20793, 
      n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, 
      n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, 
      n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, 
      n20821, n20822, n20823, n20824, n20825, n20827, n20828, n20829, n20830, 
      n20831, n20832, n20833, n20835, n20836, n20837, n20838, n20839, n20840, 
      n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, 
      n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, 
      n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, 
      n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, 
      n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, 
      n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, 
      n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, 
      n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, 
      n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, 
      n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, 
      n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, 
      n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, 
      n20950, n20951, n20953, n20954, n20955, n20956, n20957, n20958, n20959, 
      n20960, n20961, n20963, n20964, n20965, n20966, n20967, n20968, n20969, 
      n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, 
      n20979, n20980, n20982, n20983, n20984, n20985, n20986, n20987, n20988, 
      n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, 
      n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, 
      n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, 
      n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, 
      n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, 
      n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, 
      n21044, n21045, n21047, n21050, n21051, n21052, n21053, n21054, n21055, 
      n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, 
      n21065, n21066, n21067, n21068, n21069, n21071, n21072, n21073, n21074, 
      n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, 
      n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, 
      n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21101, n21102, 
      n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, 
      n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, 
      n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, 
      n21131, n21132, n21133, n21134, n21135, n21137, n21138, n21139, n21140, 
      n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, 
      n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, 
      n21159, n21161, n21162, n21163, n21165, n21166, n21167, n21168, n21169, 
      n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, 
      n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, 
      n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, 
      n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, 
      n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, 
      n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, 
      n21225, n21226, n21227, n21228, n21230, n21231, n21232, n21233, n21234, 
      n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, 
      n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, 
      n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, 
      n21262, n21263, n21265, n21266, n21267, n21268, n21269, n21270, n21271, 
      n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, 
      n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, 
      n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, 
      n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, 
      n21308, n21309, n21311, n21312, n21313, n21314, n21315, n21316, n21317, 
      n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, 
      n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, 
      n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, 
      n21345, n21346, n21347, n21348, n21349, n21351, n21352, n21353, n21354, 
      n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, 
      n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, 
      n21373, n21374, n21375, n21376, n21378, n21379, n21380, n21381, n21382, 
      n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, 
      n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, 
      n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, 
      n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, 
      n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, 
      n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, 
      n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, 
      n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, 
      n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, 
      n21465, n21467, n21469, n21470, n21471, n21472, n21473, n21474, n21475, 
      n21476, n21477, n21478, n21479, n21480, n21481, n21483, n21484, n21485, 
      n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, 
      n21495, n21496, n21497, n21499, n21500, n21501, n21503, n21504, n21505, 
      n21506, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, 
      n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, 
      n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, 
      n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, 
      n21543, n21544, n21545, n21546, n21547, n21549, n21550, n21551, n21552, 
      n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, 
      n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, 
      n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, 
      n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, 
      n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, 
      n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21607, 
      n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, 
      n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, 
      n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, 
      n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, 
      n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, 
      n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, 
      n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21671, 
      n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, 
      n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, 
      n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, 
      n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21708, 
      n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, 
      n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, 
      n21727, n21728, n21729, n21731, n21732, n21733, n21734, n21735, n21736, 
      n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, 
      n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, 
      n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, 
      n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, 
      n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, 
      n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, 
      n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, 
      n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, 
      n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, 
      n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, 
      n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, 
      n21836, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, 
      n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, 
      n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21864, 
      n21865, n21866, n21867, n21868, n21870, n21871, n21872, n21873, n21874, 
      n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, 
      n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, 
      n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, 
      n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, 
      n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, 
      n21920, n21921, n21922, n21924, n21925, n21926, n21927, n21928, n21929, 
      n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, 
      n21939, n21940, n21941, n21942, n21943, n21944, n21946, n21947, n21948, 
      n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, 
      n21958, n21959, n21960, n21961, n21962, n21963, n21966, n21967, n21968, 
      n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, 
      n21978, n21979, n21980, n21982, n21983, n21984, n21985, n21986, n21987, 
      n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, 
      n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, 
      n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, 
      n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, 
      n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, 
      n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, 
      n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, 
      n22052, n22053, n22055, n22056, n22057, n22058, n22059, n22060, n22061, 
      n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, 
      n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, 
      n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22088, n22089, 
      n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, 
      n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, 
      n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, 
      n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, 
      n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, 
      n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, 
      n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, 
      n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, 
      n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, 
      n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, 
      n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, 
      n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, 
      n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, 
      n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, 
      n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, 
      n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, 
      n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, 
      n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, 
      n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, 
      n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, 
      n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, 
      n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, 
      n22288, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, 
      n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, 
      n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, 
      n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, 
      n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, 
      n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, 
      n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, 
      n22352, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, 
      n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, 
      n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, 
      n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, 
      n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, 
      n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, 
      n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, 
      n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, 
      n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, 
      n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, 
      n22443, n22444, n22445, n22446, n22448, n22449, n22450, n22451, n22452, 
      n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, 
      n22462, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, 
      n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, 
      n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, 
      n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, 
      n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, 
      n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, 
      n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, 
      n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, 
      n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, 
      n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, 
      n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, 
      n22562, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, 
      n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, 
      n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, 
      n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, 
      n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, 
      n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, 
      n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, 
      n22626, n22627, n22628, n22629, n22630, n22631, n22633, n22634, n22635, 
      n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, 
      n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, 
      n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, 
      n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, 
      n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, 
      n22681, n22682, n22683, n22684, n22685, n22686, n22688, n22689, n22690, 
      n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, 
      n22701, n22702, n22703, n22705, n22706, n22707, n22708, n22709, n22710, 
      n22711, n22712, n22713, n22714, n22715, n22717, n22718, n22719, n22720, 
      n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, 
      n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, 
      n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, 
      n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, 
      n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, 
      n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, 
      n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, 
      n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, 
      n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, 
      n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, 
      n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, 
      n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, 
      n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, 
      n22838, n22839, n22841, n22842, n22843, n22844, n22845, n22847, n22848, 
      n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, 
      n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, 
      n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, 
      n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, 
      n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, 
      n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, 
      n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, 
      n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, 
      n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, 
      n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, 
      n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, 
      n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, 
      n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22967, 
      n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, 
      n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, 
      n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, 
      n22995, n22996, n22998, n22999, n23000, n23001, n23002, n23003, n23004, 
      n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23014, 
      n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, 
      n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, 
      n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, 
      n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, 
      n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, 
      n23060, n23061, n23062, n23063, n23065, n23066, n23067, n23068, n23069, 
      n23070, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, 
      n23080, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, 
      n23090, n23091, n23092, n23093, n23094, n23096, n23097, n23098, n23099, 
      n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, 
      n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, 
      n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, 
      n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, 
      n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, 
      n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, 
      n23155, n23156, n23157, n23159, n23161, n23162, n23163, n23164, n23165, 
      n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, 
      n23175, n23176, n23177, n23179, n23180, n23181, n23182, n23183, n23184, 
      n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, 
      n23194, n23195, n23196, n23197, n23200, n23201, n23202, n23203, n23204, 
      n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23213, n23214, 
      n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23224, 
      n23225, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23235, 
      n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, 
      n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, 
      n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, 
      n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, 
      n23272, n23273, n23274, n23276, n23277, n23278, n23279, n23280, n23281, 
      n23282, n23283, n23284, n23285, n23286, n23287, n23289, n23290, n23291, 
      n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, 
      n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, 
      n23311, n23313, n23314, n23316, n23317, n23318, n23319, n23320, n23321, 
      n23322, n23323, n23324, n23326, n23327, n23328, n23329, n23330, n23331, 
      n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, 
      n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, 
      n23350, n23351, n23352, n23353, n23355, n23356, n23357, n23358, n23359, 
      n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, 
      n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, 
      n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, 
      n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, 
      n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, 
      n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, 
      n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23422, n23423, 
      n23424, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, 
      n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, 
      n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, 
      n23452, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, 
      n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, 
      n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, 
      n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, 
      n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, 
      n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, 
      n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23516, 
      n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, 
      n23526, n23527, n23528, n23529, n23531, n23532, n23534, n23535, n23536, 
      n23537, n23538, n23539, n23540, n23541, n23542, n23545, n23546, n23547, 
      n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, 
      n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, 
      n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, 
      n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, 
      n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23593, 
      n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, 
      n23603, n23604, n23605, n23606, n23607, n23608, n23610, n23611, n23612, 
      n23613, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, 
      n23623, n23624, n23625, n23626, n23628, n23629, n23630, n23631, n23632, 
      n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, 
      n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, 
      n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, 
      n23660, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, 
      n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, 
      n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, 
      n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, 
      n23697, n23698, n23699, n23700, n23702, n23703, n23704, n23705, n23706, 
      n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, 
      n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, 
      n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, 
      n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, 
      n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23751, n23752, 
      n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, 
      n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, 
      n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, 
      n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, 
      n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, 
      n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, 
      n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23816, 
      n23817, n23818, n23819, n23820, n23821, n23822, n23825, n23827, n23829, 
      n23830, n23831, n23832, n23833, n23834, n23835, n23837, n23838, n23839, 
      n23840, n23841, n23842, n23843, n23845, n23846, n23848, n23849, n23850, 
      n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, 
      n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, 
      n23871, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, 
      n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, 
      n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, 
      n23900, n23901, n23902, n23904, n23905, n23906, n23907, n23908, n23909, 
      n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, 
      n23919, n23920, n23921, n23922, n23923, n23924, n23926, n23927, n23929, 
      n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, 
      n23939, n23940, n23941, n23942, n23944, n23945, n23946, n23947, n23948, 
      n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, 
      n23958, n23959, n23960, n23961, n23962, n23963, n23965, n23966, n23967, 
      n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, 
      n23977, n23978, n23979, n23980, n23981, n23982, n23984, n23985, n23986, 
      n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, 
      n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24006, 
      n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, 
      n24017, n24018, n24019, n24020, n24021, n24022, n24024, n24025, n24026, 
      n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, 
      n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, 
      n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, 
      n24054, n24055, n24056, n24057, n24058, n24060, n24061, n24062, n24063, 
      n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, 
      n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, 
      n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, 
      n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, 
      n24100, n24101, n24102, n24104, n24105, n24106, n24107, n24108, n24109, 
      n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, 
      n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24128, 
      n24129, n24130, n24131, n24133, n24134, n24135, n24136, n24137, n24138, 
      n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, 
      n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, 
      n24157, n24158, n24159, n24160, n24162, n24163, n24164, n24165, n24166, 
      n24167, n24168, n24169, n24170, n24171, n24173, n24174, n24175, n24176, 
      n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, 
      n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, 
      n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, 
      n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, 
      n24213, n24214, n24215, n24216, n24218, n24219, n24220, n24221, n24222, 
      n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, 
      n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, 
      n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, 
      n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, 
      n24259, n24261, n24262, n24263, n24264, n24266, n24267, n24268, n24269, 
      n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, 
      n24279, n24280, n24282, n24283, n24284, n24285, n24286, n24287, n24288, 
      n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, 
      n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, 
      n24307, n24308, n24310, n24311, n24312, n24314, n24315, n24316, n24317, 
      n24318, n24319, n24322, n24323, n24324, n24325, n24326, n24327, n24328, 
      n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, 
      n24338, n24339, n24340, n24341, n24342, n24343, n24345, n24347, n24348, 
      n24349, n24350, n24351, n24352, n24353, n24355, n24356, n24357, n24358, 
      n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, 
      n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24376, n24377, 
      n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, 
      n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, 
      n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, 
      n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, 
      n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, 
      n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24433, 
      n24434, n24435, n24436, n24437, n24439, n24440, n24441, n24442, n24443, 
      n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, 
      n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, 
      n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, 
      n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, 
      n24480, n24481, n24482, n24483, n24484, n24486, n24487, n24488, n24489, 
      n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, 
      n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, 
      n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, 
      n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, 
      n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, 
      n24535, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, 
      n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, 
      n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, 
      n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, 
      n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, 
      n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, 
      n24590, n24591, n24592, n24593, n24595, n24596, n24597, n24598, n24600, 
      n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, 
      n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, 
      n24619, n24620, n24621, n24623, n24624, n24625, n24626, n24627, n24628, 
      n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, 
      n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, 
      n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, 
      n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, 
      n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, 
      n24674, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, 
      n24684, n24685, n24686, n24687, n24688, n24690, n24691, n24692, n24693, 
      n24694, n24695, n24696, n24697, n24699, n24700, n24701, n24703, n24704, 
      n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, 
      n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, 
      n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, 
      n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, 
      n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24750, 
      n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24760, 
      n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, 
      n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, 
      n24779, n24780, n24781, n24782, n24784, n24785, n24786, n24787, n24788, 
      n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, 
      n24798, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, 
      n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24816, n24817, 
      n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, 
      n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, 
      n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, 
      n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, 
      n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, 
      n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, 
      n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, 
      n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, 
      n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, 
      n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, 
      n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, 
      n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, 
      n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, 
      n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24948, 
      n24949, n24950, n24951, n24952, n24954, n24955, n24956, n24957, n24958, 
      n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, 
      n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, 
      n24977, n24978, n24980, n24981, n24982, n24983, n24984, n24985, n24986, 
      n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, 
      n24996, n24998, n24999, n25001, n25002, n25003, n25004, n25005, n25006, 
      n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, 
      n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, 
      n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, 
      n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, 
      n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25052, 
      n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, 
      n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, 
      n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, 
      n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, 
      n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, 
      n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, 
      n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, 
      n25116, n25117, n25119, n25120, n25122, n25123, n25124, n25126, n25127, 
      n25128, n25129, n25130, n25132, n25133, n25134, n25135, n25136, n25137, 
      n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, 
      n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, 
      n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, 
      n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, 
      n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, 
      n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, 
      n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, 
      n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, 
      n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, 
      n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, 
      n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, 
      n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, 
      n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, 
      n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, 
      n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, 
      n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, 
      n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, 
      n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, 
      n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, 
      n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, 
      n25318, n25319, n25320, n25321, n25322, n25324, n25325, n25326, n25327, 
      n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, 
      n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, 
      n25346, n25347, n25348, n25349, n25351, n25352, n25353, n25354, n25355, 
      n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, 
      n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, 
      n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, 
      n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, 
      n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, 
      n25401, n25404, n25405, n25406, n25408, n25409, n25410, n25411, n25412, 
      n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25421, n25422, 
      n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, 
      n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, 
      n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, 
      n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, 
      n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, 
      n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, 
      n25478, n25479, n25480, n25481, n25482, n25483, n25485, n25486, n25487, 
      n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, 
      n25497, n25498, n25499, n25500, n25501, n25502, n25504, n25505, n25506, 
      n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, 
      n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, 
      n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, 
      n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, 
      n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, 
      n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, 
      n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, 
      n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, 
      n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, 
      n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, 
      n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, 
      n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, 
      n25615, n25616, n25617, n25618, n25621, n25622, n25623, n25624, n25625, 
      n25626, n25627, n25628, n25629, n25631, n25632, n25633, n25634, n25635, 
      n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, 
      n25645, n25646, n25647, n25649, n25650, n25651, n25652, n25653, n25654, 
      n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, 
      n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, 
      n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, 
      n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, 
      n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, 
      n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, 
      n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, 
      n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, 
      n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, 
      n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, 
      n25746, n25747, n25750, n25751, n25752, n25753, n25754, n25755, n25756, 
      n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, 
      n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, 
      n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, 
      n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, 
      n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, 
      n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, 
      n25811, n25812, n25813, n25814, n25815, n25817, n25818, n25819, n25820, 
      n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, 
      n25830, n25831, n25832, n25833, n25834, n25836, n25837, n25838, n25839, 
      n25840, n25841, n25842, n25844, n25845, n25846, n25847, n25848, n25849, 
      n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, 
      n25860, n25861, n25862, n25864, n25865, n25866, n25867, n25868, n25869, 
      n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, 
      n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, 
      n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, 
      n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, 
      n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, 
      n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, 
      n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, 
      n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, 
      n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, 
      n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, 
      n25960, n25961, n25963, n25964, n25965, n25966, n25968, n25969, n25970, 
      n25971, n25972, n25973, n25974, n25975, n25977, n25978, n25979, n25980, 
      n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, 
      n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, 
      n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, 
      n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, 
      n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, 
      n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26034, n26035, 
      n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, 
      n26045, n26046, n26047, n26048, n26049, n26050, n26052, n26053, n26054, 
      n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, 
      n26064, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, 
      n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, 
      n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, 
      n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, 
      n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, 
      n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, 
      n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, 
      n26128, n26129, n26130, n26131, n26132, n26133, n26135, n26136, n26137, 
      n26138, n26139, n26140, n26141, n26142, n26144, n26145, n26146, n26147, 
      n26148, n26151, n26153, n26154, n26157, n26158, n26159, n26160, n26161, 
      n26162, n26163, n26164, n26166, n26168, n26169, n26170, n26171, n26172, 
      n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, 
      n26182, n26183, n26184, n26185, n26186, n26187, n26189, n26190, n26191, 
      n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, 
      n26201, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, 
      n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26221, 
      n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, 
      n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, 
      n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, 
      n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, 
      n26258, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, 
      n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, 
      n26277, n26278, n26279, n26280, n26281, n26282, n26284, n26285, n26286, 
      n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, 
      n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, 
      n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, 
      n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, 
      n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26332, n26333, 
      n26334, n26335, n26336, n26337, n26338, n26339, n26341, n26342, n26343, 
      n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, 
      n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, 
      n26363, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, 
      n26373, n26374, n26376, n26377, n26378, n26379, n26380, n26381, n26382, 
      n26383, n26384, n26385, n26386, n26387, n26389, n26390, n26392, n26394, 
      n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, 
      n26404, n26406, n26408, n26409, n26410, n26412, n26413, n26414, n26415, 
      n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, 
      n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, 
      n26434, n26435, n26436, n26437, n26439, n26440, n26441, n26442, n26443, 
      n26444, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, 
      n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, 
      n26463, n26464, n26465, n26466, n26468, n26469, n26470, n26471, n26472, 
      n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, 
      n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, 
      n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26501, 
      n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, 
      n26511, n26512, n26513, n26515, n26516, n26517, n26518, n26519, n26520, 
      n26521, n26522, n26523, n26524, n26525, n26528, n26529, n26530, n26531, 
      n26532, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, 
      n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, 
      n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, 
      n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, 
      n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, 
      n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, 
      n26590, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, 
      n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26608, n26609, 
      n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, 
      n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26628, 
      n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, 
      n26639, n26640, n26641, n26643, n26644, n26645, n26646, n26648, n26649, 
      n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, 
      n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, 
      n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, 
      n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, 
      n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, 
      n26696, n26697, n26699, n26700, n26701, n26702, n26703, n26704, n26705, 
      n26706, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, 
      n26716, n26717, n26718, n26719, n26720, n26721, n26723, n26724, n26725, 
      n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, 
      n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, 
      n26744, n26746, n26747, n26748, n26749, n26751, n26752, n26753, n26754, 
      n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, 
      n26764, n26765, n26766, n26767, n26768, n26769, n26771, n26772, n26773, 
      n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, 
      n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, 
      n26792, n26793, n26795, n26796, n26797, n26798, n26799, n26800, n26801, 
      n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, 
      n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, 
      n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, 
      n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, 
      n26839, n26840, n26841, n26842, n26843, n26844, n26846, n26848, n26849, 
      n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, 
      n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, 
      n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, 
      n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, 
      n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, 
      n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, 
      n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, 
      n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, 
      n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, 
      n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, 
      n26941, n26942, n26943, n26944, n26946, n26948, n26949, n26950, n26951, 
      n26952, n26953, n26954, n26956, n26957, n26958, n26959, n26960, n26961, 
      n26962, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, 
      n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, 
      n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, 
      n26990, n26991, n26992, n26994, n26995, n26996, n26997, n26998, n26999, 
      n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, 
      n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, 
      n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, 
      n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, 
      n27036, n27037, n27038, n27039, n27041, n27043, n27044, n27045, n27046, 
      n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, 
      n27056, n27057, n27058, n27060, n27061, n27062, n27063, n27064, n27065, 
      n27066, n27067, n27069, n27070, n27071, n27072, n27073, n27074, n27075, 
      n27076, n27077, n27078, n27079, n27080, n27081, n27083, n27084, n27085, 
      n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, 
      n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, 
      n27104, n27105, n27106, n27107, n27109, n27110, n27111, n27112, n27113, 
      n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, 
      n27123, n27124, n27126, n27127, n27128, n27129, n27130, n27131, n27132, 
      n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, 
      n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, 
      n27151, n27152, n27153, n27154, n27155, n27156, n27158, n27159, n27160, 
      n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, 
      n27170, n27171, n27172, n27173, n27175, n27177, n27178, n27179, n27180, 
      n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27190, 
      n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, 
      n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, 
      n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, 
      n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, 
      n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, 
      n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, 
      n27246, n27247, n27248, n27249, n27250, n27252, n27253, n27254, n27255, 
      n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, 
      n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, 
      n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, 
      n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, 
      n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, 
      n27304, n27305, n27306, n27307, n27308, n27310, n27311, n27312, n27313, 
      n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, 
      n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, 
      n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, 
      n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, 
      n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, 
      n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, 
      n27368, n27369, n27370, n27371, n27372, n27374, n27375, n27376, n27377, 
      n27378, n27379, n27380, n27381, n27382, n27384, n27385, n27386, n27387, 
      n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, 
      n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, 
      n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, 
      n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, 
      n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, 
      n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, 
      n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, 
      n27453, n27454, n27456, n27457, n27458, n27459, n27460, n27461, n27462, 
      n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, 
      n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, 
      n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, 
      n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, 
      n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, 
      n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, 
      n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, 
      n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, 
      n27537, n27538, n27539, n27541, n27542, n27543, n27544, n27545, n27546, 
      n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, 
      n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, 
      n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, 
      n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, 
      n27583, n27584, n27585, n27586, n27588, n27589, n27590, n27591, n27592, 
      n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, 
      n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, 
      n27612, n27613, n27614, n27615, n27616, n27617, n27619, n27620, n27621, 
      n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, 
      n27631, n27632, n27633, n27634, n27636, n27637, n27638, n27639, n27640, 
      n27641, n27642, n27643, n27645, n27646, n27647, n27648, n27649, n27650, 
      n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, 
      n27660, n27661, n27662, n27663, n27664, n27666, n27668, n27669, n27670, 
      n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, 
      n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, 
      n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, 
      n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, 
      n27707, n27708, n27709, n27711, n27712, n27713, n27714, n27715, n27716, 
      n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, 
      n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, 
      n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, 
      n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27755, 
      n27757, n27758, n27759, n27760, n27761, n27762, n27764, n27765, n27766, 
      n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775, 
      n27776, n27777, n27778, n27779, n27780, n27782, n27784, n27785, n27786, 
      n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, 
      n27796, n27797, n27798, n27799, n27800, n27802, n27803, n27804, n27805, 
      n27806, n27807, n27808, n27809, n27811, n27812, n27813, n27814, n27815, 
      n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, 
      n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, 
      n27834, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, 
      n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, 
      n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, 
      n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, 
      n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, 
      n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, 
      n27889, n27890, n27891, n27892, n27893, n27894, n27898, n27899, n27900, 
      n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, 
      n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919, 
      n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928, 
      n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937, 
      n27938, n27940, n27941, n27942, n27943, n27944, n27947, n27948, n27949, 
      n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, 
      n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, 
      n27969, n27970, n27971, n27972, n27974, n27975, n27976, n27977, n27978, 
      n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, 
      n27988, n27989, n27990, n27991, n27995, n27996, n27997, n27998, n27999, 
      n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, 
      n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, 
      n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, 
      n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, 
      n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, 
      n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, 
      n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, 
      n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, 
      n28072, n28073, n28074, n28075, n28076, n28078, n28079, n28080, n28081, 
      n28083, n28084, n28086, n28087, n28088, n28089, n28090, n28091, n28092, 
      n28093, n28094, n28095, n28096, n28097, n28099, n28100, n28101, n28102, 
      n28103, n28104, n28105, n28107, n28108, n28109, n28110, n28111, n28112, 
      n28114, n28115, n28116, n28121, n28122, n28126, n28130, n28133, n28140, 
      n28142, n28143, n28144, n28147, n28149, n28155, n28157, n28161, n28162, 
      n28164, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28179, 
      n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, 
      n28191, n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, 
      n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28210, 
      n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, 
      n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, 
      n28229, n28230, n28231, n28232, n28233, n28235, n28236, n28237, n28238, 
      n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, 
      n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, 
      n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, 
      n28267, n28268, n28269, n28270, n28271, n28273, n28274, n28275, n28276, 
      n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, 
      n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28294, n28295, 
      n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28305, 
      n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, 
      n28315, n28316, n28317, n28319, n28320, n28321, n28322, n28323, n28324, 
      n28326, n28327, n28329, n28330, n28331, n28332, n28333, n28334, n28335, 
      n28336, n28337, n28339, n28340, n28341, n28343, n28344, n28345, n28347, 
      n28348, n28349, n28351, n28352, n28353, n28354, n28355, n28357, n28358, 
      n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28367, n28368, 
      n28369, n28370, n28371, n28372, n28373, n28376, n28377, n28378, n28379, 
      n28380, n28381, n28383, n28384, n28385, n28386, n28387, n28388, n28390, 
      n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, 
      n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, 
      n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, 
      n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, 
      n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, 
      n28437, n28438, n28439, n28440, n28441, n28442, n28444, n28445, n28446, 
      n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, 
      n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28465, n28466, 
      n28467, n28468, n28470, n28471, n28472, n28473, n28474, n28475, n28476, 
      n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, 
      n28486, n28487, n28488, n28489, n28491, n28492, n28493, n28494, n28495, 
      n28496, n28497, n28499, n28500, n28501, n28503, n28504, n28505, n28506, 
      n28507, n28508, n28509, n28510, n28512, n28513, n28514, n28515, n28516, 
      n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, 
      n28526, n28527, n28528, n28530, n28531, n28532, n28534, n28535, n28536, 
      n28538, n28540, n28541, n28542, n28543, n28544, n28545, n28547, n28548, 
      n28549, n28550, n28551, n28552, n28554, n28555, n28557, n28558, n28559, 
      n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, 
      n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, 
      n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, 
      n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, 
      n28596, n28597, n28598, n28600, n28601, n28602, n28603, n28604, n28605, 
      n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, 
      n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, 
      n28624, n28625, n28626, n28627, n28628, n28630, n28631, n28632, n28633, 
      n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, 
      n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, 
      n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, 
      n28661, n28662, n28663, n28665, n28666, n28667, n28668, n28669, n28670, 
      n28671, n28672, n28674, n28676, n28677, n28678, n28679, n28680, n28681, 
      n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, 
      n28691, n28692, n28693, n28694, n28695, n28696, n28698, n28699, n28701, 
      n28702, n28703, n28704, n28706, n28707, n28708, n28709, n28710, n28711, 
      n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, 
      n28721, n28722, n28723, n28725, n28726, n28727, n28728, n28729, n28730, 
      n28732, n28733, n28734, n28736, n28737, n28738, n28739, n28741, n28742, 
      n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, 
      n28752, n28753, n28754, n28756, n28757, n28759, n28761, n28762, n28763, 
      n28764, n28765, n28766, n28767, n28768, n28769, n28771, n28775, n28776, 
      n28779, n28783, n28785, n28789, n28790, n28791, n28792, n28793, n28794, 
      n28796, n28797, n28798, n28800, n28801, n28802, n28803, n28804, n28805, 
      n28806, n28807, n28808, n28810, n28811, n28812, n28813, n28814, n28815, 
      n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, 
      n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, 
      n28834, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28844, 
      n28845, n28847, n28848, n28849, n28851, n28852, n28853, n28854, n28855, 
      n28856, n28857, n28858, n28860, n28861, n28862, n28863, n28864, n28866, 
      n28867, n28869, n28871, n28872, n28874, n28875, n28876, n28877, n28878, 
      n28879, n28882, n28883, n28885, n28886, n28887, n28888, n28889, n28890, 
      n28891, n28892, n28894, n28895, n28896, n28897, n28898, n28899, n28900, 
      n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, 
      n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, 
      n28919, n28920, n28921, n28922, n28923, n28924, n28928, n28929, n28930, 
      n28931, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, 
      n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, 
      n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28958, n28960, 
      n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28969, n28970, 
      n28971, n28972, n28973, n28974, n28975, n28977, n28978, n28979, n28980, 
      n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, 
      n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28998, n28999, 
      n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, 
      n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, 
      n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, 
      n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, 
      n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, 
      n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, 
      n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, 
      n29063, n29064, n29065, n29066, n29067, n29069, n29070, n29071, n29072, 
      n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29081, n29082, 
      n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, 
      n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, 
      n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, 
      n29110, n29111, n29112, n29114, n29115, n29116, n29117, n29118, n29119, 
      n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, 
      n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, 
      n29138, n29139, n29140, n29142, n29143, n29144, n29145, n29146, n29147, 
      n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, 
      n29157, n29158, n29159, n29160, n29161, n29163, n29164, n29165, n29166, 
      n29168, n29169, n29171, n29172, n29173, n29174, n29175, n29176, n29177, 
      n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, 
      n29187, n29188, n29189, n29191, n29192, n29193, n29194, n29195, n29196, 
      n29197, n29198, n29199, n29201, n29202, n29203, n29204, n29205, n29206, 
      n29207, n29208, n29209, n29210, n29211, n29212, n29214, n29215, n29217, 
      n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, 
      n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29235, n29236, 
      n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, 
      n29246, n29247, n29248, n29249, n29251, n29253, n29255, n29256, n29257, 
      n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29268, 
      n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, 
      n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, 
      n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, 
      n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, 
      n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, 
      n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, 
      n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, 
      n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, 
      n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, 
      n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, 
      n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, 
      n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, 
      n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, 
      n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, 
      n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, 
      n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, 
      n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, 
      n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, 
      n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, 
      n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, 
      n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, 
      n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, 
      n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, 
      n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, 
      n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, 
      n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, 
      n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, 
      n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, 
      n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, 
      n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, 
      n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, 
      n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, 
      n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, 
      n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, 
      n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, 
      n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, 
      n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, 
      n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, 
      n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, 
      n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, 
      n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, 
      n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, 
      n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, 
      n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, 
      n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, 
      n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, 
      n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, 
      n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, 
      n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, 
      n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, 
      n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, 
      n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, 
      n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, 
      n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, 
      n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, 
      n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, 
      n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, 
      n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, 
      n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, 
      n29800, n29801 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n26973, A2 => n28213, ZN => n114);
   U2 : AOI22_X1 port map( A1 => n27917, A2 => n27918, B1 => n27907, B2 => 
                           n27906, ZN => n27914);
   U3 : INV_X1 port map( A => n27671, ZN => n85);
   U6 : BUF_X1 port map( A => n26652, Z => n27539);
   U7 : AND3_X1 port map( A1 => n278, A2 => n923, A3 => n921, ZN => n27877);
   U8 : INV_X1 port map( A => n3722, ZN => n27978);
   U9 : AND3_X1 port map( A1 => n4064, A2 => n2013, A3 => n4063, ZN => n25914);
   U14 : OR2_X1 port map( A1 => n23051, A2 => n24341, ZN => n1223);
   U16 : INV_X1 port map( A => n24758, ZN => n171);
   U18 : OAI21_X2 port map( B1 => n23019, B2 => n23018, A => n23017, ZN => 
                           n24688);
   U22 : OR2_X1 port map( A1 => n28460, A2 => n23078, ZN => n23838);
   U25 : OR2_X1 port map( A1 => n3940, A2 => n23825, ZN => n4483);
   U29 : OR2_X1 port map( A1 => n20858, A2 => n21159, ZN => n14);
   U30 : OR2_X1 port map( A1 => n20933, A2 => n20533, ZN => n1342);
   U32 : INV_X1 port map( A => n21495, ZN => n44);
   U33 : AND2_X1 port map( A1 => n21481, A2 => n21483, ZN => n20368);
   U34 : NOR2_X1 port map( A1 => n21481, A2 => n21574, ZN => n20849);
   U35 : INV_X1 port map( A => n21497, ZN => n7);
   U39 : BUF_X1 port map( A => n20225, Z => n20503);
   U41 : OR2_X1 port map( A1 => n17849, A2 => n18137, ZN => n18142);
   U42 : OAI211_X1 port map( C1 => n18506, C2 => n18216, A => n28763, B => 
                           n18217, ZN => n2045);
   U43 : OR2_X1 port map( A1 => n18252, A2 => n17771, ZN => n3086);
   U44 : AND2_X1 port map( A1 => n18101, A2 => n18449, ZN => n106);
   U48 : OR2_X1 port map( A1 => n5200, A2 => n18173, ZN => n1137);
   U49 : OR2_X1 port map( A1 => n18324, A2 => n18263, ZN => n18323);
   U50 : AND2_X1 port map( A1 => n18306, A2 => n17679, ZN => n17680);
   U52 : INV_X1 port map( A => n18465, ZN => n145);
   U53 : INV_X1 port map( A => n18270, ZN => n48);
   U54 : AND3_X1 port map( A1 => n17187, A2 => n17186, A3 => n17185, ZN => 
                           n18122);
   U57 : OR2_X1 port map( A1 => n18507, A2 => n29496, ZN => n18074);
   U58 : INV_X1 port map( A => n18213, ZN => n511);
   U62 : OR2_X1 port map( A1 => n16917, A2 => n16916, ZN => n186);
   U64 : OAI22_X1 port map( A1 => n17315, A2 => n17316, B1 => n4220, B2 => 
                           n17562, ZN => n792);
   U65 : NOR2_X1 port map( A1 => n17528, A2 => n17524, ZN => n17182);
   U66 : OR2_X1 port map( A1 => n16811, A2 => n16812, ZN => n3302);
   U68 : XNOR2_X1 port map( A => n15068, B => n15067, ZN => n17435);
   U69 : XNOR2_X1 port map( A => n16256, B => n15977, ZN => n16627);
   U70 : OR2_X1 port map( A1 => n15399, A2 => n13638, ZN => n6856);
   U73 : OR2_X1 port map( A1 => n15370, A2 => n15009, ZN => n3783);
   U74 : OR2_X1 port map( A1 => n5049, A2 => n15274, ZN => n217);
   U75 : AND2_X1 port map( A1 => n15046, A2 => n15342, ZN => n15229);
   U81 : OR2_X1 port map( A1 => n13766, A2 => n14481, ZN => n140);
   U83 : OR2_X1 port map( A1 => n14037, A2 => n60, ZN => n13722);
   U84 : AND2_X1 port map( A1 => n29565, A2 => n29306, ZN => n12121);
   U85 : OR2_X1 port map( A1 => n14365, A2 => n14091, ZN => n731);
   U87 : NOR2_X1 port map( A1 => n12887, A2 => n1841, ZN => n245);
   U88 : INV_X1 port map( A => n14452, ZN => n190);
   U89 : INV_X1 port map( A => n13589, ZN => n58);
   U90 : INV_X1 port map( A => n29089, ZN => n60);
   U92 : OAI21_X1 port map( B1 => n30, B2 => n14400, A => n29, ZN => n2112);
   U93 : INV_X1 port map( A => n14398, ZN => n30);
   U94 : XNOR2_X1 port map( A => n12606, B => n12605, ZN => n14292);
   U95 : AND2_X1 port map( A1 => n11985, A2 => n11986, ZN => n163);
   U96 : NAND3_X1 port map( A1 => n11697, A2 => n11696, A3 => n11695, ZN => 
                           n13484);
   U97 : OR2_X1 port map( A1 => n10900, A2 => n919, ZN => n172);
   U98 : OAI211_X1 port map( C1 => n12297, C2 => n12296, A => n12295, B => 
                           n12294, ZN => n13121);
   U99 : OR2_X1 port map( A1 => n12044, A2 => n12043, ZN => n12045);
   U103 : AND3_X1 port map( A1 => n4902, A2 => n11172, A3 => n11171, ZN => 
                           n11194);
   U105 : OR2_X1 port map( A1 => n4789, A2 => n4790, ZN => n11417);
   U106 : AND2_X1 port map( A1 => n10963, A2 => n10956, ZN => n9859);
   U108 : OAI21_X1 port map( B1 => n11289, B2 => n11290, A => n11077, ZN => 
                           n5717);
   U111 : INV_X1 port map( A => n11113, ZN => n242);
   U119 : AND3_X1 port map( A1 => n1417, A2 => n1418, A3 => n7574, ZN => n15);
   U120 : OR2_X1 port map( A1 => n8360, A2 => n9037, ZN => n6189);
   U121 : INV_X1 port map( A => n9374, ZN => n11);
   U122 : BUF_X1 port map( A => n7679, Z => n9210);
   U123 : INV_X1 port map( A => n9122, ZN => n81);
   U127 : AND3_X1 port map( A1 => n5493, A2 => n7780, A3 => n7779, ZN => n8427)
                           ;
   U128 : OAI211_X1 port map( C1 => n7425, C2 => n7426, A => n3929, B => n1358,
                           ZN => n8740);
   U129 : INV_X1 port map( A => n8215, ZN => n8212);
   U130 : BUF_X1 port map( A => n8221, Z => n7827);
   U137 : AND2_X1 port map( A1 => n29621, A2 => n26125, ZN => n26860);
   U140 : OR2_X1 port map( A1 => n1807, A2 => n29043, ZN => n24418);
   U142 : AOI22_X1 port map( A1 => n21426, A2 => n5827, B1 => n20129, B2 => 
                           n6937, ZN => n5622);
   U146 : AND2_X1 port map( A1 => n26917, A2 => n26172, ZN => n26553);
   U147 : BUF_X1 port map( A => n14630, Z => n15394);
   U149 : OR2_X1 port map( A1 => n11282, A2 => n10518, ZN => n10519);
   U150 : AND2_X1 port map( A1 => n20299, A2 => n20443, ZN => n128);
   U153 : AND2_X1 port map( A1 => n17336, A2 => n17155, ZN => n15581);
   U154 : OR2_X1 port map( A1 => n17336, A2 => n17155, ZN => n241);
   U158 : AND2_X1 port map( A1 => n27711, A2 => n27724, ZN => n27694);
   U160 : AND2_X1 port map( A1 => n20547, A2 => n20546, ZN => n19960);
   U165 : OR2_X1 port map( A1 => n24347, A2 => n24436, ZN => n24442);
   U166 : OAI21_X1 port map( B1 => n29090, B2 => n85, A => n84, ZN => n27658);
   U167 : OR2_X1 port map( A1 => n11195, A2 => n11194, ZN => n179);
   U171 : XNOR2_X1 port map( A => n18568, B => n18567, ZN => n20077);
   U172 : INV_X1 port map( A => n3315, ZN => n184);
   U173 : OR2_X1 port map( A1 => n15098, A2 => n3315, ZN => n183);
   U175 : OR3_X1 port map( A1 => n395, A2 => n26880, A3 => n27300, ZN => n26882
                           );
   U176 : OR2_X1 port map( A1 => n26166, A2 => n29054, ZN => n4399);
   U177 : OR2_X1 port map( A1 => n26410, A2 => n26797, ZN => n56);
   U179 : AND2_X1 port map( A1 => n23403, A2 => n23214, ZN => n23749);
   U181 : OR2_X1 port map( A1 => n15402, A2 => n13639, ZN => n14896);
   U185 : AOI21_X1 port map( B1 => n9202, B2 => n9199, A => n231, ZN => n2196);
   U188 : OR2_X1 port map( A1 => n2794, A2 => n27739, ZN => n1216);
   U190 : OR2_X1 port map( A1 => n26965, A2 => n27497, ZN => n225);
   U191 : OAI21_X1 port map( B1 => n17997, B2 => n17883, A => n3283, ZN => 
                           n2468);
   U193 : OR2_X1 port map( A1 => n1533, A2 => n25628, ZN => n1532);
   U195 : OR3_X1 port map( A1 => n28567, A2 => n2823, A3 => n24020, ZN => n275)
                           ;
   U196 : BUF_X1 port map( A => n27407, Z => n342);
   U199 : OAI21_X1 port map( B1 => n22970, B2 => n22969, A => n22968, ZN => 
                           n26023);
   U204 : BUF_X1 port map( A => n14358, Z => n14272);
   U205 : OAI211_X1 port map( C1 => n487, C2 => n28418, A => n23838, B => 
                           n23837, ZN => n1162);
   U206 : OR2_X1 port map( A1 => n29057, A2 => n29647, ZN => n17693);
   U209 : NAND3_X1 port map( A1 => n24447, A2 => n24756, A3 => n24218, ZN => 
                           n24219);
   U210 : AND2_X2 port map( A1 => n23561, A2 => n23560, ZN => n24447);
   U211 : NOR2_X1 port map( A1 => n14392, A2 => n1, ZN => n2207);
   U212 : INV_X1 port map( A => n14391, ZN => n1);
   U213 : NAND2_X1 port map( A1 => n6048, A2 => n15284, ZN => n14391);
   U215 : NAND2_X1 port map( A1 => n28762, A2 => n3784, ZN => n2);
   U220 : NAND2_X1 port map( A1 => n9, A2 => n6, ZN => n19832);
   U221 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n6);
   U222 : NAND2_X1 port map( A1 => n28789, A2 => n20865, ZN => n8);
   U223 : NAND2_X1 port map( A1 => n19830, A2 => n21497, ZN => n9);
   U237 : NAND3_X2 port map( A1 => n6218, A2 => n19900, A3 => n6219, ZN => 
                           n3838);
   U239 : OR2_X1 port map( A1 => n11921, A2 => n11853, ZN => n3521);
   U242 : NAND2_X1 port map( A1 => n12, A2 => n10, ZN => n8571);
   U243 : NAND2_X1 port map( A1 => n9370, A2 => n11, ZN => n10);
   U244 : NAND2_X1 port map( A1 => n8569, A2 => n8929, ZN => n9370);
   U245 : NAND2_X1 port map( A1 => n9373, A2 => n9374, ZN => n12);
   U246 : NAND3_X1 port map( A1 => n24123, A2 => n24125, A3 => n24124, ZN => 
                           n153);
   U250 : NAND3_X1 port map( A1 => n3119, A2 => n21161, A3 => n13, ZN => n22656
                           );
   U253 : NAND2_X1 port map( A1 => n8208, A2 => n7700, ZN => n7423);
   U254 : NAND2_X1 port map( A1 => n3579, A2 => n3581, ZN => n888);
   U257 : BUF_X1 port map( A => n22829, Z => n355);
   U258 : XNOR2_X1 port map( A => n9673, B => n4601, ZN => n11163);
   U267 : NAND3_X1 port map( A1 => n16, A2 => n17848, A3 => n3264, ZN => n6443)
                           ;
   U268 : NAND2_X1 port map( A1 => n2811, A2 => n17847, ZN => n16);
   U275 : NAND2_X1 port map( A1 => n6829, A2 => n16974, ZN => n17717);
   U276 : NAND2_X1 port map( A1 => n18270, A2 => n18511, ZN => n1124);
   U277 : NAND2_X1 port map( A1 => n29647, A2 => n18508, ZN => n18270);
   U278 : NAND3_X1 port map( A1 => n7871, A2 => n7053, A3 => n7960, ZN => n7055
                           );
   U280 : NAND2_X1 port map( A1 => n6679, A2 => n12050, ZN => n6678);
   U284 : NAND3_X1 port map( A1 => n19, A2 => n12240, A3 => n4617, ZN => n4616)
                           ;
   U285 : NAND2_X1 port map( A1 => n12159, A2 => n11969, ZN => n19);
   U291 : AND4_X2 port map( A1 => n5502, A2 => n5504, A3 => n24627, A4 => 
                           n24626, ZN => n27025);
   U295 : NAND2_X1 port map( A1 => n22, A2 => n11185, ZN => n11327);
   U299 : NAND3_X1 port map( A1 => n18933, A2 => n21286, A3 => n21291, ZN => 
                           n24);
   U300 : NAND2_X1 port map( A1 => n21704, A2 => n21277, ZN => n21374);
   U301 : OR2_X1 port map( A1 => n8258, A2 => n28615, ZN => n7468);
   U305 : NAND2_X1 port map( A1 => n8608, A2 => n8320, ZN => n8747);
   U306 : OR2_X1 port map( A1 => n702, A2 => n20160, ZN => n273);
   U308 : NOR2_X2 port map( A1 => n6824, A2 => n25422, ZN => n27442);
   U310 : NAND2_X1 port map( A1 => n25, A2 => n11470, ZN => n12955);
   U314 : NAND3_X1 port map( A1 => n14466, A2 => n4840, A3 => n13678, ZN => 
                           n13680);
   U315 : AND3_X2 port map( A1 => n1946, A2 => n5437, A3 => n5435, ZN => n21497
                           );
   U316 : OR2_X1 port map( A1 => n10726, A2 => n10929, ZN => n10933);
   U317 : AOI21_X1 port map( B1 => n23519, B2 => n21058, A => n23516, ZN => 
                           n21059);
   U318 : NAND2_X1 port map( A1 => n23682, A2 => n29544, ZN => n23519);
   U319 : NAND2_X1 port map( A1 => n17201, A2 => n17203, ZN => n2741);
   U320 : AND2_X1 port map( A1 => n19054, A2 => n20178, ZN => n20055);
   U324 : NAND2_X1 port map( A1 => n14400, A2 => n14399, ZN => n29);
   U325 : NAND3_X1 port map( A1 => n2890, A2 => n8849, A3 => n8850, ZN => n8854
                           );
   U326 : AND2_X2 port map( A1 => n7538, A2 => n7539, ZN => n9060);
   U327 : NAND2_X1 port map( A1 => n17430, A2 => n31, ZN => n18398);
   U329 : NAND3_X1 port map( A1 => n5025, A2 => n14897, A3 => n14896, ZN => 
                           n14898);
   U331 : NAND2_X1 port map( A1 => n5658, A2 => n21495, ZN => n5657);
   U332 : XNOR2_X2 port map( A => n7117, B => Key(8), ZN => n7164);
   U333 : NAND2_X1 port map( A1 => n35, A2 => n32, ZN => n4259);
   U334 : NAND2_X1 port map( A1 => n34, A2 => n28171, ZN => n32);
   U336 : NAND2_X1 port map( A1 => n5847, A2 => n13583, ZN => n34);
   U337 : NAND2_X1 port map( A1 => n4260, A2 => n13730, ZN => n35);
   U338 : NAND3_X1 port map( A1 => n3167, A2 => n7771, A3 => n7770, ZN => n7772
                           );
   U339 : NAND3_X1 port map( A1 => n24125, A2 => n24705, A3 => n24338, ZN => 
                           n5836);
   U341 : AND2_X2 port map( A1 => n5898, A2 => n5897, ZN => n21982);
   U343 : INV_X1 port map( A => n14738, ZN => n36);
   U344 : NAND2_X1 port map( A1 => n7716, A2 => n7717, ZN => n7720);
   U346 : NAND3_X1 port map( A1 => n11321, A2 => n11322, A3 => n11181, ZN => 
                           n37);
   U347 : NAND2_X1 port map( A1 => n11324, A2 => n29316, ZN => n39);
   U352 : NAND2_X1 port map( A1 => n3753, A2 => n18286, ZN => n40);
   U354 : NAND3_X1 port map( A1 => n8998, A2 => n9435, A3 => n8996, ZN => n41);
   U355 : NAND2_X1 port map( A1 => n42, A2 => n16942, ZN => n6643);
   U359 : NAND3_X1 port map( A1 => n11063, A2 => n1851, A3 => n10641, ZN => 
                           n2084);
   U361 : NAND2_X1 port map( A1 => n28789, A2 => n44, ZN => n43);
   U364 : INV_X1 port map( A => n7266, ZN => n7709);
   U365 : XNOR2_X1 port map( A => n16051, B => n16620, ZN => n16196);
   U366 : NOR2_X1 port map( A1 => n20293, A2 => n19815, ZN => n20122);
   U368 : NAND3_X1 port map( A1 => n3175, A2 => n6352, A3 => n3488, ZN => 
                           n14696);
   U369 : OR2_X1 port map( A1 => n18449, A2 => n18451, ZN => n1026);
   U373 : NAND3_X1 port map( A1 => n4130, A2 => n27031, A3 => n4132, ZN => 
                           n3611);
   U374 : NAND2_X1 port map( A1 => n19060, A2 => n20221, ZN => n19062);
   U375 : NAND2_X1 port map( A1 => n29587, A2 => n20222, ZN => n19060);
   U377 : NAND2_X1 port map( A1 => n48, A2 => n18271, ZN => n46);
   U380 : MUX2_X1 port map( A => n11708, B => n11648, S => n11417, Z => n11408)
                           ;
   U381 : AND2_X1 port map( A1 => n23968, A2 => n24209, ZN => n23116);
   U388 : AND2_X1 port map( A1 => n12321, A2 => n12050, ZN => n77);
   U393 : NAND2_X1 port map( A1 => n50, A2 => n1048, ZN => n12504);
   U394 : NAND2_X1 port map( A1 => n11647, A2 => n743, ZN => n50);
   U395 : NOR2_X2 port map( A1 => n162, A2 => n51, ZN => n24949);
   U397 : NAND2_X1 port map( A1 => n24475, A2 => n53, ZN => n52);
   U398 : INV_X1 port map( A => n6348, ZN => n53);
   U399 : NAND2_X1 port map( A1 => n23841, A2 => n6348, ZN => n54);
   U400 : OR2_X2 port map( A1 => n10831, A2 => n10832, ZN => n11648);
   U402 : OAI21_X1 port map( B1 => n14662, B2 => n14663, A => n55, ZN => n14665
                           );
   U403 : INV_X1 port map( A => n14660, ZN => n55);
   U405 : NAND2_X1 port map( A1 => n10808, A2 => n10544, ZN => n10805);
   U406 : NAND3_X1 port map( A1 => n461, A2 => n28415, A3 => n25008, ZN => 
                           n4141);
   U411 : MUX2_X2 port map( A => n9477, B => n13082, S => n13081, Z => n13051);
   U414 : NAND2_X1 port map( A1 => n1717, A2 => n3833, ZN => n1716);
   U418 : OR2_X2 port map( A1 => n2832, A2 => n7589, ZN => n7875);
   U421 : OAI211_X1 port map( C1 => n13720, C2 => n60, A => n59, B => n58, ZN 
                           => n57);
   U425 : OAI21_X1 port map( B1 => n6904, B2 => n21471, A => n21232, ZN => 
                           n21233);
   U428 : INV_X1 port map( A => n8187, ZN => n8936);
   U433 : NAND2_X1 port map( A1 => n28894, A2 => n20616, ZN => n20256);
   U439 : NAND3_X1 port map( A1 => n9188, A2 => n9185, A3 => n9184, ZN => n887)
                           ;
   U440 : NAND2_X1 port map( A1 => n9012, A2 => n8910, ZN => n8482);
   U443 : NAND3_X2 port map( A1 => n2676, A2 => n7412, A3 => n7414, ZN => n2677
                           );
   U446 : NAND2_X1 port map( A1 => n18171, A2 => n17780, ZN => n1563);
   U448 : BUF_X1 port map( A => n27271, Z => n27923);
   U449 : INV_X1 port map( A => n21467, ZN => n19793);
   U450 : NAND2_X1 port map( A1 => n5953, A2 => n21113, ZN => n21467);
   U452 : NAND2_X1 port map( A1 => n1436, A2 => n17447, ZN => n1468);
   U455 : OR2_X1 port map( A1 => n28796, A2 => n23408, ZN => n23748);
   U459 : NAND2_X1 port map( A1 => n14122, A2 => n14366, ZN => n14093);
   U460 : OAI21_X1 port map( B1 => n28800, B2 => n17464, A => n63, ZN => n5251)
                           ;
   U461 : NAND2_X1 port map( A1 => n17466, A2 => n4246, ZN => n63);
   U463 : NAND3_X2 port map( A1 => n64, A2 => n13765, A3 => n13766, ZN => 
                           n15207);
   U464 : NAND2_X1 port map( A1 => n6744, A2 => n13947, ZN => n64);
   U467 : NAND3_X1 port map( A1 => n66, A2 => n16152, A3 => n519, ZN => n2457);
   U470 : OAI21_X1 port map( B1 => n23192, B2 => n23193, A => n28764, ZN => 
                           n3158);
   U475 : XNOR2_X2 port map( A => n15969, B => n15970, ZN => n17277);
   U476 : OAI211_X2 port map( C1 => n14060, C2 => n4185, A => n4184, B => n4181
                           , ZN => n16232);
   U477 : AND2_X1 port map( A1 => n11033, A2 => n11248, ZN => n10525);
   U478 : NAND2_X1 port map( A1 => n69, A2 => n18180, ZN => n17792);
   U479 : NAND2_X1 port map( A1 => n17788, A2 => n17789, ZN => n69);
   U480 : NAND2_X1 port map( A1 => n4477, A2 => n4476, ZN => n17789);
   U482 : NAND2_X1 port map( A1 => n6399, A2 => n6400, ZN => n20876);
   U484 : NAND2_X1 port map( A1 => n4446, A2 => n12208, ZN => n71);
   U486 : NAND2_X1 port map( A1 => n6117, A2 => n20914, ZN => n73);
   U490 : AND2_X2 port map( A1 => n76, A2 => n75, ZN => n21291);
   U491 : NAND2_X1 port map( A1 => n18891, A2 => n18892, ZN => n75);
   U492 : NAND2_X1 port map( A1 => n5424, A2 => n3911, ZN => n76);
   U493 : NAND2_X1 port map( A1 => n566, A2 => n77, ZN => n11771);
   U497 : NOR2_X2 port map( A1 => n17682, A2 => n17681, ZN => n19637);
   U503 : MUX2_X2 port map( A => n25986, B => n25985, S => n27013, Z => n28019)
                           ;
   U504 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => n6172);
   U505 : NAND2_X1 port map( A1 => n9125, A2 => n9122, ZN => n79);
   U506 : NAND2_X1 port map( A1 => n1651, A2 => n1793, ZN => n80);
   U510 : NAND2_X1 port map( A1 => n15393, A2 => n15392, ZN => n82);
   U513 : INV_X1 port map( A => n18603, ZN => n18604);
   U514 : NAND3_X1 port map( A1 => n28142, A2 => n18600, A3 => n17989, ZN => 
                           n18603);
   U515 : NOR2_X1 port map( A1 => n28522, A2 => n24804, ZN => n24805);
   U518 : NAND2_X1 port map( A1 => n400, A2 => n27701, ZN => n27163);
   U520 : NAND2_X1 port map( A1 => n29091, A2 => n27672, ZN => n84);
   U521 : BUF_X1 port map( A => n27728, Z => n1826);
   U522 : NOR2_X1 port map( A1 => n17347, A2 => n29632, ZN => n16949);
   U532 : MUX2_X1 port map( A => n9229, B => n9232, S => n9233, Z => n7000);
   U535 : NAND2_X1 port map( A1 => n6961, A2 => n6960, ZN => n87);
   U538 : OAI21_X1 port map( B1 => n6061, B2 => n14792, A => n14970, ZN => n88)
                           ;
   U539 : INV_X1 port map( A => n12517, ZN => n12077);
   U540 : MUX2_X1 port map( A => n12271, B => n12578, S => n12517, Z => n11567)
                           ;
   U541 : NOR2_X2 port map( A1 => n11098, A2 => n11097, ZN => n12517);
   U544 : NAND2_X1 port map( A1 => n432, A2 => n89, ZN => n6165);
   U545 : NOR2_X1 port map( A1 => n5258, A2 => n10431, ZN => n89);
   U547 : INV_X1 port map( A => n28105, ZN => n91);
   U548 : NAND3_X1 port map( A1 => n13944, A2 => n13941, A3 => n15025, ZN => 
                           n13950);
   U549 : OAI21_X1 port map( B1 => n26236, B2 => n26753, A => n92, ZN => n26756
                           );
   U550 : NAND2_X1 port map( A1 => n26753, A2 => n28575, ZN => n92);
   U552 : BUF_X1 port map( A => n15165, Z => n1850);
   U555 : NAND3_X1 port map( A1 => n13651, A2 => n14303, A3 => n13817, ZN => 
                           n13650);
   U557 : NAND2_X1 port map( A1 => n27124, A2 => n27190, ZN => n26336);
   U559 : OR2_X1 port map( A1 => n26338, A2 => n26339, ZN => n96);
   U561 : NAND3_X1 port map( A1 => n19899, A2 => n20645, A3 => n19927, ZN => 
                           n6218);
   U568 : NAND3_X1 port map( A1 => n7493, A2 => n7491, A3 => n28219, ZN => 
                           n9313);
   U572 : AND3_X2 port map( A1 => n983, A2 => n3736, A3 => n7459, ZN => n8320);
   U575 : XNOR2_X2 port map( A => n100, B => n2113, ZN => n14400);
   U576 : XNOR2_X1 port map( A => n12448, B => n12449, ZN => n100);
   U582 : NAND3_X2 port map( A1 => n101, A2 => n1602, A3 => n1601, ZN => n19452
                           );
   U583 : NAND2_X1 port map( A1 => n18088, A2 => n527, ZN => n101);
   U584 : INV_X1 port map( A => n20560, ZN => n20561);
   U585 : NAND2_X1 port map( A1 => n19849, A2 => n20208, ZN => n20560);
   U586 : NAND3_X1 port map( A1 => n23182, A2 => n23181, A3 => n28765, ZN => 
                           n24241);
   U589 : NAND2_X1 port map( A1 => n948, A2 => n4913, ZN => n951);
   U591 : NAND3_X1 port map( A1 => n24016, A2 => n4639, A3 => n5799, ZN => 
                           n6215);
   U594 : AND4_X2 port map( A1 => n11286, A2 => n10381, A3 => n10380, A4 => 
                           n10379, ZN => n12176);
   U598 : NAND2_X1 port map( A1 => n15271, A2 => n5948, ZN => n15956);
   U599 : AND2_X1 port map( A1 => n17564, A2 => n17772, ZN => n17577);
   U602 : NAND3_X1 port map( A1 => n104, A2 => n5623, A3 => n4732, ZN => n17329
                           );
   U603 : NAND2_X1 port map( A1 => n18138, A2 => n18137, ZN => n104);
   U605 : NAND3_X1 port map( A1 => n1798, A2 => n1799, A3 => n6500, ZN => 
                           n18193);
   U606 : OAI21_X2 port map( B1 => n18751, B2 => n20087, A => n18750, ZN => 
                           n21000);
   U607 : NAND3_X1 port map( A1 => n8701, A2 => n8703, A3 => n105, ZN => n10231
                           );
   U610 : OAI21_X1 port map( B1 => n20793, B2 => n107, A => n21198, ZN => 
                           n20796);
   U611 : NOR2_X1 port map( A1 => n21512, A2 => n21199, ZN => n107);
   U613 : NAND2_X1 port map( A1 => n17861, A2 => n18511, ZN => n5228);
   U614 : NAND2_X1 port map( A1 => n10838, A2 => n10835, ZN => n10836);
   U625 : XNOR2_X1 port map( A => n109, B => n2509, ZN => Ciphertext(140));
   U626 : NAND3_X1 port map( A1 => n26524, A2 => n26525, A3 => n26523, ZN => 
                           n109);
   U632 : XNOR2_X2 port map( A => n16562, B => n16561, ZN => n17106);
   U645 : XNOR2_X2 port map( A => n9486, B => n9485, ZN => n11318);
   U648 : NOR2_X1 port map( A1 => n29595, A2 => n18423, ZN => n111);
   U649 : INV_X1 port map( A => n4805, ZN => n112);
   U650 : NAND2_X1 port map( A1 => n17822, A2 => n29594, ZN => n113);
   U651 : NOR3_X1 port map( A1 => n21692, A2 => n21348, A3 => n6314, ZN => 
                           n20963);
   U653 : XNOR2_X1 port map( A => n22338, B => n22717, ZN => n22519);
   U656 : NAND2_X2 port map( A1 => n1207, A2 => n8901, ZN => n10328);
   U658 : NAND3_X1 port map( A1 => n1651, A2 => n8897, A3 => n29304, ZN => 
                           n1714);
   U660 : OAI22_X1 port map( A1 => n7716, A2 => n8134, B1 => n7718, B2 => 
                           n29646, ZN => n2506);
   U662 : MUX2_X2 port map( A => n11448, B => n11447, S => n12361, Z => n13166)
                           ;
   U663 : NAND2_X1 port map( A1 => n12115, A2 => n6281, ZN => n12113);
   U667 : NAND2_X1 port map( A1 => n8861, A2 => n4585, ZN => n4584);
   U668 : NOR2_X1 port map( A1 => n8378, A2 => n9075, ZN => n8861);
   U671 : NAND3_X1 port map( A1 => n10718, A2 => n11137, A3 => n11142, ZN => 
                           n10107);
   U672 : NOR2_X1 port map( A1 => n27615, A2 => n114, ZN => n27623);
   U674 : NAND2_X1 port map( A1 => n479, A2 => n23419, ZN => n22806);
   U679 : NAND2_X1 port map( A1 => n13642, A2 => n13641, ZN => n16322);
   U681 : NAND2_X1 port map( A1 => n8536, A2 => n8734, ZN => n8542);
   U682 : NAND2_X1 port map( A1 => n3558, A2 => n12058, ZN => n11295);
   U689 : NAND3_X1 port map( A1 => n5552, A2 => n23222, A3 => n5553, ZN => 
                           n24538);
   U698 : OAI211_X1 port map( C1 => n27746, C2 => n27736, A => n119, B => n118,
                           ZN => n27738);
   U699 : NAND2_X1 port map( A1 => n27733, A2 => n27749, ZN => n118);
   U700 : NAND2_X1 port map( A1 => n27734, A2 => n27757, ZN => n119);
   U701 : NAND3_X1 port map( A1 => n8006, A2 => n120, A3 => n9099, ZN => n8005)
                           ;
   U702 : NAND2_X1 port map( A1 => n9100, A2 => n8664, ZN => n120);
   U704 : NAND3_X1 port map( A1 => n8168, A2 => n8159, A3 => n8158, ZN => n8164
                           );
   U705 : NAND2_X1 port map( A1 => n121, A2 => n14802, ZN => n3287);
   U706 : NAND2_X1 port map( A1 => n3506, A2 => n3507, ZN => n121);
   U709 : NAND3_X1 port map( A1 => n1181, A2 => n4681, A3 => n17275, ZN => 
                           n4613);
   U710 : BUF_X1 port map( A => n7198, Z => n7406);
   U720 : NAND2_X1 port map( A1 => n10549, A2 => n10492, ZN => n11112);
   U722 : INV_X1 port map( A => n18190, ZN => n122);
   U723 : INV_X1 port map( A => n18188, ZN => n123);
   U726 : NAND2_X1 port map( A1 => n11609, A2 => n4404, ZN => n125);
   U732 : NAND2_X1 port map( A1 => n29321, A2 => n8024, ZN => n8022);
   U734 : NAND2_X1 port map( A1 => n21007, A2 => n4266, ZN => n2343);
   U736 : OAI22_X1 port map( A1 => n8708, A2 => n8876, B1 => n8710, B2 => n8709
                           , ZN => n127);
   U737 : NAND2_X1 port map( A1 => n415, A2 => n128, ZN => n6840);
   U738 : NAND2_X1 port map( A1 => n7843, A2 => n8024, ZN => n7010);
   U739 : NAND3_X1 port map( A1 => n10453, A2 => n130, A3 => n287, ZN => n6330)
                           ;
   U741 : INV_X1 port map( A => n11881, ZN => n130);
   U743 : NAND3_X2 port map( A1 => n16552, A2 => n16551, A3 => n16553, ZN => 
                           n18354);
   U749 : NAND2_X1 port map( A1 => n24893, A2 => n24532, ZN => n132);
   U752 : NAND3_X1 port map( A1 => n9362, A2 => n10959, A3 => n10686, ZN => 
                           n897);
   U763 : NOR2_X1 port map( A1 => n6424, A2 => n23772, ZN => n136);
   U765 : NAND3_X1 port map( A1 => n6709, A2 => n26907, A3 => n6710, ZN => 
                           n6708);
   U767 : AND3_X2 port map( A1 => n3720, A2 => n6887, A3 => n6888, ZN => n27457
                           );
   U769 : XNOR2_X1 port map( A => n19331, B => n19408, ZN => n19119);
   U771 : NOR2_X1 port map( A1 => n22967, A2 => n137, ZN => n22968);
   U772 : NOR2_X1 port map( A1 => n6686, A2 => n23127, ZN => n137);
   U776 : NAND2_X2 port map( A1 => n2620, A2 => n138, ZN => n24347);
   U780 : NAND2_X1 port map( A1 => n8574, A2 => n8579, ZN => n8767);
   U782 : NOR2_X2 port map( A1 => n13820, A2 => n13819, ZN => n16366);
   U784 : NAND2_X1 port map( A1 => n3089, A2 => n10916, ZN => n139);
   U786 : NAND3_X1 port map( A1 => n141, A2 => n12140, A3 => n140, ZN => n15407
                           );
   U793 : NAND2_X1 port map( A1 => n21425, A2 => n5827, ZN => n21086);
   U798 : NAND2_X1 port map( A1 => n626, A2 => n8217, ZN => n8215);
   U799 : NAND2_X1 port map( A1 => n144, A2 => n143, ZN => n5492);
   U800 : AOI21_X1 port map( B1 => n18465, B2 => n6079, A => n18471, ZN => n143
                           );
   U801 : NAND2_X1 port map( A1 => n145, A2 => n17916, ZN => n144);
   U802 : OR2_X2 port map( A1 => n14588, A2 => n14587, ZN => n16257);
   U803 : NAND2_X1 port map( A1 => n148, A2 => n147, ZN => n146);
   U804 : NAND2_X1 port map( A1 => n24683, A2 => n23902, ZN => n147);
   U806 : INV_X1 port map( A => n24683, ZN => n149);
   U807 : NAND2_X1 port map( A1 => n21564, A2 => n21563, ZN => n21115);
   U808 : NAND2_X1 port map( A1 => n20756, A2 => n21565, ZN => n21563);
   U810 : AOI21_X1 port map( B1 => n17002, B2 => n17276, A => n17272, ZN => 
                           n15981);
   U812 : XNOR2_X1 port map( A => n9577, B => n9878, ZN => n10123);
   U814 : NAND2_X1 port map( A1 => n3230, A2 => n3231, ZN => n27958);
   U822 : AND2_X1 port map( A1 => n15060, A2 => n15360, ZN => n15357);
   U833 : NAND2_X1 port map( A1 => n6761, A2 => n1315, ZN => n1314);
   U837 : OR2_X2 port map( A1 => n8487, A2 => n8486, ZN => n9125);
   U839 : OR2_X1 port map( A1 => n14106, A2 => n14107, ZN => n14235);
   U843 : NAND2_X1 port map( A1 => n1003, A2 => n1004, ZN => n1002);
   U845 : AOI21_X1 port map( B1 => n208, B2 => n7943, A => n29317, ZN => n155);
   U847 : AOI22_X2 port map( A1 => n17372, A2 => n17371, B1 => n17370, B2 => 
                           n17369, ZN => n18404);
   U848 : OR2_X1 port map( A1 => n14842, A2 => n14600, ZN => n14071);
   U850 : XNOR2_X1 port map( A => n156, B => n26590, ZN => Ciphertext(48));
   U851 : NAND4_X1 port map( A1 => n5367, A2 => n5369, A3 => n26589, A4 => 
                           n26588, ZN => n156);
   U855 : NOR2_X1 port map( A1 => n23179, A2 => n157, ZN => n23182);
   U856 : NOR3_X1 port map( A1 => n1838, A2 => n23645, A3 => n23640, ZN => n157
                           );
   U858 : NAND3_X1 port map( A1 => n5035, A2 => n25453, A3 => n29100, ZN => 
                           n25470);
   U859 : NAND2_X1 port map( A1 => n2418, A2 => n2420, ZN => n9190);
   U863 : OAI21_X1 port map( B1 => n21420, B2 => n20806, A => n20805, ZN => 
                           n20807);
   U864 : NOR2_X1 port map( A1 => n5000, A2 => n20899, ZN => n21420);
   U865 : NAND2_X1 port map( A1 => n15464, A2 => n15160, ZN => n785);
   U867 : NAND2_X1 port map( A1 => n18478, A2 => n18304, ZN => n18309);
   U871 : BUF_X1 port map( A => n10534, Z => n10659);
   U873 : NAND3_X1 port map( A1 => n14385, A2 => n14382, A3 => n14381, ZN => 
                           n14383);
   U875 : XNOR2_X1 port map( A => n29580, B => n19637, ZN => n19430);
   U877 : XNOR2_X1 port map( A => n21789, B => n22094, ZN => n22689);
   U878 : AND2_X2 port map( A1 => n20927, A2 => n4566, ZN => n21789);
   U887 : OAI21_X1 port map( B1 => n21163, B2 => n4148, A => n21609, ZN => n159
                           );
   U890 : NAND3_X1 port map( A1 => n24412, A2 => n24711, A3 => n24714, ZN => 
                           n24413);
   U893 : NAND2_X1 port map( A1 => n161, A2 => n20858, ZN => n20530);
   U894 : NAND2_X1 port map( A1 => n21157, A2 => n21159, ZN => n161);
   U898 : NAND2_X2 port map( A1 => n23015, A2 => n3743, ZN => n24682);
   U899 : AOI21_X2 port map( B1 => n20489, B2 => n20488, A => n20487, ZN => 
                           n21611);
   U900 : NAND4_X2 port map( A1 => n2653, A2 => n5477, A3 => n2651, A4 => n2650
                           , ZN => n22633);
   U903 : OR2_X2 port map( A1 => n6537, A2 => n23056, ZN => n24713);
   U909 : BUF_X1 port map( A => n23010, Z => n23011);
   U913 : NAND2_X1 port map( A1 => n8930, A2 => n9147, ZN => n8935);
   U914 : XNOR2_X2 port map( A => Key(1), B => Plaintext(1), ZN => n7890);
   U915 : OR2_X1 port map( A1 => n8658, A2 => n8116, ZN => n8497);
   U916 : AND3_X2 port map( A1 => n23076, A2 => n1206, A3 => n3337, ZN => 
                           n24374);
   U918 : AOI22_X1 port map( A1 => n27001, A2 => n27045, B1 => n27003, B2 => 
                           n27002, ZN => n27009);
   U920 : NAND3_X1 port map( A1 => n5291, A2 => n23283, A3 => n6279, ZN => 
                           n5293);
   U921 : NAND2_X1 port map( A1 => n25423, A2 => n25424, ZN => n25425);
   U922 : OAI22_X1 port map( A1 => n23850, A2 => n24100, B1 => n23875, B2 => 
                           n24489, ZN => n162);
   U923 : NAND2_X1 port map( A1 => n377, A2 => n26560, ZN => n948);
   U924 : NAND3_X1 port map( A1 => n14065, A2 => n14064, A3 => n14325, ZN => 
                           n3125);
   U925 : NAND2_X1 port map( A1 => n694, A2 => n15335, ZN => n693);
   U926 : NAND2_X1 port map( A1 => n3415, A2 => n3416, ZN => n17782);
   U936 : XNOR2_X1 port map( A => n165, B => n8573, ZN => n11199);
   U937 : XNOR2_X1 port map( A => n9668, B => n9940, ZN => n165);
   U941 : NOR2_X1 port map( A1 => n6941, A2 => n167, ZN => n23065);
   U942 : NOR2_X1 port map( A1 => n23147, A2 => n1837, ZN => n167);
   U947 : NAND2_X1 port map( A1 => n14780, A2 => n15432, ZN => n168);
   U948 : NAND2_X1 port map( A1 => n14779, A2 => n15030, ZN => n169);
   U953 : AOI21_X1 port map( B1 => n170, B2 => n20618, A => n20616, ZN => 
                           n19923);
   U954 : NAND2_X1 port map( A1 => n20617, A2 => n500, ZN => n170);
   U955 : NAND3_X1 port map( A1 => n171, A2 => n24760, A3 => n378, ZN => n24763
                           );
   U958 : OAI211_X2 port map( C1 => n13908, C2 => n14051, A => n5730, B => 
                           n5386, ZN => n13922);
   U959 : XNOR2_X2 port map( A => n16584, B => n16583, ZN => n17470);
   U960 : BUF_X2 port map( A => n10939, Z => n11952);
   U961 : OAI211_X2 port map( C1 => n19778, C2 => n19777, A => n5075, B => 
                           n5074, ZN => n21140);
   U969 : OAI22_X1 port map( A1 => n17823, A2 => n512, B1 => n4802, B2 => 
                           n17824, ZN => n174);
   U978 : AND3_X2 port map( A1 => n3535, A2 => n941, A3 => n939, ZN => n18195);
   U979 : AND2_X2 port map( A1 => n6120, A2 => n6121, ZN => n25396);
   U983 : NAND2_X1 port map( A1 => n1178, A2 => n2390, ZN => n20298);
   U986 : NAND3_X1 port map( A1 => n3291, A2 => n23601, A3 => n3292, ZN => 
                           n24870);
   U987 : NAND4_X2 port map( A1 => n175, A2 => n11015, A3 => n11016, A4 => 
                           n11018, ZN => n12253);
   U988 : NAND2_X1 port map( A1 => n1999, A2 => n6108, ZN => n175);
   U989 : MUX2_X1 port map( A => n18215, B => n18506, S => n18213, Z => n17728)
                           ;
   U991 : XNOR2_X2 port map( A => n12910, B => n12909, ZN => n14287);
   U992 : NAND2_X1 port map( A1 => n12402, A2 => n12407, ZN => n11800);
   U993 : OR2_X2 port map( A1 => n4462, A2 => n4461, ZN => n12402);
   U998 : INV_X1 port map( A => n10250, ZN => n9674);
   U1003 : OAI21_X2 port map( B1 => n22448, B2 => n1740, A => n178, ZN => 
                           n24734);
   U1004 : NAND2_X1 port map( A1 => n639, A2 => n23192, ZN => n178);
   U1005 : NAND2_X1 port map( A1 => n1040, A2 => n1082, ZN => n19887);
   U1006 : NAND3_X1 port map( A1 => n15448, A2 => n15322, A3 => n15446, ZN => 
                           n15016);
   U1007 : INV_X1 port map( A => n8925, ZN => n7403);
   U1008 : NAND2_X1 port map( A1 => n9340, A2 => n6718, ZN => n8925);
   U1009 : XNOR2_X1 port map( A => n18756, B => n27225, ZN => n18704);
   U1010 : BUF_X1 port map( A => n25120, Z => n27182);
   U1011 : AOI21_X2 port map( B1 => n26402, B2 => n26401, A => n26400, ZN => 
                           n27561);
   U1012 : XNOR2_X2 port map( A => n12643, B => n12642, ZN => n14451);
   U1013 : OAI21_X2 port map( B1 => n15688, B2 => n2133, A => n15687, ZN => 
                           n18490);
   U1014 : OAI22_X1 port map( A1 => n24118, A2 => n24435, B1 => n23886, B2 => 
                           n24119, ZN => n24122);
   U1015 : NAND2_X1 port map( A1 => n5837, A2 => n179, ZN => n6850);
   U1016 : NAND2_X1 port map( A1 => n4341, A2 => n11195, ZN => n5837);
   U1020 : XNOR2_X1 port map( A => n16594, B => n16595, ZN => n180);
   U1021 : XNOR2_X1 port map( A => n181, B => n9254, ZN => n9608);
   U1022 : XNOR2_X1 port map( A => n9241, B => n9242, ZN => n181);
   U1026 : NAND2_X1 port map( A1 => n24551, A2 => n24555, ZN => n24550);
   U1028 : AND3_X2 port map( A1 => n182, A2 => n3754, A3 => n26399, ZN => 
                           n27203);
   U1029 : OAI21_X1 port map( B1 => n25122, B2 => n25123, A => n25034, ZN => 
                           n182);
   U1030 : OAI21_X1 port map( B1 => n15099, B2 => n14677, A => n183, ZN => 
                           n14682);
   U1031 : OAI211_X2 port map( C1 => n24553, C2 => n24174, A => n5510, B => 
                           n5508, ZN => n26083);
   U1032 : OAI21_X1 port map( B1 => n14170, B2 => n14169, A => n14167, ZN => 
                           n4073);
   U1038 : NAND3_X1 port map( A1 => n8492, A2 => n8630, A3 => n9100, ZN => 
                           n8493);
   U1039 : NOR2_X2 port map( A1 => n16929, A2 => n16930, ZN => n19272);
   U1040 : OAI211_X1 port map( C1 => n12159, C2 => n12241, A => n187, B => 
                           n12037, ZN => n4615);
   U1041 : NAND2_X1 port map( A1 => n188, A2 => n12241, ZN => n187);
   U1042 : INV_X1 port map( A => n12244, ZN => n188);
   U1048 : NAND2_X1 port map( A1 => n191, A2 => n190, ZN => n189);
   U1049 : NAND2_X1 port map( A1 => n14176, A2 => n14177, ZN => n191);
   U1050 : NAND2_X1 port map( A1 => n14179, A2 => n14452, ZN => n192);
   U1052 : NAND2_X1 port map( A1 => n193, A2 => n18138, ZN => n914);
   U1055 : NAND3_X1 port map( A1 => n29086, A2 => n29559, A3 => n17101, ZN => 
                           n17103);
   U1056 : NAND3_X1 port map( A1 => n11114, A2 => n29627, A3 => n28205, ZN => 
                           n2867);
   U1057 : NAND2_X2 port map( A1 => n5739, A2 => n5740, ZN => n5234);
   U1059 : NAND3_X2 port map( A1 => n2405, A2 => n8306, A3 => n8307, ZN => 
                           n8955);
   U1062 : NAND2_X1 port map( A1 => n21230, A2 => n21408, ZN => n195);
   U1064 : OAI22_X1 port map( A1 => n17693, A2 => n18516, B1 => n18270, B2 => 
                           n418, ZN => n17694);
   U1066 : NAND3_X2 port map( A1 => n6915, A2 => n2915, A3 => n9038, ZN => 
                           n10350);
   U1068 : AND3_X2 port map( A1 => n866, A2 => n275, A3 => n865, ZN => n25381);
   U1071 : NAND3_X1 port map( A1 => n9027, A2 => n9031, A3 => n9028, ZN => 
                           n9033);
   U1074 : NAND3_X1 port map( A1 => n22084, A2 => n6099, A3 => n28428, ZN => 
                           n6585);
   U1075 : NAND3_X1 port map( A1 => n197, A2 => n4924, A3 => n4919, ZN => n4918
                           );
   U1076 : NAND2_X1 port map( A1 => n27243, A2 => n27402, ZN => n197);
   U1078 : NOR2_X1 port map( A1 => n5697, A2 => n198, ZN => n5696);
   U1079 : NOR2_X1 port map( A1 => n199, A2 => n5530, ZN => n198);
   U1080 : NAND2_X1 port map( A1 => n201, A2 => n23301, ZN => n199);
   U1082 : INV_X1 port map( A => n22686, ZN => n201);
   U1085 : NOR2_X2 port map( A1 => n202, A2 => n24355, ZN => n25149);
   U1086 : OAI21_X1 port map( B1 => n24353, B2 => n28416, A => n24352, ZN => 
                           n202);
   U1089 : NAND3_X1 port map( A1 => n7010, A2 => n6299, A3 => n29106, ZN => 
                           n7014);
   U1092 : NAND2_X1 port map( A1 => n204, A2 => n7163, ZN => n2692);
   U1093 : NOR2_X1 port map( A1 => n614, A2 => n7770, ZN => n204);
   U1094 : NAND2_X1 port map( A1 => n7585, A2 => n7580, ZN => n7074);
   U1097 : NAND3_X1 port map( A1 => n17905, A2 => n3866, A3 => n17903, ZN => 
                           n3864);
   U1099 : XNOR2_X2 port map( A => n6986, B => Key(90), ZN => n7424);
   U1102 : NAND3_X1 port map( A1 => n1338, A2 => n3817, A3 => n11033, ZN => 
                           n1336);
   U1103 : AND3_X2 port map( A1 => n19009, A2 => n19008, A3 => n19007, ZN => 
                           n21287);
   U1107 : NAND2_X1 port map( A1 => n29547, A2 => n18410, ZN => n18027);
   U1113 : MUX2_X1 port map( A => n11990, B => n10863, S => n12512, Z => n10117
                           );
   U1117 : NAND2_X2 port map( A1 => n23374, A2 => n205, ZN => n25931);
   U1119 : OR2_X2 port map( A1 => n7461, A2 => n7460, ZN => n8605);
   U1120 : NAND2_X1 port map( A1 => n207, A2 => n206, ZN => n20596);
   U1121 : NAND2_X1 port map( A1 => n21591, A2 => n21322, ZN => n206);
   U1122 : NAND2_X1 port map( A1 => n20575, A2 => n20889, ZN => n207);
   U1123 : NAND2_X1 port map( A1 => n8301, A2 => n7942, ZN => n208);
   U1127 : NAND3_X1 port map( A1 => n5233, A2 => n18393, A3 => n17766, ZN => 
                           n5232);
   U1129 : NAND2_X1 port map( A1 => n4266, A2 => n20698, ZN => n19733);
   U1133 : OAI211_X1 port map( C1 => n27858, C2 => n447, A => n209, B => n4533,
                           ZN => n4535);
   U1134 : INV_X1 port map( A => n210, ZN => n209);
   U1135 : OAI22_X1 port map( A1 => n26646, A2 => n29095, B1 => n27859, B2 => 
                           n27851, ZN => n210);
   U1136 : OAI211_X1 port map( C1 => n17463, C2 => n28800, A => n528, B => 
                           n17280, ZN => n4286);
   U1137 : AOI22_X2 port map( A1 => n18338, A2 => n18339, B1 => n18336, B2 => 
                           n18337, ZN => n19384);
   U1139 : OAI22_X1 port map( A1 => n212, A2 => n211, B1 => n17057, B2 => 
                           n17542, ZN => n17059);
   U1140 : INV_X1 port map( A => n17055, ZN => n211);
   U1141 : NAND2_X1 port map( A1 => n17213, A2 => n15787, ZN => n212);
   U1144 : NAND3_X1 port map( A1 => n20628, A2 => n28186, A3 => n20623, ZN => 
                           n6883);
   U1145 : NAND2_X1 port map( A1 => n213, A2 => n3279, ZN => n7646);
   U1146 : NAND2_X1 port map( A1 => n251, A2 => n7985, ZN => n213);
   U1148 : NAND2_X1 port map( A1 => n4856, A2 => n7100, ZN => n7761);
   U1151 : AND3_X2 port map( A1 => n216, A2 => n1363, A3 => n215, ZN => n18087)
                           ;
   U1152 : NAND2_X1 port map( A1 => n16823, A2 => n17710, ZN => n215);
   U1153 : NAND2_X1 port map( A1 => n1366, A2 => n1365, ZN => n216);
   U1154 : OR2_X2 port map( A1 => n5465, A2 => n11615, ZN => n13450);
   U1157 : NAND2_X1 port map( A1 => n1909, A2 => n8058, ZN => n8352);
   U1158 : NAND3_X1 port map( A1 => n7765, A2 => n4855, A3 => n7764, ZN => 
                           n1909);
   U1161 : NAND4_X2 port map( A1 => n11745, A2 => n12360, A3 => n11744, A4 => 
                           n11743, ZN => n13039);
   U1166 : OR2_X1 port map( A1 => n7909, A2 => n8290, ZN => n2898);
   U1171 : NAND2_X1 port map( A1 => n15400, A2 => n28518, ZN => n13636);
   U1172 : OAI21_X1 port map( B1 => n1285, B2 => n10681, A => n10680, ZN => 
                           n10682);
   U1173 : NAND2_X1 port map( A1 => n1285, A2 => n28608, ZN => n10680);
   U1174 : NAND2_X1 port map( A1 => n16550, A2 => n16547, ZN => n699);
   U1176 : XNOR2_X2 port map( A => n1756, B => n1755, ZN => n20511);
   U1179 : NAND2_X1 port map( A1 => n1255, A2 => n14498, ZN => n2488);
   U1182 : AND2_X2 port map( A1 => n6527, A2 => n6531, ZN => n22271);
   U1184 : NAND2_X1 port map( A1 => n221, A2 => n220, ZN => n219);
   U1185 : NAND2_X1 port map( A1 => n4685, A2 => n5004, ZN => n221);
   U1186 : AOI21_X1 port map( B1 => n223, B2 => n15409, A => n15108, ZN => 
                           n3918);
   U1187 : INV_X1 port map( A => n3922, ZN => n223);
   U1188 : BUF_X2 port map( A => n17687, Z => n20941);
   U1195 : AND3_X2 port map( A1 => n874, A2 => n1518, A3 => n1613, ZN => n15668
                           );
   U1196 : NAND3_X1 port map( A1 => n1643, A2 => n29138, A3 => n6306, ZN => 
                           n1306);
   U1197 : NAND2_X1 port map( A1 => n26428, A2 => n26381, ZN => n26429);
   U1198 : XNOR2_X2 port map( A => n7122, B => Key(38), ZN => n8141);
   U1206 : NAND3_X1 port map( A1 => n7827, A2 => n7825, A3 => n7824, ZN => 
                           n7826);
   U1208 : NAND3_X1 port map( A1 => n5604, A2 => n5605, A3 => n225, ZN => n2380
                           );
   U1215 : NAND2_X1 port map( A1 => n226, A2 => n5956, ZN => n1020);
   U1216 : NAND2_X1 port map( A1 => n794, A2 => n13647, ZN => n226);
   U1218 : OAI21_X1 port map( B1 => n17210, B2 => n17824, A => n227, ZN => 
                           n5551);
   U1223 : NAND3_X2 port map( A1 => n5960, A2 => n8528, A3 => n5959, ZN => 
                           n9755);
   U1227 : NOR2_X1 port map( A1 => n23083, A2 => n23082, ZN => n1777);
   U1232 : NAND2_X1 port map( A1 => n4484, A2 => n229, ZN => n5080);
   U1233 : OAI21_X1 port map( B1 => n23845, B2 => n23722, A => n23721, ZN => 
                           n229);
   U1240 : NAND3_X1 port map( A1 => n7685, A2 => n7843, A3 => n7515, ZN => 
                           n7519);
   U1241 : AND2_X1 port map( A1 => n28451, A2 => n27244, ZN => n27948);
   U1244 : INV_X1 port map( A => n4880, ZN => n19283);
   U1245 : NAND2_X1 port map( A1 => n1231, A2 => n1232, ZN => n4880);
   U1246 : BUF_X1 port map( A => n8592, Z => n8978);
   U1247 : NAND2_X1 port map( A1 => n5389, A2 => n29481, ZN => n5388);
   U1249 : INV_X1 port map( A => n15071, ZN => n14639);
   U1250 : NAND4_X2 port map( A1 => n12940, A2 => n12939, A3 => n12941, A4 => 
                           n6562, ZN => n15071);
   U1251 : NAND3_X1 port map( A1 => n6479, A2 => n11486, A3 => n4744, ZN => 
                           n11306);
   U1257 : NAND3_X1 port map( A1 => n12190, A2 => n2483, A3 => n11724, ZN => 
                           n11723);
   U1258 : NAND2_X1 port map( A1 => n232, A2 => n5148, ZN => n5147);
   U1259 : NAND3_X1 port map( A1 => n7868, A2 => n7173, A3 => n7867, ZN => n232
                           );
   U1260 : BUF_X1 port map( A => n7233, Z => n7592);
   U1261 : NAND2_X1 port map( A1 => n17939, A2 => n17601, ZN => n17943);
   U1262 : OAI211_X2 port map( C1 => n16151, C2 => n16853, A => n16150, B => 
                           n3587, ZN => n17939);
   U1266 : NAND3_X1 port map( A1 => n705, A2 => n706, A3 => n12167, ZN => n233)
                           ;
   U1270 : NAND2_X2 port map( A1 => n4268, A2 => n4267, ZN => n21253);
   U1272 : XNOR2_X2 port map( A => n6979, B => Key(99), ZN => n7635);
   U1277 : AND2_X2 port map( A1 => n1469, A2 => n1471, ZN => n27340);
   U1280 : NAND3_X1 port map( A1 => n8856, A2 => n8857, A3 => n28212, ZN => 
                           n881);
   U1282 : OAI21_X1 port map( B1 => n2549, B2 => n13877, A => n235, ZN => n2607
                           );
   U1283 : NAND2_X1 port map( A1 => n13877, A2 => n14402, ZN => n235);
   U1285 : NAND2_X1 port map( A1 => n237, A2 => n17435, ZN => n4427);
   U1287 : OAI21_X1 port map( B1 => n8428, B2 => n1909, A => n238, ZN => n8432)
                           ;
   U1293 : AND2_X1 port map( A1 => n21000, A2 => n20972, ZN => n20968);
   U1295 : NAND2_X1 port map( A1 => n16774, A2 => n17016, ZN => n16865);
   U1296 : OAI211_X2 port map( C1 => n7927, C2 => n8216, A => n2556, B => n7627
                           , ZN => n9200);
   U1297 : NAND4_X2 port map( A1 => n16793, A2 => n16796, A3 => n16794, A4 => 
                           n16795, ZN => n19549);
   U1300 : AOI22_X1 port map( A1 => n28437, A2 => n27120, B1 => n26512, B2 => 
                           n402, ZN => n27122);
   U1302 : OAI22_X1 port map( A1 => n18749, A2 => n19755, B1 => n29114, B2 => 
                           n20040, ZN => n18750);
   U1303 : NAND2_X1 port map( A1 => n29104, A2 => n20090, ZN => n19755);
   U1304 : NAND2_X1 port map( A1 => n15125, A2 => n14998, ZN => n13985);
   U1311 : NAND3_X2 port map( A1 => n4619, A2 => n4620, A3 => n4622, ZN => 
                           n16377);
   U1318 : NAND2_X1 port map( A1 => n8926, A2 => n9131, ZN => n240);
   U1319 : BUF_X2 port map( A => n26374, Z => n26950);
   U1327 : NAND3_X1 port map( A1 => n11291, A2 => n11077, A3 => n11076, ZN => 
                           n4352);
   U1332 : NAND2_X1 port map( A1 => n11115, A2 => n11114, ZN => n243);
   U1335 : NAND4_X2 port map( A1 => n8697, A2 => n8694, A3 => n8695, A4 => 
                           n8696, ZN => n10232);
   U1350 : MUX2_X2 port map( A => n15524, B => n15523, S => n18478, Z => n19495
                           );
   U1351 : NAND3_X1 port map( A1 => n29475, A2 => n6419, A3 => n5188, ZN => 
                           n26317);
   U1352 : XNOR2_X2 port map( A => n4961, B => n12918, ZN => n14285);
   U1355 : NAND2_X1 port map( A1 => n14761, A2 => n14762, ZN => n14765);
   U1356 : OAI211_X2 port map( C1 => n21129, C2 => n21497, A => n21128, B => 
                           n244, ZN => n22409);
   U1357 : NAND3_X1 port map( A1 => n21126, A2 => n21127, A3 => n21497, ZN => 
                           n244);
   U1360 : NAND3_X1 port map( A1 => n530, A2 => n29636, A3 => n17379, ZN => 
                           n16876);
   U1363 : AOI21_X1 port map( B1 => n28761, B2 => n28200, A => n245, ZN => 
                           n2295);
   U1365 : NAND3_X2 port map( A1 => n248, A2 => n8423, A3 => n8424, ZN => 
                           n12202);
   U1368 : OAI21_X1 port map( B1 => n250, B2 => n8223, A => n249, ZN => n8226);
   U1369 : NAND2_X1 port map( A1 => n8223, A2 => n8224, ZN => n249);
   U1370 : INV_X1 port map( A => n8225, ZN => n250);
   U1371 : OAI21_X1 port map( B1 => n15102, B2 => n15105, A => n14936, ZN => 
                           n6022);
   U1373 : NAND2_X1 port map( A1 => n5838, A2 => n11622, ZN => n6705);
   U1374 : NAND3_X1 port map( A1 => n4926, A2 => n4925, A3 => n26820, ZN => 
                           n3263);
   U1376 : NAND2_X1 port map( A1 => n7191, A2 => n7641, ZN => n251);
   U1379 : OAI21_X1 port map( B1 => n4100, B2 => n16911, A => n252, ZN => 
                           n15848);
   U1380 : NAND2_X1 port map( A1 => n4099, A2 => n16911, ZN => n252);
   U1382 : OR2_X1 port map( A1 => n11330, A2 => n10821, ZN => n5366);
   U1385 : OR2_X2 port map( A1 => n6485, A2 => n5732, ZN => n18353);
   U1386 : OR2_X2 port map( A1 => n10845, A2 => n10846, ZN => n4617);
   U1387 : XNOR2_X1 port map( A => n253, B => n11575, ZN => n11577);
   U1395 : OAI211_X1 port map( C1 => n26603, C2 => n6859, A => n2053, B => n255
                           , ZN => n6858);
   U1396 : NAND2_X1 port map( A1 => n28026, A2 => n28030, ZN => n255);
   U1401 : NAND2_X1 port map( A1 => n1599, A2 => n14471, ZN => n1598);
   U1403 : NAND2_X1 port map( A1 => n3914, A2 => n17197, ZN => n18414);
   U1404 : AND2_X2 port map( A1 => n2705, A2 => n2704, ZN => n19511);
   U1406 : NAND2_X1 port map( A1 => n19981, A2 => n29066, ZN => n702);
   U1408 : MUX2_X2 port map( A => n25596, B => n25595, S => n29482, Z => n28035
                           );
   U1412 : XNOR2_X1 port map( A => n9754, B => n9992, ZN => n10376);
   U1414 : BUF_X1 port map( A => n26322, Z => n26992);
   U1417 : NAND2_X1 port map( A1 => n257, A2 => n24750, ZN => n2880);
   U1418 : OAI21_X1 port map( B1 => n24746, B2 => n28550, A => n4980, ZN => 
                           n257);
   U1421 : NAND2_X1 port map( A1 => n1527, A2 => n8760, ZN => n8759);
   U1425 : NAND3_X1 port map( A1 => n15315, A2 => n15319, A3 => n15308, ZN => 
                           n14855);
   U1428 : NAND2_X2 port map( A1 => n649, A2 => n19979, ZN => n4937);
   U1429 : NAND3_X2 port map( A1 => n14857, A2 => n1067, A3 => n14858, ZN => 
                           n16165);
   U1430 : NAND2_X1 port map( A1 => n398, A2 => n27041, ZN => n4487);
   U1433 : AOI22_X1 port map( A1 => n27886, A2 => n27885, B1 => n27884, B2 => 
                           n27923, ZN => n27888);
   U1436 : NOR2_X2 port map( A1 => n15590, A2 => n15589, ZN => n18292);
   U1439 : BUF_X1 port map( A => n15239, Z => n15234);
   U1440 : NAND3_X1 port map( A1 => n24531, A2 => n24894, A3 => n24530, ZN => 
                           n24537);
   U1441 : OR2_X1 port map( A1 => n7231, A2 => n441, ZN => n7871);
   U1443 : OAI21_X1 port map( B1 => n8899, B2 => n1793, A => n610, ZN => n1792)
                           ;
   U1444 : OAI211_X1 port map( C1 => n8908, C2 => n1770, A => n9016, B => n1769
                           , ZN => n1771);
   U1445 : OR2_X1 port map( A1 => n8752, A2 => n9529, ZN => n749);
   U1446 : NOR2_X1 port map( A1 => n8908, A2 => n9014, ZN => n8662);
   U1447 : AOI22_X1 port map( A1 => n8092, A2 => n9047, B1 => n5945, B2 => 
                           n8091, ZN => n9577);
   U1449 : XNOR2_X1 port map( A => n9749, B => n748, ZN => n9946);
   U1450 : AND2_X1 port map( A1 => n6779, A2 => n11004, ZN => n1380);
   U1451 : XNOR2_X1 port map( A => n1396, B => n1397, ZN => n11227);
   U1458 : XNOR2_X1 port map( A => n16131, B => n15854, ZN => n16267);
   U1459 : OR2_X1 port map( A1 => n28775, A2 => n17374, ZN => n4652);
   U1460 : AND2_X1 port map( A1 => n18493, A2 => n28633, ZN => n18495);
   U1461 : INV_X1 port map( A => n21047, ZN => n21412);
   U1464 : AND2_X1 port map( A1 => n23338, A2 => n29108, ZN => n1263);
   U1465 : XNOR2_X1 port map( A => n271, B => n22432, ZN => n23469);
   U1467 : OR2_X1 port map( A1 => n24765, A2 => n24767, ZN => n3054);
   U1469 : OR2_X1 port map( A1 => n6198, A2 => n630, ZN => n1301);
   U1471 : XNOR2_X1 port map( A => n277, B => n25212, ZN => n26480);
   U1472 : OR2_X1 port map( A1 => n26476, A2 => n26186, ZN => n24204);
   U1474 : INV_X1 port map( A => n29538, ZN => n27372);
   U1475 : AND3_X1 port map( A1 => n631, A2 => n8270, A3 => n7485, ZN => n258);
   U1476 : XOR2_X1 port map( A => n16603, B => n16476, Z => n259);
   U1477 : XOR2_X1 port map( A => n9505, B => n653, Z => n260);
   U1478 : AND3_X1 port map( A1 => n7765, A2 => n4855, A3 => n7764, ZN => n261)
                           ;
   U1479 : BUF_X1 port map( A => n10793, Z => n12155);
   U1481 : BUF_X1 port map( A => n17206, Z => n18129);
   U1482 : XNOR2_X1 port map( A => n25223, B => n25222, ZN => n26727);
   U1484 : AND3_X1 port map( A1 => n11069, A2 => n1851, A3 => n11243, ZN => 
                           n262);
   U1485 : NAND2_X2 port map( A1 => n5089, A2 => n10115, ZN => n12507);
   U1486 : AND2_X2 port map( A1 => n3941, A2 => n3942, ZN => n3946);
   U1489 : OR2_X1 port map( A1 => n13310, A2 => n13309, ZN => n263);
   U1494 : AND2_X1 port map( A1 => n14144, A2 => n2974, ZN => n265);
   U1495 : XOR2_X1 port map( A => n16313, B => n634, Z => n266);
   U1496 : NOR2_X2 port map( A1 => n13792, A2 => n13791, ZN => n15070);
   U1501 : AND2_X2 port map( A1 => n17036, A2 => n17035, ZN => n18332);
   U1502 : XOR2_X1 port map( A => n19622, B => n3728, Z => n267);
   U1504 : OR2_X1 port map( A1 => n20121, A2 => n20302, ZN => n268);
   U1506 : OR3_X1 port map( A1 => n21587, A2 => n21586, A3 => n21585, ZN => 
                           n269);
   U1507 : OR3_X1 port map( A1 => n22142, A2 => n21624, A3 => n22141, ZN => 
                           n270);
   U1509 : XOR2_X1 port map( A => n22430, B => n22429, Z => n271);
   U1511 : XOR2_X1 port map( A => n28450, B => n3622, Z => n272);
   U1512 : XOR2_X1 port map( A => n21947, B => n1538, Z => n274);
   U1514 : OR3_X1 port map( A1 => n23897, A2 => n25006, A3 => n25005, ZN => 
                           n276);
   U1515 : XOR2_X1 port map( A => n25211, B => n25467, Z => n277);
   U1517 : OR2_X1 port map( A1 => n28228, A2 => n925, ZN => n278);
   U1521 : XNOR2_X1 port map( A => n9546, B => n9545, ZN => n11037);
   U1523 : XNOR2_X1 port map( A => n24360, B => n24359, ZN => n26466);
   U1528 : XNOR2_X1 port map( A => n25292, B => n25291, ZN => n26717);
   U1539 : NAND4_X2 port map( A1 => n8567, A2 => n8568, A3 => n8566, A4 => 
                           n8565, ZN => n10436);
   U1542 : AOI22_X2 port map( A1 => n16921, A2 => n17414, B1 => n15811, B2 => 
                           n15522, ZN => n17679);
   U1551 : NOR2_X2 port map( A1 => n5967, A2 => n16769, ZN => n18109);
   U1552 : BUF_X1 port map( A => n23448, Z => n292);
   U1553 : XNOR2_X1 port map( A => n22739, B => n22738, ZN => n23448);
   U1557 : AND2_X1 port map( A1 => n11782, A2 => n11778, ZN => n11784);
   U1561 : OR2_X1 port map( A1 => n16807, A2 => n29574, ZN => n16672);
   U1564 : BUF_X1 port map( A => n27378, Z => n294);
   U1566 : OAI21_X1 port map( B1 => n5582, B2 => n26485, A => n26199, ZN => 
                           n27378);
   U1570 : XNOR2_X1 port map( A => n18965, B => n18964, ZN => n20224);
   U1575 : BUF_X2 port map( A => n26090, Z => n300);
   U1576 : INV_X1 port map( A => n26865, ZN => n401);
   U1578 : OAI211_X1 port map( C1 => n8795, C2 => n9034, A => n8794, B => n8793
                           , ZN => n10222);
   U1580 : XNOR2_X2 port map( A => n4531, B => n16007, ZN => n16977);
   U1582 : NAND2_X2 port map( A1 => n24563, A2 => n24562, ZN => n25947);
   U1584 : BUF_X1 port map( A => n12226, Z => n303);
   U1593 : BUF_X1 port map( A => n27028, Z => n307);
   U1594 : OAI22_X1 port map( A1 => n26925, A2 => n28711, B1 => n23864, B2 => 
                           n29552, ZN => n27028);
   U1595 : BUF_X2 port map( A => n14122, Z => n308);
   U1596 : XNOR2_X1 port map( A => n12959, B => n12958, ZN => n14122);
   U1598 : NAND3_X2 port map( A1 => n14503, A2 => n264, A3 => n14502, ZN => 
                           n16558);
   U1599 : XNOR2_X2 port map( A => n7086, B => Key(3), ZN => n7315);
   U1602 : AND3_X2 port map( A1 => n2709, A2 => n2710, A3 => n3553, ZN => 
                           n13445);
   U1606 : OR2_X1 port map( A1 => n29541, A2 => n27364, ZN => n799);
   U1607 : OR2_X1 port map( A1 => n27074, A2 => n29622, ZN => n3771);
   U1617 : OAI211_X1 port map( C1 => n14284, C2 => n14081, A => n13823, B => 
                           n13822, ZN => n14981);
   U1621 : XNOR2_X1 port map( A => n3582, B => n16169, ZN => n17466);
   U1623 : XNOR2_X2 port map( A => n21828, B => n21827, ZN => n23768);
   U1624 : AND2_X2 port map( A1 => n21725, A2 => n21724, ZN => n24747);
   U1626 : BUF_X1 port map( A => n16289, Z => n320);
   U1627 : OAI211_X1 port map( C1 => n4514, C2 => n4515, A => n5016, B => n4512
                           , ZN => n16289);
   U1628 : AND2_X1 port map( A1 => n26731, A2 => n26480, ZN => n26485);
   U1629 : NOR2_X2 port map( A1 => n6601, A2 => n5441, ZN => n22896);
   U1636 : BUF_X1 port map( A => n27718, Z => n326);
   U1637 : AOI21_X1 port map( B1 => n27690, B2 => n27688, A => n27687, ZN => 
                           n27718);
   U1640 : XNOR2_X2 port map( A => n1609, B => Key(25), ZN => n7792);
   U1641 : OAI22_X1 port map( A1 => n15032, A2 => n14825, B1 => n1644, B2 => 
                           n14826, ZN => n14780);
   U1646 : OAI21_X2 port map( B1 => n24136, B2 => n24135, A => n24134, ZN => 
                           n5275);
   U1649 : XNOR2_X1 port map( A => n24402, B => n24401, ZN => n26458);
   U1651 : XNOR2_X2 port map( A => n15672, B => n15671, ZN => n4218);
   U1652 : NAND2_X2 port map( A1 => n10909, A2 => n10910, ZN => n13414);
   U1654 : XNOR2_X2 port map( A => n4600, B => n9933, ZN => n11113);
   U1661 : AOI21_X2 port map( B1 => n15378, B2 => n15377, A => n15376, ZN => 
                           n16081);
   U1665 : AND3_X2 port map( A1 => n1477, A2 => n1479, A3 => n1476, ZN => 
                           n26029);
   U1666 : AOI21_X2 port map( B1 => n20775, B2 => n20774, A => n20773, ZN => 
                           n22219);
   U1671 : MUX2_X2 port map( A => n23237, B => n23236, S => n23716, Z => n24653
                           );
   U1674 : BUF_X1 port map( A => n337, Z => n336);
   U1675 : OAI21_X2 port map( B1 => n24083, B2 => n23506, A => n23505, ZN => 
                           n25751);
   U1681 : BUF_X2 port map( A => n23777, Z => n339);
   U1682 : NOR2_X2 port map( A1 => n18084, A2 => n6228, ZN => n19717);
   U1685 : BUF_X1 port map( A => n8269, Z => n341);
   U1686 : XNOR2_X1 port map( A => Key(147), B => Plaintext(147), ZN => n8269);
   U1687 : NAND3_X2 port map( A1 => n1392, A2 => n5614, A3 => n1393, ZN => 
                           n16563);
   U1689 : AOI22_X2 port map( A1 => n23495, A2 => n23323, B1 => n23321, B2 => 
                           n23322, ZN => n24672);
   U1691 : NOR3_X1 port map( A1 => n25612, A2 => n25611, A3 => n25610, ZN => 
                           n27407);
   U1695 : NOR2_X2 port map( A1 => n19759, A2 => n19758, ZN => n22143);
   U1700 : NOR2_X1 port map( A1 => n470, A2 => n23946, ZN => n1483);
   U1701 : AND2_X1 port map( A1 => n20609, A2 => n29508, ZN => n899);
   U1703 : OAI211_X2 port map( C1 => n4374, C2 => n4373, A => n4372, B => n4371
                           , ZN => n19669);
   U1705 : OAI211_X2 port map( C1 => n14100, C2 => n14099, A => n3750, B => 
                           n3749, ZN => n15217);
   U1709 : OR2_X1 port map( A1 => n4088, A2 => n13060, ZN => n14350);
   U1711 : NOR2_X2 port map( A1 => n17755, A2 => n5688, ZN => n19045);
   U1725 : XNOR2_X2 port map( A => Key(35), B => Plaintext(35), ZN => n8161);
   U1727 : XNOR2_X2 port map( A => n7115, B => Key(6), ZN => n7116);
   U1731 : NOR2_X2 port map( A1 => n17946, A2 => n17945, ZN => n19267);
   U1733 : NOR2_X2 port map( A1 => n17126, A2 => n17125, ZN => n18136);
   U1739 : BUF_X1 port map( A => n7369, Z => n370);
   U1740 : XNOR2_X1 port map( A => Key(89), B => Plaintext(89), ZN => n7369);
   U1751 : NOR2_X2 port map( A1 => n4648, A2 => n4602, ZN => n24668);
   U1758 : XNOR2_X2 port map( A => n26009, B => n26010, ZN => n27155);
   U1759 : OAI22_X1 port map( A1 => n27795, A2 => n27821, B1 => n29469, B2 => 
                           n27819, ZN => n27823);
   U1761 : INV_X1 port map( A => n28025, ZN => n376);
   U1766 : INV_X1 port map( A => n26459, ZN => n377);
   U1768 : INV_X1 port map( A => n24215, ZN => n378);
   U1769 : CLKBUF_X1 port map( A => n22935, Z => n23449);
   U1770 : INV_X1 port map( A => n23266, ZN => n379);
   U1771 : INV_X1 port map( A => n23587, ZN => n380);
   U1774 : OAI21_X1 port map( B1 => n3953, B2 => n3952, A => n3951, ZN => 
                           n21530);
   U1775 : INV_X1 port map( A => n21000, ZN => n381);
   U1776 : INV_X1 port map( A => n20477, ZN => n382);
   U1779 : INV_X1 port map( A => n20488, ZN => n384);
   U1780 : INV_X1 port map( A => n20166, ZN => n385);
   U1781 : INV_X1 port map( A => n20601, ZN => n386);
   U1784 : INV_X1 port map( A => n16879, ZN => n17382);
   U1785 : XNOR2_X1 port map( A => n16089, B => n16088, ZN => n17456);
   U1786 : INV_X1 port map( A => n17463, ZN => n387);
   U1788 : NAND4_X1 port map( A1 => n14859, A2 => n14862, A3 => n14860, A4 => 
                           n14861, ZN => n16313);
   U1789 : BUF_X1 port map( A => n15323, Z => n546);
   U1790 : INV_X1 port map( A => n13789, ZN => n388);
   U1792 : XNOR2_X1 port map( A => n11670, B => n5805, ZN => n14479);
   U1793 : INV_X1 port map( A => n14016, ZN => n389);
   U1795 : NAND2_X1 port map( A1 => n12188, A2 => n12187, ZN => n12128);
   U1798 : INV_X1 port map( A => n11004, ZN => n10997);
   U1799 : INV_X1 port map( A => n10963, ZN => n10780);
   U1802 : INV_X1 port map( A => n10948, ZN => n391);
   U1805 : CLKBUF_X1 port map( A => n7101, Z => n8179);
   U1811 : CLKBUF_X1 port map( A => Key(25), Z => n1175);
   U1812 : CLKBUF_X1 port map( A => Key(35), Z => n3116);
   U1813 : CLKBUF_X1 port map( A => Key(46), Z => n2325);
   U1815 : CLKBUF_X1 port map( A => Key(56), Z => n3029);
   U1816 : CLKBUF_X1 port map( A => Key(123), Z => n3380);
   U1818 : CLKBUF_X1 port map( A => Key(147), Z => n21537);
   U1819 : CLKBUF_X1 port map( A => Key(188), Z => n3751);
   U1820 : CLKBUF_X1 port map( A => Key(52), Z => n3635);
   U1821 : CLKBUF_X1 port map( A => Key(38), Z => n2984);
   U1822 : CLKBUF_X1 port map( A => Key(17), Z => n3317);
   U1823 : CLKBUF_X1 port map( A => Key(57), Z => n3686);
   U1824 : CLKBUF_X1 port map( A => Key(132), Z => n2522);
   U1825 : CLKBUF_X1 port map( A => Key(145), Z => n3154);
   U1827 : CLKBUF_X1 port map( A => Key(41), Z => n3528);
   U1828 : CLKBUF_X1 port map( A => Key(54), Z => n1179);
   U1830 : CLKBUF_X1 port map( A => Key(65), Z => n1246);
   U1831 : CLKBUF_X1 port map( A => Key(191), Z => n3607);
   U1834 : CLKBUF_X1 port map( A => Key(2), Z => n3586);
   U1835 : CLKBUF_X1 port map( A => Key(64), Z => n1887);
   U1836 : CLKBUF_X1 port map( A => Key(107), Z => n3662);
   U1837 : AOI21_X1 port map( B1 => n802, B2 => n27366, A => n29387, ZN => n801
                           );
   U1838 : INV_X1 port map( A => n6568, ZN => n393);
   U1841 : INV_X1 port map( A => n27549, ZN => n394);
   U1843 : INV_X1 port map( A => n27308, ZN => n395);
   U1845 : OR2_X1 port map( A1 => n1427, A2 => n1622, ZN => n5582);
   U1850 : OAI21_X1 port map( B1 => n26482, B2 => n1622, A => n29501, ZN => 
                           n1470);
   U1851 : INV_X1 port map( A => n29054, ZN => n1279);
   U1852 : OR2_X1 port map( A1 => n4678, A2 => n26426, ZN => n2033);
   U1853 : NOR3_X1 port map( A1 => n26927, A2 => n26926, A3 => n26581, ZN => 
                           n24823);
   U1854 : AND2_X1 port map( A1 => n26995, A2 => n29481, ZN => n26735);
   U1855 : OR3_X1 port map( A1 => n28532, A2 => n26632, A3 => n29481, ZN => 
                           n25971);
   U1856 : INV_X1 port map( A => n28783, ZN => n398);
   U1857 : CLKBUF_X1 port map( A => n25666, Z => n26475);
   U1858 : CLKBUF_X1 port map( A => n25119, Z => n26357);
   U1860 : INV_X1 port map( A => n27052, ZN => n399);
   U1861 : INV_X1 port map( A => n27700, ZN => n400);
   U1862 : INV_X1 port map( A => n26835, ZN => n402);
   U1863 : XNOR2_X1 port map( A => n25261, B => n25366, ZN => n1254);
   U1865 : OAI21_X1 port map( B1 => n24506, B2 => n24263, A => n24262, ZN => 
                           n26090);
   U1867 : OAI22_X1 port map( A1 => n24506, A2 => n28523, B1 => n24505, B2 => 
                           n24806, ZN => n25844);
   U1868 : OR2_X1 port map( A1 => n24258, A2 => n23467, ZN => n1250);
   U1870 : NAND2_X1 port map( A1 => n28415, A2 => n25008, ZN => n1522);
   U1872 : OR2_X1 port map( A1 => n24484, A2 => n24046, ZN => n966);
   U1873 : AND3_X1 port map( A1 => n3723, A2 => n4254, A3 => n6822, ZN => n1955
                           );
   U1874 : CLKBUF_X1 port map( A => n23962, Z => n24468);
   U1875 : OR2_X1 port map( A1 => n23045, A2 => n477, ZN => n1805);
   U1876 : INV_X1 port map( A => n24435, ZN => n403);
   U1877 : OAI211_X1 port map( C1 => n23061, C2 => n23344, A => n4137, B => 
                           n4138, ZN => n23867);
   U1878 : INV_X1 port map( A => n24672, ZN => n404);
   U1881 : OR2_X1 port map( A1 => n481, A2 => n22531, ZN => n1531);
   U1882 : MUX2_X1 port map( A => n480, B => n23062, S => n23417, Z => n23063);
   U1884 : INV_X1 port map( A => n960, ZN => n23622);
   U1885 : INV_X1 port map( A => n4231, ZN => n405);
   U1886 : INV_X1 port map( A => n23612, ZN => n406);
   U1887 : CLKBUF_X1 port map( A => n23825, Z => n23829);
   U1891 : INV_X1 port map( A => n23820, ZN => n407);
   U1896 : INV_X1 port map( A => n23432, ZN => n408);
   U1897 : INV_X1 port map( A => n23250, ZN => n409);
   U1898 : XNOR2_X1 port map( A => n22684, B => n1818, ZN => n23773);
   U1899 : XNOR2_X1 port map( A => n22459, B => n621, ZN => n22382);
   U1900 : AND2_X1 port map( A1 => n5014, A2 => n5013, ZN => n22320);
   U1902 : AOI22_X1 port map( A1 => n21556, A2 => n21555, B1 => n21554, B2 => 
                           n21553, ZN => n22829);
   U1905 : OR2_X1 port map( A1 => n20886, A2 => n21322, ZN => n21590);
   U1909 : INV_X1 port map( A => n1925, ZN => n1924);
   U1911 : INV_X1 port map( A => n21679, ZN => n412);
   U1912 : OAI22_X1 port map( A1 => n821, A2 => n20474, B1 => n2062, B2 => n382
                           , ZN => n21328);
   U1914 : NAND2_X1 port map( A1 => n20134, A2 => n507, ZN => n6770);
   U1915 : AOI21_X1 port map( B1 => n19920, B2 => n20619, A => n500, ZN => 
                           n1565);
   U1917 : NAND2_X1 port map( A1 => n20586, A2 => n20587, ZN => n1429);
   U1918 : INV_X1 port map( A => n19949, ZN => n20587);
   U1919 : OAI21_X1 port map( B1 => n502, B2 => n20109, A => n703, ZN => n20111
                           );
   U1920 : INV_X1 port map( A => n20049, ZN => n413);
   U1921 : INV_X1 port map( A => n20282, ZN => n19808);
   U1923 : OR2_X1 port map( A1 => n505, A2 => n20549, ZN => n5982);
   U1924 : XNOR2_X1 port map( A => n19037, B => n19038, ZN => n20477);
   U1925 : XNOR2_X1 port map( A => n18953, B => n18952, ZN => n20166);
   U1927 : INV_X1 port map( A => n20088, ZN => n414);
   U1929 : XNOR2_X1 port map( A => n16982, B => n16983, ZN => n20549);
   U1930 : INV_X1 port map( A => n19947, ZN => n416);
   U1931 : XNOR2_X1 port map( A => n19504, B => n19503, ZN => n6843);
   U1932 : XNOR2_X1 port map( A => n19191, B => n19452, ZN => n19540);
   U1936 : OR2_X1 port map( A1 => n18466, A2 => n1384, ZN => n1383);
   U1937 : OR2_X1 port map( A1 => n17875, A2 => n525, ZN => n1034);
   U1938 : OR2_X1 port map( A1 => n18449, A2 => n18198, ZN => n18452);
   U1940 : AND2_X1 port map( A1 => n510, A2 => n18507, ZN => n1125);
   U1941 : AND2_X1 port map( A1 => n17618, A2 => n17617, ZN => n17825);
   U1942 : AND2_X1 port map( A1 => n29044, A2 => n527, ZN => n18189);
   U1944 : INV_X1 port map( A => n18411, ZN => n417);
   U1945 : OR2_X1 port map( A1 => n18242, A2 => n522, ZN => n2786);
   U1946 : INV_X1 port map( A => n18507, ZN => n418);
   U1948 : INV_X1 port map( A => n18148, ZN => n420);
   U1949 : OAI21_X1 port map( B1 => n926, B2 => n533, A => n17394, ZN => n1367)
                           ;
   U1950 : AOI21_X1 port map( B1 => n17281, B2 => n528, A => n784, ZN => n783);
   U1952 : NAND2_X1 port map( A1 => n16067, A2 => n1464, ZN => n17941);
   U1953 : OAI211_X1 port map( C1 => n29373, C2 => n17492, A => n4314, B => 
                           n1153, ZN => n4313);
   U1954 : INV_X1 port map( A => n6371, ZN => n1090);
   U1955 : INV_X1 port map( A => n16812, ZN => n421);
   U1958 : INV_X1 port map( A => n17259, ZN => n422);
   U1959 : INV_X1 port map( A => n17571, ZN => n423);
   U1961 : XNOR2_X1 port map( A => n16624, B => n16623, ZN => n16803);
   U1964 : OAI21_X1 port map( B1 => n14788, B2 => n552, A => n14787, ZN => 
                           n16077);
   U1966 : AND3_X1 port map( A1 => n1571, A2 => n552, A3 => n1570, ZN => n13820
                           );
   U1968 : NAND3_X1 port map( A1 => n5197, A2 => n15153, A3 => n5196, ZN => 
                           n16434);
   U1969 : OAI211_X1 port map( C1 => n15518, C2 => n15519, A => n15517, B => 
                           n15516, ZN => n15928);
   U1971 : INV_X1 port map( A => n15323, ZN => n1926);
   U1973 : INV_X1 port map( A => n15343, ZN => n425);
   U1975 : NAND2_X1 port map( A1 => n13810, A2 => n13809, ZN => n15182);
   U1977 : INV_X1 port map( A => n15370, ZN => n426);
   U1978 : OAI21_X1 port map( B1 => n14150, B2 => n557, A => n713, ZN => n14151
                           );
   U1979 : OAI211_X1 port map( C1 => n13934, C2 => n14158, A => n646, B => n558
                           , ZN => n645);
   U1981 : INV_X1 port map( A => n14358, ZN => n13829);
   U1986 : OR2_X1 port map( A1 => n14061, A2 => n13652, ZN => n14322);
   U1988 : INV_X1 port map( A => n14293, ZN => n428);
   U1992 : INV_X1 port map( A => n13069, ZN => n429);
   U1994 : OR2_X1 port map( A1 => n11930, A2 => n568, ZN => n1489);
   U1995 : INV_X1 port map( A => n11951, ZN => n11862);
   U1997 : NAND2_X1 port map( A1 => n29137, A2 => n11778, ZN => n11552);
   U1998 : NAND3_X1 port map( A1 => n11051, A2 => n11050, A3 => n11049, ZN => 
                           n12266);
   U2000 : INV_X1 port map( A => n12150, ZN => n430);
   U2001 : INV_X1 port map( A => n10939, ZN => n11945);
   U2002 : NAND2_X1 port map( A1 => n9292, A2 => n9291, ZN => n13086);
   U2003 : NOR2_X1 port map( A1 => n1375, A2 => n9654, ZN => n9692);
   U2004 : AOI21_X1 port map( B1 => n10923, B2 => n10922, A => n10921, ZN => 
                           n10939);
   U2009 : OAI21_X1 port map( B1 => n1359, B2 => n391, A => n6366, ZN => n11984
                           );
   U2010 : NOR2_X1 port map( A1 => n391, A2 => n10972, ZN => n10969);
   U2011 : OR2_X1 port map( A1 => n595, A2 => n11210, ZN => n11082);
   U2012 : AND2_X1 port map( A1 => n11210, A2 => n595, ZN => n6604);
   U2016 : INV_X1 port map( A => n11207, ZN => n432);
   U2017 : XNOR2_X1 port map( A => n9571, B => n9926, ZN => n1338);
   U2019 : INV_X1 port map( A => n11337, ZN => n434);
   U2020 : XNOR2_X1 port map( A => n10349, B => n1855, ZN => n1854);
   U2022 : INV_X1 port map( A => n11218, ZN => n435);
   U2023 : OAI21_X1 port map( B1 => n606, B2 => n7328, A => n7327, ZN => n10007
                           );
   U2025 : OAI211_X1 port map( C1 => n8379, C2 => n882, A => n881, B => n880, 
                           ZN => n10207);
   U2026 : OR2_X1 port map( A1 => n937, A2 => n7714, ZN => n2915);
   U2027 : INV_X1 port map( A => n8617, ZN => n882);
   U2028 : OR2_X1 port map( A1 => n8617, A2 => n28212, ZN => n880);
   U2033 : INV_X1 port map( A => n8983, ZN => n436);
   U2034 : OAI211_X1 port map( C1 => n7659, C2 => n29317, A => n7402, B => 
                           n7401, ZN => n9134);
   U2037 : OR2_X1 port map( A1 => n7690, A2 => n7817, ZN => n7501);
   U2039 : NOR2_X1 port map( A1 => n7089, A2 => n29112, ZN => n3188);
   U2040 : INV_X1 port map( A => n7997, ZN => n437);
   U2041 : INV_X1 port map( A => n7775, ZN => n438);
   U2042 : XNOR2_X1 port map( A => n7136, B => Key(51), ZN => n7742);
   U2044 : CLKBUF_X1 port map( A => Key(174), Z => n3462);
   U2046 : CLKBUF_X1 port map( A => Key(93), Z => n1172);
   U2047 : CLKBUF_X1 port map( A => Key(49), Z => n1928);
   U2048 : CLKBUF_X1 port map( A => Key(159), Z => n1927);
   U2049 : CLKBUF_X1 port map( A => Key(20), Z => n3770);
   U2050 : CLKBUF_X1 port map( A => Key(10), Z => n2402);
   U2051 : CLKBUF_X1 port map( A => Key(86), Z => n2511);
   U2054 : CLKBUF_X1 port map( A => Key(149), Z => n3180);
   U2055 : CLKBUF_X1 port map( A => Key(142), Z => n3386);
   U2056 : CLKBUF_X1 port map( A => Key(110), Z => n1193);
   U2057 : CLKBUF_X1 port map( A => Key(50), Z => n3697);
   U2058 : CLKBUF_X1 port map( A => Key(27), Z => n3493);
   U2059 : CLKBUF_X1 port map( A => Key(23), Z => n3622);
   U2060 : CLKBUF_X1 port map( A => Key(72), Z => n3212);
   U2061 : CLKBUF_X1 port map( A => Key(103), Z => n2505);
   U2062 : CLKBUF_X1 port map( A => Key(96), Z => n3374);
   U2064 : CLKBUF_X1 port map( A => Key(13), Z => n5059);
   U2065 : CLKBUF_X1 port map( A => Key(94), Z => n1119);
   U2066 : CLKBUF_X1 port map( A => Key(81), Z => n2476);
   U2067 : CLKBUF_X1 port map( A => Key(179), Z => n1247);
   U2068 : CLKBUF_X1 port map( A => Key(104), Z => n3625);
   U2069 : CLKBUF_X1 port map( A => Key(146), Z => n2577);
   U2070 : CLKBUF_X1 port map( A => Key(16), Z => n730);
   U2071 : CLKBUF_X1 port map( A => Key(3), Z => n1187);
   U2072 : CLKBUF_X1 port map( A => Key(37), Z => n1248);
   U2073 : CLKBUF_X1 port map( A => Key(67), Z => n2441);
   U2074 : CLKBUF_X1 port map( A => Key(88), Z => n3114);
   U2075 : CLKBUF_X1 port map( A => Key(74), Z => n22489);
   U2076 : CLKBUF_X1 port map( A => Key(128), Z => n3211);
   U2077 : CLKBUF_X1 port map( A => Key(8), Z => n2973);
   U2078 : CLKBUF_X1 port map( A => Key(97), Z => n2509);
   U2079 : CLKBUF_X1 port map( A => Key(160), Z => n1046);
   U2080 : CLKBUF_X1 port map( A => Key(121), Z => n1184);
   U2082 : CLKBUF_X1 port map( A => Key(181), Z => n2385);
   U2083 : CLKBUF_X1 port map( A => Key(60), Z => n2541);
   U2084 : CLKBUF_X1 port map( A => Key(85), Z => n3067);
   U2085 : CLKBUF_X1 port map( A => Key(18), Z => n2381);
   U2086 : CLKBUF_X1 port map( A => Key(11), Z => n21865);
   U2087 : INV_X1 port map( A => n7369, ZN => n439);
   U2088 : CLKBUF_X1 port map( A => Key(90), Z => n3035);
   U2089 : CLKBUF_X1 port map( A => Key(135), Z => n3457);
   U2090 : CLKBUF_X1 port map( A => Key(173), Z => n24897);
   U2092 : CLKBUF_X1 port map( A => Key(106), Z => n3244);
   U2093 : CLKBUF_X1 port map( A => Key(51), Z => n22072);
   U2094 : CLKBUF_X1 port map( A => Key(140), Z => n3109);
   U2095 : CLKBUF_X1 port map( A => Key(24), Z => n1196);
   U2098 : CLKBUF_X1 port map( A => Key(9), Z => n3606);
   U2100 : CLKBUF_X1 port map( A => Key(168), Z => n3508);
   U2101 : CLKBUF_X1 port map( A => Key(78), Z => n857);
   U2103 : CLKBUF_X1 port map( A => Key(118), Z => n3232);
   U2105 : CLKBUF_X1 port map( A => Key(114), Z => n3336);
   U2106 : CLKBUF_X1 port map( A => Key(34), Z => n2602);
   U2107 : CLKBUF_X1 port map( A => Key(69), Z => n3321);
   U2109 : CLKBUF_X1 port map( A => Key(22), Z => n2446);
   U2110 : INV_X1 port map( A => n3029, ZN => n440);
   U2111 : CLKBUF_X1 port map( A => Key(21), Z => n1133);
   U2112 : CLKBUF_X1 port map( A => Key(156), Z => n2353);
   U2114 : CLKBUF_X1 port map( A => Key(58), Z => n2544);
   U2115 : CLKBUF_X1 port map( A => Key(42), Z => n2306);
   U2116 : CLKBUF_X1 port map( A => Key(43), Z => n3378);
   U2117 : CLKBUF_X1 port map( A => Key(163), Z => n3191);
   U2118 : CLKBUF_X1 port map( A => Key(115), Z => n2912);
   U2119 : CLKBUF_X1 port map( A => Key(75), Z => n3372);
   U2120 : CLKBUF_X1 port map( A => Key(61), Z => n1062);
   U2121 : CLKBUF_X1 port map( A => Key(155), Z => n27956);
   U2122 : CLKBUF_X1 port map( A => Key(178), Z => n3463);
   U2123 : CLKBUF_X1 port map( A => Key(87), Z => n3482);
   U2124 : CLKBUF_X1 port map( A => Key(184), Z => n3323);
   U2126 : CLKBUF_X1 port map( A => Key(136), Z => n2996);
   U2128 : CLKBUF_X1 port map( A => Key(177), Z => n2889);
   U2129 : CLKBUF_X1 port map( A => Key(80), Z => n3660);
   U2130 : CLKBUF_X1 port map( A => Key(190), Z => n1923);
   U2131 : CLKBUF_X1 port map( A => Key(82), Z => n3516);
   U2132 : CLKBUF_X1 port map( A => Key(157), Z => n900);
   U2133 : CLKBUF_X1 port map( A => Key(164), Z => n3728);
   U2134 : CLKBUF_X1 port map( A => Key(176), Z => n27231);
   U2135 : CLKBUF_X1 port map( A => Key(170), Z => n1123);
   U2136 : CLKBUF_X1 port map( A => Key(108), Z => n26531);
   U2137 : CLKBUF_X1 port map( A => Key(12), Z => n2411);
   U2139 : CLKBUF_X1 port map( A => Key(55), Z => n2982);
   U2141 : CLKBUF_X1 port map( A => Key(113), Z => n3451);
   U2142 : CLKBUF_X1 port map( A => Key(109), Z => n2404);
   U2145 : CLKBUF_X1 port map( A => Key(169), Z => n3369);
   U2146 : CLKBUF_X1 port map( A => Key(63), Z => n3334);
   U2147 : CLKBUF_X1 port map( A => Key(40), Z => n891);
   U2149 : CLKBUF_X1 port map( A => Key(120), Z => n2274);
   U2150 : CLKBUF_X1 port map( A => Key(14), Z => n2894);
   U2151 : CLKBUF_X1 port map( A => Key(33), Z => n3633);
   U2153 : CLKBUF_X1 port map( A => Key(127), Z => n2981);
   U2154 : CLKBUF_X1 port map( A => Key(141), Z => n3752);
   U2155 : CLKBUF_X1 port map( A => Key(28), Z => n2995);
   U2156 : CLKBUF_X1 port map( A => Key(76), Z => n2598);
   U2158 : CLKBUF_X1 port map( A => Key(148), Z => n1161);
   U2159 : CLKBUF_X1 port map( A => Key(137), Z => n3742);
   U2161 : OR2_X1 port map( A1 => n26145, A2 => n27727, ZN => n26147);
   U2162 : OR2_X1 port map( A1 => n28005, A2 => n28006, ZN => n1546);
   U2164 : AOI22_X1 port map( A1 => n28027, A2 => n376, B1 => n25601, B2 => 
                           n28035, ZN => n26664);
   U2165 : NOR2_X1 port map( A1 => n27586, A2 => n27585, ZN => n931);
   U2166 : INV_X1 port map( A => n1548, ZN => n28000);
   U2167 : INV_X1 port map( A => n27862, ZN => n27873);
   U2168 : AOI211_X1 port map( C1 => n27431, C2 => n27430, A => n1821, B => 
                           n1820, ZN => n1819);
   U2169 : OAI21_X1 port map( B1 => n27387, B2 => n27408, A => n26960, ZN => 
                           n27403);
   U2170 : AND2_X1 port map( A1 => n27387, A2 => n25629, ZN => n27409);
   U2171 : INV_X1 port map( A => n25629, ZN => n27400);
   U2172 : OR2_X1 port map( A1 => n397, A2 => n27759, ZN => n2794);
   U2173 : INV_X1 port map( A => n6095, ZN => n27526);
   U2175 : NOR3_X1 port map( A1 => n27429, A2 => n27426, A3 => n27425, ZN => 
                           n1821);
   U2176 : INV_X1 port map( A => n27573, ZN => n27553);
   U2177 : NOR2_X1 port map( A1 => n29056, A2 => n28111, ZN => n1691);
   U2178 : NOR2_X1 port map( A1 => n28089, A2 => n28111, ZN => n28109);
   U2179 : NOR2_X1 port map( A1 => n27830, A2 => n27829, ZN => n27100);
   U2180 : OR2_X1 port map( A1 => n27938, A2 => n27244, ZN => n1011);
   U2181 : OR2_X1 port map( A1 => n28016, A2 => n28017, ZN => n1548);
   U2182 : NOR2_X1 port map( A1 => n27855, A2 => n26641, ZN => n26696);
   U2184 : INV_X1 port map( A => n27362, ZN => n27370);
   U2185 : INV_X1 port map( A => n28179, ZN => n930);
   U2187 : INV_X1 port map( A => n27588, ZN => n933);
   U2188 : NOR2_X1 port map( A1 => n27582, A2 => n27590, ZN => n27589);
   U2189 : INV_X1 port map( A => n27439, ZN => n26829);
   U2190 : NOR2_X1 port map( A1 => n26069, A2 => n26068, ZN => n27728);
   U2191 : AND3_X1 port map( A1 => n27429, A2 => n27428, A3 => n27427, ZN => 
                           n1820);
   U2192 : AND3_X1 port map( A1 => n5735, A2 => n24825, A3 => n24824, ZN => 
                           n6568);
   U2194 : NOR2_X1 port map( A1 => n25201, A2 => n25200, ZN => n27549);
   U2195 : NOR2_X1 port map( A1 => n27547, A2 => n26652, ZN => n27200);
   U2196 : INV_X1 port map( A => n27630, ZN => n442);
   U2197 : OAI211_X1 port map( C1 => n26361, C2 => n1076, A => n2033, B => 
                           n1075, ZN => n27614);
   U2198 : INV_X1 port map( A => n28019, ZN => n443);
   U2199 : INV_X1 port map( A => n27301, ZN => n444);
   U2200 : INV_X1 port map( A => n28016, ZN => n445);
   U2203 : AND2_X1 port map( A1 => n3703, A2 => n3702, ZN => n27286);
   U2204 : NOR2_X1 port map( A1 => n1968, A2 => n26262, ZN => n27597);
   U2205 : INV_X1 port map( A => n27213, ZN => n446);
   U2208 : INV_X1 port map( A => n27863, ZN => n27871);
   U2209 : NAND3_X1 port map( A1 => n798, A2 => n29055, A3 => n4173, ZN => 
                           n27362);
   U2210 : INV_X1 port map( A => n27859, ZN => n447);
   U2213 : NOR2_X1 port map( A1 => n26743, A2 => n26744, ZN => n28090);
   U2215 : INV_X1 port map( A => n27465, ZN => n449);
   U2218 : MUX2_X1 port map( A => n26509, B => n26508, S => n27084, Z => n26639
                           );
   U2220 : OAI21_X1 port map( B1 => n27122, B2 => n26516, A => n26515, ZN => 
                           n27854);
   U2221 : NOR2_X1 port map( A1 => n26635, A2 => n26634, ZN => n27972);
   U2222 : OAI21_X1 port map( B1 => n26301, B2 => n27904, A => n25953, ZN => 
                           n27863);
   U2223 : AOI21_X1 port map( B1 => n27151, B2 => n401, A => n27152, ZN => 
                           n3590);
   U2224 : NOR2_X1 port map( A1 => n26356, A2 => n28650, ZN => n27186);
   U2225 : AND2_X1 port map( A1 => n28575, A2 => n26761, ZN => n1169);
   U2226 : NAND2_X1 port map( A1 => n27012, A2 => n399, ZN => n1535);
   U2228 : INV_X1 port map( A => n1622, ZN => n1472);
   U2229 : AND2_X1 port map( A1 => n26727, A2 => n26480, ZN => n1533);
   U2231 : NOR2_X1 port map( A1 => n26241, A2 => n26753, ZN => n25650);
   U2232 : BUF_X1 port map( A => n26729, Z => n26482);
   U2233 : NOR2_X1 port map( A1 => n26200, A2 => n26235, ZN => n26741);
   U2234 : OAI21_X1 port map( B1 => n26461, B2 => n26457, A => n28578, ZN => 
                           n949);
   U2235 : AOI21_X1 port map( B1 => n28504, B2 => n27161, A => n27701, ZN => 
                           n5994);
   U2236 : OR2_X1 port map( A1 => n27124, A2 => n28513, ZN => n5486);
   U2237 : OR3_X1 port map( A1 => n26426, A2 => n26382, A3 => n26381, ZN => 
                           n26383);
   U2238 : INV_X1 port map( A => n26736, ZN => n826);
   U2240 : INV_X1 port map( A => n25406, ZN => n26469);
   U2241 : INV_X1 port map( A => n27067, ZN => n922);
   U2244 : XNOR2_X1 port map( A => n6436, B => n25064, ZN => n4820);
   U2245 : OR2_X1 port map( A1 => n26997, A2 => n26733, ZN => n26736);
   U2247 : XNOR2_X1 port map( A => n23941, B => n23940, ZN => n26448);
   U2250 : BUF_X1 port map( A => n25676, Z => n27041);
   U2253 : XNOR2_X1 port map( A => n24988, B => n24989, ZN => n27169);
   U2254 : INV_X1 port map( A => n26727, ZN => n1622);
   U2256 : INV_X1 port map( A => n25365, ZN => n26928);
   U2261 : XNOR2_X1 port map( A => n25742, B => n25741, ZN => n5263);
   U2264 : XNOR2_X1 port map( A => n25804, B => n25805, ZN => n26841);
   U2267 : INV_X1 port map( A => n26919, ZN => n454);
   U2269 : XNOR2_X1 port map( A => n24695, B => n24696, ZN => n25365);
   U2270 : XNOR2_X1 port map( A => n4084, B => n4082, ZN => n26740);
   U2271 : INV_X1 port map( A => n27704, ZN => n455);
   U2272 : INV_X1 port map( A => n26941, ZN => n456);
   U2273 : XNOR2_X1 port map( A => n25587, B => n25586, ZN => n26995);
   U2274 : INV_X1 port map( A => n26917, ZN => n457);
   U2276 : XNOR2_X1 port map( A => n23893, B => n23892, ZN => n26179);
   U2278 : NOR2_X1 port map( A1 => n24981, A2 => n24980, ZN => n25411);
   U2279 : XNOR2_X1 port map( A => n1303, B => n25891, ZN => n1302);
   U2280 : XNOR2_X1 port map( A => n25262, B => n26070, ZN => n25081);
   U2282 : INV_X1 port map( A => n24870, ZN => n25944);
   U2283 : XNOR2_X1 port map( A => n25703, B => n5146, ZN => n26101);
   U2284 : AND3_X1 port map( A1 => n4691, A2 => n4694, A3 => n4690, ZN => 
                           n25369);
   U2285 : NOR2_X1 port map( A1 => n24615, A2 => n5136, ZN => n25876);
   U2287 : NOR2_X1 port map( A1 => n3567, A2 => n24122, ZN => n25268);
   U2288 : NOR2_X1 port map( A1 => n22871, A2 => n22872, ZN => n25293);
   U2289 : OR2_X1 port map( A1 => n820, A2 => n3654, ZN => n1458);
   U2295 : AND4_X1 port map( A1 => n276, A2 => n1517, A3 => n25007, A4 => n1515
                           , ZN => n1514);
   U2296 : OAI211_X1 port map( C1 => n24442, C2 => n24441, A => n24440, B => 
                           n24439, ZN => n25564);
   U2297 : OR2_X1 port map( A1 => n1283, A2 => n24589, ZN => n1282);
   U2300 : OR2_X1 port map( A1 => n24649, A2 => n672, ZN => n24660);
   U2302 : INV_X1 port map( A => n966, ZN => n24482);
   U2303 : OAI22_X1 port map( A1 => n24083, A2 => n24408, B1 => n6266, B2 => 
                           n24405, ZN => n24407);
   U2304 : AND2_X1 port map( A1 => n23971, A2 => n24479, ZN => n1655);
   U2305 : NOR2_X1 port map( A1 => n24806, A2 => n803, ZN => n24263);
   U2308 : INV_X1 port map( A => n24454, ZN => n458);
   U2309 : INV_X1 port map( A => n29555, ZN => n1274);
   U2311 : NOR2_X1 port map( A1 => n24467, A2 => n24582, ZN => n1203);
   U2312 : INV_X1 port map( A => n24278, ZN => n24590);
   U2313 : INV_X1 port map( A => n1808, ZN => n24338);
   U2314 : NOR2_X1 port map( A1 => n25793, A2 => n25794, ZN => n25800);
   U2315 : AND2_X1 port map( A1 => n24745, A2 => n24751, ZN => n24616);
   U2316 : INV_X1 port map( A => n24612, ZN => n459);
   U2317 : INV_X1 port map( A => n23389, ZN => n811);
   U2318 : OR2_X1 port map( A1 => n831, A2 => n24592, ZN => n2586);
   U2319 : AND2_X1 port map( A1 => n24739, A2 => n24735, ZN => n24604);
   U2320 : NOR2_X1 port map( A1 => n22867, A2 => n22866, ZN => n24173);
   U2321 : INV_X1 port map( A => n24706, ZN => n24417);
   U2322 : NAND2_X1 port map( A1 => n24339, A2 => n24340, ZN => n3731);
   U2323 : OR2_X1 port map( A1 => n24388, A2 => n24077, ZN => n24135);
   U2324 : AND2_X1 port map( A1 => n4849, A2 => n2557, ZN => n1856);
   U2325 : INV_X1 port map( A => n831, ZN => n4693);
   U2326 : AND2_X1 port map( A1 => n25008, A2 => n24138, ZN => n1516);
   U2327 : INV_X1 port map( A => n24804, ZN => n24162);
   U2328 : OR2_X1 port map( A1 => n24241, A2 => n24559, ZN => n1726);
   U2330 : OR2_X1 port map( A1 => n24133, A2 => n24081, ZN => n1617);
   U2332 : INV_X1 port map( A => n3061, ZN => n673);
   U2334 : INV_X1 port map( A => n29695, ZN => n460);
   U2335 : OR2_X1 port map( A1 => n24629, A2 => n4364, ZN => n24531);
   U2336 : OR2_X1 port map( A1 => n23897, A2 => n25008, ZN => n1515);
   U2337 : INV_X1 port map( A => n24747, ZN => n1631);
   U2338 : INV_X1 port map( A => n24457, ZN => n1426);
   U2339 : INV_X1 port map( A => n29309, ZN => n24775);
   U2340 : INV_X1 port map( A => n24369, ZN => n461);
   U2341 : INV_X1 port map( A => n24745, ZN => n462);
   U2342 : AND2_X1 port map( A1 => n24891, A2 => n24631, ZN => n23982);
   U2347 : OR2_X1 port map( A1 => n25008, A2 => n24138, ZN => n1448);
   U2348 : INV_X1 port map( A => n23945, ZN => n463);
   U2349 : INV_X1 port map( A => n1955, ZN => n464);
   U2350 : AND2_X1 port map( A1 => n5696, A2 => n5698, ZN => n24555);
   U2354 : INV_X1 port map( A => n24635, ZN => n465);
   U2355 : OAI211_X1 port map( C1 => n23741, C2 => n23383, A => n1638, B => 
                           n1637, ZN => n24133);
   U2356 : OAI21_X1 port map( B1 => n23444, B2 => n4794, A => n2169, ZN => 
                           n1498);
   U2358 : NOR2_X1 port map( A1 => n21929, A2 => n6310, ZN => n6309);
   U2359 : OAI21_X1 port map( B1 => n23424, B2 => n23426, A => n23115, ZN => 
                           n24483);
   U2360 : INV_X1 port map( A => n24310, ZN => n466);
   U2362 : OR2_X1 port map( A1 => n24367, A2 => n24138, ZN => n1551);
   U2364 : INV_X1 port map( A => n24972, ZN => n468);
   U2366 : NAND2_X1 port map( A1 => n5080, A2 => n24093, ZN => n24489);
   U2367 : AND2_X1 port map( A1 => n23805, A2 => n22742, ZN => n1240);
   U2368 : AND3_X1 port map( A1 => n6609, A2 => n6608, A3 => n6607, ZN => 
                           n24337);
   U2369 : INV_X1 port map( A => n24211, ZN => n469);
   U2370 : AOI21_X1 port map( B1 => n1531, B2 => n22863, A => n23835, ZN => 
                           n22867);
   U2371 : AOI22_X1 port map( A1 => n23690, A2 => n23802, B1 => n23689, B2 => 
                           n23688, ZN => n24205);
   U2372 : INV_X1 port map( A => n24779, ZN => n470);
   U2376 : OR2_X1 port map( A1 => n23440, A2 => n23441, ZN => n1228);
   U2378 : INV_X1 port map( A => n24509, ZN => n471);
   U2380 : AND2_X1 port map( A1 => n23189, A2 => n1286, ZN => n23757);
   U2381 : OR2_X1 port map( A1 => n23253, A2 => n23252, ZN => n867);
   U2382 : OAI22_X1 port map( A1 => n6054, A2 => n2141, B1 => n943, B2 => 
                           n23735, ZN => n22009);
   U2383 : OR2_X1 port map( A1 => n2066, A2 => n23558, ZN => n1556);
   U2384 : OR3_X1 port map( A1 => n23180, A2 => n23645, A3 => n23643, ZN => 
                           n23181);
   U2385 : OAI21_X1 port map( B1 => n808, B2 => n23787, A => n23036, ZN => 
                           n1642);
   U2386 : OR2_X1 port map( A1 => n23395, A2 => n23396, ZN => n907);
   U2387 : AND2_X1 port map( A1 => n754, A2 => n755, ZN => n23402);
   U2388 : OR2_X1 port map( A1 => n23384, A2 => n23385, ZN => n1637);
   U2389 : AND2_X1 port map( A1 => n23442, A2 => n23370, ZN => n23444);
   U2390 : NOR2_X1 port map( A1 => n23626, A2 => n23566, ZN => n23274);
   U2391 : NOR2_X1 port map( A1 => n23074, A2 => n28653, ZN => n23811);
   U2392 : OR2_X1 port map( A1 => n23538, A2 => n1913, ZN => n712);
   U2393 : AND3_X1 port map( A1 => n28594, A2 => n23807, A3 => n29102, ZN => 
                           n23814);
   U2394 : AND2_X1 port map( A1 => n22451, A2 => n22452, ZN => n23704);
   U2395 : NAND2_X1 port map( A1 => n23787, A2 => n23786, ZN => n1641);
   U2396 : AND2_X1 port map( A1 => n23305, A2 => n22686, ZN => n23303);
   U2397 : OR2_X1 port map( A1 => n23808, A2 => n29102, ZN => n1284);
   U2398 : OR2_X1 port map( A1 => n23073, A2 => n23099, ZN => n2400);
   U2399 : INV_X1 port map( A => n23615, ZN => n760);
   U2401 : OR2_X1 port map( A1 => n23829, A2 => n23382, ZN => n23383);
   U2405 : OR2_X1 port map( A1 => n23735, A2 => n23736, ZN => n755);
   U2406 : XNOR2_X1 port map( A => n21782, B => n21781, ZN => n23767);
   U2407 : XNOR2_X1 port map( A => n4228, B => n22924, ZN => n23461);
   U2409 : INV_X1 port map( A => n23784, ZN => n473);
   U2410 : XNOR2_X1 port map( A => n22203, B => n22202, ZN => n23612);
   U2411 : INV_X1 port map( A => n23679, ZN => n474);
   U2412 : INV_X1 port map( A => n23825, ZN => n885);
   U2415 : XNOR2_X1 port map( A => n22276, B => n2393, ZN => n23633);
   U2416 : INV_X1 port map( A => n23787, ZN => n475);
   U2417 : XNOR2_X1 port map( A => n22324, B => n22323, ZN => n23762);
   U2418 : INV_X1 port map( A => n379, ZN => n476);
   U2419 : INV_X1 port map( A => n23557, ZN => n477);
   U2421 : XNOR2_X1 port map( A => n22816, B => n22817, ZN => n23820);
   U2423 : INV_X1 port map( A => n23647, ZN => n641);
   U2425 : CLKBUF_X1 port map( A => n23258, Z => n23398);
   U2426 : INV_X1 port map( A => n22979, ZN => n23405);
   U2429 : INV_X1 port map( A => n22946, ZN => n23385);
   U2430 : INV_X1 port map( A => n23416, ZN => n479);
   U2431 : OR2_X1 port map( A1 => n23733, A2 => n23258, ZN => n754);
   U2432 : INV_X1 port map( A => n23099, ZN => n480);
   U2433 : INV_X1 port map( A => n23077, ZN => n481);
   U2434 : INV_X1 port map( A => n23382, ZN => n482);
   U2436 : INV_X1 port map( A => n23419, ZN => n483);
   U2437 : INV_X1 port map( A => n28164, ZN => n484);
   U2439 : INV_X1 port map( A => n23418, ZN => n485);
   U2440 : INV_X1 port map( A => n23360, ZN => n486);
   U2441 : XNOR2_X1 port map( A => n22425, B => n22424, ZN => n23647);
   U2443 : INV_X1 port map( A => n28460, ZN => n487);
   U2447 : XNOR2_X1 port map( A => n21835, B => n21834, ZN => n23777);
   U2448 : XNOR2_X1 port map( A => n22390, B => n1451, ZN => n23618);
   U2449 : XNOR2_X1 port map( A => n1500, B => n22711, ZN => n1055);
   U2450 : XNOR2_X1 port map( A => n22610, B => n22007, ZN => n4968);
   U2451 : XNOR2_X1 port map( A => n22156, B => n22155, ZN => n23587);
   U2454 : XNOR2_X1 port map( A => n22522, B => n3372, ZN => n1538);
   U2455 : XNOR2_X1 port map( A => n22912, B => n21990, ZN => n22533);
   U2456 : XNOR2_X1 port map( A => n22923, B => n1501, ZN => n1500);
   U2457 : INV_X1 port map( A => n22710, ZN => n1501);
   U2460 : XNOR2_X1 port map( A => n21982, B => n22110, ZN => n22395);
   U2461 : XNOR2_X1 port map( A => n22245, B => n3635, ZN => n6389);
   U2462 : XNOR2_X1 port map( A => n22830, B => n22525, ZN => n21847);
   U2464 : INV_X1 port map( A => n22690, ZN => n22169);
   U2468 : AND2_X1 port map( A1 => n20991, A2 => n20990, ZN => n22006);
   U2470 : INV_X1 port map( A => n22099, ZN => n22098);
   U2471 : AND2_X1 port map( A1 => n20185, A2 => n5018, ZN => n22132);
   U2472 : NAND3_X1 port map( A1 => n270, A2 => n3889, A3 => n3891, ZN => n1271
                           );
   U2476 : OAI211_X1 port map( C1 => n21619, C2 => n21618, A => n21617, B => 
                           n21616, ZN => n22813);
   U2478 : AND3_X1 port map( A1 => n1289, A2 => n269, A3 => n1288, ZN => n3486)
                           ;
   U2479 : OR2_X1 port map( A1 => n19859, A2 => n4467, ZN => n4466);
   U2480 : OAI211_X1 port map( C1 => n21619, C2 => n20906, A => n20524, B => 
                           n20523, ZN => n22609);
   U2482 : AND3_X1 port map( A1 => n650, A2 => n648, A3 => n647, ZN => n3578);
   U2486 : OR2_X1 port map( A1 => n21748, A2 => n20658, ZN => n1327);
   U2487 : AOI22_X1 port map( A1 => n1621, A2 => n21550, B1 => n21553, B2 => 
                           n21547, ZN => n21181);
   U2488 : AND2_X1 port map( A1 => n21178, A2 => n21179, ZN => n879);
   U2489 : OAI21_X1 port map( B1 => n21015, B2 => n21016, A => n22404, ZN => 
                           n1720);
   U2490 : AOI21_X1 port map( B1 => n21236, B2 => n21237, A => n21748, ZN => 
                           n952);
   U2491 : OAI21_X1 port map( B1 => n20844, B2 => n1814, A => n21125, ZN => 
                           n1083);
   U2493 : AND2_X1 port map( A1 => n20848, A2 => n21481, ZN => n854);
   U2494 : OR2_X1 port map( A1 => n28791, A2 => n21334, ZN => n4776);
   U2495 : OR2_X1 port map( A1 => n4960, A2 => n20744, ZN => n3119);
   U2497 : AND2_X1 port map( A1 => n21306, A2 => n21311, ZN => n906);
   U2498 : INV_X1 port map( A => n21171, ZN => n21409);
   U2499 : NOR2_X1 port map( A1 => n20688, A2 => n20689, ZN => n21716);
   U2500 : INV_X1 port map( A => n21090, ZN => n701);
   U2501 : INV_X1 port map( A => n21530, ZN => n1543);
   U2502 : INV_X1 port map( A => n21532, ZN => n1540);
   U2504 : OR2_X1 port map( A1 => n20886, A2 => n21587, ZN => n1288);
   U2505 : INV_X1 port map( A => n20786, ZN => n21930);
   U2507 : NOR2_X1 port map( A1 => n22286, A2 => n22290, ZN => n1693);
   U2508 : INV_X1 port map( A => n21221, ZN => n20703);
   U2509 : OR2_X1 port map( A1 => n21113, A2 => n21464, ZN => n4224);
   U2511 : INV_X1 port map( A => n20988, ZN => n20914);
   U2516 : OR2_X1 port map( A1 => n20854, A2 => n21145, ZN => n2427);
   U2517 : INV_X1 port map( A => n21213, ZN => n489);
   U2518 : INV_X1 port map( A => n21574, ZN => n21485);
   U2519 : INV_X1 port map( A => n20783, ZN => n21550);
   U2520 : AND2_X1 port map( A1 => n21014, A2 => n21429, ZN => n21016);
   U2521 : INV_X1 port map( A => n21736, ZN => n21471);
   U2524 : NOR2_X1 port map( A1 => n20878, A2 => n20877, ZN => n20879);
   U2525 : INV_X1 port map( A => n21119, ZN => n21117);
   U2527 : INV_X1 port map( A => n21408, ZN => n490);
   U2529 : INV_X1 port map( A => n20393, ZN => n21541);
   U2530 : AND2_X1 port map( A1 => n21599, A2 => n21600, ZN => n20905);
   U2531 : AND2_X1 port map( A1 => n6771, A2 => n6770, ZN => n20899);
   U2532 : AND2_X1 port map( A1 => n21679, A2 => n21674, ZN => n21449);
   U2534 : OR2_X1 port map( A1 => n19980, A2 => n6114, ZN => n649);
   U2535 : OR2_X1 port map( A1 => n21118, A2 => n21145, ZN => n21141);
   U2537 : INV_X1 port map( A => n21078, ZN => n491);
   U2545 : OR2_X1 port map( A1 => n6577, A2 => n19994, ZN => n1462);
   U2546 : INV_X1 port map( A => n21143, ZN => n492);
   U2548 : INV_X1 port map( A => n21473, ZN => n493);
   U2549 : OR2_X1 port map( A1 => n20045, A2 => n19985, ZN => n18884);
   U2550 : NOR2_X1 port map( A1 => n20328, A2 => n28491, ZN => n1335);
   U2551 : INV_X1 port map( A => n20744, ZN => n494);
   U2552 : AND2_X1 port map( A1 => n681, A2 => n680, ZN => n20139);
   U2555 : INV_X1 port map( A => n20533, ZN => n495);
   U2556 : OAI211_X1 port map( C1 => n20198, C2 => n20588, A => n1428, B => 
                           n1429, ZN => n21679);
   U2560 : OR2_X1 port map( A1 => n18848, A2 => n836, ZN => n835);
   U2561 : INV_X1 port map( A => n21704, ZN => n496);
   U2562 : INV_X1 port map( A => n21400, ZN => n497);
   U2563 : AOI21_X1 port map( B1 => n19808, B2 => n20284, A => n20283, ZN => 
                           n680);
   U2568 : INV_X1 port map( A => n21362, ZN => n19458);
   U2569 : INV_X1 port map( A => n6840, ZN => n21248);
   U2572 : INV_X1 port map( A => n20248, ZN => n20636);
   U2573 : NOR2_X1 port map( A1 => n20354, A2 => n20478, ZN => n20474);
   U2574 : AND2_X1 port map( A1 => n20162, A2 => n29066, ZN => n19872);
   U2575 : AND2_X1 port map( A1 => n384, A2 => n20486, ZN => n869);
   U2576 : AND2_X1 port map( A1 => n19765, A2 => n20049, ZN => n18848);
   U2577 : INV_X1 port map( A => n21353, ZN => n20517);
   U2579 : OR2_X1 port map( A1 => n4657, A2 => n19973, ZN => n4656);
   U2581 : OR2_X1 port map( A1 => n20607, A2 => n20441, ZN => n20612);
   U2582 : INV_X1 port map( A => n19993, ZN => n20222);
   U2583 : INV_X1 port map( A => n20549, ZN => n1781);
   U2584 : XNOR2_X1 port map( A => n19674, B => n19673, ZN => n20137);
   U2586 : INV_X1 port map( A => n20504, ZN => n1626);
   U2587 : BUF_X1 port map( A => n18699, Z => n20379);
   U2589 : INV_X1 port map( A => n20637, ZN => n498);
   U2591 : OR2_X1 port map( A1 => n20299, A2 => n20130, ZN => n1178);
   U2592 : XNOR2_X1 port map( A => n19545, B => n19544, ZN => n19554);
   U2593 : XNOR2_X1 port map( A => n19319, B => n19318, ZN => n1881);
   U2594 : AND2_X1 port map( A1 => n20209, A2 => n19851, ZN => n20397);
   U2595 : OR2_X1 port map( A1 => n19993, A2 => n20166, ZN => n20221);
   U2596 : INV_X1 port map( A => n20209, ZN => n20394);
   U2597 : XNOR2_X1 port map( A => n19352, B => n19353, ZN => n19920);
   U2598 : OR2_X1 port map( A1 => n20458, A2 => n4569, ZN => n20275);
   U2599 : INV_X1 port map( A => n20182, ZN => n499);
   U2600 : INV_X1 port map( A => n20431, ZN => n500);
   U2601 : XNOR2_X1 port map( A => n18623, B => n19690, ZN => n20567);
   U2602 : XNOR2_X1 port map( A => n18911, B => n18910, ZN => n20144);
   U2604 : XNOR2_X1 port map( A => n1757, B => n19617, ZN => n1755);
   U2607 : INV_X1 port map( A => n21355, ZN => n501);
   U2609 : BUF_X1 port map( A => n19093, Z => n20239);
   U2610 : XNOR2_X1 port map( A => n774, B => n773, ZN => n20618);
   U2611 : INV_X1 port map( A => n28140, ZN => n503);
   U2612 : XNOR2_X1 port map( A => n17655, B => n17656, ZN => n20580);
   U2613 : XNOR2_X1 port map( A => n17606, B => n17605, ZN => n20414);
   U2615 : XNOR2_X1 port map( A => n18678, B => n18679, ZN => n20375);
   U2616 : INV_X1 port map( A => n20178, ZN => n504);
   U2619 : XNOR2_X1 port map( A => n5211, B => n18721, ZN => n20088);
   U2621 : XNOR2_X1 port map( A => n5161, B => n19484, ZN => n19315);
   U2622 : XNOR2_X1 port map( A => n18116, B => n18115, ZN => n19947);
   U2623 : XNOR2_X1 port map( A => n19591, B => n775, ZN => n774);
   U2624 : INV_X1 port map( A => n19855, ZN => n505);
   U2625 : INV_X1 port map( A => n20284, ZN => n506);
   U2626 : XNOR2_X1 port map( A => n19225, B => n3087, ZN => n1757);
   U2627 : XNOR2_X1 port map( A => n1823, B => n1822, ZN => n20130);
   U2628 : INV_X1 port map( A => n19270, ZN => n1054);
   U2631 : XNOR2_X1 port map( A => n18804, B => n18805, ZN => n20098);
   U2632 : XNOR2_X1 port map( A => n18985, B => n18986, ZN => n20173);
   U2633 : INV_X1 port map( A => n6843, ZN => n507);
   U2634 : XNOR2_X1 port map( A => n1504, B => n19349, ZN => n19445);
   U2635 : XNOR2_X1 port map( A => n1825, B => n1824, ZN => n1822);
   U2636 : XNOR2_X1 port map( A => n19330, B => n267, ZN => n773);
   U2637 : XNOR2_X1 port map( A => n18782, B => n19332, ZN => n19175);
   U2638 : NOR2_X1 port map( A1 => n18594, A2 => n2341, ZN => n19300);
   U2640 : INV_X1 port map( A => n1733, ZN => n1783);
   U2642 : XNOR2_X1 port map( A => n19481, B => n19483, ZN => n1825);
   U2644 : XNOR2_X1 port map( A => n1733, B => n19207, ZN => n19528);
   U2645 : XNOR2_X1 port map( A => n19192, B => n1741, ZN => n19356);
   U2646 : INV_X1 port map( A => n19086, ZN => n18906);
   U2647 : XNOR2_X1 port map( A => n19206, B => n18695, ZN => n19330);
   U2648 : INV_X1 port map( A => n19490, ZN => n18085);
   U2649 : NAND2_X1 port map( A1 => n2150, A2 => n2147, ZN => n19475);
   U2650 : INV_X1 port map( A => n19246, ZN => n19616);
   U2651 : INV_X1 port map( A => n19349, ZN => n1505);
   U2653 : INV_X1 port map( A => n19228, ZN => n1503);
   U2655 : XNOR2_X1 port map( A => n19482, B => n22072, ZN => n1824);
   U2661 : OR2_X1 port map( A1 => n1455, A2 => n17602, ZN => n19490);
   U2663 : AND3_X1 port map( A1 => n1506, A2 => n18066, A3 => n18065, ZN => 
                           n19349);
   U2664 : NAND2_X1 port map( A1 => n16981, A2 => n3544, ZN => n19483);
   U2666 : NOR2_X1 port map( A1 => n5178, A2 => n17936, ZN => n19323);
   U2672 : NOR2_X1 port map( A1 => n17591, A2 => n17590, ZN => n18725);
   U2673 : AND3_X1 port map( A1 => n2045, A2 => n5857, A3 => n5985, ZN => 
                           n19122);
   U2676 : AND3_X1 port map( A1 => n2770, A2 => n2771, A3 => n17757, ZN => 
                           n19273);
   U2678 : AND2_X1 port map( A1 => n17638, A2 => n6930, ZN => n19305);
   U2682 : AND2_X1 port map( A1 => n18181, A2 => n18444, ZN => n18448);
   U2683 : INV_X1 port map( A => n18100, ZN => n18199);
   U2686 : MUX2_X1 port map( A => n18219, B => n18218, S => n18217, Z => n18877
                           );
   U2687 : OAI21_X1 port map( B1 => n17652, B2 => n17653, A => n17651, ZN => 
                           n18773);
   U2688 : INV_X1 port map( A => n3439, ZN => n1731);
   U2689 : OR2_X1 port map( A1 => n18098, A2 => n18444, ZN => n1304);
   U2691 : INV_X1 port map( A => n18173, ZN => n1708);
   U2692 : AND2_X1 port map( A1 => n17942, A2 => n17941, ZN => n1433);
   U2694 : AND2_X1 port map( A1 => n18304, A2 => n18306, ZN => n17933);
   U2695 : INV_X1 port map( A => n17793, ZN => n671);
   U2696 : OR2_X1 port map( A1 => n18333, A2 => n817, ZN => n17652);
   U2697 : OR2_X1 port map( A1 => n18195, A2 => n18449, ZN => n18100);
   U2698 : AND2_X1 port map( A1 => n15734, A2 => n18490, ZN => n18016);
   U2699 : AND2_X1 port map( A1 => n17858, A2 => n18285, ZN => n18521);
   U2700 : INV_X1 port map( A => n420, ZN => n1758);
   U2701 : AND2_X1 port map( A1 => n18261, A2 => n18263, ZN => n697);
   U2702 : AND2_X1 port map( A1 => n17842, A2 => n18242, ZN => n2787);
   U2704 : AND2_X1 port map( A1 => n17564, A2 => n17771, ZN => n1378);
   U2705 : INV_X1 port map( A => n18706, ZN => n876);
   U2706 : NOR2_X1 port map( A1 => n18333, A2 => n18334, ZN => n1180);
   U2707 : OR2_X1 port map( A1 => n18402, A2 => n18232, ZN => n1524);
   U2708 : AND2_X1 port map( A1 => n18268, A2 => n18326, ZN => n1717);
   U2709 : INV_X1 port map( A => n18422, ZN => n1530);
   U2711 : OR2_X1 port map( A1 => n17132, A2 => n17131, ZN => n18137);
   U2712 : NAND2_X1 port map( A1 => n6643, A2 => n6642, ZN => n18537);
   U2713 : INV_X1 port map( A => n18342, ZN => n17906);
   U2714 : AND2_X1 port map( A1 => n15892, A2 => n18299, ZN => n18061);
   U2715 : OAI21_X1 port map( B1 => n17717, B2 => n17431, A => n5329, ZN => 
                           n18522);
   U2716 : INV_X1 port map( A => n817, ZN => n4412);
   U2720 : OR2_X1 port map( A1 => n17939, A2 => n17872, ZN => n1436);
   U2722 : INV_X1 port map( A => n18040, ZN => n17824);
   U2723 : AND2_X1 port map( A1 => n18421, A2 => n17802, ZN => n1577);
   U2724 : AND2_X1 port map( A1 => n18040, A2 => n18421, ZN => n1576);
   U2725 : INV_X1 port map( A => n17864, ZN => n509);
   U2726 : NAND4_X1 port map( A1 => n679, A2 => n16893, A3 => n16892, A4 => 
                           n16894, ZN => n18511);
   U2727 : OAI211_X1 port map( C1 => n16825, C2 => n4571, A => n4113, B => 
                           n4112, ZN => n18476);
   U2728 : OAI21_X1 port map( B1 => n1509, B2 => n17037, A => n1508, ZN => 
                           n18299);
   U2729 : INV_X1 port map( A => n1384, ZN => n17916);
   U2730 : INV_X1 port map( A => n18508, ZN => n510);
   U2733 : INV_X1 port map( A => n18441, ZN => n513);
   U2736 : OAI21_X1 port map( B1 => n17513, B2 => n4273, A => n4705, ZN => 
                           n17696);
   U2737 : INV_X1 port map( A => n18506, ZN => n515);
   U2738 : AND2_X1 port map( A1 => n18251, A2 => n18017, ZN => n17961);
   U2739 : AND2_X1 port map( A1 => n18020, A2 => n18017, ZN => n17959);
   U2741 : NOR2_X1 port map( A1 => n17021, A2 => n17020, ZN => n17854);
   U2742 : INV_X1 port map( A => n18172, ZN => n516);
   U2743 : AND2_X1 port map( A1 => n1665, A2 => n1667, ZN => n17781);
   U2745 : INV_X1 port map( A => n17601, ZN => n517);
   U2746 : INV_X1 port map( A => n19560, ZN => n18188);
   U2748 : OR2_X1 port map( A1 => n17059, A2 => n17058, ZN => n817);
   U2751 : OAI211_X1 port map( C1 => n387, C2 => n1666, A => n4286, B => n4285,
                           ZN => n17872);
   U2752 : INV_X1 port map( A => n17939, ZN => n519);
   U2753 : AND2_X1 port map( A1 => n17008, A2 => n2827, ZN => n17715);
   U2754 : INV_X1 port map( A => n17667, ZN => n824);
   U2755 : OR2_X1 port map( A1 => n2819, A2 => n17710, ZN => n1363);
   U2758 : INV_X1 port map( A => n18402, ZN => n521);
   U2759 : INV_X1 port map( A => n18236, ZN => n522);
   U2760 : OAI21_X1 port map( B1 => n17467, B2 => n4246, A => n1481, ZN => 
                           n16674);
   U2761 : INV_X1 port map( A => n18178, ZN => n523);
   U2762 : AND3_X1 port map( A1 => n4900, A2 => n4901, A3 => n16700, ZN => 
                           n5814);
   U2763 : OAI21_X1 port map( B1 => n422, B2 => n16782, A => n16781, ZN => 
                           n17902);
   U2764 : INV_X1 port map( A => n17941, ZN => n525);
   U2767 : NAND3_X1 port map( A1 => n1387, A2 => n17436, A3 => n16828, ZN => 
                           n19560);
   U2768 : AND2_X1 port map( A1 => n1253, A2 => n1252, ZN => n17292);
   U2770 : OR2_X1 port map( A1 => n16906, A2 => n17566, ZN => n15892);
   U2771 : OR2_X1 port map( A1 => n16787, A2 => n2826, ZN => n1226);
   U2772 : AND2_X1 port map( A1 => n29513, A2 => n17570, ZN => n17318);
   U2773 : OR2_X1 port map( A1 => n17361, A2 => n17365, ZN => n15717);
   U2774 : NOR3_X1 port map( A1 => n17512, A2 => n4273, A3 => n17830, ZN => 
                           n4272);
   U2776 : INV_X1 port map( A => n6465, ZN => n1181);
   U2777 : INV_X1 port map( A => n16883, ZN => n17526);
   U2779 : AND2_X1 port map( A1 => n17467, A2 => n4246, ZN => n784);
   U2780 : OR2_X1 port map( A1 => n16543, A2 => n17120, ZN => n17462);
   U2781 : OR2_X1 port map( A1 => n2768, A2 => n17229, ZN => n1307);
   U2782 : NOR2_X1 port map( A1 => n17279, A2 => n17278, ZN => n779);
   U2784 : AND2_X1 port map( A1 => n2122, A2 => n17552, ZN => n17051);
   U2785 : XNOR2_X1 port map( A => n16402, B => n16403, ZN => n16883);
   U2786 : OR2_X1 port map( A1 => n17396, A2 => n14871, ZN => n16825);
   U2787 : INV_X1 port map( A => n17262, ZN => n1657);
   U2789 : NOR2_X1 port map( A1 => n424, A2 => n16879, ZN => n17384);
   U2790 : INV_X1 port map( A => n4246, ZN => n528);
   U2791 : OR2_X1 port map( A1 => n17293, A2 => n17393, ZN => n1253);
   U2793 : OR2_X1 port map( A1 => n17830, A2 => n17829, ZN => n16547);
   U2795 : AOI21_X1 port map( B1 => n29559, B2 => n1466, A => n16860, ZN => 
                           n1465);
   U2796 : AND2_X1 port map( A1 => n17569, A2 => n29138, ZN => n4317);
   U2797 : NOR2_X1 port map( A1 => n17229, A2 => n17569, ZN => n1507);
   U2798 : INV_X1 port map( A => n17106, ZN => n796);
   U2801 : INV_X1 port map( A => n6002, ZN => n16790);
   U2802 : AND3_X1 port map( A1 => n17275, A2 => n17277, A3 => n17276, ZN => 
                           n780);
   U2803 : AOI21_X1 port map( B1 => n29737, B2 => n1482, A => n17464, ZN => 
                           n17094);
   U2804 : OR2_X1 port map( A1 => n17258, A2 => n1438, ZN => n1437);
   U2805 : OR2_X1 port map( A1 => n16541, A2 => n16810, ZN => n16543);
   U2807 : OR2_X1 port map( A1 => n4316, A2 => n17566, ZN => n6417);
   U2808 : INV_X1 port map( A => n17437, ZN => n529);
   U2809 : INV_X1 port map( A => n17396, ZN => n17294);
   U2811 : INV_X1 port map( A => n17528, ZN => n17158);
   U2812 : INV_X1 port map( A => n17375, ZN => n530);
   U2813 : XNOR2_X1 port map( A => n6650, B => n6649, ZN => n17542);
   U2818 : INV_X1 port map( A => n16706, ZN => n531);
   U2820 : BUF_X1 port map( A => n16736, Z => n17488);
   U2821 : INV_X1 port map( A => n17315, ZN => n532);
   U2826 : XNOR2_X1 port map( A => n16507, B => n16508, ZN => n17452);
   U2827 : INV_X1 port map( A => n17277, ZN => n17001);
   U2828 : INV_X1 port map( A => n17124, ZN => n1816);
   U2829 : INV_X1 port map( A => n17467, ZN => n1482);
   U2832 : CLKBUF_X1 port map( A => n16668, Z => n17258);
   U2833 : XNOR2_X1 port map( A => n16142, B => n1575, ZN => n1438);
   U2834 : XNOR2_X1 port map( A => n14914, B => n14913, ZN => n17397);
   U2835 : XNOR2_X1 port map( A => n15653, B => n15652, ZN => n17552);
   U2837 : XNOR2_X1 port map( A => n16420, B => n16419, ZN => n17528);
   U2838 : INV_X1 port map( A => n17393, ZN => n533);
   U2840 : INV_X1 port map( A => n16803, ZN => n534);
   U2841 : INV_X1 port map( A => n15731, ZN => n535);
   U2843 : XNOR2_X1 port map( A => n16064, B => n16063, ZN => n17097);
   U2844 : INV_X1 port map( A => n17062, ZN => n536);
   U2846 : XNOR2_X1 port map( A => n15564, B => n6929, ZN => n16937);
   U2847 : XNOR2_X1 port map( A => n1778, B => n1348, ZN => n17356);
   U2849 : XNOR2_X1 port map( A => n15794, B => n15793, ZN => n17545);
   U2851 : XNOR2_X1 port map( A => n6160, B => n6158, ZN => n17137);
   U2852 : XNOR2_X1 port map( A => n15778, B => n15777, ZN => n6649);
   U2854 : XNOR2_X1 port map( A => n16163, B => n16164, ZN => n17463);
   U2857 : INV_X1 port map( A => n29632, ZN => n542);
   U2858 : XNOR2_X1 port map( A => n16434, B => n4323, ZN => n16050);
   U2859 : XNOR2_X1 port map( A => n15982, B => n15940, ZN => n16201);
   U2860 : XNOR2_X1 port map( A => n16233, B => n1259, ZN => n1258);
   U2861 : XNOR2_X1 port map( A => n14719, B => n16422, ZN => n16145);
   U2862 : INV_X1 port map( A => n16278, ZN => n16281);
   U2863 : XNOR2_X1 port map( A => n1310, B => n15668, ZN => n16278);
   U2864 : NAND2_X1 port map( A1 => n14866, A2 => n4324, ZN => n4323);
   U2865 : INV_X1 port map( A => n16232, ZN => n769);
   U2867 : XNOR2_X1 port map( A => n15900, B => n16023, ZN => n16302);
   U2868 : AND2_X1 port map( A1 => n14800, A2 => n2190, ZN => n15760);
   U2869 : INV_X1 port map( A => n16304, ZN => n16131);
   U2870 : XNOR2_X1 port map( A => n16230, B => n16090, ZN => n1259);
   U2873 : XNOR2_X1 port map( A => n16084, B => n2116, ZN => n16205);
   U2874 : AND2_X1 port map( A1 => n6760, A2 => n6758, ZN => n16585);
   U2876 : NAND2_X1 port map( A1 => n14911, A2 => n14910, ZN => n16070);
   U2880 : AND3_X1 port map( A1 => n6090, A2 => n6089, A3 => n6088, ZN => 
                           n15992);
   U2882 : NOR2_X1 port map( A1 => n14528, A2 => n14527, ZN => n16024);
   U2883 : NOR2_X1 port map( A1 => n2208, A2 => n2207, ZN => n15565);
   U2884 : NAND3_X1 port map( A1 => n14673, A2 => n14674, A3 => n2699, ZN => 
                           n2700);
   U2887 : OAI21_X1 port map( B1 => n4955, B2 => n4957, A => n14110, ZN => 
                           n16332);
   U2889 : OAI211_X1 port map( C1 => n14532, C2 => n14533, A => n14531, B => 
                           n14530, ZN => n16052);
   U2890 : OR2_X1 port map( A1 => n15131, A2 => n15132, ZN => n1597);
   U2892 : OAI211_X1 port map( C1 => n14940, C2 => n15406, A => n14939, B => 
                           n14938, ZN => n16241);
   U2893 : OAI21_X1 port map( B1 => n15227, B2 => n1149, A => n1148, ZN => 
                           n3923);
   U2894 : OR2_X1 port map( A1 => n756, A2 => n15288, ZN => n4184);
   U2895 : INV_X1 port map( A => n16172, ZN => n543);
   U2896 : AND2_X1 port map( A1 => n14855, A2 => n14856, ZN => n1067);
   U2897 : AND2_X1 port map( A1 => n15373, A2 => n15374, ZN => n1662);
   U2899 : OAI22_X1 port map( A1 => n15353, A2 => n5238, B1 => n14191, B2 => 
                           n15228, ZN => n16176);
   U2901 : INV_X1 port map( A => n15458, ZN => n1701);
   U2902 : BUF_X1 port map( A => n14882, Z => n14884);
   U2903 : INV_X1 port map( A => n15185, ZN => n972);
   U2904 : MUX2_X1 port map( A => n15187, B => n13818, S => n15190, Z => n13819
                           );
   U2905 : AND2_X1 port map( A1 => n15310, A2 => n15272, ZN => n1095);
   U2906 : NAND3_X1 port map( A1 => n4259, A2 => n13732, A3 => n14070, ZN => 
                           n15373);
   U2907 : OAI21_X1 port map( B1 => n14737, B2 => n15009, A => n837, ZN => 
                           n14738);
   U2909 : OAI211_X1 port map( C1 => n15275, C2 => n15274, A => n15514, B => 
                           n1328, ZN => n1518);
   U2910 : OR2_X1 port map( A1 => n14220, A2 => n15047, ZN => n3615);
   U2912 : OR2_X1 port map( A1 => n15371, A2 => n15370, ZN => n683);
   U2914 : AND2_X1 port map( A1 => n15290, A2 => n15292, ZN => n15040);
   U2916 : INV_X1 port map( A => n15115, ZN => n544);
   U2917 : OR2_X1 port map( A1 => n29380, A2 => n15394, ZN => n1326);
   U2919 : INV_X1 port map( A => n15001, ZN => n1745);
   U2922 : AND2_X1 port map( A1 => n14835, A2 => n2456, ZN => n2455);
   U2923 : INV_X1 port map( A => n15447, ZN => n15322);
   U2924 : INV_X1 port map( A => n15117, ZN => n1001);
   U2925 : INV_X1 port map( A => n15190, ZN => n14785);
   U2926 : OR2_X1 port map( A1 => n15456, A2 => n28803, ZN => n3079);
   U2928 : INV_X1 port map( A => n15160, ZN => n545);
   U2930 : INV_X1 port map( A => n15119, ZN => n1005);
   U2931 : INV_X1 port map( A => n15190, ZN => n547);
   U2933 : AND2_X1 port map( A1 => n5666, A2 => n2304, ZN => n15155);
   U2936 : INV_X1 port map( A => n15444, ZN => n548);
   U2939 : AND2_X1 port map( A1 => n14550, A2 => n14549, ZN => n1809);
   U2941 : NAND3_X1 port map( A1 => n14441, A2 => n14442, A3 => n14443, ZN => 
                           n14923);
   U2942 : INV_X1 port map( A => n15127, ZN => n1744);
   U2945 : INV_X1 port map( A => n15102, ZN => n549);
   U2946 : BUF_X1 port map( A => n14153, Z => n15360);
   U2947 : AND3_X1 port map( A1 => n14904, A2 => n14905, A3 => n14906, ZN => 
                           n14908);
   U2948 : INV_X1 port map( A => n15152, ZN => n5198);
   U2949 : INV_X1 port map( A => n15222, ZN => n550);
   U2950 : INV_X1 port map( A => n15123, ZN => n551);
   U2952 : NAND4_X1 port map( A1 => n4435, A2 => n4432, A3 => n13688, A4 => 
                           n4431, ZN => n14992);
   U2953 : AOI21_X1 port map( B1 => n13773, B2 => n13774, A => n13772, ZN => 
                           n14963);
   U2956 : AND2_X1 port map( A1 => n1628, A2 => n1629, ZN => n1627);
   U2957 : OAI21_X1 port map( B1 => n13793, B2 => n13217, A => n13216, ZN => 
                           n15085);
   U2958 : INV_X1 port map( A => n15182, ZN => n552);
   U2960 : OR2_X1 port map( A1 => n13797, A2 => n13796, ZN => n1569);
   U2962 : AND2_X1 port map( A1 => n13709, A2 => n13708, ZN => n15246);
   U2963 : BUF_X1 port map( A => n14115, Z => n15248);
   U2964 : NAND2_X1 port map( A1 => n14139, A2 => n14140, ZN => n4992);
   U2966 : OAI21_X1 port map( B1 => n14770, B2 => n14771, A => n14769, ZN => 
                           n14713);
   U2967 : INV_X1 port map( A => n15456, ZN => n553);
   U2970 : AOI21_X1 port map( B1 => n830, B2 => n14273, A => n4666, ZN => 
                           n15513);
   U2971 : OAI21_X1 port map( B1 => n815, B2 => n13903, A => n814, ZN => n13904
                           );
   U2972 : NOR2_X1 port map( A1 => n13751, A2 => n13750, ZN => n15151);
   U2976 : OR2_X1 port map( A1 => n4074, A2 => n14168, ZN => n998);
   U2977 : OR2_X1 port map( A1 => n5409, A2 => n14437, ZN => n727);
   U2979 : OR2_X1 port map( A1 => n4837, A2 => n28986, ZN => n5015);
   U2982 : INV_X1 port map( A => n4666, ZN => n829);
   U2984 : AND2_X1 port map( A1 => n11372, A2 => n1580, ZN => n1776);
   U2988 : NAND3_X1 port map( A1 => n14429, A2 => n14428, A3 => n28199, ZN => 
                           n14430);
   U2989 : INV_X1 port map( A => n4893, ZN => n14355);
   U2990 : CLKBUF_X1 port map( A => n13257, Z => n14320);
   U2991 : AND2_X1 port map( A1 => n14244, A2 => n28172, ZN => n956);
   U2992 : AOI21_X1 port map( B1 => n13903, B2 => n389, A => n1661, ZN => n1660
                           );
   U2993 : OR2_X1 port map( A1 => n1320, A2 => n14452, ZN => n1322);
   U2994 : BUF_X1 port map( A => n13775, Z => n14250);
   U2995 : INV_X1 port map( A => n1742, ZN => n13614);
   U2996 : INV_X1 port map( A => n28804, ZN => n4012);
   U2997 : AND2_X1 port map( A1 => n29589, A2 => n4425, ZN => n815);
   U2998 : OR2_X1 port map( A1 => n13999, A2 => n14038, ZN => n1016);
   U2999 : AND2_X1 port map( A1 => n14480, A2 => n13936, ZN => n644);
   U3002 : XNOR2_X1 port map( A => n13225, B => n4041, ZN => n14043);
   U3003 : INV_X1 port map( A => n13595, ZN => n14146);
   U3004 : INV_X1 port map( A => n13716, ZN => n13903);
   U3005 : INV_X1 port map( A => n14158, ZN => n14474);
   U3006 : AND2_X1 port map( A1 => n29589, A2 => n13902, ZN => n1661);
   U3007 : OR3_X1 port map( A1 => n14285, A2 => n14083, A3 => n14084, ZN => 
                           n14283);
   U3008 : INV_X1 port map( A => n14217, ZN => n555);
   U3011 : INV_X1 port map( A => n14322, ZN => n1346);
   U3013 : INV_X1 port map( A => n14327, ZN => n14323);
   U3014 : INV_X1 port map( A => n5531, ZN => n6351);
   U3015 : AND2_X1 port map( A1 => n14593, A2 => n14101, ZN => n12938);
   U3016 : XNOR2_X1 port map( A => n13276, B => n13275, ZN => n14053);
   U3017 : INV_X1 port map( A => n13837, ZN => n556);
   U3018 : INV_X1 port map( A => n14381, ZN => n557);
   U3019 : INV_X1 port map( A => n14479, ZN => n558);
   U3020 : XNOR2_X1 port map( A => n12526, B => n12525, ZN => n13874);
   U3021 : XNOR2_X1 port map( A => n13041, B => n1956, ZN => n14126);
   U3022 : INV_X1 port map( A => n14122, ZN => n559);
   U3023 : XNOR2_X1 port map( A => n12710, B => n12709, ZN => n14200);
   U3024 : INV_X1 port map( A => n14309, ZN => n560);
   U3025 : XNOR2_X1 port map( A => n3624, B => n13011, ZN => n4166);
   U3026 : INV_X1 port map( A => n1368, ZN => n13901);
   U3027 : INV_X1 port map( A => n14083, ZN => n561);
   U3029 : XNOR2_X1 port map( A => n13498, B => n13499, ZN => n13589);
   U3030 : XNOR2_X1 port map( A => n11370, B => n11369, ZN => n14101);
   U3032 : INV_X1 port map( A => n14435, ZN => n562);
   U3033 : XNOR2_X1 port map( A => n12439, B => n12438, ZN => n14399);
   U3035 : XNOR2_X1 port map( A => n13367, B => n13368, ZN => n13716);
   U3038 : XNOR2_X1 port map( A => n12821, B => n12820, ZN => n13953);
   U3039 : XNOR2_X1 port map( A => n12694, B => n12695, ZN => n14455);
   U3040 : INV_X1 port map( A => n14238, ZN => n563);
   U3041 : XNOR2_X1 port map( A => n13268, B => n13267, ZN => n13816);
   U3042 : XNOR2_X1 port map( A => n11410, B => n3687, ZN => n13943);
   U3043 : XNOR2_X1 port map( A => n12873, B => n12874, ZN => n12878);
   U3045 : XNOR2_X1 port map( A => n12832, B => n12829, ZN => n1085);
   U3046 : XNOR2_X1 port map( A => n12901, B => n1780, ZN => n12902);
   U3047 : INV_X1 port map( A => n14123, ZN => n564);
   U3049 : XNOR2_X1 port map( A => n12884, B => n12885, ZN => n4041);
   U3051 : XNOR2_X1 port map( A => n13101, B => n13348, ZN => n13246);
   U3052 : INV_X1 port map( A => n12461, ZN => n13298);
   U3053 : XNOR2_X1 port map( A => n12504, B => n12813, ZN => n13521);
   U3054 : AND2_X1 port map( A1 => n5468, A2 => n5467, ZN => n13227);
   U3055 : XNOR2_X1 port map( A => n13297, B => n1664, ZN => n13501);
   U3057 : OR2_X1 port map( A1 => n6645, A2 => n15576, ZN => n961);
   U3058 : INV_X1 port map( A => n6645, ZN => n962);
   U3059 : XNOR2_X1 port map( A => n12799, B => n1293, ZN => n13346);
   U3060 : NOR2_X1 port map( A1 => n11407, A2 => n5076, ZN => n12747);
   U3061 : NAND2_X1 port map( A1 => n11931, A2 => n1491, ZN => n1293);
   U3065 : BUF_X1 port map( A => n12608, Z => n13359);
   U3066 : AND2_X1 port map( A1 => n4017, A2 => n11956, ZN => n860);
   U3067 : NAND3_X1 port map( A1 => n2604, A2 => n12002, A3 => n2603, ZN => 
                           n12879);
   U3068 : AND2_X1 port map( A1 => n4102, A2 => n12130, ZN => n13538);
   U3071 : INV_X1 port map( A => n12529, ZN => n565);
   U3077 : OAI211_X1 port map( C1 => n12256, C2 => n11598, A => n11597, B => 
                           n11596, ZN => n13504);
   U3078 : NAND2_X1 port map( A1 => n11691, A2 => n11690, ZN => n13043);
   U3079 : AND4_X1 port map( A1 => n10955, A2 => n10954, A3 => n10953, A4 => 
                           n10952, ZN => n13069);
   U3082 : OR2_X1 port map( A1 => n12280, A2 => n4105, ZN => n12284);
   U3090 : OR2_X1 port map( A1 => n12103, A2 => n12164, ZN => n705);
   U3091 : OR2_X1 port map( A1 => n375, A2 => n776, ZN => n11541);
   U3092 : OR2_X1 port map( A1 => n12027, A2 => n1291, ZN => n1107);
   U3093 : AOI22_X1 port map( A1 => n11862, A2 => n11861, B1 => n11860, B2 => 
                           n11947, ZN => n1526);
   U3094 : INV_X1 port map( A => n12288, ZN => n1103);
   U3095 : INV_X1 port map( A => n11844, ZN => n706);
   U3096 : OAI21_X1 port map( B1 => n12177, B2 => n11413, A => n11412, ZN => 
                           n12788);
   U3097 : AND2_X1 port map( A1 => n1484, A2 => n11715, ZN => n11650);
   U3099 : OR2_X1 port map( A1 => n11703, A2 => n12205, ZN => n11439);
   U3101 : AND2_X1 port map( A1 => n13086, A2 => n13081, ZN => n11812);
   U3103 : INV_X1 port map( A => n9692, ZN => n12210);
   U3104 : INV_X1 port map( A => n11648, ZN => n1706);
   U3105 : OR2_X1 port map( A1 => n11417, A2 => n11648, ZN => n11714);
   U3106 : AND2_X1 port map( A1 => n12354, A2 => n12352, ZN => n1371);
   U3107 : CLKBUF_X1 port map( A => n12293, Z => n12061);
   U3108 : OR2_X1 port map( A1 => n1890, A2 => n12177, ZN => n1318);
   U3109 : INV_X1 port map( A => n12508, ZN => n1746);
   U3110 : INV_X1 port map( A => n11505, ZN => n12280);
   U3111 : INV_X1 port map( A => n12315, ZN => n566);
   U3113 : INV_X1 port map( A => n11551, ZN => n1453);
   U3115 : INV_X1 port map( A => n11867, ZN => n11360);
   U3117 : OR2_X1 port map( A1 => n5905, A2 => n10935, ZN => n11947);
   U3118 : OAI21_X1 port map( B1 => n10911, B2 => n10452, A => n10451, ZN => 
                           n11876);
   U3119 : INV_X1 port map( A => n11852, ZN => n11547);
   U3122 : INV_X1 port map( A => n11715, ZN => n1485);
   U3123 : NOR2_X1 port map( A1 => n12337, A2 => n11473, ZN => n1292);
   U3128 : INV_X1 port map( A => n12266, ZN => n568);
   U3129 : AND2_X1 port map( A1 => n12508, A2 => n12507, ZN => n11616);
   U3130 : OR2_X1 port map( A1 => n11980, A2 => n12226, ZN => n11981);
   U3132 : AND4_X2 port map( A1 => n10107, A2 => n10104, A3 => n10106, A4 => 
                           n10105, ZN => n12508);
   U3133 : AOI22_X1 port map( A1 => n11107, A2 => n11106, B1 => n11217, B2 => 
                           n11105, ZN => n12577);
   U3135 : OAI21_X1 port map( B1 => n11143, B2 => n11142, A => n1452, ZN => 
                           n11780);
   U3137 : NAND2_X1 port map( A1 => n6720, A2 => n3570, ZN => n11969);
   U3139 : INV_X1 port map( A => n12181, ZN => n570);
   U3142 : INV_X1 port map( A => n12132, ZN => n12265);
   U3144 : INV_X1 port map( A => n11536, ZN => n572);
   U3145 : INV_X1 port map( A => n12146, ZN => n573);
   U3146 : INV_X1 port map( A => n11855, ZN => n574);
   U3148 : INV_X1 port map( A => n11574, ZN => n575);
   U3150 : INV_X1 port map( A => n10863, ZN => n577);
   U3152 : INV_X1 port map( A => n12050, ZN => n12316);
   U3153 : OAI211_X1 port map( C1 => n10844, C2 => n10523, A => n11039, B => 
                           n4145, ZN => n12328);
   U3155 : OR2_X1 port map( A1 => n10542, A2 => n10541, ZN => n989);
   U3156 : OAI211_X1 port map( C1 => n1975, C2 => n2143, A => n1399, B => n1400
                           , ZN => n12163);
   U3157 : AND2_X1 port map( A1 => n10755, A2 => n10756, ZN => n11672);
   U3159 : INV_X1 port map( A => n11463, ZN => n578);
   U3160 : INV_X1 port map( A => n11856, ZN => n579);
   U3161 : AND4_X1 port map( A1 => n2086, A2 => n10642, A3 => n2085, A4 => 
                           n2084, ZN => n11962);
   U3162 : OR2_X1 port map( A1 => n10996, A2 => n10995, ZN => n1786);
   U3165 : NAND2_X1 port map( A1 => n10652, A2 => n10884, ZN => n1261);
   U3166 : INV_X1 port map( A => n11901, ZN => n580);
   U3167 : OR2_X1 port map( A1 => n3801, A2 => n10694, ZN => n12194);
   U3168 : OR2_X1 port map( A1 => n10963, A2 => n10956, ZN => n3413);
   U3169 : INV_X1 port map( A => n10726, ZN => n10928);
   U3171 : AND2_X1 port map( A1 => n10893, A2 => n11290, ZN => n1736);
   U3172 : OR2_X1 port map( A1 => n11082, A2 => n11083, ZN => n1399);
   U3173 : CLKBUF_X1 port map( A => n11323, Z => n11328);
   U3174 : OR2_X1 port map( A1 => n1703, A2 => n1338, ZN => n10526);
   U3176 : OR2_X1 port map( A1 => n10520, A2 => n10884, ZN => n1260);
   U3177 : OR2_X1 port map( A1 => n11241, A2 => n11244, ZN => n787);
   U3178 : INV_X1 port map( A => n28624, ZN => n1357);
   U3179 : AND2_X1 port map( A1 => n11121, A2 => n11119, ZN => n10506);
   U3180 : NOR2_X1 port map( A1 => n969, A2 => n10806, ZN => n10741);
   U3181 : INV_X1 port map( A => n11209, ZN => n11213);
   U3182 : INV_X1 port map( A => n1338, ZN => n1704);
   U3183 : NOR2_X1 port map( A1 => n433, A2 => n11210, ZN => n1975);
   U3190 : INV_X1 port map( A => n28407, ZN => n10998);
   U3193 : OR2_X1 port map( A1 => n11064, A2 => n11067, ZN => n11068);
   U3194 : INV_X1 port map( A => n11199, ZN => n581);
   U3195 : XNOR2_X1 port map( A => n10416, B => n10415, ZN => n11207);
   U3196 : INV_X1 port map( A => n11196, ZN => n3585);
   U3197 : CLKBUF_X1 port map( A => n10882, Z => n11211);
   U3198 : INV_X1 port map( A => n11064, ZN => n11244);
   U3199 : XNOR2_X1 port map( A => n9809, B => n9808, ZN => n10786);
   U3203 : XNOR2_X1 port map( A => n8376, B => n8377, ZN => n11166);
   U3204 : INV_X1 port map( A => n10970, ZN => n1285);
   U3206 : INV_X1 port map( A => n2690, ZN => n11255);
   U3207 : OR2_X1 port map( A1 => n11243, A2 => n11240, ZN => n1760);
   U3208 : OR2_X1 port map( A1 => n11315, A2 => n2690, ZN => n1537);
   U3209 : CLKBUF_X1 port map( A => n10524, Z => n11248);
   U3210 : XNOR2_X1 port map( A => n10301, B => n10300, ZN => n11294);
   U3212 : XNOR2_X1 port map( A => n8775, B => n8774, ZN => n11337);
   U3213 : INV_X1 port map( A => n11149, ZN => n582);
   U3218 : XNOR2_X1 port map( A => n9302, B => n9915, ZN => n10300);
   U3219 : INV_X1 port map( A => n11282, ZN => n584);
   U3221 : INV_X1 port map( A => n11084, ZN => n10883);
   U3222 : INV_X1 port map( A => n1854, ZN => n585);
   U3223 : XNOR2_X1 port map( A => n9968, B => n9967, ZN => n10502);
   U3224 : XNOR2_X1 port map( A => n8620, B => n8621, ZN => n11196);
   U3225 : INV_X1 port map( A => n11033, ZN => n586);
   U3227 : INV_X1 port map( A => n11093, ZN => n587);
   U3229 : XNOR2_X1 port map( A => n9720, B => n9719, ZN => n11226);
   U3231 : INV_X1 port map( A => n10930, ZN => n588);
   U3232 : INV_X1 port map( A => n10984, ZN => n589);
   U3234 : XNOR2_X1 port map( A => n10389, B => n10390, ZN => n11094);
   U3235 : INV_X1 port map( A => n10932, ZN => n590);
   U3236 : XNOR2_X1 port map( A => n10213, B => n10214, ZN => n11066);
   U3237 : INV_X1 port map( A => n10976, ZN => n591);
   U3238 : XNOR2_X1 port map( A => n1761, B => n10187, ZN => n11243);
   U3241 : XNOR2_X1 port map( A => n9629, B => n9379, ZN => n9721);
   U3243 : INV_X1 port map( A => n10752, ZN => n593);
   U3244 : INV_X1 port map( A => n11253, ZN => n594);
   U3246 : INV_X1 port map( A => n11084, ZN => n595);
   U3249 : XNOR2_X1 port map( A => n654, B => n10207, ZN => n9590);
   U3250 : XNOR2_X1 port map( A => n10322, B => n9295, ZN => n9977);
   U3251 : XNOR2_X1 port map( A => n655, B => n10310, ZN => n9956);
   U3253 : AND2_X1 port map( A1 => n2596, A2 => n2597, ZN => n10228);
   U3256 : XNOR2_X1 port map( A => n4479, B => n10353, ZN => n10433);
   U3257 : OR2_X1 port map( A1 => n8606, A2 => n963, ZN => n10246);
   U3259 : INV_X1 port map( A => n9648, ZN => n9900);
   U3262 : XNOR2_X1 port map( A => n9696, B => n10171, ZN => n9596);
   U3269 : AND2_X1 port map( A1 => n2290, A2 => n5330, ZN => n10359);
   U3271 : XNOR2_X1 port map( A => n9426, B => n10357, ZN => n9722);
   U3273 : INV_X1 port map( A => n9505, ZN => n654);
   U3275 : AND2_X1 port map( A1 => n10233, A2 => n8724, ZN => n8606);
   U3277 : AND2_X1 port map( A1 => n843, A2 => n842, ZN => n10064);
   U3281 : NAND4_X1 port map( A1 => n4728, A2 => n8689, A3 => n8690, A4 => 
                           n9024, ZN => n9899);
   U3285 : OR2_X1 port map( A1 => n7575, A2 => n8537, ZN => n1355);
   U3288 : OAI21_X1 port map( B1 => n970, B2 => n8355, A => n8354, ZN => n971);
   U3290 : NAND4_X1 port map( A1 => n9049, A2 => n4730, A3 => n4731, A4 => 
                           n8691, ZN => n10227);
   U3292 : NAND3_X1 port map( A1 => n8417, A2 => n8416, A3 => n8415, ZN => 
                           n10073);
   U3293 : OR2_X1 port map( A1 => n7575, A2 => n8537, ZN => n1416);
   U3294 : MUX2_X1 port map( A => n8960, B => n8959, S => n8958, Z => n9613);
   U3295 : OAI21_X1 port map( B1 => n744, B2 => n8120, A => n5449, ZN => n9992)
                           ;
   U3296 : OAI22_X1 port map( A1 => n9340, A2 => n8755, B1 => n1934, B2 => 
                           n8754, ZN => n8756);
   U3297 : MUX2_X1 port map( A => n7001, B => n7000, S => n9045, Z => n9732);
   U3298 : INV_X1 port map( A => n8993, ZN => n1047);
   U3299 : AND3_X1 port map( A1 => n2861, A2 => n2860, A3 => n2863, ZN => 
                           n10302);
   U3300 : OR2_X1 port map( A1 => n8483, A2 => n440, ZN => n1710);
   U3301 : OR2_X1 port map( A1 => n1788, A2 => n8760, ZN => n1790);
   U3302 : OAI21_X1 port map( B1 => n8426, B2 => n8427, A => n8078, ZN => n8120
                           );
   U3305 : OR2_X1 port map( A1 => n9049, A2 => n9235, ZN => n1117);
   U3306 : NOR2_X1 port map( A1 => n844, A2 => n9137, ZN => n843);
   U3307 : AOI21_X1 port map( B1 => n8920, B2 => n8919, A => n8918, ZN => n9647
                           );
   U3308 : OR2_X1 port map( A1 => n8610, A2 => n9530, ZN => n714);
   U3310 : AND2_X1 port map( A1 => n9135, A2 => n9134, ZN => n844);
   U3311 : AND2_X1 port map( A1 => n6747, A2 => n9374, ZN => n8570);
   U3312 : NOR2_X1 port map( A1 => n9140, A2 => n638, ZN => n637);
   U3313 : OR2_X1 port map( A1 => n5568, A2 => n5945, ZN => n9238);
   U3314 : NOR2_X1 port map( A1 => n8819, A2 => n8594, ZN => n8823);
   U3315 : INV_X1 port map( A => n8058, ZN => n8426);
   U3316 : NOR2_X1 port map( A1 => n9438, A2 => n8777, ZN => n8993);
   U3317 : OR2_X1 port map( A1 => n8931, A2 => n9148, ZN => n8761);
   U3318 : MUX2_X1 port map( A => n8661, B => n8482, S => n9016, Z => n8483);
   U3319 : AND2_X1 port map( A1 => n8961, A2 => n9171, ZN => n9173);
   U3320 : OR2_X1 port map( A1 => n8827, A2 => n8586, ZN => n8465);
   U3321 : INV_X1 port map( A => n8699, ZN => n8403);
   U3322 : OAI211_X1 port map( C1 => n9140, C2 => n8562, A => n8561, B => n1803
                           , ZN => n2336);
   U3323 : OR2_X1 port map( A1 => n1934, A2 => n9133, ZN => n1670);
   U3324 : OR2_X1 port map( A1 => n8764, A2 => n8763, ZN => n9564);
   U3326 : OR2_X1 port map( A1 => n9013, A2 => n9014, ZN => n1615);
   U3327 : AND2_X1 port map( A1 => n4938, A2 => n7091, ZN => n1839);
   U3328 : OAI21_X1 port map( B1 => n8924, B2 => n6718, A => n1934, ZN => n8552
                           );
   U3329 : INV_X1 port map( A => n9037, ZN => n1634);
   U3330 : OR2_X1 port map( A1 => n8782, A2 => n9186, ZN => n8784);
   U3331 : OR2_X1 port map( A1 => n9148, A2 => n8929, ZN => n1528);
   U3332 : OR2_X1 port map( A1 => n8983, A2 => n8981, ZN => n8408);
   U3335 : AND2_X1 port map( A1 => n9125, A2 => n8899, ZN => n1794);
   U3336 : AND2_X1 port map( A1 => n8500, A2 => n8652, ZN => n7906);
   U3337 : INV_X1 port map( A => n1910, ZN => n8430);
   U3338 : INV_X1 port map( A => n9122, ZN => n1793);
   U3339 : CLKBUF_X1 port map( A => n8777, Z => n9208);
   U3340 : OAI21_X1 port map( B1 => n8353, B2 => n8077, A => n8427, ZN => n745)
                           ;
   U3341 : INV_X1 port map( A => n8963, ZN => n9170);
   U3344 : OR2_X1 port map( A1 => n8183, A2 => n8182, ZN => n8980);
   U3345 : INV_X1 port map( A => n9144, ZN => n638);
   U3347 : INV_X1 port map( A => n8981, ZN => n596);
   U3350 : INV_X1 port map( A => n9228, ZN => n597);
   U3351 : OR2_X1 port map( A1 => n7476, A2 => n7475, ZN => n8848);
   U3352 : INV_X1 port map( A => n9139, ZN => n598);
   U3353 : INV_X1 port map( A => n8562, ZN => n599);
   U3355 : AOI21_X1 port map( B1 => n1586, B2 => n1587, A => n1589, ZN => n8326
                           );
   U3356 : INV_X1 port map( A => n8792, ZN => n9035);
   U3357 : INV_X1 port map( A => n9132, ZN => n600);
   U3358 : INV_X1 port map( A => n9134, ZN => n601);
   U3360 : INV_X1 port map( A => n8977, ZN => n602);
   U3362 : OAI211_X1 port map( C1 => n7725, C2 => n8043, A => n7724, B => n7723
                           , ZN => n9007);
   U3363 : INV_X1 port map( A => n8579, ZN => n603);
   U3365 : INV_X1 port map( A => n9171, ZN => n605);
   U3368 : OR2_X1 port map( A1 => n7217, A2 => n742, ZN => n3301);
   U3369 : OAI21_X1 port map( B1 => n5911, B2 => n8247, A => n5910, ZN => n8966
                           );
   U3370 : NAND3_X1 port map( A1 => n1352, A2 => n1351, A3 => n1349, ZN => 
                           n8384);
   U3371 : INV_X1 port map( A => n9421, ZN => n606);
   U3373 : INV_X1 port map( A => n1589, ZN => n1585);
   U3374 : OR2_X1 port map( A1 => n7317, A2 => n7775, ZN => n1586);
   U3375 : INV_X1 port map( A => n8819, ZN => n607);
   U3376 : AOI21_X1 port map( B1 => n1568, B2 => n5256, A => n5255, ZN => n7973
                           );
   U3377 : INV_X1 port map( A => n9016, ZN => n608);
   U3378 : NAND4_X1 port map( A1 => n7182, A2 => n7183, A3 => n7181, A4 => 
                           n7180, ZN => n8733);
   U3380 : OAI211_X1 port map( C1 => n7704, C2 => n7840, A => n7702, B => n7703
                           , ZN => n8792);
   U3382 : AOI22_X1 port map( A1 => n7209, A2 => n7208, B1 => n7207, B2 => 
                           n7206, ZN => n8525);
   U3383 : OR2_X1 port map( A1 => n7766, A2 => n4856, ZN => n4855);
   U3385 : AOI22_X1 port map( A1 => n8052, A2 => n8132, B1 => n8051, B2 => 
                           n8050, ZN => n9363);
   U3386 : INV_X1 port map( A => n9396, ZN => n609);
   U3390 : OR2_X1 port map( A1 => n7385, A2 => n6748, ZN => n9374);
   U3391 : NOR2_X1 port map( A1 => n7316, A2 => n1700, ZN => n1589);
   U3392 : INV_X1 port map( A => n3654, ZN => n771);
   U3393 : AND3_X1 port map( A1 => n7381, A2 => n7380, A3 => n7379, ZN => n8929
                           );
   U3394 : OAI21_X1 port map( B1 => n7864, B2 => n7172, A => n5149, ZN => n5148
                           );
   U3395 : AND2_X1 port map( A1 => n7290, A2 => n7759, ZN => n2630);
   U3396 : OR2_X1 port map( A1 => n8260, A2 => n28614, ZN => n1198);
   U3398 : AND2_X1 port map( A1 => n8044, A2 => n7722, ZN => n889);
   U3399 : INV_X1 port map( A => n1354, ZN => n1350);
   U3400 : BUF_X1 port map( A => n7399, Z => n8304);
   U3401 : BUF_X1 port map( A => n7400, Z => n8305);
   U3404 : AND2_X1 port map( A1 => n7368, A2 => n439, ZN => n1295);
   U3405 : OR2_X1 port map( A1 => n7456, A2 => n7040, ZN => n7645);
   U3406 : OR2_X1 port map( A1 => n7793, A2 => n7150, ZN => n2545);
   U3407 : INV_X1 port map( A => n7283, ZN => n8150);
   U3409 : INV_X1 port map( A => n7742, ZN => n7744);
   U3410 : BUF_X1 port map( A => n7283, Z => n7542);
   U3411 : INV_X1 port map( A => n7793, ZN => n3810);
   U3413 : CLKBUF_X1 port map( A => n7405, Z => n8276);
   U3415 : INV_X1 port map( A => n2804, ZN => n1911);
   U3416 : INV_X1 port map( A => n7456, ZN => n612);
   U3417 : XNOR2_X1 port map( A => n7038, B => Key(154), ZN => n7641);
   U3418 : INV_X1 port map( A => n7349, ZN => n8168);
   U3419 : INV_X1 port map( A => n27742, ZN => n5633);
   U3421 : BUF_X1 port map( A => n7488, Z => n8264);
   U3422 : INV_X1 port map( A => n8173, ZN => n613);
   U3423 : INV_X1 port map( A => n3083, ZN => n653);
   U3424 : BUF_X1 port map( A => n7082, Z => n7303);
   U3425 : XNOR2_X1 port map( A => n7109, B => Key(190), ZN => n7897);
   U3428 : INV_X1 port map( A => n2511, ZN => n1782);
   U3429 : INV_X1 port map( A => n7164, ZN => n614);
   U3430 : INV_X1 port map( A => n7089, ZN => n1354);
   U3431 : CLKBUF_X1 port map( A => n7466, Z => n7946);
   U3432 : CLKBUF_X1 port map( A => n7589, Z => n7960);
   U3433 : INV_X1 port map( A => n8131, ZN => n615);
   U3434 : INV_X1 port map( A => n3482, ZN => n1412);
   U3436 : INV_X1 port map( A => n7839, ZN => n7367);
   U3437 : INV_X1 port map( A => n7817, ZN => n616);
   U3438 : XNOR2_X1 port map( A => n7154, B => Key(30), ZN => n7348);
   U3439 : INV_X1 port map( A => n3752, ZN => n1229);
   U3441 : INV_X1 port map( A => n2350, ZN => n927);
   U3442 : CLKBUF_X1 port map( A => n7150, Z => n7541);
   U3443 : INV_X1 port map( A => n7250, ZN => n617);
   U3444 : XNOR2_X1 port map( A => n6996, B => Key(121), ZN => n7912);
   U3445 : INV_X1 port map( A => n7268, ZN => n618);
   U3447 : CLKBUF_X1 port map( A => Key(73), Z => n2523);
   U3448 : CLKBUF_X1 port map( A => Key(83), Z => n27452);
   U3452 : XNOR2_X1 port map( A => Key(77), B => Plaintext(77), ZN => n7851);
   U3453 : CLKBUF_X1 port map( A => Key(180), Z => n2987);
   U3454 : CLKBUF_X1 port map( A => Key(187), Z => n26825);
   U3455 : INV_X1 port map( A => n7836, ZN => n619);
   U3457 : INV_X1 port map( A => Plaintext(25), ZN => n1609);
   U3458 : INV_X1 port map( A => n3219, ZN => n621);
   U3459 : INV_X1 port map( A => n1179, ZN => n622);
   U3460 : CLKBUF_X1 port map( A => Key(68), Z => n26680);
   U3461 : CLKBUF_X1 port map( A => Key(129), Z => n3276);
   U3464 : INV_X1 port map( A => n3751, ZN => n623);
   U3468 : CLKBUF_X1 port map( A => Key(139), Z => n3501);
   U3469 : CLKBUF_X1 port map( A => Key(48), Z => n3650);
   U3470 : INV_X1 port map( A => n3528, ZN => n625);
   U3471 : INV_X1 port map( A => n7924, ZN => n626);
   U3472 : INV_X1 port map( A => n7626, ZN => n627);
   U3473 : INV_X1 port map( A => n3686, ZN => n628);
   U3474 : CLKBUF_X1 port map( A => Key(32), Z => n3003);
   U3475 : INV_X1 port map( A => n3697, ZN => n629);
   U3479 : CLKBUF_X1 port map( A => Key(98), Z => n3666);
   U3480 : INV_X1 port map( A => n26665, ZN => n630);
   U3481 : INV_X1 port map( A => n8269, ZN => n631);
   U3482 : CLKBUF_X1 port map( A => Key(182), Z => n3710);
   U3487 : CLKBUF_X1 port map( A => Key(130), Z => n26032);
   U3489 : CLKBUF_X1 port map( A => Key(119), Z => n27298);
   U3490 : INV_X1 port map( A => n3423, ZN => n632);
   U3491 : CLKBUF_X1 port map( A => Key(91), Z => n3134);
   U3492 : INV_X1 port map( A => n3742, ZN => n633);
   U3494 : INV_X1 port map( A => n1175, ZN => n634);
   U3495 : INV_X1 port map( A => n2325, ZN => n635);
   U3498 : NAND2_X1 port map( A1 => n9140, A2 => n638, ZN => n2928);
   U3499 : NAND2_X1 port map( A1 => n8561, A2 => n636, ZN => n8567);
   U3500 : NOR2_X1 port map( A1 => n9140, A2 => n599, ZN => n636);
   U3501 : NAND2_X1 port map( A1 => n599, A2 => n637, ZN => n8189);
   U3503 : NAND2_X1 port map( A1 => n641, A2 => n28391, ZN => n23048);
   U3504 : OAI21_X1 port map( B1 => n641, B2 => n23470, A => n23469, ZN => 
                           n23471);
   U3505 : INV_X1 port map( A => n640, ZN => n639);
   U3506 : OAI211_X1 port map( C1 => n661, C2 => n641, A => n23193, B => n640, 
                           ZN => n660);
   U3508 : NAND2_X1 port map( A1 => n14474, A2 => n644, ZN => n643);
   U3509 : XNOR2_X2 port map( A => n11735, B => n11734, ZN => n14158);
   U3510 : NAND2_X1 port map( A1 => n13934, A2 => n14480, ZN => n646);
   U3511 : NAND3_X1 port map( A1 => n21410, A2 => n21408, A3 => n21412, ZN => 
                           n647);
   U3513 : NAND3_X1 port map( A1 => n20663, A2 => n21047, A3 => n4937, ZN => 
                           n648);
   U3514 : NAND2_X1 port map( A1 => n490, A2 => n651, ZN => n650);
   U3515 : NOR2_X1 port map( A1 => n21171, A2 => n21047, ZN => n651);
   U3517 : NAND2_X1 port map( A1 => n652, A2 => n10523, ZN => n11041);
   U3520 : XNOR2_X1 port map( A => n654, B => n9941, ZN => n8835);
   U3521 : XNOR2_X1 port map( A => n654, B => n10271, ZN => n10274);
   U3522 : OAI21_X2 port map( B1 => n8983, B2 => n8411, A => n8410, ZN => n655)
                           ;
   U3523 : XNOR2_X1 port map( A => n655, B => n1187, ZN => n9484);
   U3524 : XNOR2_X1 port map( A => n655, B => n10073, ZN => n8418);
   U3525 : XNOR2_X1 port map( A => n10272, B => n655, ZN => n8844);
   U3526 : XNOR2_X1 port map( A => n655, B => n10353, ZN => n10354);
   U3527 : NAND2_X1 port map( A1 => n21143, A2 => n21117, ZN => n21146);
   U3528 : AOI21_X1 port map( B1 => n21145, B2 => n492, A => n21119, ZN => n657
                           );
   U3529 : NAND2_X1 port map( A1 => n657, A2 => n21141, ZN => n656);
   U3530 : OAI21_X2 port map( B1 => n19781, B2 => n20081, A => n19780, ZN => 
                           n21143);
   U3531 : NAND2_X1 port map( A1 => n492, A2 => n20852, ZN => n658);
   U3533 : NAND2_X1 port map( A1 => n659, A2 => n21314, ZN => n3531);
   U3534 : NAND2_X1 port map( A1 => n659, A2 => n21138, ZN => n21139);
   U3535 : NAND2_X1 port map( A1 => n20723, A2 => n20724, ZN => n659);
   U3536 : NAND2_X1 port map( A1 => n24324, A2 => n24677, ZN => n3480);
   U3537 : NAND2_X1 port map( A1 => n24397, A2 => n24678, ZN => n24324);
   U3538 : NAND3_X2 port map( A1 => n660, A2 => n2046, A3 => n662, ZN => n24678
                           );
   U3539 : INV_X1 port map( A => n23318, ZN => n661);
   U3540 : NAND2_X1 port map( A1 => n1740, A2 => n23654, ZN => n662);
   U3542 : NAND2_X1 port map( A1 => n26734, A2 => n26995, ZN => n663);
   U3543 : NAND2_X1 port map( A1 => n29486, A2 => n25972, ZN => n664);
   U3544 : OAI21_X1 port map( B1 => n11782, B2 => n11550, A => n11785, ZN => 
                           n666);
   U3546 : NAND2_X1 port map( A1 => n11786, A2 => n11502, ZN => n667);
   U3547 : NAND2_X1 port map( A1 => n17793, A2 => n513, ZN => n668);
   U3549 : NAND2_X1 port map( A1 => n17739, A2 => n17740, ZN => n669);
   U3550 : NAND2_X1 port map( A1 => n17738, A2 => n671, ZN => n670);
   U3551 : NAND2_X1 port map( A1 => n510, A2 => n18072, ZN => n18076);
   U3553 : AOI21_X1 port map( B1 => n24029, B2 => n24651, A => n673, ZN => 
                           n6664);
   U3554 : NAND2_X1 port map( A1 => n3061, A2 => n629, ZN => n672);
   U3556 : NAND3_X1 port map( A1 => n24657, A2 => n24656, A3 => n673, ZN => 
                           n24658);
   U3557 : NAND2_X1 port map( A1 => n17658, A2 => n17657, ZN => n993);
   U3559 : OR2_X1 port map( A1 => n17436, A2 => n17437, ZN => n4988);
   U3560 : NAND2_X1 port map( A1 => n15489, A2 => n15485, ZN => n5644);
   U3561 : NAND3_X1 port map( A1 => n1541, A2 => n1540, A3 => n21535, ZN => 
                           n1539);
   U3563 : NAND3_X1 port map( A1 => n23271, A2 => n23272, A3 => n23273, ZN => 
                           n674);
   U3564 : XNOR2_X1 port map( A => n675, B => n26003, ZN => Ciphertext(6));
   U3565 : NAND3_X1 port map( A1 => n26002, A2 => n26000, A3 => n26001, ZN => 
                           n675);
   U3567 : NOR2_X1 port map( A1 => n26180, A2 => n24204, ZN => n25611);
   U3568 : NAND2_X1 port map( A1 => n1480, A2 => n18340, ZN => n18347);
   U3574 : NAND3_X1 port map( A1 => n7765, A2 => n4855, A3 => n7764, ZN => 
                           n1910);
   U3575 : OAI21_X1 port map( B1 => n23486, B2 => n23154, A => n23155, ZN => 
                           n1390);
   U3576 : NAND3_X1 port map( A1 => n678, A2 => n11529, A3 => n13087, ZN => 
                           n11530);
   U3577 : NAND2_X1 port map( A1 => n13084, A2 => n11980, ZN => n678);
   U3579 : NAND2_X1 port map( A1 => n16890, A2 => n17078, ZN => n679);
   U3580 : NAND3_X1 port map( A1 => n2216, A2 => n18600, A3 => n2215, ZN => 
                           n2214);
   U3582 : NAND2_X1 port map( A1 => n26817, A2 => n27025, ZN => n26816);
   U3583 : INV_X1 port map( A => n17838, ZN => n17839);
   U3586 : NAND2_X1 port map( A1 => n17715, A2 => n17431, ZN => n5329);
   U3587 : NAND3_X1 port map( A1 => n6686, A2 => n24547, A3 => n23126, ZN => 
                           n865);
   U3588 : NAND2_X1 port map( A1 => n19938, A2 => n506, ZN => n681);
   U3591 : NAND2_X1 port map( A1 => n17663, A2 => n17947, ZN => n757);
   U3592 : NAND3_X1 port map( A1 => n17596, A2 => n686, A3 => n29024, ZN => 
                           n17594);
   U3595 : NAND2_X1 port map( A1 => n13872, A2 => n13703, ZN => n4837);
   U3597 : OAI211_X2 port map( C1 => n14884, C2 => n14585, A => n14584, B => 
                           n688, ZN => n16256);
   U3598 : NAND2_X1 port map( A1 => n14884, A2 => n14582, ZN => n688);
   U3599 : INV_X1 port map( A => n690, ZN => n689);
   U3602 : NAND2_X1 port map( A1 => n691, A2 => n14275, ZN => n14834);
   U3603 : NAND2_X1 port map( A1 => n14361, A2 => n28507, ZN => n691);
   U3604 : OAI21_X2 port map( B1 => n4656, B2 => n19517, A => n19516, ZN => 
                           n21806);
   U3605 : NAND3_X1 port map( A1 => n17416, A2 => n3234, A3 => n15811, ZN => 
                           n17417);
   U3606 : INV_X1 port map( A => n8790, ZN => n7606);
   U3607 : NAND2_X1 port map( A1 => n8414, A2 => n8788, ZN => n8790);
   U3610 : INV_X1 port map( A => n15047, ZN => n694);
   U3611 : NAND2_X1 port map( A1 => n15336, A2 => n15047, ZN => n695);
   U3612 : OAI21_X1 port map( B1 => n18441, B2 => n523, A => n696, ZN => n18098
                           );
   U3613 : NAND2_X1 port map( A1 => n18441, A2 => n18179, ZN => n696);
   U3614 : NOR2_X2 port map( A1 => n19012, A2 => n19011, ZN => n21292);
   U3618 : NAND2_X1 port map( A1 => n21090, A2 => n5817, ZN => n20801);
   U3620 : AND2_X1 port map( A1 => n20790, A2 => n20791, ZN => n698);
   U3621 : OAI21_X1 port map( B1 => n28203, B2 => n12206, A => n1221, ZN => 
                           n11833);
   U3622 : NAND2_X1 port map( A1 => n699, A2 => n4270, ZN => n5791);
   U3623 : NAND2_X1 port map( A1 => n2296, A2 => n700, ZN => n20789);
   U3624 : NAND2_X1 port map( A1 => n20802, A2 => n701, ZN => n700);
   U3625 : NAND2_X1 port map( A1 => n20109, A2 => n20322, ZN => n703);
   U3626 : NAND2_X1 port map( A1 => n15253, A2 => n707, ZN => n15254);
   U3627 : NAND3_X1 port map( A1 => n15251, A2 => n15250, A3 => n15252, ZN => 
                           n707);
   U3628 : NAND3_X2 port map( A1 => n3765, A2 => n708, A3 => n2288, ZN => 
                           n12760);
   U3629 : NAND3_X1 port map( A1 => n1061, A2 => n12400, A3 => n11800, ZN => 
                           n708);
   U3630 : XNOR2_X1 port map( A => n18608, B => n19299, ZN => n19683);
   U3632 : NOR2_X1 port map( A1 => n26505, A2 => n26506, ZN => n26638);
   U3633 : NOR2_X1 port map( A1 => n24846, A2 => n709, ZN => n24857);
   U3634 : NOR2_X1 port map( A1 => n26361, A2 => n26425, ZN => n709);
   U3635 : XNOR2_X1 port map( A => n710, B => n21573, ZN => n21584);
   U3636 : XNOR2_X1 port map( A => n21566, B => n22271, ZN => n710);
   U3640 : NAND2_X1 port map( A1 => n14150, A2 => n14382, ZN => n713);
   U3643 : XNOR2_X1 port map( A => n22315, B => n22077, ZN => n21341);
   U3644 : XNOR2_X1 port map( A => n22596, B => n21325, ZN => n22315);
   U3645 : NAND2_X1 port map( A1 => n26648, A2 => n29532, ZN => n26979);
   U3647 : NAND2_X1 port map( A1 => n2708, A2 => n22084, ZN => n1635);
   U3648 : OR2_X1 port map( A1 => n7640, A2 => n612, ZN => n983);
   U3650 : OR3_X1 port map( A1 => n14380, A2 => n13837, A3 => n14381, ZN => 
                           n6105);
   U3651 : INV_X1 port map( A => n24616, ZN => n1262);
   U3653 : NAND2_X1 port map( A1 => n16895, A2 => n16896, ZN => n715);
   U3656 : NAND2_X1 port map( A1 => n6072, A2 => n8760, ZN => n8930);
   U3657 : INV_X1 port map( A => n15010, ZN => n14865);
   U3658 : NAND2_X1 port map( A1 => n14863, A2 => n15370, ZN => n15010);
   U3659 : AND2_X1 port map( A1 => n11308, A2 => n11053, ZN => n10852);
   U3660 : OAI21_X1 port map( B1 => n2132, B2 => n24322, A => n24324, ZN => 
                           n2131);
   U3661 : OAI21_X1 port map( B1 => n20639, B2 => n717, A => n20638, ZN => 
                           n20640);
   U3662 : OAI21_X1 port map( B1 => n20633, B2 => n28538, A => n20632, ZN => 
                           n717);
   U3663 : NAND3_X1 port map( A1 => n20202, A2 => n20302, A3 => n20304, ZN => 
                           n19948);
   U3664 : NAND2_X1 port map( A1 => n719, A2 => n3717, ZN => n3716);
   U3665 : NAND2_X1 port map( A1 => n810, A2 => n3954, ZN => n719);
   U3666 : MUX2_X2 port map( A => n24393, B => n24394, S => n24683, Z => n25689
                           );
   U3667 : NAND2_X1 port map( A1 => n1744, A2 => n15004, ZN => n14746);
   U3668 : NAND2_X1 port map( A1 => n23369, A2 => n23368, ZN => n24316);
   U3669 : NAND2_X1 port map( A1 => n2508, A2 => n720, ZN => n18667);
   U3670 : NAND3_X1 port map( A1 => n1523, A2 => n18234, A3 => n1524, ZN => 
                           n720);
   U3671 : OR2_X1 port map( A1 => n5817, A2 => n21089, ZN => n20186);
   U3672 : NAND3_X1 port map( A1 => n4355, A2 => n2064, A3 => n4354, ZN => 
                           n4353);
   U3674 : OR3_X1 port map( A1 => n24140, A2 => n25009, A3 => n24139, ZN => 
                           n2153);
   U3675 : NAND2_X1 port map( A1 => n3207, A2 => n721, ZN => n19192);
   U3676 : OAI21_X1 port map( B1 => n18377, B2 => n18378, A => n3283, ZN => 
                           n721);
   U3677 : OAI21_X1 port map( B1 => n11460, B2 => n11459, A => n390, ZN => n722
                           );
   U3678 : NAND2_X1 port map( A1 => n6403, A2 => n18327, ZN => n3757);
   U3679 : NAND3_X1 port map( A1 => n836, A2 => n19762, A3 => n20063, ZN => 
                           n1699);
   U3680 : NAND2_X1 port map( A1 => n18765, A2 => n19761, ZN => n836);
   U3683 : NAND2_X1 port map( A1 => n15072, A2 => n15071, ZN => n14641);
   U3684 : NAND2_X1 port map( A1 => n20553, A2 => n20406, ZN => n20407);
   U3686 : NAND2_X1 port map( A1 => n22391, A2 => n23567, ZN => n724);
   U3688 : INV_X1 port map( A => n23567, ZN => n726);
   U3689 : NAND3_X2 port map( A1 => n728, A2 => n727, A3 => n4300, ZN => n15389
                           );
   U3690 : NAND2_X1 port map( A1 => n3851, A2 => n14432, ZN => n728);
   U3691 : INV_X1 port map( A => n7906, ZN => n944);
   U3692 : XNOR2_X1 port map( A => n729, B => n25361, ZN => Ciphertext(10));
   U3693 : OAI211_X1 port map( C1 => n6806, C2 => n29387, A => n3623, B => 
                           n5359, ZN => n729);
   U3694 : INV_X1 port map( A => n17844, ZN => n17607);
   U3695 : NAND2_X1 port map( A1 => n18242, A2 => n17969, ZN => n17844);
   U3696 : NAND3_X1 port map( A1 => n19837, A2 => n19750, A3 => n29143, ZN => 
                           n5100);
   U3697 : NOR2_X1 port map( A1 => n14000, A2 => n14036, ZN => n1019);
   U3698 : INV_X1 port map( A => n22977, ZN => n23252);
   U3700 : AOI21_X1 port map( B1 => n26990, B2 => n28521, A => n29622, ZN => 
                           n26994);
   U3702 : NOR2_X1 port map( A1 => n780, A2 => n779, ZN => n778);
   U3703 : NOR2_X1 port map( A1 => n19345, A2 => n19890, ZN => n19369);
   U3704 : NAND2_X1 port map( A1 => n14370, A2 => n731, ZN => n5796);
   U3705 : AOI21_X1 port map( B1 => n7735, B2 => n7736, A => n7734, ZN => n732)
                           ;
   U3706 : INV_X1 port map( A => n893, ZN => n14832);
   U3707 : NAND2_X1 port map( A1 => n733, A2 => n564, ZN => n893);
   U3708 : NAND2_X1 port map( A1 => n14092, A2 => n14093, ZN => n733);
   U3710 : NAND2_X1 port map( A1 => n12928, A2 => n561, ZN => n734);
   U3711 : NAND2_X1 port map( A1 => n12927, A2 => n14083, ZN => n735);
   U3712 : AND2_X2 port map( A1 => n737, A2 => n736, ZN => n22671);
   U3713 : NAND2_X1 port map( A1 => n19460, A2 => n21717, ZN => n736);
   U3714 : NAND2_X1 port map( A1 => n738, A2 => n19461, ZN => n737);
   U3715 : NAND2_X1 port map( A1 => n19419, A2 => n19418, ZN => n738);
   U3717 : AOI21_X1 port map( B1 => n29547, B2 => n17818, A => n18122, ZN => 
                           n739);
   U3718 : XNOR2_X2 port map( A => n19031, B => n19030, ZN => n20480);
   U3719 : NAND2_X1 port map( A1 => n740, A2 => n1779, ZN => n17360);
   U3720 : NAND2_X1 port map( A1 => n28793, A2 => n17356, ZN => n740);
   U3721 : NAND2_X1 port map( A1 => n28175, A2 => n28559, ZN => n10754);
   U3722 : XNOR2_X1 port map( A => n10078, B => n10077, ZN => n10556);
   U3724 : NAND2_X1 port map( A1 => n742, A2 => n8284, ZN => n7673);
   U3725 : NAND2_X1 port map( A1 => n742, A2 => n8280, ZN => n7669);
   U3726 : NAND2_X1 port map( A1 => n742, A2 => n8276, ZN => n8277);
   U3727 : NAND3_X1 port map( A1 => n8282, A2 => n8281, A3 => n742, ZN => n8283
                           );
   U3728 : NAND2_X1 port map( A1 => n7215, A2 => n742, ZN => n7216);
   U3730 : OAI21_X1 port map( B1 => n743, B2 => n1485, A => n12143, ZN => 
                           n12148);
   U3731 : NAND2_X1 port map( A1 => n573, A2 => n11712, ZN => n743);
   U3732 : NOR2_X1 port map( A1 => n1910, A2 => n745, ZN => n744);
   U3733 : INV_X1 port map( A => n7312, ZN => n7804);
   U3735 : NAND2_X1 port map( A1 => n7804, A2 => n7898, ZN => n746);
   U3736 : NAND2_X1 port map( A1 => n7805, A2 => n7804, ZN => n747);
   U3737 : XNOR2_X1 port map( A => n748, B => n10228, ZN => n9724);
   U3738 : XNOR2_X1 port map( A => n748, B => n1895, ZN => n9988);
   U3740 : NAND2_X1 port map( A1 => n4858, A2 => n4860, ZN => n750);
   U3741 : NAND3_X1 port map( A1 => n750, A2 => n820, A3 => n3654, ZN => n772);
   U3742 : NAND2_X1 port map( A1 => n750, A2 => n820, ZN => n1459);
   U3743 : AND2_X2 port map( A1 => n751, A2 => n753, ZN => n24369);
   U3746 : NAND2_X1 port map( A1 => n23259, A2 => n23735, ZN => n753);
   U3747 : NAND2_X1 port map( A1 => n14600, A2 => n15284, ZN => n756);
   U3748 : NAND2_X1 port map( A1 => n17665, A2 => n757, ZN => n4191);
   U3749 : INV_X1 port map( A => n7231, ZN => n758);
   U3750 : NAND2_X1 port map( A1 => n758, A2 => n7589, ZN => n3740);
   U3751 : NAND2_X1 port map( A1 => n758, A2 => n441, ZN => n5120);
   U3752 : NAND3_X1 port map( A1 => n7592, A2 => n7591, A3 => n758, ZN => n7593
                           );
   U3753 : NAND3_X1 port map( A1 => n7873, A2 => n7957, A3 => n758, ZN => n7054
                           );
   U3755 : NAND3_X1 port map( A1 => n10929, A2 => n762, A3 => n761, ZN => n763)
                           ;
   U3756 : NAND2_X1 port map( A1 => n590, A2 => n10726, ZN => n761);
   U3757 : NAND2_X1 port map( A1 => n588, A2 => n10932, ZN => n762);
   U3758 : XNOR2_X2 port map( A => n9474, B => n9473, ZN => n10726);
   U3759 : NAND2_X1 port map( A1 => n765, A2 => n763, ZN => n11878);
   U3761 : NAND2_X1 port map( A1 => n10460, A2 => n10927, ZN => n765);
   U3762 : NAND3_X1 port map( A1 => n17392, A2 => n766, A3 => n5021, ZN => 
                           n17391);
   U3763 : NAND2_X1 port map( A1 => n18248, A2 => n18709, ZN => n766);
   U3764 : NAND2_X1 port map( A1 => n5023, A2 => n18706, ZN => n17392);
   U3765 : NAND2_X1 port map( A1 => n26735, A2 => n26736, ZN => n767);
   U3766 : NAND2_X1 port map( A1 => n26734, A2 => n28532, ZN => n28100);
   U3767 : NAND3_X1 port map( A1 => n2094, A2 => n26736, A3 => n29486, ZN => 
                           n768);
   U3768 : XNOR2_X1 port map( A => n16232, B => n622, ZN => n14602);
   U3769 : XNOR2_X1 port map( A => n543, B => n16232, ZN => n15991);
   U3770 : XNOR2_X1 port map( A => n769, B => n16400, ZN => n15619);
   U3771 : NAND3_X1 port map( A1 => n4858, A2 => n4860, A3 => n771, ZN => n770)
                           ;
   U3773 : XNOR2_X1 port map( A => n1733, B => n19332, ZN => n775);
   U3774 : INV_X1 port map( A => n375, ZN => n777);
   U3776 : NAND3_X1 port map( A1 => n4349, A2 => n12235, A3 => n777, ZN => 
                           n11681);
   U3777 : NAND2_X1 port map( A1 => n17274, A2 => n6465, ZN => n781);
   U3778 : NAND2_X1 port map( A1 => n17273, A2 => n1181, ZN => n782);
   U3779 : AOI21_X1 port map( B1 => n4734, B2 => n785, A => n15462, ZN => 
                           n15468);
   U3781 : NAND2_X1 port map( A1 => n18503, A2 => n515, ZN => n17866);
   U3782 : NAND2_X1 port map( A1 => n18502, A2 => n515, ZN => n5985);
   U3783 : OAI211_X2 port map( C1 => n788, C2 => n1851, A => n787, B => n786, 
                           ZN => n12050);
   U3784 : NAND2_X1 port map( A1 => n11245, A2 => n11244, ZN => n786);
   U3785 : MUX2_X1 port map( A => n1900, B => n11240, S => n11244, Z => n788);
   U3787 : INV_X1 port map( A => n4220, ZN => n790);
   U3788 : XNOR2_X2 port map( A => n15759, B => n15758, ZN => n4220);
   U3789 : OR2_X1 port map( A1 => n14301, A2 => n13816, ZN => n794);
   U3790 : NAND2_X1 port map( A1 => n13816, A2 => n14053, ZN => n13647);
   U3791 : NAND2_X1 port map( A1 => n17520, A2 => n795, ZN => n16743);
   U3792 : NOR2_X1 port map( A1 => n17106, A2 => n29406, ZN => n795);
   U3793 : NAND2_X1 port map( A1 => n17473, A2 => n796, ZN => n3812);
   U3794 : OAI21_X1 port map( B1 => n29364, B2 => n22286, A => n21187, ZN => 
                           n797);
   U3795 : NAND2_X1 port map( A1 => n22023, A2 => n22290, ZN => n21187);
   U3797 : NAND2_X1 port map( A1 => n797, A2 => n22288, ZN => n3857);
   U3798 : NAND2_X1 port map( A1 => n800, A2 => n799, ZN => n26809);
   U3799 : NAND2_X1 port map( A1 => n27362, A2 => n27366, ZN => n800);
   U3800 : AOI21_X1 port map( B1 => n26809, B2 => n28562, A => n801, ZN => 
                           n26810);
   U3801 : NAND2_X1 port map( A1 => n27362, A2 => n29538, ZN => n802);
   U3803 : INV_X1 port map( A => n24804, ZN => n803);
   U3804 : OAI21_X2 port map( B1 => n23788, B2 => n807, A => n804, ZN => n24806
                           );
   U3805 : NAND2_X1 port map( A1 => n24027, A2 => n24263, ZN => n2807);
   U3806 : NAND2_X1 port map( A1 => n805, A2 => n23788, ZN => n804);
   U3807 : OAI21_X1 port map( B1 => n23785, B2 => n475, A => n806, ZN => n805);
   U3808 : NAND2_X1 port map( A1 => n23785, A2 => n23786, ZN => n806);
   U3809 : MUX2_X1 port map( A => n808, B => n473, S => n23036, Z => n807);
   U3810 : INV_X1 port map( A => n23783, ZN => n808);
   U3811 : OAI21_X2 port map( B1 => n23757, B2 => n23034, A => n3192, ZN => 
                           n24804);
   U3812 : NAND2_X1 port map( A1 => n20946, A2 => n28185, ZN => n2724);
   U3813 : AND2_X1 port map( A1 => n21501, A2 => n20944, ZN => n20946);
   U3814 : INV_X1 port map( A => n24341, ZN => n5571);
   U3815 : NAND2_X1 port map( A1 => n24708, A2 => n24341, ZN => n24125);
   U3818 : OR2_X1 port map( A1 => n1908, A2 => n810, ZN => n825);
   U3819 : NAND2_X1 port map( A1 => n20456, A2 => n810, ZN => n3953);
   U3820 : NAND2_X1 port map( A1 => n20636, A2 => n20635, ZN => n810);
   U3821 : NAND2_X1 port map( A1 => n29470, A2 => n24386, ZN => n813);
   U3822 : NAND3_X1 port map( A1 => n24133, A2 => n24386, A3 => n29470, ZN => 
                           n812);
   U3823 : NAND2_X1 port map( A1 => n5307, A2 => n813, ZN => n24134);
   U3824 : INV_X1 port map( A => n2874, ZN => n814);
   U3825 : NAND2_X1 port map( A1 => n18334, A2 => n817, ZN => n18331);
   U3827 : NAND2_X1 port map( A1 => n18370, A2 => n817, ZN => n4213);
   U3828 : NAND2_X1 port map( A1 => n17652, A2 => n816, ZN => n18002);
   U3829 : NAND2_X1 port map( A1 => n817, A2 => n18332, ZN => n816);
   U3831 : OAI211_X1 port map( C1 => n5728, C2 => n29470, A => n24081, B => 
                           n24135, ZN => n818);
   U3832 : NAND3_X1 port map( A1 => n616, A2 => n7017, A3 => n7692, ZN => n3637
                           );
   U3833 : XNOR2_X2 port map( A => Plaintext(83), B => Key(83), ZN => n7692);
   U3834 : XNOR2_X2 port map( A => n819, B => Key(78), ZN => n7817);
   U3835 : INV_X1 port map( A => Plaintext(78), ZN => n819);
   U3836 : NAND2_X1 port map( A1 => n4857, A2 => n23911, ZN => n820);
   U3837 : NAND2_X1 port map( A1 => n822, A2 => n382, ZN => n821);
   U3838 : NAND2_X1 port map( A1 => n383, A2 => n20476, ZN => n822);
   U3839 : NAND3_X1 port map( A1 => n5310, A2 => n28527, A3 => n823, ZN => 
                           n23407);
   U3840 : NAND2_X1 port map( A1 => n23405, A2 => n2239, ZN => n823);
   U3842 : NAND3_X1 port map( A1 => n2746, A2 => n20456, A3 => n825, ZN => 
                           n21532);
   U3843 : OAI211_X1 port map( C1 => n28102, C2 => n826, A => n28101, B => 
                           n28100, ZN => n28104);
   U3845 : NAND2_X1 port map( A1 => n14272, A2 => n14359, ZN => n827);
   U3846 : NAND2_X1 port map( A1 => n14271, A2 => n4166, ZN => n14361);
   U3849 : NAND2_X1 port map( A1 => n831, A2 => n24141, ZN => n3541);
   U3851 : NAND2_X1 port map( A1 => n24277, A2 => n831, ZN => n5094);
   U3852 : NOR2_X1 port map( A1 => n24590, A2 => n831, ZN => n23855);
   U3853 : OAI21_X1 port map( B1 => n24277, B2 => n831, A => n24592, ZN => 
                           n23856);
   U3854 : NAND2_X1 port map( A1 => n24279, A2 => n831, ZN => n5118);
   U3855 : OAI22_X1 port map( A1 => n24593, A2 => n4692, B1 => n4966, B2 => 
                           n831, ZN => n4152);
   U3857 : NAND2_X1 port map( A1 => n23854, A2 => n831, ZN => n840);
   U3858 : NAND2_X1 port map( A1 => n3251, A2 => n831, ZN => n5117);
   U3859 : NAND2_X1 port map( A1 => n832, A2 => n20522, ZN => n21334);
   U3860 : NAND2_X1 port map( A1 => n1200, A2 => n1199, ZN => n832);
   U3861 : OAI21_X1 port map( B1 => n8786, B2 => n8717, A => n8716, ZN => n8791
                           );
   U3862 : NAND2_X1 port map( A1 => n834, A2 => n8788, ZN => n8716);
   U3863 : INV_X1 port map( A => n8414, ZN => n834);
   U3864 : INV_X1 port map( A => n8414, ZN => n8720);
   U3865 : NAND2_X1 port map( A1 => n8791, A2 => n8790, ZN => n1294);
   U3867 : NAND3_X1 port map( A1 => n15009, A2 => n15372, A3 => n14863, ZN => 
                           n837);
   U3868 : OAI211_X2 port map( C1 => n14374, C2 => n13594, A => n4330, B => 
                           n13727, ZN => n14863);
   U3869 : NAND2_X1 port map( A1 => n15370, A2 => n15371, ZN => n14737);
   U3870 : OAI21_X1 port map( B1 => n24474, B2 => n24471, A => n53, ZN => n6123
                           );
   U3872 : MUX2_X1 port map( A => n23876, B => n23875, S => n6348, Z => n23877)
                           ;
   U3873 : NAND2_X1 port map( A1 => n20483, A2 => n20485, ZN => n20241);
   U3874 : XNOR2_X2 port map( A => n22708, B => n22709, ZN => n23442);
   U3875 : INV_X1 port map( A => n17565, ZN => n1166);
   U3876 : OAI22_X1 port map( A1 => n8343, A2 => n9133, B1 => n1670, B2 => n600
                           , ZN => n839);
   U3877 : INV_X1 port map( A => n20598, ZN => n20273);
   U3880 : NAND2_X1 port map( A1 => n23855, A2 => n24593, ZN => n841);
   U3881 : NAND2_X1 port map( A1 => n9136, A2 => n601, ZN => n842);
   U3882 : NAND2_X1 port map( A1 => n846, A2 => n28567, ZN => n866);
   U3884 : NAND2_X1 port map( A1 => n24019, A2 => n24541, ZN => n846);
   U3885 : XNOR2_X1 port map( A => n847, B => n26601, ZN => Ciphertext(144));
   U3886 : NAND4_X1 port map( A1 => n26600, A2 => n26598, A3 => n26597, A4 => 
                           n26599, ZN => n847);
   U3887 : NAND2_X1 port map( A1 => n5514, A2 => n15419, ZN => n3705);
   U3889 : AOI21_X2 port map( B1 => n11418, B2 => n12146, A => n848, ZN => 
                           n12595);
   U3890 : AOI21_X1 port map( B1 => n11416, B2 => n11417, A => n11645, ZN => 
                           n848);
   U3891 : INV_X1 port map( A => n1287, ZN => n23060);
   U3892 : NAND2_X1 port map( A1 => n23343, A2 => n23338, ZN => n1287);
   U3894 : NAND3_X1 port map( A1 => n14204, A2 => n2959, A3 => n14459, ZN => 
                           n12704);
   U3899 : NAND3_X1 port map( A1 => n4547, A2 => n4548, A3 => n14575, ZN => 
                           n2731);
   U3901 : OAI21_X1 port map( B1 => n16779, B2 => n17262, A => n17258, ZN => 
                           n16151);
   U3902 : OAI22_X1 port map( A1 => n18430, A2 => n850, B1 => n17814, B2 => 
                           n18148, ZN => n17817);
   U3903 : NAND2_X1 port map( A1 => n18431, A2 => n18433, ZN => n850);
   U3904 : NAND2_X1 port map( A1 => n17517, A2 => n17518, ZN => n17472);
   U3905 : NAND2_X1 port map( A1 => n23336, A2 => n851, ZN => n25761);
   U3907 : OAI21_X2 port map( B1 => n24190, B2 => n24191, A => n24189, ZN => 
                           n25440);
   U3908 : OAI22_X1 port map( A1 => n25669, A2 => n25670, B1 => n26474, B2 => 
                           n26181, ZN => n852);
   U3911 : NAND2_X1 port map( A1 => n3830, A2 => n13582, ZN => n13645);
   U3914 : AND2_X1 port map( A1 => n20351, A2 => n20783, ZN => n20931);
   U3915 : NAND2_X1 port map( A1 => n20847, A2 => n854, ZN => n5942);
   U3916 : NAND2_X1 port map( A1 => n21485, A2 => n20749, ZN => n20847);
   U3917 : OAI21_X1 port map( B1 => n28225, B2 => n406, A => n855, ZN => n23001
                           );
   U3918 : NAND2_X1 port map( A1 => n28225, A2 => n379, ZN => n855);
   U3919 : NOR3_X1 port map( A1 => n24617, A2 => n28550, A3 => n1631, ZN => 
                           n24620);
   U3922 : XNOR2_X1 port map( A => n10029, B => n9934, ZN => n10287);
   U3923 : OR2_X1 port map( A1 => n11594, A2 => n11932, ZN => n11597);
   U3924 : AOI22_X1 port map( A1 => n18508, A2 => n18271, B1 => n18273, B2 => 
                           n29057, ZN => n856);
   U3926 : NAND2_X1 port map( A1 => n8963, A2 => n605, ZN => n2289);
   U3927 : XNOR2_X1 port map( A => n858, B => n10391, ZN => n9357);
   U3928 : INV_X1 port map( A => n9447, ZN => n858);
   U3929 : NAND2_X1 port map( A1 => n18297, A2 => n28745, ZN => n2459);
   U3930 : AND2_X2 port map( A1 => n7360, A2 => n7361, ZN => n9148);
   U3931 : XNOR2_X1 port map( A => n859, B => n8940, ZN => n10472);
   U3932 : XNOR2_X1 port map( A => n8952, B => n9523, ZN => n859);
   U3934 : OR2_X1 port map( A1 => n20972, A2 => n20966, ZN => n21215);
   U3935 : NAND2_X1 port map( A1 => n10853, A2 => n10851, ZN => n11162);
   U3936 : NAND2_X1 port map( A1 => n861, A2 => n18248, ZN => n1784);
   U3937 : NAND2_X1 port map( A1 => n863, A2 => n862, ZN => n861);
   U3938 : NAND2_X1 port map( A1 => n18707, A2 => n17353, ZN => n862);
   U3940 : OR2_X1 port map( A1 => n13888, A2 => n14317, ZN => n12585);
   U3941 : INV_X1 port map( A => n15223, ZN => n15227);
   U3942 : XNOR2_X1 port map( A => n16871, B => n16870, ZN => n20405);
   U3944 : OAI22_X1 port map( A1 => n20548, A2 => n19857, B1 => n5982, B2 => 
                           n6315, ZN => n21696);
   U3945 : XNOR2_X1 port map( A => n864, B => n10285, ZN => n5562);
   U3946 : XNOR2_X1 port map( A => n10284, B => n10283, ZN => n864);
   U3947 : OAI21_X1 port map( B1 => n1736, B2 => n1735, A => n11077, ZN => 
                           n1734);
   U3949 : OR2_X1 port map( A1 => n9140, A2 => n598, ZN => n1127);
   U3950 : NAND2_X1 port map( A1 => n27191, A2 => n27190, ZN => n26290);
   U3951 : NOR2_X1 port map( A1 => n23254, A2 => n867, ZN => n23255);
   U3952 : NAND2_X1 port map( A1 => n27645, A2 => n868, ZN => n26672);
   U3953 : NAND2_X1 port map( A1 => n27641, A2 => n27639, ZN => n868);
   U3954 : NAND2_X1 port map( A1 => n20001, A2 => n869, ZN => n6137);
   U3955 : XNOR2_X1 port map( A => n16377, B => n3856, ZN => n16121);
   U3956 : OR2_X1 port map( A1 => n29585, A2 => n27191, ZN => n26138);
   U3957 : NAND2_X1 port map( A1 => n18231, A2 => n18398, ZN => n18397);
   U3958 : OAI21_X1 port map( B1 => n12363, B2 => n12361, A => n870, ZN => 
                           n10899);
   U3961 : NOR2_X1 port map( A1 => n15036, A2 => n15290, ZN => n4955);
   U3962 : OAI211_X1 port map( C1 => n21692, C2 => n21242, A => n6311, B => 
                           n21348, ZN => n6312);
   U3963 : NAND2_X1 port map( A1 => n1165, A2 => n1167, ZN => n871);
   U3964 : INV_X1 port map( A => n21645, ZN => n21042);
   U3965 : NAND2_X1 port map( A1 => n10110, A2 => n10704, ZN => n10708);
   U3967 : NAND2_X1 port map( A1 => n1673, A2 => n1674, ZN => n872);
   U3969 : NAND2_X2 port map( A1 => n5970, A2 => n5969, ZN => n15900);
   U3970 : XNOR2_X1 port map( A => n22357, B => n22600, ZN => n22361);
   U3971 : NAND2_X1 port map( A1 => n5349, A2 => n24435, ZN => n873);
   U3972 : NAND2_X1 port map( A1 => n6293, A2 => n14605, ZN => n874);
   U3973 : OAI21_X1 port map( B1 => n18707, B2 => n876, A => n875, ZN => n18250
                           );
   U3974 : NAND2_X1 port map( A1 => n18707, A2 => n18404, ZN => n875);
   U3975 : NAND2_X1 port map( A1 => n2690, A2 => n11022, ZN => n11316);
   U3976 : INV_X1 port map( A => n21511, ZN => n20463);
   U3977 : NAND2_X1 port map( A1 => n21532, A2 => n21534, ZN => n21511);
   U3978 : XOR2_X1 port map( A => n16482, B => n16478, Z => n1094);
   U3979 : NAND3_X1 port map( A1 => n877, A2 => n3342, A3 => n3343, ZN => 
                           n18305);
   U3980 : NAND2_X1 port map( A1 => n14694, A2 => n29600, ZN => n877);
   U3982 : OAI21_X1 port map( B1 => n23556, B2 => n23636, A => n5143, ZN => 
                           n878);
   U3983 : MUX2_X1 port map( A => n24068, B => n24067, S => n24677, Z => n24069
                           );
   U3984 : AOI22_X1 port map( A1 => n26483, A2 => n1623, B1 => n29501, B2 => 
                           n26484, ZN => n26487);
   U3985 : INV_X1 port map( A => n22514, ZN => n21182);
   U3986 : INV_X1 port map( A => n21549, ZN => n1621);
   U3987 : INV_X1 port map( A => n18333, ZN => n1650);
   U3988 : NAND2_X1 port map( A1 => n883, A2 => n8569, ZN => n7387);
   U3989 : OAI21_X1 port map( B1 => n9150, B2 => n8929, A => n9374, ZN => n883)
                           ;
   U3991 : OAI211_X1 port map( C1 => n28181, C2 => n23741, A => n886, B => n885
                           , ZN => n884);
   U3992 : NAND2_X1 port map( A1 => n23741, A2 => n482, ZN => n886);
   U3995 : NAND2_X1 port map( A1 => n6832, A2 => n12513, ZN => n3382);
   U3996 : NOR2_X2 port map( A1 => n12715, A2 => n888, ZN => n15420);
   U3997 : NAND2_X1 port map( A1 => n25617, A2 => n27395, ZN => n25621);
   U3998 : NAND2_X1 port map( A1 => n17164, A2 => n28775, ZN => n4293);
   U3999 : NAND2_X1 port map( A1 => n890, A2 => n889, ZN => n7724);
   U4000 : NAND2_X1 port map( A1 => n7721, A2 => n7336, ZN => n890);
   U4003 : NAND2_X1 port map( A1 => n18382, A2 => n17881, ZN => n18350);
   U4004 : NAND2_X1 port map( A1 => n903, A2 => n905, ZN => n23754);
   U4005 : NAND2_X1 port map( A1 => n12510, A2 => n11990, ZN => n6833);
   U4006 : NAND2_X1 port map( A1 => n8740, A2 => n9073, ZN => n9072);
   U4008 : AOI21_X1 port map( B1 => n23796, B2 => n23321, A => n23039, ZN => 
                           n24336);
   U4009 : XNOR2_X1 port map( A => n892, B => n19356, ZN => n19358);
   U4010 : XNOR2_X1 port map( A => n19355, B => n19354, ZN => n892);
   U4011 : AND2_X1 port map( A1 => n4478, A2 => n17361, ZN => n17047);
   U4012 : NAND2_X1 port map( A1 => n12206, A2 => n4037, ZN => n4446);
   U4013 : AOI22_X1 port map( A1 => n11851, A2 => n11853, B1 => n11852, B2 => 
                           n11921, ZN => n11854);
   U4014 : OR2_X1 port map( A1 => n14665, A2 => n14666, ZN => n1053);
   U4015 : NAND3_X1 port map( A1 => n5529, A2 => n20230, A3 => n4557, ZN => 
                           n5528);
   U4018 : NAND2_X1 port map( A1 => n1354, A2 => n29112, ZN => n7088);
   U4019 : NAND3_X1 port map( A1 => n24996, A2 => n24995, A3 => n894, ZN => 
                           n24998);
   U4021 : NAND2_X1 port map( A1 => n897, A2 => n895, ZN => n10968);
   U4022 : NAND2_X1 port map( A1 => n10687, A2 => n10961, ZN => n895);
   U4023 : INV_X1 port map( A => n10959, ZN => n896);
   U4025 : NOR2_X1 port map( A1 => n11070, A2 => n262, ZN => n898);
   U4026 : NAND2_X1 port map( A1 => n20614, A2 => n899, ZN => n1082);
   U4027 : AOI22_X1 port map( A1 => n28036, A2 => n28037, B1 => n28034, B2 => 
                           n28035, ZN => n28042);
   U4028 : NAND2_X1 port map( A1 => n26661, A2 => n26662, ZN => n28036);
   U4029 : AND3_X2 port map( A1 => n23092, A2 => n23091, A3 => n3990, ZN => 
                           n24380);
   U4030 : NAND3_X1 port map( A1 => n9436, A2 => n9210, A3 => n8996, ZN => 
                           n7680);
   U4031 : NAND2_X1 port map( A1 => n7662, A2 => n8271, ZN => n901);
   U4034 : NAND2_X1 port map( A1 => n23744, A2 => n24514, ZN => n905);
   U4035 : OR2_X1 port map( A1 => n20479, A2 => n20480, ZN => n4556);
   U4036 : NAND2_X1 port map( A1 => n20298, A2 => n5933, ZN => n20301);
   U4038 : NAND2_X1 port map( A1 => n23848, A2 => n23845, ZN => n908);
   U4039 : OAI21_X1 port map( B1 => n909, B2 => n29227, A => n21706, ZN => 
                           n21711);
   U4040 : AOI21_X1 port map( B1 => n21702, B2 => n21705, A => n496, ZN => n909
                           );
   U4041 : NAND3_X1 port map( A1 => n23911, A2 => n23389, A3 => n24077, ZN => 
                           n23410);
   U4042 : OR2_X1 port map( A1 => n21443, A2 => n21656, ZN => n1109);
   U4043 : NAND2_X1 port map( A1 => n14284, A2 => n14283, ZN => n14290);
   U4044 : NAND2_X1 port map( A1 => n7909, A2 => n8287, ZN => n7474);
   U4046 : OAI211_X1 port map( C1 => n23415, C2 => n23417, A => n2435, B => 
                           n23419, ZN => n910);
   U4048 : OAI22_X1 port map( A1 => n23807, A2 => n29102, B1 => n28594, B2 => 
                           n28653, ZN => n22745);
   U4050 : NAND2_X1 port map( A1 => n14079, A2 => n13744, ZN => n912);
   U4052 : NAND2_X1 port map( A1 => n914, A2 => n17846, ZN => n913);
   U4053 : NAND2_X1 port map( A1 => n917, A2 => n18144, ZN => n916);
   U4054 : NAND2_X1 port map( A1 => n918, A2 => n18143, ZN => n917);
   U4055 : NAND2_X1 port map( A1 => n2811, A2 => n18137, ZN => n918);
   U4057 : OAI211_X1 port map( C1 => n17526, C2 => n17157, A => n920, B => 
                           n17181, ZN => n5919);
   U4058 : NAND2_X1 port map( A1 => n17157, A2 => n17528, ZN => n920);
   U4059 : NAND2_X1 port map( A1 => n27865, A2 => n27877, ZN => n27866);
   U4060 : NAND2_X1 port map( A1 => n25720, A2 => n922, ZN => n921);
   U4061 : NAND3_X1 port map( A1 => n924, A2 => n3332, A3 => n27069, ZN => n923
                           );
   U4062 : NAND2_X1 port map( A1 => n29076, A2 => n29520, ZN => n924);
   U4063 : NAND2_X1 port map( A1 => n28545, A2 => n29520, ZN => n925);
   U4064 : INV_X1 port map( A => n14871, ZN => n17400);
   U4065 : INV_X1 port map( A => n16825, ZN => n926);
   U4066 : XNOR2_X1 port map( A => n928, B => n927, ZN => Ciphertext(87));
   U4067 : NAND3_X1 port map( A1 => n936, A2 => n932, A3 => n929, ZN => n928);
   U4068 : NAND2_X1 port map( A1 => n931, A2 => n930, ZN => n929);
   U4069 : INV_X1 port map( A => n27591, ZN => n27585);
   U4070 : NAND2_X1 port map( A1 => n934, A2 => n933, ZN => n932);
   U4071 : NOR2_X1 port map( A1 => n27589, A2 => n935, ZN => n934);
   U4072 : AND2_X1 port map( A1 => n27591, A2 => n27590, ZN => n935);
   U4073 : NAND2_X1 port map( A1 => n27592, A2 => n1901, ZN => n936);
   U4074 : AND2_X1 port map( A1 => n2502, A2 => n937, ZN => n938);
   U4075 : NAND2_X1 port map( A1 => n8433, A2 => n9029, ZN => n937);
   U4076 : INV_X1 port map( A => n17159, ZN => n940);
   U4077 : NAND2_X1 port map( A1 => n940, A2 => n424, ZN => n939);
   U4078 : NAND2_X1 port map( A1 => n17384, A2 => n18069, ZN => n941);
   U4079 : XNOR2_X1 port map( A => n942, B => n18145, ZN => n18167);
   U4080 : XNOR2_X1 port map( A => n19469, B => n942, ZN => n19470);
   U4081 : XNOR2_X1 port map( A => n942, B => n19017, ZN => n19018);
   U4082 : XNOR2_X1 port map( A => n19370, B => n18134, ZN => n942);
   U4083 : NAND2_X1 port map( A1 => n2141, A2 => n23258, ZN => n943);
   U4084 : NAND4_X2 port map( A1 => n8636, A2 => n8638, A3 => n8637, A4 => n944
                           , ZN => n10160);
   U4085 : NAND2_X1 port map( A1 => n945, A2 => n2325, ZN => n947);
   U4087 : NAND3_X1 port map( A1 => n24587, A2 => n6055, A3 => n635, ZN => n946
                           );
   U4088 : XNOR2_X1 port map( A => n945, B => n3232, ZN => n24925);
   U4089 : XNOR2_X1 port map( A => n945, B => n3516, ZN => n25168);
   U4090 : XNOR2_X1 port map( A => n945, B => n3114, ZN => n25576);
   U4091 : XNOR2_X1 port map( A => n945, B => n3635, ZN => n25938);
   U4092 : XNOR2_X1 port map( A => n25785, B => n945, ZN => n25467);
   U4093 : NAND2_X1 port map( A1 => n951, A2 => n949, ZN => n25362);
   U4095 : XNOR2_X2 port map( A => n24574, B => n24573, ZN => n26560);
   U4096 : NAND2_X1 port map( A1 => n954, A2 => n953, ZN => n15301);
   U4097 : NAND2_X1 port map( A1 => n14172, A2 => n957, ZN => n953);
   U4098 : NAND3_X1 port map( A1 => n14244, A2 => n957, A3 => n28172, ZN => 
                           n954);
   U4099 : OAI21_X2 port map( B1 => n956, B2 => n14172, A => n957, ZN => n15436
                           );
   U4100 : NAND2_X1 port map( A1 => n6573, A2 => n958, ZN => n957);
   U4101 : OR2_X1 port map( A1 => n13943, A2 => n15194, ZN => n958);
   U4102 : AND2_X1 port map( A1 => n14239, A2 => n14240, ZN => n6573);
   U4103 : NAND2_X1 port map( A1 => n23618, A2 => n960, ZN => n23626);
   U4104 : NOR2_X1 port map( A1 => n23566, A2 => n960, ZN => n22986);
   U4105 : NAND3_X1 port map( A1 => n23566, A2 => n23621, A3 => n960, ZN => 
                           n23272);
   U4106 : OAI21_X1 port map( B1 => n23570, B2 => n23571, A => n960, ZN => 
                           n23572);
   U4107 : OAI211_X1 port map( C1 => n6646, C2 => n962, A => n1947, B => n961, 
                           ZN => n13222);
   U4108 : NAND3_X1 port map( A1 => n581, A2 => n3585, A3 => n10563, ZN => 
                           n10511);
   U4109 : NAND2_X1 port map( A1 => n20299, A2 => n20443, ZN => n19924);
   U4111 : NAND2_X1 port map( A1 => n10237, A2 => n3116, ZN => n963);
   U4112 : XNOR2_X1 port map( A => n25933, B => n26100, ZN => n25112);
   U4113 : NAND3_X1 port map( A1 => n965, A2 => n966, A3 => n24486, ZN => n964)
                           ;
   U4114 : OR2_X1 port map( A1 => n24481, A2 => n24480, ZN => n965);
   U4115 : NAND2_X1 port map( A1 => n968, A2 => n6539, ZN => n6538);
   U4116 : NOR2_X1 port map( A1 => n17015, A2 => n968, ZN => n17021);
   U4117 : NAND2_X1 port map( A1 => n10808, A2 => n28627, ZN => n969);
   U4119 : NAND2_X1 port map( A1 => n261, A2 => n8427, ZN => n8354);
   U4120 : INV_X1 port map( A => n8352, ZN => n970);
   U4122 : NAND2_X1 port map( A1 => n547, A2 => n15185, ZN => n1570);
   U4123 : OAI21_X1 port map( B1 => n14784, B2 => n972, A => n15182, ZN => 
                           n14532);
   U4124 : NAND2_X1 port map( A1 => n15186, A2 => n972, ZN => n1571);
   U4125 : OAI211_X1 port map( C1 => n15190, C2 => n15183, A => n15186, B => 
                           n972, ZN => n14800);
   U4126 : NAND2_X1 port map( A1 => n13801, A2 => n13802, ZN => n973);
   U4127 : NAND2_X1 port map( A1 => n13800, A2 => n14312, ZN => n974);
   U4128 : NAND2_X1 port map( A1 => n18071, A2 => n18070, ZN => n975);
   U4129 : NOR2_X1 port map( A1 => n29496, A2 => n2032, ZN => n18075);
   U4130 : NOR2_X2 port map( A1 => n975, A2 => n5814, ZN => n18510);
   U4132 : NAND2_X1 port map( A1 => n626, A2 => n977, ZN => n7436);
   U4133 : INV_X1 port map( A => n8217, ZN => n977);
   U4134 : NAND2_X1 port map( A1 => n14934, A2 => n14935, ZN => n6286);
   U4138 : NAND2_X1 port map( A1 => n24071, A2 => n24316, ZN => n980);
   U4141 : MUX2_X1 port map( A => n11549, B => n11922, S => n11852, Z => n10095
                           );
   U4142 : AND2_X2 port map( A1 => n6151, A2 => n10004, ZN => n11852);
   U4143 : NAND2_X1 port map( A1 => n3580, A2 => n427, ZN => n981);
   U4148 : NAND2_X1 port map( A1 => n23885, A2 => n24437, ZN => n5349);
   U4149 : NAND2_X1 port map( A1 => n24436, A2 => n24347, ZN => n23885);
   U4150 : NOR2_X1 port map( A1 => n23154, A2 => n23482, ZN => n984);
   U4153 : NAND2_X1 port map( A1 => n987, A2 => n15115, ZN => n986);
   U4154 : NAND2_X1 port map( A1 => n14740, A2 => n15117, ZN => n987);
   U4155 : NAND2_X1 port map( A1 => n1003, A2 => n544, ZN => n988);
   U4156 : NAND2_X1 port map( A1 => n990, A2 => n989, ZN => n11536);
   U4157 : NAND2_X1 port map( A1 => n10540, A2 => n10760, ZN => n990);
   U4158 : NAND2_X1 port map( A1 => n13586, A2 => n13602, ZN => n13592);
   U4159 : NAND2_X1 port map( A1 => n2248, A2 => n8350, ZN => n2247);
   U4161 : AOI21_X1 port map( B1 => n19880, B2 => n19881, A => n20028, ZN => 
                           n19885);
   U4164 : NAND3_X2 port map( A1 => n3070, A2 => n3069, A3 => n3068, ZN => 
                           n19440);
   U4165 : NAND2_X1 port map( A1 => n14076, A2 => n14253, ZN => n14096);
   U4166 : NAND2_X1 port map( A1 => n991, A2 => n2824, ZN => n2821);
   U4167 : NAND2_X1 port map( A1 => n2822, A2 => n28567, ZN => n991);
   U4168 : INV_X1 port map( A => n1650, ZN => n1087);
   U4169 : OAI211_X2 port map( C1 => n493, C2 => n21391, A => n21390, B => n992
                           , ZN => n22326);
   U4170 : NAND2_X1 port map( A1 => n21388, A2 => n21387, ZN => n992);
   U4172 : NOR2_X2 port map( A1 => n994, A2 => n993, ZN => n19123);
   U4175 : XNOR2_X1 port map( A => n22922, B => n272, ZN => n21996);
   U4177 : NAND2_X1 port map( A1 => n997, A2 => n996, ZN => n8058);
   U4178 : NAND2_X1 port map( A1 => n7806, A2 => n7805, ZN => n996);
   U4179 : INV_X1 port map( A => n20441, ZN => n1081);
   U4180 : NAND2_X1 port map( A1 => n11183, A2 => n11323, ZN => n11186);
   U4181 : NAND2_X1 port map( A1 => n8605, A2 => n9081, ZN => n8850);
   U4182 : NAND2_X1 port map( A1 => n4072, A2 => n998, ZN => n15342);
   U4184 : INV_X1 port map( A => n24240, ZN => n25794);
   U4185 : NAND2_X1 port map( A1 => n999, A2 => n23186, ZN => n24240);
   U4186 : NAND2_X1 port map( A1 => n23184, A2 => n23566, ZN => n999);
   U4187 : NAND2_X1 port map( A1 => n17221, A2 => n29142, ZN => n15847);
   U4188 : NAND2_X1 port map( A1 => n5179, A2 => n5561, ZN => n5178);
   U4189 : NOR2_X1 port map( A1 => n12260, A2 => n11622, ZN => n11581);
   U4191 : NAND2_X1 port map( A1 => n1002, A2 => n1001, ZN => n1000);
   U4192 : NAND2_X1 port map( A1 => n15113, A2 => n15119, ZN => n1003);
   U4193 : NAND2_X1 port map( A1 => n15114, A2 => n1005, ZN => n1004);
   U4194 : NAND2_X1 port map( A1 => n15118, A2 => n15117, ZN => n1006);
   U4195 : XNOR2_X1 port map( A => n9352, B => n10335, ZN => n9242);
   U4196 : NOR2_X1 port map( A1 => n3155, A2 => n258, ZN => n1007);
   U4197 : NAND3_X1 port map( A1 => n17173, A2 => n29635, A3 => n16874, ZN => 
                           n1799);
   U4199 : NAND2_X1 port map( A1 => n1009, A2 => n17858, ZN => n3540);
   U4200 : NAND3_X1 port map( A1 => n17718, A2 => n5329, A3 => n17719, ZN => 
                           n1009);
   U4203 : AOI22_X2 port map( A1 => n7249, A2 => n8135, B1 => n1010, B2 => n615
                           , ZN => n8553);
   U4205 : OAI211_X1 port map( C1 => n4998, C2 => n27926, A => n27950, B => 
                           n1011, ZN => n4999);
   U4206 : INV_X1 port map( A => n29082, ZN => n6615);
   U4209 : NAND2_X1 port map( A1 => n3833, A2 => n3834, ZN => n3832);
   U4210 : AND2_X1 port map( A1 => n20483, A2 => n20484, ZN => n19791);
   U4211 : NAND2_X1 port map( A1 => n4058, A2 => n4059, ZN => n18265);
   U4212 : INV_X1 port map( A => n18263, ZN => n18262);
   U4215 : AND2_X1 port map( A1 => n1166, A2 => n29098, ZN => n1723);
   U4216 : INV_X1 port map( A => n17439, ZN => n16962);
   U4217 : INV_X1 port map( A => n11780, ZN => n11421);
   U4218 : INV_X1 port map( A => n18042, ZN => n16862);
   U4219 : XNOR2_X1 port map( A => n10196, B => n10197, ZN => n11064);
   U4220 : INV_X1 port map( A => n21705, ZN => n21373);
   U4222 : XNOR2_X1 port map( A => n15742, B => n15743, ZN => n16837);
   U4224 : AOI21_X1 port map( B1 => n1013, B2 => n1012, A => n24405, ZN => 
                           n23910);
   U4225 : NAND2_X1 port map( A1 => n3797, A2 => n24085, ZN => n1012);
   U4226 : NAND2_X1 port map( A1 => n6265, A2 => n24404, ZN => n1013);
   U4227 : XNOR2_X2 port map( A => n1015, B => n19281, ZN => n19985);
   U4228 : XNOR2_X1 port map( A => n3659, B => n18876, ZN => n1015);
   U4230 : NAND2_X1 port map( A1 => n20020, A2 => n19795, ZN => n20518);
   U4231 : NAND2_X1 port map( A1 => n6465, A2 => n17275, ZN => n1017);
   U4232 : NAND2_X1 port map( A1 => n16844, A2 => n539, ZN => n1018);
   U4234 : OAI21_X1 port map( B1 => n8579, B2 => n606, A => n604, ZN => n8771);
   U4235 : NAND3_X1 port map( A1 => n7585, A2 => n7584, A3 => n7884, ZN => 
                           n7304);
   U4236 : NAND2_X1 port map( A1 => n1930, A2 => n21471, ZN => n21475);
   U4237 : NAND2_X1 port map( A1 => n1021, A2 => n5625, ZN => n5624);
   U4239 : OR2_X1 port map( A1 => n28478, A2 => n13646, ZN => n5341);
   U4240 : OAI211_X1 port map( C1 => n18153, C2 => n18154, A => n18158, B => 
                           n1022, ZN => n1232);
   U4241 : NAND2_X1 port map( A1 => n17825, A2 => n18154, ZN => n1022);
   U4242 : NAND2_X1 port map( A1 => n1309, A2 => n1023, ZN => n15011);
   U4243 : INV_X1 port map( A => n1024, ZN => n1023);
   U4244 : AOI21_X1 port map( B1 => n14614, B2 => n14615, A => n632, ZN => 
                           n1024);
   U4245 : NAND2_X1 port map( A1 => n15302, A2 => n15436, ZN => n13944);
   U4246 : NAND2_X1 port map( A1 => n1026, A2 => n1025, ZN => n17810);
   U4248 : XNOR2_X2 port map( A => n7030, B => Key(63), ZN => n7266);
   U4249 : NAND2_X1 port map( A1 => n1028, A2 => n7915, ZN => n1797);
   U4250 : OAI21_X1 port map( B1 => n29568, B2 => n7909, A => n7474, ZN => 
                           n1028);
   U4251 : NAND3_X1 port map( A1 => n15131, A2 => n14999, A3 => n15132, ZN => 
                           n5866);
   U4252 : NAND2_X1 port map( A1 => n14998, A2 => n15123, ZN => n15131);
   U4253 : NAND2_X1 port map( A1 => n26380, A2 => n1076, ZN => n1029);
   U4254 : INV_X1 port map( A => n26425, ZN => n1030);
   U4256 : NAND2_X1 port map( A1 => n29321, A2 => n7846, ZN => n6299);
   U4258 : NAND2_X1 port map( A1 => n7522, A2 => n7268, ZN => n1033);
   U4261 : OAI211_X1 port map( C1 => n3440, C2 => n623, A => n1730, B => n1729,
                           ZN => n19433);
   U4262 : NAND3_X1 port map( A1 => n2318, A2 => n2838, A3 => n2317, ZN => 
                           n18867);
   U4263 : NAND2_X1 port map( A1 => n1035, A2 => n20136, ZN => n20138);
   U4264 : NAND2_X1 port map( A1 => n19896, A2 => n2152, ZN => n1035);
   U4267 : AND2_X2 port map( A1 => n12624, A2 => n12625, ZN => n3315);
   U4269 : NAND2_X1 port map( A1 => n3737, A2 => n3739, ZN => n18466);
   U4270 : OAI21_X1 port map( B1 => n28015, B2 => n445, A => n1037, ZN => 
                           n28012);
   U4271 : NAND2_X1 port map( A1 => n28015, A2 => n28017, ZN => n1037);
   U4273 : NOR2_X1 port map( A1 => n28104, A2 => n28103, ZN => n1690);
   U4275 : INV_X1 port map( A => n4617, ZN => n12037);
   U4276 : XNOR2_X1 port map( A => n10045, B => n10411, ZN => n1572);
   U4277 : AOI21_X2 port map( B1 => n15354, B2 => n15353, A => n15352, ZN => 
                           n16279);
   U4278 : XNOR2_X1 port map( A => n9930, B => n3073, ZN => n9743);
   U4280 : NAND3_X1 port map( A1 => n15434, A2 => n15431, A3 => n15432, ZN => 
                           n14022);
   U4284 : NAND2_X1 port map( A1 => n18136, A2 => n17846, ZN => n17849);
   U4287 : OR2_X1 port map( A1 => n18311, A2 => n17920, ZN => n4629);
   U4288 : NAND3_X1 port map( A1 => n24412, A2 => n24714, A3 => n28524, ZN => 
                           n24411);
   U4290 : NOR2_X1 port map( A1 => n21653, A2 => n6275, ZN => n20244);
   U4291 : NAND2_X1 port map( A1 => n17972, A2 => n17973, ZN => n19409);
   U4292 : NAND3_X1 port map( A1 => n20607, A2 => n1081, A3 => n20611, ZN => 
                           n1040);
   U4294 : AOI21_X1 port map( B1 => n5303, B2 => n20494, A => n6834, ZN => 
                           n1041);
   U4295 : NAND2_X1 port map( A1 => n2514, A2 => n2516, ZN => n1042);
   U4296 : INV_X1 port map( A => n20938, ZN => n21309);
   U4297 : NAND2_X1 port map( A1 => n1043, A2 => n20938, ZN => n1315);
   U4298 : NAND3_X1 port map( A1 => n20308, A2 => n20307, A3 => n20309, ZN => 
                           n20938);
   U4299 : INV_X1 port map( A => n21306, ZN => n1043);
   U4301 : OAI21_X1 port map( B1 => n20055, B2 => n1044, A => n2555, ZN => 
                           n20058);
   U4302 : AOI21_X1 port map( B1 => n20054, B2 => n20172, A => n6114, ZN => 
                           n1044);
   U4303 : NAND2_X1 port map( A1 => n20917, A2 => n21287, ZN => n20918);
   U4304 : NOR2_X1 port map( A1 => n20986, A2 => n21288, ZN => n20917);
   U4306 : AND2_X1 port map( A1 => n1938, A2 => n7675, ZN => n7678);
   U4309 : INV_X1 port map( A => n18421, ZN => n4805);
   U4310 : OAI22_X1 port map( A1 => n1456, A2 => n525, B1 => n17762, B2 => 
                           n17943, ZN => n1455);
   U4313 : NAND2_X1 port map( A1 => n13803, A2 => n14292, ZN => n13804);
   U4316 : NAND3_X1 port map( A1 => n5129, A2 => n5594, A3 => n8579, ZN => 
                           n1045);
   U4318 : NAND2_X1 port map( A1 => n11714, A2 => n11650, ZN => n1048);
   U4319 : INV_X1 port map( A => n16815, ZN => n1091);
   U4320 : OAI22_X1 port map( A1 => n21893, A2 => n28444, B1 => n23689, B2 => 
                           n23537, ZN => n23690);
   U4321 : NOR2_X2 port map( A1 => n23528, A2 => n1049, ZN => n24765);
   U4322 : NOR3_X1 port map( A1 => n23527, A2 => n23662, A3 => n23526, ZN => 
                           n1049);
   U4324 : NAND2_X1 port map( A1 => n3936, A2 => n21562, ZN => n1050);
   U4325 : NAND2_X1 port map( A1 => n15434, A2 => n15030, ZN => n5407);
   U4326 : NAND2_X1 port map( A1 => n27340, A2 => n29052, ZN => n27348);
   U4327 : NAND2_X1 port map( A1 => n1052, A2 => n1051, ZN => n1256);
   U4328 : NAND2_X1 port map( A1 => n1622, A2 => n29579, ZN => n1051);
   U4329 : NAND2_X1 port map( A1 => n26726, A2 => n26727, ZN => n1052);
   U4331 : NAND2_X1 port map( A1 => n23600, A2 => n23467, ZN => n23601);
   U4332 : NAND2_X1 port map( A1 => n2656, A2 => n6526, ZN => n17990);
   U4333 : NAND2_X1 port map( A1 => n14664, A2 => n1053, ZN => n15304);
   U4334 : XNOR2_X1 port map( A => n19271, B => n1054, ZN => n20272);
   U4336 : OR2_X1 port map( A1 => n8265, A2 => n341, ZN => n2472);
   U4338 : OAI21_X1 port map( B1 => n22878, B2 => n4385, A => n22743, ZN => 
                           n22744);
   U4339 : AOI21_X1 port map( B1 => n8459, B2 => n8524, A => n8680, ZN => n1056
                           );
   U4340 : XNOR2_X1 port map( A => n19315, B => n1057, ZN => n18694);
   U4341 : XNOR2_X1 port map( A => n18689, B => n18880, ZN => n1057);
   U4342 : NAND2_X1 port map( A1 => n1059, A2 => n1058, ZN => n8577);
   U4343 : NAND2_X1 port map( A1 => n8576, A2 => n29395, ZN => n1058);
   U4344 : NAND2_X1 port map( A1 => n1060, A2 => n8749, ZN => n1059);
   U4345 : NAND2_X1 port map( A1 => n9532, A2 => n9530, ZN => n1060);
   U4346 : NAND2_X1 port map( A1 => n1256, A2 => n1532, ZN => n25629);
   U4348 : NAND2_X1 port map( A1 => n2167, A2 => n12281, ZN => n1061);
   U4352 : NAND2_X1 port map( A1 => n1063, A2 => n12231, ZN => n11987);
   U4353 : NAND2_X1 port map( A1 => n9433, A2 => n11981, ZN => n1063);
   U4354 : NAND2_X1 port map( A1 => n13083, A2 => n303, ZN => n9433);
   U4356 : XOR2_X1 port map( A => n13543, B => n440, Z => n6270);
   U4358 : OR2_X1 port map( A1 => n2228, A2 => n10871, ZN => n1163);
   U4361 : NAND2_X1 port map( A1 => n18144, A2 => n526, ZN => n17845);
   U4362 : OAI211_X1 port map( C1 => n28206, C2 => n10742, A => n28876, B => 
                           n1064, ZN => n10744);
   U4364 : NAND2_X1 port map( A1 => n1066, A2 => n1065, ZN => n14524);
   U4365 : NAND2_X1 port map( A1 => n425, A2 => n15046, ZN => n1065);
   U4366 : NAND2_X1 port map( A1 => n15227, A2 => n15343, ZN => n1066);
   U4369 : OAI21_X1 port map( B1 => n27954, B2 => n27965, A => n28636, ZN => 
                           n1068);
   U4370 : NAND2_X1 port map( A1 => n1069, A2 => n20322, ZN => n3341);
   U4371 : OAI22_X1 port map( A1 => n19956, A2 => n20319, B1 => n20324, B2 => 
                           n20323, ZN => n1069);
   U4372 : NAND2_X1 port map( A1 => n11782, A2 => n11502, ZN => n11420);
   U4373 : OAI211_X1 port map( C1 => n1292, C2 => n12343, A => n1070, B => 
                           n11474, ZN => n11475);
   U4374 : NAND2_X1 port map( A1 => n1290, A2 => n431, ZN => n1070);
   U4375 : NAND2_X1 port map( A1 => n1071, A2 => n11253, ZN => n4649);
   U4376 : NAND2_X1 port map( A1 => n11258, A2 => n11318, ZN => n1071);
   U4377 : NAND3_X1 port map( A1 => n15434, A2 => n15030, A3 => n14821, ZN => 
                           n14023);
   U4379 : OR2_X1 port map( A1 => n17277, A2 => n17276, ZN => n17004);
   U4380 : INV_X1 port map( A => n1073, ZN => n22875);
   U4383 : NAND2_X1 port map( A1 => n26432, A2 => n26361, ZN => n1075);
   U4384 : INV_X1 port map( A => n26425, ZN => n1076);
   U4385 : XNOR2_X1 port map( A => n19267, B => n6319, ZN => n17974);
   U4386 : INV_X1 port map( A => n12677, ZN => n1511);
   U4388 : NAND2_X1 port map( A1 => n12239, A2 => n11514, ZN => n4140);
   U4389 : NAND2_X1 port map( A1 => n1450, A2 => n4141, ZN => n1449);
   U4392 : AOI21_X1 port map( B1 => n2246, B2 => n24461, A => n24809, ZN => 
                           n23951);
   U4395 : NAND3_X1 port map( A1 => n1220, A2 => n1219, A3 => n10989, ZN => 
                           n1080);
   U4396 : NAND2_X1 port map( A1 => n11551, A2 => n11784, ZN => n1140);
   U4398 : NAND2_X1 port map( A1 => n1198, A2 => n7388, ZN => n7392);
   U4399 : NAND2_X1 port map( A1 => n21570, A2 => n21567, ZN => n1084);
   U4400 : XNOR2_X2 port map( A => n1085, B => n2293, ZN => n14393);
   U4401 : OAI211_X1 port map( C1 => n27326, C2 => n28641, A => n27325, B => 
                           n1086, ZN => Ciphertext(148));
   U4402 : NAND4_X1 port map( A1 => n27323, A2 => n27320, A3 => n27322, A4 => 
                           n27321, ZN => n1086);
   U4407 : XOR2_X1 port map( A => n22589, B => n2522, Z => n1773);
   U4408 : OAI21_X1 port map( B1 => n18001, B2 => n18334, A => n1087, ZN => 
                           n1649);
   U4409 : NAND3_X1 port map( A1 => n4586, A2 => n13724, A3 => n4331, ZN => 
                           n4330);
   U4410 : OAI211_X1 port map( C1 => n29086, C2 => n1091, A => n1090, B => 
                           n1089, ZN => n1088);
   U4411 : NAND2_X1 port map( A1 => n29086, A2 => n1466, ZN => n1089);
   U4412 : NAND3_X1 port map( A1 => n15434, A2 => n15432, A3 => n15030, ZN => 
                           n15034);
   U4413 : NOR2_X2 port map( A1 => n18030, A2 => n1092, ZN => n18981);
   U4414 : OAI22_X1 port map( A1 => n18027, A2 => n417, B1 => n29547, B2 => 
                           n18029, ZN => n1092);
   U4416 : NAND2_X1 port map( A1 => n7706, A2 => n7853, ZN => n2590);
   U4417 : NAND2_X1 port map( A1 => n7496, A2 => n7494, ZN => n7706);
   U4420 : INV_X1 port map( A => n4270, ZN => n17512);
   U4422 : XNOR2_X2 port map( A => n1094, B => n5784, ZN => n4270);
   U4424 : NAND2_X1 port map( A1 => n15271, A2 => n1095, ZN => n14615);
   U4425 : XOR2_X1 port map( A => n16246, B => n15639, Z => n1348);
   U4430 : NAND2_X1 port map( A1 => n8874, A2 => n8699, ZN => n8710);
   U4431 : OAI21_X1 port map( B1 => n1334, B2 => n20517, A => n20329, ZN => 
                           n1099);
   U4432 : NAND3_X1 port map( A1 => n14190, A2 => n14189, A3 => n14188, ZN => 
                           n15223);
   U4433 : INV_X1 port map( A => n17954, ZN => n20314);
   U4434 : OAI211_X1 port map( C1 => n11280, C2 => n584, A => n1100, B => n585,
                           ZN => n3018);
   U4435 : NAND2_X1 port map( A1 => n11280, A2 => n11281, ZN => n1100);
   U4437 : NAND2_X1 port map( A1 => n12079, A2 => n12296, ZN => n1101);
   U4438 : NAND3_X1 port map( A1 => n1104, A2 => n11482, A3 => n1103, ZN => 
                           n1102);
   U4439 : INV_X1 port map( A => n11796, ZN => n1104);
   U4440 : NAND2_X1 port map( A1 => n618, A2 => n7266, ZN => n8027);
   U4441 : XNOR2_X2 port map( A => n7027, B => Key(65), ZN => n7268);
   U4442 : XNOR2_X1 port map( A => n28566, B => n22641, ZN => n22565);
   U4443 : NAND2_X1 port map( A1 => n2619, A2 => n24437, ZN => n24120);
   U4444 : INV_X1 port map( A => n19923, ZN => n1105);
   U4445 : NAND2_X1 port map( A1 => n1106, A2 => n13976, ZN => n13977);
   U4447 : NAND2_X1 port map( A1 => n1108, A2 => n2256, ZN => n9292);
   U4448 : NAND2_X1 port map( A1 => n2255, A2 => n10946, ZN => n1108);
   U4449 : NAND2_X1 port map( A1 => n18415, A2 => n18416, ZN => n18417);
   U4452 : NAND2_X1 port map( A1 => n21660, A2 => n21656, ZN => n1110);
   U4453 : NAND2_X1 port map( A1 => n8304, A2 => n7942, ZN => n7659);
   U4454 : NAND3_X1 port map( A1 => n13857, A2 => n13858, A3 => n29036, ZN => 
                           n13860);
   U4456 : NAND2_X1 port map( A1 => n15557, A2 => n542, ZN => n1591);
   U4458 : NAND2_X1 port map( A1 => n13585, A2 => n13645, ZN => n1111);
   U4459 : NOR2_X2 port map( A1 => n11667, A2 => n11668, ZN => n13048);
   U4460 : MUX2_X1 port map( A => n1883, B => n24372, S => n24373, Z => n24381)
                           ;
   U4462 : NAND2_X1 port map( A1 => n15395, A2 => n1112, ZN => n1164);
   U4463 : NAND2_X1 port map( A1 => n14723, A2 => n15144, ZN => n1112);
   U4465 : NAND2_X1 port map( A1 => n1594, A2 => n17348, ZN => n1593);
   U4468 : NAND2_X1 port map( A1 => n7920, A2 => n7619, ZN => n7921);
   U4469 : OAI21_X1 port map( B1 => n8228, B2 => n8227, A => n8226, ZN => n8230
                           );
   U4470 : NAND2_X1 port map( A1 => n18124, A2 => n18589, ZN => n5475);
   U4471 : NAND2_X1 port map( A1 => n1115, A2 => n2944, ZN => n7537);
   U4472 : NAND2_X1 port map( A1 => n8162, A2 => n7349, ZN => n1115);
   U4473 : OAI21_X1 port map( B1 => n11318, B2 => n594, A => n1116, ZN => 
                           n11259);
   U4474 : NAND2_X1 port map( A1 => n11318, A2 => n2690, ZN => n1116);
   U4477 : NAND2_X1 port map( A1 => n9046, A2 => n5945, ZN => n1118);
   U4479 : NAND4_X2 port map( A1 => n2635, A2 => n18142, A3 => n2633, A4 => 
                           n18139, ZN => n18852);
   U4480 : OR2_X1 port map( A1 => n4188, A2 => n17259, ZN => n1374);
   U4482 : INV_X1 port map( A => n17025, ZN => n1121);
   U4483 : NAND2_X1 port map( A1 => n17026, A2 => n17025, ZN => n1122);
   U4484 : NAND3_X2 port map( A1 => n5525, A2 => n5524, A3 => n11808, ZN => 
                           n12776);
   U4485 : NAND2_X1 port map( A1 => n4799, A2 => n14429, ZN => n14199);
   U4486 : OAI21_X1 port map( B1 => n1125, B2 => n18511, A => n1124, ZN => 
                           n18274);
   U4487 : NAND3_X1 port map( A1 => n5931, A2 => n15284, A3 => n2893, ZN => 
                           n5930);
   U4489 : NAND2_X1 port map( A1 => n1127, A2 => n1126, ZN => n9145);
   U4490 : NAND2_X1 port map( A1 => n599, A2 => n9140, ZN => n1126);
   U4491 : NAND2_X1 port map( A1 => n13308, A2 => n263, ZN => n15083);
   U4493 : OR2_X1 port map( A1 => n24082, A2 => n24081, ZN => n1128);
   U4495 : NAND2_X1 port map( A1 => n1131, A2 => n1130, ZN => n1129);
   U4496 : AOI21_X1 port map( B1 => n17157, B2 => n16706, A => n17181, ZN => 
                           n1130);
   U4497 : NAND2_X1 port map( A1 => n17526, A2 => n531, ZN => n1131);
   U4499 : NAND2_X1 port map( A1 => n1625, A2 => n6605, ZN => n1132);
   U4500 : NAND2_X1 port map( A1 => n24998, A2 => n24999, ZN => n25052);
   U4501 : NAND2_X1 port map( A1 => n1135, A2 => n1134, ZN => n15332);
   U4502 : NAND2_X1 port map( A1 => n16968, A2 => n17421, ZN => n1134);
   U4503 : NAND2_X1 port map( A1 => n17305, A2 => n17012, ZN => n1135);
   U4506 : AND2_X1 port map( A1 => n13803, A2 => n13699, ZN => n12614);
   U4507 : NAND2_X1 port map( A1 => n1561, A2 => n1137, ZN => n6342);
   U4508 : XNOR2_X1 port map( A => n22710, B => n22923, ZN => n5841);
   U4509 : INV_X1 port map( A => n15184, ZN => n15186);
   U4510 : INV_X1 port map( A => n10287, ZN => n9311);
   U4512 : NOR2_X1 port map( A1 => n11000, A2 => n10997, ZN => n10683);
   U4513 : NAND2_X1 port map( A1 => n11233, A2 => n11234, ZN => n3442);
   U4514 : AOI21_X1 port map( B1 => n23221, B2 => n23222, A => n23220, ZN => 
                           n23225);
   U4515 : NAND2_X1 port map( A1 => n2708, A2 => n23700, ZN => n23221);
   U4516 : NAND2_X1 port map( A1 => n28810, A2 => n7935, ZN => n7609);
   U4519 : NAND2_X1 port map( A1 => n23740, A2 => n23741, ZN => n23742);
   U4520 : NAND2_X1 port map( A1 => n2911, A2 => n21624, ZN => n3227);
   U4521 : NAND2_X1 port map( A1 => n20381, A2 => n20567, ZN => n18624);
   U4522 : XNOR2_X2 port map( A => n12397, B => n12398, ZN => n5584);
   U4524 : NAND2_X1 port map( A1 => n1620, A2 => n7837, ZN => n1139);
   U4526 : XNOR2_X1 port map( A => n9627, B => n10079, ZN => n1141);
   U4527 : OAI21_X1 port map( B1 => n27603, B2 => n27604, A => n1142, ZN => 
                           n27606);
   U4528 : OAI21_X1 port map( B1 => n27602, B2 => n27607, A => n27617, ZN => 
                           n1142);
   U4529 : XOR2_X1 port map( A => n16616, B => n16141, Z => n1575);
   U4530 : XOR2_X1 port map( A => n22000, B => n22204, Z => n1640);
   U4531 : NAND2_X1 port map( A1 => n6663, A2 => n18197, ZN => n1143);
   U4532 : OAI21_X1 port map( B1 => n24243, B2 => n24242, A => n1144, ZN => 
                           n24244);
   U4533 : NAND2_X1 port map( A1 => n1217, A2 => n1145, ZN => n1144);
   U4534 : AND2_X1 port map( A1 => n24240, A2 => n24241, ZN => n1145);
   U4535 : INV_X1 port map( A => n4295, ZN => n1801);
   U4536 : NAND2_X1 port map( A1 => n9232, A2 => n9229, ZN => n8544);
   U4537 : OAI21_X2 port map( B1 => n6994, B2 => n6993, A => n6992, ZN => n9232
                           );
   U4539 : NAND2_X1 port map( A1 => n11065, A2 => n11242, ZN => n1146);
   U4541 : NAND2_X1 port map( A1 => n3924, A2 => n15343, ZN => n1148);
   U4542 : NAND2_X1 port map( A1 => n550, A2 => n425, ZN => n1149);
   U4544 : NAND2_X1 port map( A1 => n1808, A2 => n24341, ZN => n5795);
   U4547 : NAND2_X1 port map( A1 => n8663, A2 => n284, ZN => n1789);
   U4549 : NAND2_X1 port map( A1 => n24590, A2 => n24141, ZN => n24144);
   U4552 : NAND2_X1 port map( A1 => n23075, A2 => n23285, ZN => n1150);
   U4553 : NAND2_X1 port map( A1 => n23808, A2 => n23810, ZN => n1151);
   U4554 : NAND2_X1 port map( A1 => n2416, A2 => n15484, ZN => n16921);
   U4557 : NAND2_X1 port map( A1 => n17492, A2 => n536, ZN => n1153);
   U4558 : NAND2_X1 port map( A1 => n10778, A2 => n10958, ZN => n10779);
   U4559 : NAND3_X1 port map( A1 => n15733, A2 => n15732, A3 => n17236, ZN => 
                           n18488);
   U4560 : NAND2_X1 port map( A1 => n1154, A2 => n21547, ZN => n20932);
   U4561 : NAND2_X1 port map( A1 => n21553, A2 => n21519, ZN => n1154);
   U4562 : OAI21_X1 port map( B1 => n27715, B2 => n26126, A => n1155, ZN => 
                           n27696);
   U4563 : INV_X1 port map( A => n26889, ZN => n1155);
   U4564 : NAND2_X1 port map( A1 => n4980, A2 => n1156, ZN => n21727);
   U4565 : NAND2_X1 port map( A1 => n28223, A2 => n462, ZN => n1156);
   U4570 : NAND2_X1 port map( A1 => n1158, A2 => n442, ZN => n2414);
   U4571 : NAND2_X1 port map( A1 => n27627, A2 => n27632, ZN => n1158);
   U4573 : NAND2_X1 port map( A1 => n1159, A2 => n760, ZN => n23218);
   U4574 : NAND2_X1 port map( A1 => n23217, A2 => n476, ZN => n1159);
   U4575 : NAND2_X2 port map( A1 => n1160, A2 => n6146, ZN => n13226);
   U4576 : NAND2_X1 port map( A1 => n6145, A2 => n6658, ZN => n1160);
   U4577 : NAND2_X1 port map( A1 => n18034, A2 => n18033, ZN => n17621);
   U4579 : OR2_X1 port map( A1 => n8221, A2 => n7371, ZN => n1358);
   U4580 : AOI22_X1 port map( A1 => n26793, A2 => n28710, B1 => n26575, B2 => 
                           n26576, ZN => n26925);
   U4582 : NAND2_X1 port map( A1 => n1245, A2 => n5926, ZN => n22298);
   U4584 : NOR3_X1 port map( A1 => n25231, A2 => n25230, A3 => n26485, ZN => 
                           n25238);
   U4586 : NAND2_X1 port map( A1 => n19871, A2 => n3400, ZN => n19879);
   U4587 : XOR2_X1 port map( A => n16495, B => n15855, Z => n1234);
   U4588 : OAI21_X1 port map( B1 => n4557, B2 => n20474, A => n5528, ZN => 
                           n20739);
   U4589 : XNOR2_X1 port map( A => n22712, B => n20923, ZN => n1502);
   U4590 : AOI21_X1 port map( B1 => n5761, B2 => n26748, A => n5035, ZN => 
                           n26634);
   U4591 : NAND2_X1 port map( A1 => n27169, A2 => n28573, ZN => n24990);
   U4592 : XNOR2_X1 port map( A => n25412, B => n1302, ZN => n24982);
   U4594 : NAND2_X1 port map( A1 => n1166, A2 => n17227, ZN => n1165);
   U4595 : NAND2_X1 port map( A1 => n4717, A2 => n29138, ZN => n1167);
   U4596 : XNOR2_X2 port map( A => n12591, B => n12592, ZN => n13803);
   U4599 : NAND2_X1 port map( A1 => n17219, A2 => n17220, ZN => n17223);
   U4600 : OR2_X1 port map( A1 => n10517, A2 => n1854, ZN => n10520);
   U4601 : OR2_X1 port map( A1 => n7715, A2 => n6860, ZN => n8793);
   U4602 : AND2_X1 port map( A1 => n11113, A2 => n10461, ZN => n1494);
   U4604 : NOR2_X1 port map( A1 => n25650, A2 => n1169, ZN => n25276);
   U4605 : NAND3_X1 port map( A1 => n28494, A2 => n6621, A3 => n27372, ZN => 
                           n6620);
   U4606 : NAND2_X1 port map( A1 => n17205, A2 => n17818, ZN => n1170);
   U4607 : NAND4_X2 port map( A1 => n6192, A2 => n6189, A3 => n6190, A4 => 
                           n6191, ZN => n10384);
   U4608 : NAND2_X1 port map( A1 => n8362, A2 => n8361, ZN => n1171);
   U4609 : NAND2_X1 port map( A1 => n9012, A2 => n9016, ZN => n5676);
   U4611 : NAND2_X1 port map( A1 => n17232, A2 => n17361, ZN => n17236);
   U4612 : INV_X1 port map( A => n17263, ZN => n16991);
   U4613 : NAND2_X1 port map( A1 => n18136, A2 => n526, ZN => n2719);
   U4614 : NAND2_X1 port map( A1 => n24303, A2 => n24369, ZN => n1450);
   U4615 : NAND2_X1 port map( A1 => n16725, A2 => n17481, ZN => n4368);
   U4617 : NAND3_X1 port map( A1 => n598, A2 => n9140, A3 => n8185, ZN => n9141
                           );
   U4619 : OAI21_X1 port map( B1 => n4815, B2 => n11319, A => n11318, ZN => 
                           n1174);
   U4620 : NAND2_X1 port map( A1 => n8147, A2 => n7792, ZN => n7794);
   U4622 : NAND2_X1 port map( A1 => n18174, A2 => n18171, ZN => n1395);
   U4623 : AND3_X1 port map( A1 => n23678, A2 => n23676, A3 => n23131, ZN => 
                           n23365);
   U4624 : INV_X1 port map( A => n23469, ZN => n23649);
   U4625 : NAND2_X1 port map( A1 => n23469, A2 => n23647, ZN => n22433);
   U4626 : NAND2_X1 port map( A1 => n1441, A2 => n1443, ZN => n17946);
   U4627 : NAND2_X1 port map( A1 => n8360, A2 => n8433, ZN => n8362);
   U4629 : NAND2_X1 port map( A1 => n23684, A2 => n29544, ZN => n1176);
   U4630 : NAND2_X1 port map( A1 => n23685, A2 => n28457, ZN => n1177);
   U4631 : NAND2_X1 port map( A1 => n18087, A2 => n16985, ZN => n16843);
   U4632 : NAND3_X1 port map( A1 => n1546, A2 => n1547, A3 => n28004, ZN => 
                           n1545);
   U4633 : NAND2_X1 port map( A1 => n18332, A2 => n1180, ZN => n1973);
   U4634 : INV_X1 port map( A => n7840, ZN => n7420);
   U4635 : NAND2_X1 port map( A1 => n7835, A2 => n7840, ZN => n3112);
   U4636 : XNOR2_X2 port map( A => Key(87), B => Plaintext(87), ZN => n7840);
   U4637 : XOR2_X1 port map( A => n21855, B => n6364, Z => n1818);
   U4638 : AOI21_X1 port map( B1 => n17710, B2 => n17572, A => n423, ZN => 
                           n1366);
   U4639 : XNOR2_X1 port map( A => n10252, B => n1713, ZN => n10254);
   U4640 : NOR2_X2 port map( A1 => n21648, A2 => n1182, ZN => n22067);
   U4641 : OAI21_X1 port map( B1 => n21647, B2 => n21749, A => n21646, ZN => 
                           n1182);
   U4643 : XNOR2_X1 port map( A => n19650, B => n1183, ZN => n19282);
   U4644 : XNOR2_X1 port map( A => n19279, B => n19280, ZN => n1183);
   U4645 : NAND2_X1 port map( A1 => n21458, A2 => n21457, ZN => n20846);
   U4647 : XNOR2_X1 port map( A => n1185, B => n26106, ZN => n2902);
   U4648 : INV_X1 port map( A => n26107, ZN => n1185);
   U4649 : NAND2_X1 port map( A1 => n7912, A2 => n7628, ZN => n8291);
   U4650 : AOI21_X1 port map( B1 => n27630, B2 => n27616, A => n1186, ZN => 
                           n27622);
   U4652 : NAND3_X1 port map( A1 => n29600, A2 => n29299, A3 => n17263, ZN => 
                           n3878);
   U4653 : NAND2_X1 port map( A1 => n14516, A2 => n1904, ZN => n13668);
   U4654 : NAND2_X1 port map( A1 => n13979, A2 => n14743, ZN => n14516);
   U4655 : NAND3_X1 port map( A1 => n1353, A2 => n1700, A3 => n7888, ZN => 
                           n1352);
   U4656 : NAND2_X1 port map( A1 => n1413, A2 => n20165, ZN => n1188);
   U4657 : NAND2_X1 port map( A1 => n1415, A2 => n19993, ZN => n1189);
   U4658 : NAND2_X1 port map( A1 => n8371, A2 => n8372, ZN => n8373);
   U4659 : OR2_X1 port map( A1 => n11168, A2 => n11166, ZN => n10823);
   U4660 : OAI211_X1 port map( C1 => n11336, C2 => n11338, A => n1190, B => 
                           n10558, ZN => n2521);
   U4662 : NOR2_X1 port map( A1 => n18468, A2 => n1191, ZN => n6077);
   U4663 : NAND2_X1 port map( A1 => n18472, A2 => n18469, ZN => n1191);
   U4665 : NAND2_X1 port map( A1 => n9231, A2 => n6590, ZN => n5158);
   U4666 : NAND2_X1 port map( A1 => n21213, A2 => n21211, ZN => n21020);
   U4667 : NAND2_X1 port map( A1 => n4217, A2 => n17421, ZN => n16791);
   U4668 : NAND2_X1 port map( A1 => n1737, A2 => n16789, ZN => n4217);
   U4671 : NAND2_X1 port map( A1 => n504, A2 => n29584, ZN => n2555);
   U4672 : OAI21_X1 port map( B1 => n24677, B2 => n24678, A => n1194, ZN => 
                           n24399);
   U4673 : NAND2_X1 port map( A1 => n24677, A2 => n24395, ZN => n1194);
   U4674 : INV_X1 port map( A => n5714, ZN => n1738);
   U4675 : NAND2_X1 port map( A1 => n5645, A2 => n5644, ZN => n1244);
   U4676 : NOR2_X2 port map( A1 => n1356, A2 => n14606, ZN => n15309);
   U4679 : NAND2_X1 port map( A1 => n21680, A2 => n21675, ZN => n21672);
   U4680 : NAND2_X1 port map( A1 => n10586, A2 => n11468, ZN => n2589);
   U4681 : NAND2_X1 port map( A1 => n3700, A2 => n3699, ZN => n3698);
   U4682 : NAND3_X1 port map( A1 => n21401, A2 => n21749, A3 => n20658, ZN => 
                           n4647);
   U4685 : NAND2_X1 port map( A1 => n20518, A2 => n501, ZN => n1199);
   U4686 : NAND2_X1 port map( A1 => n1201, A2 => n28126, ZN => n1200);
   U4687 : NAND2_X1 port map( A1 => n20520, A2 => n20517, ZN => n1201);
   U4689 : NAND2_X1 port map( A1 => n1204, A2 => n1203, ZN => n1202);
   U4692 : NAND2_X1 port map( A1 => n6451, A2 => n6452, ZN => n21283);
   U4693 : OR2_X1 port map( A1 => n14468, A2 => n4840, ZN => n1628);
   U4694 : OR2_X1 port map( A1 => n18068, A2 => n18067, ZN => n1506);
   U4695 : NAND2_X1 port map( A1 => n7802, A2 => n7803, ZN => n7806);
   U4696 : NAND2_X1 port map( A1 => n23805, A2 => n28594, ZN => n1206);
   U4697 : INV_X1 port map( A => n15491, ZN => n14703);
   U4698 : XNOR2_X1 port map( A => n1505, B => n19243, ZN => n19020);
   U4699 : XNOR2_X2 port map( A => Key(41), B => Plaintext(41), ZN => n7336);
   U4702 : AOI21_X1 port map( B1 => n27097, B2 => n27531, A => n1208, ZN => 
                           n27098);
   U4703 : OAI22_X1 port map( A1 => n27509, A2 => n27527, B1 => n27531, B2 => 
                           n27221, ZN => n1208);
   U4704 : XNOR2_X1 port map( A => n1209, B => n9917, ZN => n9920);
   U4705 : XNOR2_X1 port map( A => n9918, B => n1920, ZN => n1209);
   U4706 : NAND3_X1 port map( A1 => n8905, A2 => n6147, A3 => n9013, ZN => 
                           n8907);
   U4707 : NAND2_X1 port map( A1 => n1596, A2 => n29632, ZN => n1592);
   U4708 : NAND2_X1 port map( A1 => n1593, A2 => n1595, ZN => n1596);
   U4709 : NAND2_X1 port map( A1 => n16687, A2 => n6380, ZN => n6379);
   U4711 : AOI21_X1 port map( B1 => n6469, B2 => n28822, A => n26949, ZN => 
                           n1210);
   U4712 : NAND2_X1 port map( A1 => n5903, A2 => n5904, ZN => n3089);
   U4713 : NAND2_X1 port map( A1 => n3147, A2 => n23771, ZN => n6543);
   U4714 : NAND2_X1 port map( A1 => n1211, A2 => n7835, ZN => n7842);
   U4715 : NAND2_X1 port map( A1 => n619, A2 => n7369, ZN => n1211);
   U4716 : AND2_X2 port map( A1 => n1213, A2 => n1212, ZN => n16586);
   U4717 : NAND2_X1 port map( A1 => n14809, A2 => n14810, ZN => n1212);
   U4718 : NAND2_X1 port map( A1 => n14811, A2 => n14812, ZN => n1213);
   U4719 : NAND2_X1 port map( A1 => n14715, A2 => n13922, ZN => n14811);
   U4721 : MUX2_X1 port map( A => n11286, B => n11285, S => n11284, Z => n1214)
                           ;
   U4722 : OAI22_X1 port map( A1 => n4423, A2 => n2974, B1 => n13903, B2 => 
                           n13902, ZN => n14020);
   U4724 : NAND2_X1 port map( A1 => n17481, A2 => n17476, ZN => n3171);
   U4726 : INV_X1 port map( A => n24559, ZN => n1217);
   U4727 : NAND3_X1 port map( A1 => n17663, A2 => n18343, A3 => n17906, ZN => 
                           n4075);
   U4728 : NAND2_X1 port map( A1 => n2769, A2 => n17569, ZN => n2768);
   U4729 : XNOR2_X1 port map( A => n1218, B => n22413, ZN => n22417);
   U4730 : XNOR2_X1 port map( A => n22412, B => n22411, ZN => n1218);
   U4731 : NAND2_X1 port map( A1 => n6636, A2 => n21465, ZN => n3936);
   U4734 : NAND2_X1 port map( A1 => n10985, A2 => n589, ZN => n1219);
   U4735 : NAND2_X1 port map( A1 => n3804, A2 => n10984, ZN => n1220);
   U4736 : OAI21_X1 port map( B1 => n14045, B2 => n13906, A => n14049, ZN => 
                           n14052);
   U4737 : NAND2_X1 port map( A1 => n12206, A2 => n12111, ZN => n1221);
   U4738 : XNOR2_X2 port map( A => n3663, B => n10300, ZN => n10972);
   U4739 : OAI21_X1 port map( B1 => n17815, B2 => n18045, A => n1224, ZN => 
                           n17816);
   U4740 : NAND3_X1 port map( A1 => n1894, A2 => n18148, A3 => n18430, ZN => 
                           n1224);
   U4743 : MUX2_X1 port map( A => n27551, B => n27571, S => n27573, Z => n27219
                           );
   U4746 : XNOR2_X1 port map( A => n1230, B => n1229, ZN => Ciphertext(64));
   U4747 : NAND3_X1 port map( A1 => n27284, A2 => n5331, A3 => n27283, ZN => 
                           n1230);
   U4748 : OR2_X1 port map( A1 => n1914, A2 => n28444, ZN => n23024);
   U4749 : INV_X1 port map( A => n17827, ZN => n1231);
   U4750 : NAND2_X1 port map( A1 => n27088, A2 => n27084, ZN => n27020);
   U4751 : XNOR2_X1 port map( A => n1234, B => n16627, ZN => n1233);
   U4752 : INV_X1 port map( A => n7967, ZN => n1568);
   U4755 : NAND3_X1 port map( A1 => n4348, A2 => n4347, A3 => n17673, ZN => 
                           n18520);
   U4756 : XNOR2_X1 port map( A => n10251, B => n1709, ZN => n1713);
   U4758 : AOI21_X1 port map( B1 => n7281, B2 => n7282, A => n8150, ZN => n1237
                           );
   U4760 : NAND2_X1 port map( A1 => n1238, A2 => n12300, ZN => n2219);
   U4762 : NAND2_X1 port map( A1 => n23813, A2 => n1239, ZN => n24472);
   U4763 : NOR2_X1 port map( A1 => n1240, A2 => n23814, ZN => n1239);
   U4765 : OAI22_X1 port map( A1 => n15847, A2 => n17553, B1 => n17224, B2 => 
                           n17556, ZN => n1241);
   U4768 : OR2_X2 port map( A1 => n1242, A2 => n7588, ZN => n8718);
   U4769 : NAND2_X1 port map( A1 => n2236, A2 => n2237, ZN => n1242);
   U4771 : NAND2_X1 port map( A1 => n1244, A2 => n15268, ZN => n1243);
   U4773 : NAND2_X1 port map( A1 => n24100, A2 => n29051, ZN => n23875);
   U4775 : OAI211_X1 port map( C1 => n24973, C2 => n24258, A => n471, B => n468
                           , ZN => n24259);
   U4777 : NAND2_X1 port map( A1 => n468, A2 => n23467, ZN => n1249);
   U4780 : MUX2_X1 port map( A => n468, B => n23467, S => n24976, Z => n24014);
   U4781 : OAI21_X2 port map( B1 => n17292, B2 => n28729, A => n6524, ZN => 
                           n6526);
   U4782 : NAND2_X1 port map( A1 => n17400, A2 => n17397, ZN => n1252);
   U4783 : XNOR2_X1 port map( A => n1254, B => n25728, ZN => n25733);
   U4784 : XNOR2_X1 port map( A => n1254, B => n25015, ZN => n24170);
   U4785 : XNOR2_X1 port map( A => n1254, B => n25432, ZN => n25433);
   U4787 : INV_X1 port map( A => n29037, ZN => n1255);
   U4790 : XNOR2_X1 port map( A => n16093, B => n16091, ZN => n1257);
   U4791 : NAND2_X1 port map( A1 => n1261, A2 => n1260, ZN => n10654);
   U4794 : NAND2_X1 port map( A1 => n1265, A2 => n1817, ZN => n1264);
   U4795 : NAND2_X1 port map( A1 => n1419, A2 => n16803, ZN => n1265);
   U4796 : NAND2_X1 port map( A1 => n17477, A2 => n3883, ZN => n1419);
   U4797 : XNOR2_X1 port map( A => n1266, B => n1271, ZN => n1270);
   U4799 : OR2_X1 port map( A1 => n3237, A2 => n628, ZN => n1268);
   U4800 : NAND2_X1 port map( A1 => n3237, A2 => n21088, ZN => n22394);
   U4801 : OR2_X1 port map( A1 => n21088, A2 => n628, ZN => n1269);
   U4802 : INV_X1 port map( A => n1271, ZN => n22773);
   U4803 : XNOR2_X1 port map( A => n1270, B => n22395, ZN => n3338);
   U4804 : NAND2_X1 port map( A1 => n5505, A2 => n26489, ZN => n1280);
   U4805 : NOR2_X1 port map( A1 => n24678, A2 => n29555, ZN => n24673);
   U4806 : NAND3_X1 port map( A1 => n6406, A2 => n24674, A3 => n1272, ZN => 
                           n24680);
   U4807 : NAND2_X1 port map( A1 => n1274, A2 => n1273, ZN => n1272);
   U4808 : NOR2_X1 port map( A1 => n24678, A2 => n404, ZN => n1273);
   U4809 : AOI21_X1 port map( B1 => n29054, B2 => n26928, A => n26927, ZN => 
                           n1281);
   U4810 : NAND2_X1 port map( A1 => n1276, A2 => n1275, ZN => n26712);
   U4811 : NAND2_X1 port map( A1 => n27433, A2 => n27439, ZN => n1275);
   U4812 : NAND2_X1 port map( A1 => n26829, A2 => n27434, ZN => n1276);
   U4813 : OAI211_X2 port map( C1 => n1279, C2 => n26166, A => n1278, B => 
                           n1277, ZN => n27439);
   U4814 : NAND2_X1 port map( A1 => n1280, A2 => n1281, ZN => n1278);
   U4817 : NAND2_X1 port map( A1 => n23074, A2 => n23285, ZN => n22878);
   U4818 : NAND2_X1 port map( A1 => n5265, A2 => n1285, ZN => n4171);
   U4819 : NAND2_X1 port map( A1 => n10723, A2 => n1285, ZN => n10725);
   U4820 : NAND2_X1 port map( A1 => n5743, A2 => n1286, ZN => n5742);
   U4821 : NAND2_X1 port map( A1 => n23474, A2 => n29620, ZN => n1286);
   U4822 : NAND2_X1 port map( A1 => n4546, A2 => n17977, ZN => n17976);
   U4823 : NAND2_X1 port map( A1 => n1287, A2 => n23428, ZN => n23424);
   U4824 : NAND3_X1 port map( A1 => n21591, A2 => n5983, A3 => n1921, ZN => 
                           n4962);
   U4825 : NAND2_X1 port map( A1 => n21588, A2 => n29569, ZN => n1289);
   U4826 : AOI21_X1 port map( B1 => n21323, B2 => n21588, A => n1921, ZN => 
                           n21324);
   U4827 : NOR2_X1 port map( A1 => n1291, A2 => n12337, ZN => n1290);
   U4828 : INV_X1 port map( A => n12026, ZN => n1291);
   U4829 : INV_X1 port map( A => n20354, ZN => n19032);
   U4831 : XNOR2_X1 port map( A => n1293, B => n13556, ZN => n13152);
   U4832 : XNOR2_X1 port map( A => n1293, B => n12854, ZN => n11939);
   U4833 : XNOR2_X1 port map( A => n13263, B => n1293, ZN => n12435);
   U4834 : XNOR2_X1 port map( A => n13244, B => n1293, ZN => n12538);
   U4835 : NAND2_X1 port map( A1 => n1296, A2 => n1295, ZN => n1297);
   U4836 : NAND2_X1 port map( A1 => n7367, A2 => n7840, ZN => n1296);
   U4837 : NAND2_X1 port map( A1 => n7370, A2 => n370, ZN => n1298);
   U4838 : NAND3_X1 port map( A1 => n23075, A2 => n23074, A3 => n29102, ZN => 
                           n22743);
   U4839 : OAI21_X1 port map( B1 => n23074, B2 => n23806, A => n23810, ZN => 
                           n22638);
   U4840 : NAND2_X1 port map( A1 => n24263, A2 => n28522, ZN => n1299);
   U4842 : OAI21_X1 port map( B1 => n24298, B2 => n1301, A => n1300, ZN => 
                           n1303);
   U4843 : OAI21_X1 port map( B1 => n24298, B2 => n6198, A => n630, ZN => n1300
                           );
   U4844 : NOR2_X2 port map( A1 => n18096, A2 => n18091, ZN => n17793);
   U4845 : NAND2_X1 port map( A1 => n1308, A2 => n10937, ZN => n9417);
   U4846 : AND2_X1 port map( A1 => n1308, A2 => n10936, ZN => n11005);
   U4847 : NAND2_X1 port map( A1 => n11002, A2 => n28407, ZN => n3640);
   U4848 : NOR2_X1 port map( A1 => n11002, A2 => n28407, ZN => n10684);
   U4849 : OAI21_X1 port map( B1 => n10999, B2 => n10936, A => n1308, ZN => 
                           n9693);
   U4850 : NAND3_X1 port map( A1 => n11002, A2 => n5573, A3 => n28407, ZN => 
                           n11007);
   U4851 : NAND3_X1 port map( A1 => n14614, A2 => n14615, A3 => n632, ZN => 
                           n1309);
   U4852 : XNOR2_X1 port map( A => n1310, B => n857, ZN => n16046);
   U4853 : XNOR2_X1 port map( A => n15070, B => n1310, ZN => n15796);
   U4854 : XNOR2_X1 port map( A => n9645, B => n9746, ZN => n9687);
   U4856 : NAND3_X1 port map( A1 => n8961, A2 => n8963, A3 => n9171, ZN => 
                           n1311);
   U4858 : OAI21_X1 port map( B1 => n21269, B2 => n20818, A => n20711, ZN => 
                           n1312);
   U4859 : NAND2_X1 port map( A1 => n21266, A2 => n20816, ZN => n20818);
   U4860 : NOR2_X2 port map( A1 => n20876, A2 => n20877, ZN => n21269);
   U4862 : NAND2_X1 port map( A1 => n6362, A2 => n1314, ZN => n6363);
   U4863 : NAND2_X1 port map( A1 => n1314, A2 => n21150, ZN => n21151);
   U4864 : NAND3_X1 port map( A1 => n1318, A2 => n12181, A3 => n1319, ZN => 
                           n1317);
   U4866 : NAND2_X1 port map( A1 => n10441, A2 => n570, ZN => n1316);
   U4867 : NAND2_X1 port map( A1 => n1890, A2 => n12124, ZN => n1319);
   U4868 : INV_X1 port map( A => n14177, ZN => n1320);
   U4870 : NAND2_X1 port map( A1 => n13850, A2 => n1322, ZN => n1321);
   U4871 : NAND2_X1 port map( A1 => n1324, A2 => n1323, ZN => n4299);
   U4872 : NAND2_X1 port map( A1 => n14991, A2 => n15389, ZN => n1323);
   U4873 : NAND2_X1 port map( A1 => n1326, A2 => n15145, ZN => n1324);
   U4875 : AOI21_X1 port map( B1 => n21644, B2 => n1327, A => n21643, ZN => 
                           n21648);
   U4876 : NAND2_X1 port map( A1 => n15275, A2 => n15513, ZN => n1328);
   U4877 : NAND3_X2 port map( A1 => n1748, A2 => n1749, A3 => n6511, ZN => 
                           n15274);
   U4879 : AOI21_X1 port map( B1 => n2930, B2 => n2931, A => n20567, ZN => 
                           n1329);
   U4880 : OAI21_X1 port map( B1 => n6237, B2 => n97, A => n6236, ZN => n1330);
   U4883 : NAND2_X1 port map( A1 => n17458, A2 => n421, ZN => n1332);
   U4884 : NAND3_X1 port map( A1 => n17116, A2 => n16812, A3 => n17118, ZN => 
                           n1333);
   U4885 : NAND2_X1 port map( A1 => n29083, A2 => n29539, ZN => n17458);
   U4887 : AND2_X1 port map( A1 => n415, A2 => n6843, ZN => n5934);
   U4888 : NAND2_X1 port map( A1 => n6840, A2 => n507, ZN => n6839);
   U4889 : NAND2_X1 port map( A1 => n19505, A2 => n507, ZN => n6838);
   U4890 : NAND2_X1 port map( A1 => n19796, A2 => n28126, ZN => n1334);
   U4891 : OAI211_X2 port map( C1 => n2843, C2 => n1337, A => n1521, B => n1336
                           , ZN => n12132);
   U4892 : INV_X1 port map( A => n1704, ZN => n1337);
   U4893 : NAND2_X1 port map( A1 => n3820, A2 => n1338, ZN => n10838);
   U4894 : NAND2_X1 port map( A1 => n3817, A2 => n1338, ZN => n1440);
   U4897 : OAI22_X1 port map( A1 => n1340, A2 => n22011, B1 => n20762, B2 => 
                           n4828, ZN => n1339);
   U4899 : NAND2_X1 port map( A1 => n21823, A2 => n4828, ZN => n1340);
   U4900 : AOI21_X1 port map( B1 => n21077, B2 => n1342, A => n21823, ZN => 
                           n22014);
   U4901 : XNOR2_X2 port map( A => n13149, B => n13148, ZN => n14327);
   U4903 : OAI211_X1 port map( C1 => n14324, C2 => n13653, A => n14322, B => 
                           n14323, ZN => n1344);
   U4904 : NAND2_X1 port map( A1 => n1346, A2 => n14328, ZN => n1345);
   U4906 : NAND3_X1 port map( A1 => n3731, A2 => n6506, A3 => n1808, ZN => 
                           n2460);
   U4907 : NAND3_X1 port map( A1 => n7774, A2 => n1350, A3 => n438, ZN => n1349
                           );
   U4908 : NAND2_X1 port map( A1 => n3188, A2 => n438, ZN => n1351);
   U4909 : NAND2_X1 port map( A1 => n7774, A2 => n7777, ZN => n1353);
   U4910 : XNOR2_X1 port map( A => n10019, B => n1884, ZN => n8883);
   U4911 : NAND2_X1 port map( A1 => n8739, A2 => n8369, ZN => n1417);
   U4912 : NAND3_X1 port map( A1 => n11213, A2 => n11212, A3 => n1357, ZN => 
                           n11214);
   U4913 : AOI21_X1 port map( B1 => n1358, B2 => n7696, A => n7695, ZN => n7699
                           );
   U4914 : OR2_X1 port map( A1 => n10680, A2 => n29577, ZN => n11983);
   U4915 : NAND2_X1 port map( A1 => n11984, A2 => n11983, ZN => n12231);
   U4916 : AND2_X1 port map( A1 => n5265, A2 => n10970, ZN => n1359);
   U4919 : OAI21_X1 port map( B1 => n17562, B2 => n532, A => n4220, ZN => n1361
                           );
   U4920 : NAND2_X1 port map( A1 => n4873, A2 => n17561, ZN => n1362);
   U4921 : NAND2_X1 port map( A1 => n4220, A2 => n17315, ZN => n17561);
   U4922 : OR2_X1 port map( A1 => n17313, A2 => n17312, ZN => n4873);
   U4923 : NAND2_X1 port map( A1 => n423, A2 => n17570, ZN => n2819);
   U4924 : NAND2_X1 port map( A1 => n17320, A2 => n17707, ZN => n1365);
   U4926 : NAND3_X1 port map( A1 => n389, A2 => n1368, A3 => n4425, ZN => n3741
                           );
   U4927 : OR2_X1 port map( A1 => n14144, A2 => n1368, ZN => n6924);
   U4928 : NAND2_X1 port map( A1 => n4423, A2 => n1368, ZN => n14018);
   U4929 : NAND2_X1 port map( A1 => n265, A2 => n13901, ZN => n4421);
   U4930 : OAI21_X1 port map( B1 => n389, B2 => n1368, A => n14141, ZN => 
                           n14145);
   U4931 : NAND2_X1 port map( A1 => n1368, A2 => n2974, ZN => n14141);
   U4932 : NAND3_X1 port map( A1 => n12355, A2 => n1370, A3 => n1369, ZN => 
                           n12461);
   U4933 : NAND2_X1 port map( A1 => n10586, A2 => n1371, ZN => n1370);
   U4935 : NAND3_X1 port map( A1 => n4085, A2 => n1374, A3 => n17262, ZN => 
                           n1373);
   U4936 : NOR2_X1 port map( A1 => n12207, A2 => n12210, ZN => n12209);
   U4937 : NAND2_X1 port map( A1 => n9653, A2 => n11043, ZN => n1375);
   U4938 : OAI21_X1 port map( B1 => n28370, B2 => n17582, A => n1377, ZN => 
                           n1376);
   U4939 : NAND2_X1 port map( A1 => n524, A2 => n17771, ZN => n6912);
   U4940 : NAND2_X1 port map( A1 => n524, A2 => n1378, ZN => n1377);
   U4941 : NAND2_X1 port map( A1 => n7373, A2 => n1379, ZN => n7374);
   U4942 : NAND3_X1 port map( A1 => n8227, A2 => n28721, A3 => n8221, ZN => 
                           n1379);
   U4943 : INV_X1 port map( A => n6988, ZN => n8227);
   U4944 : NAND2_X1 port map( A1 => n592, A2 => n1380, ZN => n2554);
   U4946 : XNOR2_X1 port map( A => n9745, B => n9744, ZN => n11010);
   U4947 : INV_X1 port map( A => n11010, ZN => n1381);
   U4948 : OAI21_X1 port map( B1 => n10628, B2 => n11235, A => n11012, ZN => 
                           n10579);
   U4949 : NAND2_X1 port map( A1 => n1381, A2 => n11235, ZN => n11012);
   U4950 : INV_X1 port map( A => n11010, ZN => n6108);
   U4951 : NOR2_X1 port map( A1 => n16338, A2 => n1382, ZN => n16493);
   U4952 : AND2_X1 port map( A1 => n6079, A2 => n1384, ZN => n1382);
   U4953 : NAND2_X1 port map( A1 => n1384, A2 => n18466, ZN => n18472);
   U4954 : AND2_X1 port map( A1 => n18467, A2 => n1384, ZN => n18314);
   U4955 : AOI21_X1 port map( B1 => n17915, B2 => n1384, A => n18006, ZN => 
                           n18010);
   U4956 : NAND2_X1 port map( A1 => n16442, A2 => n1383, ZN => n16492);
   U4958 : NAND2_X1 port map( A1 => n603, A2 => n1386, ZN => n9580);
   U4959 : NAND2_X1 port map( A1 => n7912, A2 => n8290, ZN => n7913);
   U4960 : NAND2_X1 port map( A1 => n1388, A2 => n1961, ZN => n14969);
   U4961 : NAND2_X1 port map( A1 => n13470, A2 => n13469, ZN => n1388);
   U4962 : OAI211_X1 port map( C1 => n8914, C2 => n9107, A => n8071, B => n8669
                           , ZN => n8072);
   U4963 : NAND2_X1 port map( A1 => n8071, A2 => n8669, ZN => n8916);
   U4965 : NAND2_X1 port map( A1 => n23155, A2 => n1641, ZN => n1391);
   U4966 : MUX2_X1 port map( A => n17535, B => n17536, S => n18242, Z => n17538
                           );
   U4967 : NAND3_X1 port map( A1 => n14696, A2 => n14845, A3 => n14695, ZN => 
                           n1393);
   U4968 : NAND2_X1 port map( A1 => n28198, A2 => n14842, ZN => n1394);
   U4969 : NAND2_X1 port map( A1 => n1395, A2 => n18170, ZN => n2591);
   U4970 : NAND2_X1 port map( A1 => n18169, A2 => n1395, ZN => n18177);
   U4971 : NOR2_X1 port map( A1 => n10622, A2 => n11227, ZN => n10624);
   U4972 : XNOR2_X1 port map( A => n9956, B => n260, ZN => n1396);
   U4973 : XNOR2_X1 port map( A => n9722, B => n9721, ZN => n1397);
   U4974 : NAND2_X1 port map( A1 => n436, A2 => n1398, ZN => n8988);
   U4975 : NOR2_X1 port map( A1 => n609, A2 => n8981, ZN => n1398);
   U4976 : NAND3_X1 port map( A1 => n10883, A2 => n11209, A3 => n11085, ZN => 
                           n1400);
   U4978 : OAI21_X1 port map( B1 => n12429, B2 => n12428, A => n5134, ZN => 
                           n1401);
   U4979 : OR2_X1 port map( A1 => n12354, A2 => n580, ZN => n5134);
   U4980 : OR2_X1 port map( A1 => n7088, A2 => n438, ZN => n1404);
   U4981 : NAND2_X1 port map( A1 => n1403, A2 => n1402, ZN => n4938);
   U4982 : NAND2_X1 port map( A1 => n7088, A2 => n1700, ZN => n1402);
   U4983 : NAND2_X1 port map( A1 => n4939, A2 => n438, ZN => n1403);
   U4985 : OAI21_X1 port map( B1 => n17316, B2 => n790, A => n1406, ZN => n1405
                           );
   U4986 : OR2_X1 port map( A1 => n4220, A2 => n17315, ZN => n1406);
   U4988 : NAND3_X1 port map( A1 => n27301, A2 => n6150, A3 => n395, ZN => 
                           n1407);
   U4989 : XNOR2_X1 port map( A => n1410, B => n1412, ZN => Ciphertext(70));
   U4990 : NAND3_X1 port map( A1 => n5425, A2 => n29493, A3 => n444, ZN => 
                           n1411);
   U4992 : NAND2_X1 port map( A1 => n20223, A2 => n297, ZN => n1415);
   U4993 : NAND2_X1 port map( A1 => n6578, A2 => n20219, ZN => n20223);
   U4994 : NAND2_X1 port map( A1 => n6901, A2 => n8734, ZN => n1418);
   U4995 : NOR2_X1 port map( A1 => n1419, A2 => n16723, ZN => n17667);
   U4997 : INV_X1 port map( A => n29307, ZN => n1420);
   U5000 : NAND2_X1 port map( A1 => n1425, A2 => n1423, ZN => n1422);
   U5001 : NAND2_X1 port map( A1 => n29309, A2 => n23945, ZN => n1423);
   U5002 : NAND3_X1 port map( A1 => n470, A2 => n463, A3 => n29309, ZN => n1424
                           );
   U5003 : OR2_X1 port map( A1 => n1427, A2 => n1470, ZN => n1469);
   U5004 : NOR2_X1 port map( A1 => n26484, A2 => n26731, ZN => n1427);
   U5005 : NAND2_X1 port map( A1 => n20197, A2 => n20589, ZN => n1428);
   U5007 : INV_X1 port map( A => n13802, ZN => n1430);
   U5008 : NAND2_X1 port map( A1 => n14319, A2 => n14317, ZN => n13802);
   U5009 : OR2_X1 port map( A1 => n13802, A2 => n560, ZN => n13712);
   U5010 : OAI21_X1 port map( B1 => n13258, B2 => n1430, A => n560, ZN => n2331
                           );
   U5012 : NAND2_X1 port map( A1 => n28191, A2 => n17941, ZN => n17763);
   U5013 : NAND2_X1 port map( A1 => n28191, A2 => n1433, ZN => n17944);
   U5014 : NOR2_X1 port map( A1 => n1434, A2 => n17942, ZN => n17602);
   U5015 : NAND2_X1 port map( A1 => n525, A2 => n17762, ZN => n1434);
   U5016 : NAND3_X1 port map( A1 => n17937, A2 => n17939, A3 => n28191, ZN => 
                           n16189);
   U5017 : INV_X1 port map( A => n1438, ZN => n1574);
   U5018 : NAND2_X1 port map( A1 => n1657, A2 => n1438, ZN => n16852);
   U5019 : NAND3_X1 port map( A1 => n1658, A2 => n1657, A3 => n1437, ZN => 
                           n1656);
   U5020 : OAI21_X1 port map( B1 => n16780, B2 => n16850, A => n1438, ZN => 
                           n16781);
   U5021 : NAND2_X1 port map( A1 => n501, A2 => n20261, ZN => n19794);
   U5022 : NAND3_X1 port map( A1 => n501, A2 => n20261, A3 => n28133, ZN => 
                           n21362);
   U5023 : NAND2_X1 port map( A1 => n1439, A2 => n5716, ZN => n12080);
   U5024 : OAI22_X1 port map( A1 => n11251, A2 => n11250, B1 => n29149, B2 => 
                           n586, ZN => n1439);
   U5025 : NAND2_X1 port map( A1 => n1440, A2 => n3818, ZN => n11251);
   U5026 : XNOR2_X2 port map( A => n9578, B => n9933, ZN => n11033);
   U5027 : NAND2_X1 port map( A1 => n1442, A2 => n17941, ZN => n1463);
   U5028 : NAND2_X1 port map( A1 => n1442, A2 => n17939, ZN => n1441);
   U5029 : NAND2_X1 port map( A1 => n17940, A2 => n519, ZN => n1443);
   U5030 : XNOR2_X1 port map( A => n22334, B => n21955, ZN => n22809);
   U5032 : NAND2_X1 port map( A1 => n21450, A2 => n21675, ZN => n1445);
   U5033 : INV_X1 port map( A => n1617, ZN => n6111);
   U5034 : OAI211_X1 port map( C1 => n28431, C2 => n22084, A => n1635, B => 
                           n6099, ZN => n1446);
   U5035 : XNOR2_X1 port map( A => n25508, B => n2602, ZN => n24306);
   U5036 : NOR2_X2 port map( A1 => n1449, A2 => n1447, ZN => n25508);
   U5037 : AOI21_X1 port map( B1 => n1448, B2 => n24305, A => n23897, ZN => 
                           n1447);
   U5038 : XNOR2_X1 port map( A => n2532, B => n22389, ZN => n1451);
   U5039 : NAND2_X1 port map( A1 => n1453, A2 => n29137, ZN => n1668);
   U5041 : NOR2_X1 port map( A1 => n15132, A2 => n15127, ZN => n1454);
   U5043 : NAND2_X1 port map( A1 => n1454, A2 => n13632, ZN => n13635);
   U5044 : NAND2_X1 port map( A1 => n17943, A2 => n1457, ZN => n1456);
   U5045 : NAND2_X1 port map( A1 => n517, A2 => n28656, ZN => n1457);
   U5046 : XNOR2_X1 port map( A => n1459, B => n27894, ZN => n25837);
   U5047 : XNOR2_X1 port map( A => n1459, B => n25351, ZN => n25082);
   U5048 : NAND2_X1 port map( A1 => n21230, A2 => n21409, ZN => n4632);
   U5050 : NAND2_X1 port map( A1 => n1467, A2 => n1465, ZN => n1464);
   U5051 : INV_X1 port map( A => n16679, ZN => n1466);
   U5052 : NAND2_X1 port map( A1 => n16814, A2 => n17282, ZN => n1467);
   U5053 : AOI22_X1 port map( A1 => n25641, A2 => n29579, B1 => n1473, B2 => 
                           n1472, ZN => n1471);
   U5054 : NOR2_X1 port map( A1 => n26480, A2 => n29579, ZN => n1473);
   U5056 : XNOR2_X1 port map( A => n26029, B => n4263, ZN => n25507);
   U5057 : NAND2_X1 port map( A1 => n23502, A2 => n23945, ZN => n1476);
   U5058 : NAND2_X1 port map( A1 => n1478, A2 => n458, ZN => n1477);
   U5059 : AOI21_X1 port map( B1 => n24780, B2 => n23946, A => n23945, ZN => 
                           n1478);
   U5060 : NAND2_X1 port map( A1 => n24454, A2 => n24775, ZN => n1479);
   U5062 : NAND2_X1 port map( A1 => n17280, A2 => n4246, ZN => n1481);
   U5064 : NAND2_X1 port map( A1 => n1485, A2 => n11708, ZN => n11709);
   U5065 : NAND2_X1 port map( A1 => n11648, A2 => n12145, ZN => n1484);
   U5066 : NAND2_X1 port map( A1 => n15286, A2 => n14696, ZN => n15287);
   U5068 : AND2_X1 port map( A1 => n14842, A2 => n28996, ZN => n15286);
   U5071 : NAND2_X1 port map( A1 => n11645, A2 => n1487, ZN => n3143);
   U5072 : NOR2_X1 port map( A1 => n573, A2 => n11715, ZN => n1487);
   U5075 : NAND2_X1 port map( A1 => n11437, A2 => n12265, ZN => n1490);
   U5077 : NAND2_X1 port map( A1 => n1493, A2 => n11552, ZN => n11554);
   U5078 : NAND2_X1 port map( A1 => n1669, A2 => n1493, ZN => n11504);
   U5079 : NAND2_X1 port map( A1 => n11115, A2 => n11113, ZN => n4128);
   U5080 : NAND2_X1 port map( A1 => n11115, A2 => n1494, ZN => n4630);
   U5082 : NAND3_X1 port map( A1 => n24484, A2 => n1496, A3 => n1497, ZN => 
                           n1495);
   U5083 : NAND2_X1 port map( A1 => n29597, A2 => n24209, ZN => n1496);
   U5084 : NAND2_X1 port map( A1 => n24480, A2 => n24479, ZN => n1497);
   U5086 : INV_X1 port map( A => n19229, ZN => n1504);
   U5087 : XNOR2_X1 port map( A => n19349, B => n1503, ZN => n19518);
   U5088 : NOR2_X1 port map( A1 => n4317, A2 => n1507, ZN => n1509);
   U5089 : NAND2_X1 port map( A1 => n15884, A2 => n17037, ZN => n1508);
   U5090 : XNOR2_X1 port map( A => n12677, B => n1510, ZN => n13177);
   U5091 : INV_X1 port map( A => n13175, ZN => n1510);
   U5092 : XNOR2_X1 port map( A => n1511, B => n13380, ZN => n13383);
   U5093 : XNOR2_X1 port map( A => n22459, B => n633, ZN => n21779);
   U5094 : NAND3_X1 port map( A1 => n1513, A2 => n7796, A3 => n7794, ZN => 
                           n1512);
   U5095 : NAND2_X1 port map( A1 => n7541, A2 => n7793, ZN => n1513);
   U5096 : XNOR2_X2 port map( A => n7149, B => Key(24), ZN => n7793);
   U5097 : NAND2_X1 port map( A1 => n1516, A2 => n28528, ZN => n25007);
   U5098 : NAND2_X1 port map( A1 => n25009, A2 => n28528, ZN => n1517);
   U5099 : INV_X1 port map( A => n15514, ZN => n15510);
   U5100 : AND2_X1 port map( A1 => n1519, A2 => n14438, ZN => n3851);
   U5101 : INV_X1 port map( A => n1876, ZN => n1519);
   U5102 : OR2_X1 port map( A1 => n14438, A2 => n1841, ZN => n13959);
   U5103 : OAI21_X1 port map( B1 => n13957, B2 => n13671, A => n28200, ZN => 
                           n4300);
   U5104 : OAI21_X2 port map( B1 => n28200, B2 => n13849, A => n13848, ZN => 
                           n15168);
   U5105 : NAND3_X1 port map( A1 => n586, A2 => n11248, A3 => n29148, ZN => 
                           n1521);
   U5107 : INV_X1 port map( A => n18232, ZN => n18401);
   U5108 : NAND2_X1 port map( A1 => n18399, A2 => n18232, ZN => n1523);
   U5109 : NAND2_X1 port map( A1 => n390, A2 => n11867, ZN => n6304);
   U5110 : NAND2_X1 port map( A1 => n4126, A2 => n11116, ZN => n1525);
   U5112 : XNOR2_X2 port map( A => n25266, B => n25265, ZN => n26753);
   U5115 : XNOR2_X1 port map( A => n22592, B => n6938, ZN => n23825);
   U5116 : OAI21_X2 port map( B1 => n21297, B2 => n21296, A => n21295, ZN => 
                           n22644);
   U5119 : NAND2_X1 port map( A1 => n9146, A2 => n8929, ZN => n1529);
   U5120 : OR2_X2 port map( A1 => n7374, A2 => n7375, ZN => n9146);
   U5121 : AOI21_X1 port map( B1 => n1530, B2 => n18042, A => n29595, ZN => 
                           n18044);
   U5122 : AND2_X2 port map( A1 => n16855, A2 => n16854, ZN => n18042);
   U5123 : INV_X1 port map( A => n22531, ZN => n23833);
   U5124 : INV_X1 port map( A => n1534, ZN => n27941);
   U5125 : OAI211_X1 port map( C1 => n27016, C2 => n27017, A => n1536, B => 
                           n1535, ZN => n1534);
   U5126 : NAND2_X1 port map( A1 => n28441, A2 => n28451, ZN => n1775);
   U5127 : NAND2_X1 port map( A1 => n27011, A2 => n28446, ZN => n1536);
   U5128 : INV_X1 port map( A => n11315, ZN => n2689);
   U5129 : NAND2_X1 port map( A1 => n4327, A2 => n1537, ZN => n4329);
   U5130 : AOI21_X1 port map( B1 => n2094, B2 => n29486, A => n26735, ZN => 
                           n28102);
   U5132 : NAND2_X1 port map( A1 => n21533, A2 => n21534, ZN => n1541);
   U5133 : NAND3_X1 port map( A1 => n1544, A2 => n21536, A3 => n1543, ZN => 
                           n1542);
   U5134 : INV_X1 port map( A => n21531, ZN => n1544);
   U5135 : XNOR2_X1 port map( A => n1545, B => n28007, ZN => Ciphertext(171));
   U5136 : NAND3_X1 port map( A1 => n1548, A2 => n28002, A3 => n443, ZN => 
                           n1547);
   U5137 : NAND3_X1 port map( A1 => n23897, A2 => n25006, A3 => n28415, ZN => 
                           n1549);
   U5138 : NAND2_X1 port map( A1 => n1550, A2 => n1549, ZN => n4558);
   U5139 : NAND2_X1 port map( A1 => n4559, A2 => n1551, ZN => n1550);
   U5140 : NAND2_X1 port map( A1 => n12321, A2 => n12050, ZN => n1552);
   U5141 : NAND3_X1 port map( A1 => n12318, A2 => n12319, A3 => n1552, ZN => 
                           n2979);
   U5142 : NAND2_X1 port map( A1 => n428, A2 => n14295, ZN => n13805);
   U5143 : NAND2_X1 port map( A1 => n13806, A2 => n428, ZN => n13702);
   U5144 : NAND2_X1 port map( A1 => n17712, A2 => n18263, ZN => n3834);
   U5146 : NAND2_X1 port map( A1 => n16919, A2 => n790, ZN => n1553);
   U5147 : NAND2_X1 port map( A1 => n16920, A2 => n17317, ZN => n1554);
   U5150 : NAND2_X1 port map( A1 => n23555, A2 => n477, ZN => n1555);
   U5151 : MUX2_X1 port map( A => n24635, B => n24634, S => n24633, Z => n25793
                           );
   U5152 : NAND2_X1 port map( A1 => n23187, A2 => n23557, ZN => n1558);
   U5155 : NAND2_X1 port map( A1 => n1562, A2 => n1563, ZN => n1561);
   U5156 : NAND2_X1 port map( A1 => n18173, A2 => n18170, ZN => n1562);
   U5157 : NAND2_X1 port map( A1 => n20432, A2 => n1565, ZN => n1564);
   U5159 : INV_X1 port map( A => n19920, ZN => n20255);
   U5164 : OAI21_X1 port map( B1 => n7678, B2 => n4697, A => n1567, ZN => n6540
                           );
   U5165 : NAND2_X1 port map( A1 => n7676, A2 => n4697, ZN => n1567);
   U5166 : NAND3_X2 port map( A1 => n1569, A2 => n4251, A3 => n4252, ZN => 
                           n15190);
   U5167 : XNOR2_X1 port map( A => n1572, B => n10188, ZN => n1761);
   U5168 : XNOR2_X1 port map( A => n1572, B => n9518, ZN => n9522);
   U5169 : XNOR2_X1 port map( A => n9805, B => n1572, ZN => n9809);
   U5170 : AOI21_X1 port map( B1 => n17262, B2 => n1574, A => n17260, ZN => 
                           n16782);
   U5173 : NAND2_X1 port map( A1 => n16850, A2 => n1574, ZN => n16150);
   U5179 : INV_X1 port map( A => n12938, ZN => n1580);
   U5181 : MUX2_X1 port map( A => n16995, B => n16992, S => n17263, Z => n1581)
                           ;
   U5182 : NAND2_X1 port map( A1 => n28176, A2 => n1865, ZN => n6542);
   U5186 : NAND2_X1 port map( A1 => n1584, A2 => n1585, ZN => n8574);
   U5187 : NAND2_X1 port map( A1 => n1586, A2 => n1587, ZN => n1584);
   U5188 : OAI21_X1 port map( B1 => n7777, B2 => n7890, A => n1354, ZN => n1588
                           );
   U5189 : NAND2_X1 port map( A1 => n7317, A2 => n1588, ZN => n1587);
   U5190 : NAND2_X1 port map( A1 => n1590, A2 => n14264, ZN => n13615);
   U5191 : NAND2_X1 port map( A1 => n14267, A2 => n1742, ZN => n1590);
   U5192 : NAND2_X1 port map( A1 => n1743, A2 => n14260, ZN => n1742);
   U5194 : NAND2_X1 port map( A1 => n14099, A2 => n14259, ZN => n14267);
   U5197 : INV_X1 port map( A => n17025, ZN => n1594);
   U5198 : NAND2_X1 port map( A1 => n5420, A2 => n17025, ZN => n1595);
   U5200 : NAND2_X1 port map( A1 => n14659, A2 => n14658, ZN => n15018);
   U5201 : NAND2_X1 port map( A1 => n1598, A2 => n14467, ZN => n14659);
   U5202 : NAND2_X1 port map( A1 => n14185, A2 => n13933, ZN => n1599);
   U5203 : NAND2_X1 port map( A1 => n14466, A2 => n1600, ZN => n14658);
   U5204 : NAND2_X1 port map( A1 => n13933, A2 => n3843, ZN => n1600);
   U5205 : OR2_X1 port map( A1 => n14469, A2 => n14464, ZN => n3843);
   U5206 : NAND3_X1 port map( A1 => n527, A2 => n29044, A3 => n18087, ZN => 
                           n1601);
   U5207 : NAND3_X1 port map( A1 => n16843, A2 => n29125, A3 => n1603, ZN => 
                           n1602);
   U5208 : OR2_X1 port map( A1 => n18087, A2 => n18188, ZN => n1603);
   U5209 : NOR2_X1 port map( A1 => n19561, A2 => n18190, ZN => n18088);
   U5212 : NAND3_X1 port map( A1 => n7792, A2 => n1607, A3 => n7796, ZN => 
                           n1606);
   U5213 : INV_X1 port map( A => n7542, ZN => n1607);
   U5214 : OAI21_X1 port map( B1 => n7792, B2 => n7541, A => n8150, ZN => n1608
                           );
   U5215 : OAI211_X1 port map( C1 => n12063, C2 => n12289, A => n12062, B => 
                           n1610, ZN => n12697);
   U5216 : NAND3_X1 port map( A1 => n12060, A2 => n29498, A3 => n1611, ZN => 
                           n1610);
   U5217 : NAND3_X1 port map( A1 => n12058, A2 => n12061, A3 => n12290, ZN => 
                           n1611);
   U5219 : NAND3_X1 port map( A1 => n7839, A2 => n370, A3 => n7840, ZN => n1612
                           );
   U5220 : NAND2_X1 port map( A1 => n14604, A2 => n15515, ZN => n1613);
   U5221 : AOI21_X1 port map( B1 => n1616, B2 => n1615, A => n608, ZN => n1614)
                           ;
   U5222 : NAND2_X1 port map( A1 => n6147, A2 => n9014, ZN => n1616);
   U5223 : NAND2_X1 port map( A1 => n1617, A2 => n28401, ZN => n4860);
   U5225 : NAND2_X1 port map( A1 => n15731, A2 => n17232, ZN => n17045);
   U5226 : INV_X1 port map( A => n17362, ZN => n17232);
   U5228 : XNOR2_X1 port map( A => n19540, B => n18639, ZN => n1619);
   U5229 : NAND2_X1 port map( A1 => n8210, A2 => n8211, ZN => n1620);
   U5230 : OR2_X1 port map( A1 => n7836, A2 => n7839, ZN => n8211);
   U5231 : NAND3_X1 port map( A1 => n21551, A2 => n1621, A3 => n21177, ZN => 
                           n20930);
   U5232 : NAND2_X1 port map( A1 => n21552, A2 => n1621, ZN => n21522);
   U5233 : MUX2_X1 port map( A => n20351, B => n21551, S => n21549, Z => n20784
                           );
   U5236 : INV_X1 port map( A => n26480, ZN => n1623);
   U5237 : NOR2_X1 port map( A1 => n1624, A2 => n20504, ZN => n1625);
   U5238 : INV_X1 port map( A => n20506, ZN => n1624);
   U5240 : OAI21_X1 port map( B1 => n6605, B2 => n29601, A => n1626, ZN => 
                           n19150);
   U5241 : NAND3_X1 port map( A1 => n11963, A2 => n12219, A3 => n2846, ZN => 
                           n11535);
   U5242 : NAND2_X1 port map( A1 => n11963, A2 => n12219, ZN => n11697);
   U5243 : NAND3_X1 port map( A1 => n14466, A2 => n4840, A3 => n14467, ZN => 
                           n1629);
   U5245 : NOR2_X1 port map( A1 => n19791, A2 => n20486, ZN => n1804);
   U5248 : NAND2_X1 port map( A1 => n24746, A2 => n1632, ZN => n24266);
   U5249 : NAND2_X1 port map( A1 => n24617, A2 => n24747, ZN => n1632);
   U5250 : MUX2_X2 port map( A => n21726, B => n21727, S => n24747, Z => n25901
                           );
   U5251 : NAND3_X1 port map( A1 => n9034, A2 => n9035, A3 => n1634, ZN => 
                           n2502);
   U5253 : NAND3_X1 port map( A1 => n6472, A2 => n23739, A3 => n6474, ZN => 
                           n1638);
   U5255 : XNOR2_X1 port map( A => n22777, B => n1640, ZN => n21742);
   U5256 : OR2_X1 port map( A1 => n6081, A2 => n1642, ZN => n24687);
   U5257 : NAND2_X1 port map( A1 => n4118, A2 => n17569, ZN => n1643);
   U5258 : XNOR2_X2 port map( A => n15868, B => n16237, ZN => n17569);
   U5259 : AND2_X2 port map( A1 => n1646, A2 => n1645, ZN => n1644);
   U5260 : INV_X2 port map( A => n1644, ZN => n15434);
   U5261 : NAND2_X1 port map( A1 => n15027, A2 => n1644, ZN => n15028);
   U5262 : NAND2_X1 port map( A1 => n1644, A2 => n14821, ZN => n14683);
   U5263 : NAND3_X1 port map( A1 => n15032, A2 => n1644, A3 => n15031, ZN => 
                           n15033);
   U5264 : MUX2_X1 port map( A => n14823, B => n14822, S => n1644, Z => n14829)
                           ;
   U5265 : INV_X1 port map( A => n14014, ZN => n1645);
   U5266 : NAND2_X1 port map( A1 => n14015, A2 => n14351, ZN => n1646);
   U5267 : NAND2_X1 port map( A1 => n1648, A2 => n1647, ZN => n18373);
   U5268 : NAND2_X1 port map( A1 => n4412, A2 => n18333, ZN => n1647);
   U5269 : NAND2_X1 port map( A1 => n18371, A2 => n1650, ZN => n1648);
   U5270 : MUX2_X1 port map( A => n1650, B => n18370, S => n18337, Z => n18374)
                           ;
   U5271 : NAND2_X1 port map( A1 => n1649, A2 => n17061, ZN => n19096);
   U5272 : MUX2_X1 port map( A => n1651, B => n8485, S => n81, Z => n8489);
   U5273 : NAND3_X1 port map( A1 => n24457, A2 => n24777, A3 => n24775, ZN => 
                           n1654);
   U5274 : NAND2_X1 port map( A1 => n24212, A2 => n29597, ZN => n1652);
   U5275 : NAND2_X1 port map( A1 => n1655, A2 => n24480, ZN => n1653);
   U5276 : INV_X1 port map( A => n24211, ZN => n24480);
   U5277 : NAND2_X1 port map( A1 => n17258, A2 => n17259, ZN => n1658);
   U5278 : NAND2_X1 port map( A1 => n13717, A2 => n13900, ZN => n1659);
   U5279 : XNOR2_X1 port map( A => n6647, B => n1664, ZN => n12707);
   U5281 : AND3_X1 port map( A1 => n11971, A2 => n11972, A3 => n11973, ZN => 
                           n1663);
   U5282 : XNOR2_X1 port map( A => n12644, B => n1664, ZN => n12588);
   U5283 : XNOR2_X1 port map( A => n11975, B => n1664, ZN => n11988);
   U5284 : NAND2_X1 port map( A1 => n20368, A2 => n21581, ZN => n6694);
   U5285 : AOI21_X1 port map( B1 => n29737, B2 => n387, A => n1666, ZN => n1665
                           );
   U5286 : INV_X1 port map( A => n17464, ZN => n1666);
   U5287 : NAND2_X1 port map( A1 => n528, A2 => n17280, ZN => n1667);
   U5288 : NAND2_X1 port map( A1 => n11420, A2 => n1668, ZN => n1669);
   U5289 : NAND2_X1 port map( A1 => n1669, A2 => n3900, ZN => n11425);
   U5290 : NAND2_X1 port map( A1 => n8342, A2 => n9132, ZN => n8755);
   U5291 : INV_X1 port map( A => n1934, ZN => n8342);
   U5293 : OAI22_X1 port map( A1 => n14400, A2 => n28804, B1 => n13963, B2 => 
                           n29628, ZN => n1671);
   U5295 : NAND2_X1 port map( A1 => n21212, A2 => n28790, ZN => n1673);
   U5296 : NAND2_X1 port map( A1 => n5855, A2 => n22023, ZN => n1674);
   U5297 : XNOR2_X1 port map( A => n22783, B => n3317, ZN => n22785);
   U5298 : NAND3_X1 port map( A1 => n479, A2 => n28626, A3 => n483, ZN => n1675
                           );
   U5302 : AND2_X1 port map( A1 => n24204, A2 => n1679, ZN => n25321);
   U5303 : NAND2_X1 port map( A1 => n28561, A2 => n28547, ZN => n1679);
   U5306 : OAI21_X1 port map( B1 => n1683, B2 => n26498, A => n27372, ZN => 
                           n1681);
   U5308 : NOR2_X1 port map( A1 => n26497, A2 => n27364, ZN => n1683);
   U5309 : INV_X1 port map( A => n25995, ZN => n1684);
   U5310 : XNOR2_X1 port map( A => n16596, B => n16393, ZN => n16116);
   U5311 : OAI211_X2 port map( C1 => n14739, C2 => n5198, A => n5815, B => 
                           n1685, ZN => n16596);
   U5312 : NAND3_X1 port map( A1 => n15379, A2 => n15384, A3 => n2203, ZN => 
                           n1685);
   U5313 : INV_X1 port map( A => n12420, ZN => n12980);
   U5314 : XNOR2_X1 port map( A => n11432, B => n1686, ZN => n11445);
   U5315 : XNOR2_X1 port map( A => n1687, B => n12420, ZN => n1686);
   U5316 : INV_X1 port map( A => n13179, ZN => n1687);
   U5317 : XNOR2_X1 port map( A => n1688, B => n28108, ZN => Ciphertext(190));
   U5321 : NAND2_X1 port map( A1 => n1693, A2 => n489, ZN => n1692);
   U5322 : NAND2_X1 port map( A1 => n1695, A2 => n28790, ZN => n1694);
   U5323 : MUX2_X1 port map( A => n22286, B => n22290, S => n21211, Z => n1695)
                           ;
   U5325 : NAND2_X1 port map( A1 => n29294, A2 => n17179, ZN => n1697);
   U5328 : AOI21_X1 port map( B1 => n1698, B2 => n7628, A => n7914, ZN => n6999
                           );
   U5329 : NAND2_X1 port map( A1 => n7396, A2 => n1698, ZN => n1796);
   U5330 : NAND2_X1 port map( A1 => n7912, A2 => n7911, ZN => n1698);
   U5331 : INV_X1 port map( A => n28692, ZN => n1700);
   U5332 : OR2_X1 port map( A1 => n28608, A2 => n591, ZN => n10678);
   U5333 : NAND3_X1 port map( A1 => n5267, A2 => n5265, A3 => n391, ZN => 
                           n10950);
   U5334 : NAND3_X1 port map( A1 => n6368, A2 => n6367, A3 => n391, ZN => n6366
                           );
   U5336 : NAND3_X1 port map( A1 => n553, A2 => n15180, A3 => n15459, ZN => 
                           n1702);
   U5337 : INV_X1 port map( A => n15180, ZN => n15457);
   U5338 : NAND2_X1 port map( A1 => n1934, A2 => n9134, ZN => n8343);
   U5339 : NAND2_X1 port map( A1 => n1934, A2 => n9133, ZN => n9131);
   U5340 : NAND2_X1 port map( A1 => n8753, A2 => n1934, ZN => n7411);
   U5341 : NAND2_X1 port map( A1 => n7397, A2 => n1934, ZN => n7414);
   U5342 : NAND2_X1 port map( A1 => n11248, A2 => n29666, ZN => n1703);
   U5343 : NAND2_X1 port map( A1 => n3819, A2 => n1704, ZN => n3814);
   U5344 : NAND2_X1 port map( A1 => n1706, A2 => n12145, ZN => n11711);
   U5345 : AOI21_X1 port map( B1 => n1706, B2 => n11645, A => n11715, ZN => 
                           n11647);
   U5346 : OAI21_X1 port map( B1 => n12144, B2 => n1706, A => n1705, ZN => 
                           n5636);
   U5347 : NAND2_X1 port map( A1 => n12147, A2 => n1706, ZN => n1705);
   U5348 : NAND2_X1 port map( A1 => n1707, A2 => n11322, ZN => n6510);
   U5349 : NAND2_X1 port map( A1 => n11184, A2 => n1707, ZN => n8992);
   U5350 : NAND3_X1 port map( A1 => n11181, A2 => n10473, A3 => n1707, ZN => 
                           n3906);
   U5351 : INV_X1 port map( A => n10810, ZN => n1707);
   U5352 : AND2_X1 port map( A1 => n516, A2 => n18173, ZN => n5223);
   U5354 : OAI21_X1 port map( B1 => n17689, B2 => n4884, A => n1708, ZN => 
                           n16821);
   U5356 : OR2_X1 port map( A1 => n8484, A2 => n440, ZN => n1711);
   U5357 : NAND3_X1 port map( A1 => n1710, A2 => n1711, A3 => n1712, ZN => 
                           n1709);
   U5358 : NAND3_X1 port map( A1 => n8483, A2 => n8484, A3 => n440, ZN => n1712
                           );
   U5359 : NAND2_X1 port map( A1 => n4060, A2 => n610, ZN => n1715);
   U5360 : XNOR2_X1 port map( A => n10328, B => n625, ZN => n8902);
   U5361 : NAND2_X1 port map( A1 => n17896, A2 => n18322, ZN => n1718);
   U5362 : NAND2_X2 port map( A1 => n1721, A2 => n5999, ZN => n18261);
   U5364 : NAND2_X1 port map( A1 => n6417, A2 => n29138, ZN => n16906);
   U5366 : OAI22_X1 port map( A1 => n27758, A2 => n1724, B1 => n27740, B2 => 
                           n27741, ZN => n27743);
   U5367 : INV_X1 port map( A => n27229, ZN => n1724);
   U5368 : OR2_X1 port map( A1 => n27732, A2 => n27759, ZN => n27229);
   U5370 : NAND2_X1 port map( A1 => n1725, A2 => n14667, ZN => n14668);
   U5371 : INV_X1 port map( A => n15020, ZN => n1725);
   U5372 : AND2_X1 port map( A1 => n465, A2 => n24559, ZN => n23989);
   U5373 : OAI21_X1 port map( B1 => n24242, B2 => n1727, A => n1726, ZN => 
                           n24194);
   U5374 : INV_X1 port map( A => n24633, ZN => n1727);
   U5375 : NAND2_X1 port map( A1 => n402, A2 => n26837, ZN => n1728);
   U5377 : OAI211_X1 port map( C1 => n28631, C2 => n402, A => n27120, B => 
                           n1728, ZN => n2270);
   U5378 : NAND2_X1 port map( A1 => n3440, A2 => n3439, ZN => n1733);
   U5380 : NAND2_X1 port map( A1 => n1731, A2 => n3751, ZN => n1730);
   U5381 : XNOR2_X1 port map( A => n1783, B => n1732, ZN => n19036);
   U5382 : INV_X1 port map( A => n19320, ZN => n1732);
   U5383 : NAND2_X1 port map( A1 => n5563, A2 => n1734, ZN => n10533);
   U5384 : NOR2_X1 port map( A1 => n11290, A2 => n29116, ZN => n1735);
   U5385 : INV_X1 port map( A => n14240, ZN => n2714);
   U5386 : NAND2_X1 port map( A1 => n17615, A2 => n4217, ZN => n3250);
   U5387 : NAND2_X1 port map( A1 => n1738, A2 => n6002, ZN => n1737);
   U5389 : NAND2_X1 port map( A1 => n1739, A2 => n26228, ZN => n26233);
   U5390 : NAND2_X1 port map( A1 => n1740, A2 => n23648, ZN => n5555);
   U5391 : XNOR2_X1 port map( A => n1741, B => n3516, ZN => n18666);
   U5392 : XNOR2_X1 port map( A => n18912, B => n1741, ZN => n16696);
   U5393 : XNOR2_X1 port map( A => n18913, B => n1741, ZN => n19133);
   U5394 : INV_X1 port map( A => n14260, ZN => n13611);
   U5395 : INV_X1 port map( A => n14267, ZN => n13613);
   U5396 : INV_X1 port map( A => n14268, ZN => n1743);
   U5397 : NOR2_X1 port map( A1 => n1744, A2 => n14998, ZN => n15126);
   U5398 : NOR2_X1 port map( A1 => n1745, A2 => n15127, ZN => n13986);
   U5399 : NAND2_X1 port map( A1 => n1745, A2 => n15004, ZN => n14685);
   U5400 : NAND2_X1 port map( A1 => n14686, A2 => n1745, ZN => n14687);
   U5401 : NAND2_X1 port map( A1 => n1746, A2 => n12507, ZN => n10864);
   U5402 : NOR2_X1 port map( A1 => n577, A2 => n12508, ZN => n11989);
   U5404 : NAND3_X1 port map( A1 => n12512, A2 => n577, A3 => n1746, ZN => 
                           n11992);
   U5405 : NAND3_X1 port map( A1 => n1747, A2 => n10165, A3 => n10166, ZN => 
                           n10168);
   U5406 : NAND2_X1 port map( A1 => n10572, A2 => n10883, ZN => n1747);
   U5407 : NAND2_X1 port map( A1 => n15511, A2 => n15274, ZN => n15509);
   U5408 : MUX2_X1 port map( A => n14356, B => n14357, S => n4893, Z => n1749);
   U5410 : MUX2_X1 port map( A => n9243, B => n9041, S => n9247, Z => n1750);
   U5411 : XNOR2_X1 port map( A => n1751, B => n21847, ZN => n21852);
   U5412 : XNOR2_X1 port map( A => n21849, B => n21848, ZN => n1751);
   U5414 : NAND2_X1 port map( A1 => n1753, A2 => n1752, ZN => n5023);
   U5416 : NAND2_X1 port map( A1 => n17360, A2 => n17359, ZN => n1753);
   U5417 : XNOR2_X1 port map( A => n19231, B => n19227, ZN => n1756);
   U5419 : MUX2_X1 port map( A => n2853, B => n18430, S => n18431, Z => n1759);
   U5420 : AND2_X1 port map( A1 => n11068, A2 => n1760, ZN => n5063);
   U5421 : INV_X1 port map( A => n11067, ZN => n10880);
   U5422 : NAND2_X1 port map( A1 => n3189, A2 => n1762, ZN => n6049);
   U5423 : AOI21_X1 port map( B1 => n23680, B2 => n474, A => n28457, ZN => 
                           n1762);
   U5424 : INV_X1 port map( A => n12166, ZN => n12102);
   U5426 : NAND2_X1 port map( A1 => n21033, A2 => n21473, ZN => n1763);
   U5427 : NAND2_X1 port map( A1 => n1765, A2 => n493, ZN => n1764);
   U5428 : NAND2_X1 port map( A1 => n1766, A2 => n21472, ZN => n1765);
   U5429 : NAND2_X1 port map( A1 => n29314, A2 => n21736, ZN => n1766);
   U5430 : AND3_X2 port map( A1 => n3341, A2 => n2956, A3 => n19957, ZN => 
                           n21736);
   U5431 : NOR2_X1 port map( A1 => n9247, A2 => n28211, ZN => n6344);
   U5432 : NAND3_X1 port map( A1 => n9248, A2 => n28211, A3 => n1768, ZN => 
                           n9249);
   U5433 : INV_X1 port map( A => n9247, ZN => n1768);
   U5434 : INV_X1 port map( A => n9014, ZN => n1770);
   U5435 : NAND2_X1 port map( A1 => n9015, A2 => n9014, ZN => n1769);
   U5436 : OAI211_X2 port map( C1 => n9019, C2 => n5674, A => n9017, B => n1771
                           , ZN => n10362);
   U5437 : XNOR2_X1 port map( A => n22651, B => n1773, ZN => n1772);
   U5438 : OAI21_X1 port map( B1 => n1775, B2 => n27925, A => n1774, ZN => 
                           n27022);
   U5439 : NAND3_X1 port map( A1 => n27925, A2 => n27944, A3 => n27938, ZN => 
                           n1774);
   U5440 : AOI21_X2 port map( B1 => n1776, B2 => n11371, A => n1969, ZN => 
                           n14893);
   U5442 : XNOR2_X1 port map( A => n15975, B => n266, ZN => n1778);
   U5443 : NAND2_X1 port map( A1 => n17354, A2 => n17355, ZN => n1779);
   U5444 : XNOR2_X1 port map( A => n12420, B => n565, ZN => n1780);
   U5445 : NOR2_X1 port map( A1 => n505, A2 => n1781, ZN => n19963);
   U5446 : XNOR2_X1 port map( A => n18959, B => n1782, ZN => n18577);
   U5447 : XNOR2_X1 port map( A => n18959, B => n624, ZN => n18977);
   U5448 : XNOR2_X1 port map( A => n1783, B => n18959, ZN => n17982);
   U5449 : OAI21_X1 port map( B1 => n23604, B2 => n23606, A => n1785, ZN => 
                           n23249);
   U5450 : NAND2_X1 port map( A1 => n23607, A2 => n23606, ZN => n1785);
   U5452 : NAND2_X1 port map( A1 => n3455, A2 => n3453, ZN => n1787);
   U5453 : NAND2_X1 port map( A1 => n12251, A2 => n12252, ZN => n11934);
   U5454 : INV_X1 port map( A => n11934, ZN => n11020);
   U5455 : INV_X1 port map( A => n8760, ZN => n8569);
   U5456 : NAND3_X1 port map( A1 => n6747, A2 => n9374, A3 => n6072, ZN => 
                           n1791);
   U5457 : NAND2_X1 port map( A1 => n9148, A2 => n9149, ZN => n1788);
   U5459 : XNOR2_X2 port map( A => n13071, B => n13072, ZN => n4893);
   U5462 : AND2_X2 port map( A1 => n1797, A2 => n1796, ZN => n1934);
   U5463 : INV_X1 port map( A => n18101, ZN => n16717);
   U5464 : NAND2_X1 port map( A1 => n18193, A2 => n16718, ZN => n18101);
   U5466 : NAND2_X1 port map( A1 => n530, A2 => n29635, ZN => n1800);
   U5467 : NAND2_X1 port map( A1 => n16874, A2 => n17375, ZN => n1802);
   U5468 : NAND2_X1 port map( A1 => n8562, A2 => n9139, ZN => n1803);
   U5469 : NAND2_X1 port map( A1 => n29526, A2 => n21705, ZN => n19187);
   U5470 : OAI22_X2 port map( A1 => n1804, A2 => n20482, B1 => n20238, B2 => 
                           n19092, ZN => n21705);
   U5471 : NAND2_X1 port map( A1 => n5571, A2 => n1808, ZN => n24415);
   U5472 : OAI21_X1 port map( B1 => n24709, B2 => n1808, A => n24417, ZN => 
                           n1807);
   U5473 : NAND2_X1 port map( A1 => n24710, A2 => n1808, ZN => n5749);
   U5474 : AND2_X1 port map( A1 => n1809, A2 => n15171, ZN => n6925);
   U5475 : NAND2_X1 port map( A1 => n1810, A2 => n20276, ZN => n22657);
   U5476 : NAND2_X1 port map( A1 => n2666, A2 => n1810, ZN => n2665);
   U5478 : NAND2_X1 port map( A1 => n8242, A2 => n616, ZN => n3655);
   U5479 : OR2_X1 port map( A1 => n11038, A2 => n28612, ZN => n10671);
   U5480 : MUX2_X1 port map( A => n11273, B => n28147, S => n11038, Z => n10673
                           );
   U5481 : NOR2_X1 port map( A1 => n11039, A2 => n1811, ZN => n10846);
   U5482 : INV_X1 port map( A => n11038, ZN => n1811);
   U5484 : NAND3_X1 port map( A1 => n607, A2 => n602, A3 => n8594, ZN => n1813)
                           ;
   U5485 : INV_X1 port map( A => n21124, ZN => n1814);
   U5486 : AND2_X1 port map( A1 => n20842, A2 => n3838, ZN => n20844);
   U5487 : NAND2_X1 port map( A1 => n439, A2 => n7835, ZN => n8210);
   U5488 : MUX2_X1 port map( A => n15896, B => n15897, S => n15434, Z => n15898
                           );
   U5491 : NAND2_X1 port map( A1 => n16690, A2 => n534, ZN => n1817);
   U5492 : INV_X1 port map( A => n11085, ZN => n11212);
   U5493 : XNOR2_X1 port map( A => n1819, B => n2476, ZN => Ciphertext(28));
   U5494 : NAND2_X1 port map( A1 => n1622, A2 => n26485, ZN => n26486);
   U5496 : XNOR2_X1 port map( A => n19308, B => n4976, ZN => n1823);
   U5497 : XNOR2_X1 port map( A => n7068, B => Key(175), ZN => n7584);
   U5499 : XNOR2_X1 port map( A => n22647, B => n22648, ZN => n1829);
   U5500 : XNOR2_X1 port map( A => n22647, B => n22648, ZN => n23430);
   U5501 : INV_X1 port map( A => n14331, ZN => n1830);
   U5502 : OR2_X1 port map( A1 => n10546, A2 => n10545, ZN => n1831);
   U5504 : XNOR2_X1 port map( A => n9982, B => n9983, ZN => n1834);
   U5505 : INV_X1 port map( A => n20109, ZN => n1835);
   U5506 : INV_X1 port map( A => n578, ZN => n1836);
   U5507 : XNOR2_X1 port map( A => n5862, B => n22885, ZN => n1837);
   U5508 : NAND2_X1 port map( A1 => n19826, A2 => n19825, ZN => n20865);
   U5509 : AOI21_X1 port map( B1 => n10503, B2 => n10502, A => n3458, ZN => 
                           n11463);
   U5510 : XNOR2_X1 port map( A => n5862, B => n22885, ZN => n23145);
   U5512 : XNOR2_X1 port map( A => n22244, B => n22243, ZN => n1838);
   U5513 : XNOR2_X1 port map( A => n22244, B => n22243, ZN => n22992);
   U5514 : OAI211_X1 port map( C1 => n8761, C2 => n8760, A => n8759, B => n8758
                           , ZN => n10151);
   U5515 : INV_X1 port map( A => n21016, ZN => n1840);
   U5516 : INV_X1 port map( A => n14435, ZN => n1841);
   U5517 : NAND2_X1 port map( A1 => n7821, A2 => n7424, ZN => n1842);
   U5518 : AND2_X1 port map( A1 => n14834, A2 => n14833, ZN => n2456);
   U5519 : NAND2_X1 port map( A1 => n20016, A2 => n1844, ZN => n1845);
   U5520 : NAND2_X1 port map( A1 => n20015, A2 => n20014, ZN => n1846);
   U5521 : NAND2_X1 port map( A1 => n1845, A2 => n1846, ZN => n20669);
   U5522 : INV_X1 port map( A => n20014, ZN => n1844);
   U5525 : XNOR2_X1 port map( A => n2805, B => n21825, ZN => n22582);
   U5527 : INV_X1 port map( A => n15165, ZN => n1848);
   U5528 : AND2_X1 port map( A1 => n3844, A2 => n3846, ZN => n1849);
   U5531 : OAI211_X1 port map( C1 => n8882, C2 => n8881, A => n8880, B => n8879
                           , ZN => n1853);
   U5533 : XOR2_X1 port map( A => n10347, B => n10348, Z => n1855);
   U5537 : NAND2_X1 port map( A1 => n11713, A2 => n3174, ZN => n1857);
   U5538 : NAND2_X1 port map( A1 => n3407, A2 => n20692, ZN => n1858);
   U5539 : NAND2_X1 port map( A1 => n3407, A2 => n20692, ZN => n1859);
   U5541 : NAND2_X1 port map( A1 => n11713, A2 => n3174, ZN => n13269);
   U5544 : XOR2_X1 port map( A => n13005, B => n13260, Z => n12389);
   U5547 : OR2_X1 port map( A1 => n18061, A2 => n17931, ZN => n1863);
   U5549 : NAND4_X1 port map( A1 => n15933, A2 => n15932, A3 => n15934, A4 => 
                           n17404, ZN => n18057);
   U5550 : XNOR2_X1 port map( A => n4967, B => n4968, ZN => n23733);
   U5551 : OR2_X1 port map( A1 => n26419, A2 => n26914, ZN => n1864);
   U5552 : XNOR2_X1 port map( A => n3141, B => n5195, ZN => n1865);
   U5553 : OAI211_X1 port map( C1 => n8939, C2 => n9144, A => n8938, B => n8937
                           , ZN => n1868);
   U5556 : AOI21_X1 port map( B1 => n24004, B2 => n24547, A => n24003, ZN => 
                           n1871);
   U5557 : XNOR2_X1 port map( A => n6071, B => n25390, ZN => n1872);
   U5558 : XNOR2_X2 port map( A => n25400, B => n25401, ZN => n26914);
   U5559 : XNOR2_X1 port map( A => n3141, B => n5195, ZN => n10940);
   U5560 : OAI211_X1 port map( C1 => n8939, C2 => n9144, A => n8938, B => n8937
                           , ZN => n9894);
   U5562 : XNOR2_X1 port map( A => n6071, B => n25390, ZN => n26565);
   U5563 : INV_X1 port map( A => n23138, ZN => n1873);
   U5564 : AND2_X1 port map( A1 => n25597, A2 => n25654, ZN => n26742);
   U5565 : XNOR2_X1 port map( A => n25338, B => n25339, ZN => n1874);
   U5566 : OR2_X1 port map( A1 => n20337, A2 => n3144, ZN => n1875);
   U5567 : XNOR2_X1 port map( A => n12878, B => n12877, ZN => n1876);
   U5568 : AOI21_X1 port map( B1 => n8582, B2 => n8583, A => n8581, ZN => n1877
                           );
   U5569 : AOI21_X1 port map( B1 => n8582, B2 => n8583, A => n8581, ZN => n1878
                           );
   U5570 : XNOR2_X1 port map( A => n9445, B => n9444, ZN => n1879);
   U5571 : XNOR2_X1 port map( A => n12878, B => n12877, ZN => n14434);
   U5572 : AOI21_X1 port map( B1 => n8582, B2 => n8583, A => n8581, ZN => n9517
                           );
   U5573 : XNOR2_X1 port map( A => n19319, B => n19318, ZN => n20630);
   U5575 : NAND2_X1 port map( A1 => n6579, A2 => n5940, ZN => n1883);
   U5576 : OAI21_X1 port map( B1 => n9868, B2 => n12186, A => n9867, ZN => 
                           n1885);
   U5577 : NAND2_X1 port map( A1 => n6579, A2 => n5940, ZN => n23995);
   U5578 : AND2_X1 port map( A1 => n15691, A2 => n323, ZN => n1886);
   U5579 : BUF_X1 port map( A => n11247, Z => n12321);
   U5581 : XOR2_X1 port map( A => n18520, B => n19427, Z => n19234);
   U5582 : NAND3_X1 port map( A1 => n4623, A2 => n17550, A3 => n17551, ZN => 
                           n1888);
   U5585 : OAI211_X1 port map( C1 => n9065, C2 => n9064, A => n5537, B => n5536
                           , ZN => n1891);
   U5586 : OAI211_X1 port map( C1 => n9065, C2 => n9064, A => n5537, B => n5536
                           , ZN => n1892);
   U5587 : OAI211_X1 port map( C1 => n9065, C2 => n9064, A => n5537, B => n5536
                           , ZN => n9661);
   U5588 : AOI22_X1 port map( A1 => n6610, A2 => n23390, B1 => n6279, B2 => 
                           n23837, ZN => n1893);
   U5589 : INV_X1 port map( A => n18433, ZN => n1894);
   U5591 : XNOR2_X1 port map( A => n13253, B => n13252, ZN => n1896);
   U5592 : OR2_X1 port map( A1 => n6635, A2 => n19801, ZN => n1897);
   U5593 : XNOR2_X1 port map( A => n8706, B => n8707, ZN => n1898);
   U5594 : XNOR2_X1 port map( A => Key(21), B => Plaintext(21), ZN => n1899);
   U5595 : AOI22_X1 port map( A1 => n6610, A2 => n23390, B1 => n6279, B2 => 
                           n23837, ZN => n23393);
   U5596 : XNOR2_X1 port map( A => n8706, B => n8707, ZN => n10828);
   U5599 : XNOR2_X1 port map( A => n10175, B => n10174, ZN => n1900);
   U5600 : OR2_X1 port map( A1 => n1968, A2 => n26262, ZN => n1901);
   U5601 : NAND4_X1 port map( A1 => n7187, A2 => n7186, A3 => n7185, A4 => 
                           n7184, ZN => n1902);
   U5603 : NAND4_X1 port map( A1 => n13658, A2 => n13659, A3 => n13702, A4 => 
                           n13657, ZN => n1904);
   U5604 : NOR2_X1 port map( A1 => n11110, A2 => n11109, ZN => n1905);
   U5605 : NOR2_X1 port map( A1 => n11110, A2 => n11109, ZN => n1906);
   U5607 : INV_X1 port map( A => n498, ZN => n1908);
   U5608 : NAND4_X1 port map( A1 => n7187, A2 => n7186, A3 => n7185, A4 => 
                           n7184, ZN => n9542);
   U5609 : NAND4_X1 port map( A1 => n13658, A2 => n13659, A3 => n13702, A4 => 
                           n13657, ZN => n15119);
   U5610 : XNOR2_X1 port map( A => n24971, B => n24970, ZN => n26386);
   U5611 : XNOR2_X1 port map( A => n19401, B => n19400, ZN => n20637);
   U5613 : INV_X1 port map( A => n1914, ZN => n1913);
   U5615 : XNOR2_X1 port map( A => n19271, B => n19270, ZN => n1915);
   U5616 : XNOR2_X1 port map( A => n19271, B => n19270, ZN => n1916);
   U5617 : OAI21_X1 port map( B1 => n9155, B2 => n9154, A => n9153, ZN => n1917
                           );
   U5618 : OAI21_X1 port map( B1 => n9155, B2 => n9154, A => n9153, ZN => n1918
                           );
   U5619 : INV_X1 port map( A => n4861, ZN => n1919);
   U5620 : NOR2_X1 port map( A1 => n26355, A2 => n26354, ZN => n27629);
   U5621 : XNOR2_X1 port map( A => n21874, B => n21873, ZN => n4726);
   U5622 : OAI21_X1 port map( B1 => n9155, B2 => n9154, A => n9153, ZN => 
                           n10412);
   U5624 : INV_X1 port map( A => n20886, ZN => n1921);
   U5625 : OAI21_X1 port map( B1 => n23879, B2 => n23878, A => n23877, ZN => 
                           n1922);
   U5627 : OAI21_X1 port map( B1 => n23879, B2 => n23878, A => n23877, ZN => 
                           n25107);
   U5629 : XNOR2_X1 port map( A => n6717, B => n19018, ZN => n20354);
   U5631 : XNOR2_X1 port map( A => n9982, B => n9983, ZN => n10498);
   U5635 : XNOR2_X1 port map( A => n9667, B => n9666, ZN => n10853);
   U5637 : XNOR2_X1 port map( A => n13253, B => n13252, ZN => n14047);
   U5638 : XNOR2_X1 port map( A => n24088, B => n24089, ZN => n26186);
   U5639 : OR2_X1 port map( A1 => n8033, A2 => n8032, ZN => n4061);
   U5640 : AOI21_X1 port map( B1 => n7424, B2 => n7697, A => n7824, ZN => n7698
                           );
   U5641 : OR2_X1 port map( A1 => n4552, A2 => n7827, ZN => n4550);
   U5642 : OR2_X1 port map( A1 => n7856, A2 => n617, ZN => n7857);
   U5643 : INV_X1 port map( A => n8910, ZN => n5674);
   U5644 : XNOR2_X1 port map( A => n10137, B => n10294, ZN => n9736);
   U5646 : XNOR2_X1 port map( A => n10382, B => n5896, ZN => n5895);
   U5647 : AND2_X1 port map( A1 => n10860, A2 => n10859, ZN => n3570);
   U5648 : AOI22_X1 port map( A1 => n5753, A2 => n2680, B1 => n4591, B2 => 
                           n11165, ZN => n2678);
   U5649 : AND2_X1 port map( A1 => n5526, A2 => n11806, ZN => n5525);
   U5651 : XNOR2_X1 port map( A => n13291, B => n12776, ZN => n13513);
   U5652 : XNOR2_X1 port map( A => n13218, B => n6821, ZN => n6819);
   U5653 : XNOR2_X1 port map( A => n13219, B => n1196, ZN => n6821);
   U5654 : INV_X1 port map( A => n13674, ZN => n14492);
   U5655 : INV_X1 port map( A => n14434, ZN => n14437);
   U5656 : XNOR2_X1 port map( A => n13194, B => n13193, ZN => n13793);
   U5657 : INV_X1 port map( A => n13943, ZN => n15199);
   U5658 : OR2_X1 port map( A1 => n14070, A2 => n3798, ZN => n3175);
   U5659 : INV_X1 port map( A => n14616, ZN => n6797);
   U5660 : OR2_X1 port map( A1 => n5678, A2 => n14916, ZN => n14502);
   U5661 : NOR2_X1 port map( A1 => n17259, A2 => n29574, ZN => n16853);
   U5662 : INV_X1 port map( A => n17659, ZN => n18317);
   U5663 : NOR2_X1 port map( A1 => n18313, A2 => n18314, ZN => n18318);
   U5664 : OR2_X1 port map( A1 => n524, A2 => n2558, ZN => n17777);
   U5665 : OAI211_X1 port map( C1 => n18490, C2 => n18491, A => n18487, B => 
                           n3826, ZN => n3825);
   U5666 : XNOR2_X1 port map( A => n3222, B => n22697, ZN => n21826);
   U5667 : OAI211_X1 port map( C1 => n7165, C2 => n7279, A => n5282, B => n2692
                           , ZN => n7175);
   U5669 : OR2_X1 port map( A1 => n7533, A2 => n8014, ZN => n8018);
   U5670 : XNOR2_X1 port map( A => n6977, B => Key(101), ZN => n7830);
   U5671 : NOR2_X1 port map( A1 => n7657, A2 => n8304, ZN => n7207);
   U5672 : INV_X1 port map( A => n29317, ZN => n8297);
   U5673 : INV_X1 port map( A => n7692, ZN => n8243);
   U5674 : OR2_X1 port map( A1 => n7690, A2 => n7376, ZN => n3511);
   U5676 : OR2_X1 port map( A1 => n8927, A2 => n9132, ZN => n3101);
   U5678 : XNOR2_X1 port map( A => n4508, B => n4507, ZN => n4505);
   U5679 : XNOR2_X1 port map( A => n9714, B => n6916, ZN => n10620);
   U5680 : OR2_X1 port map( A1 => n6272, A2 => n11198, ZN => n4710);
   U5682 : AND3_X1 port map( A1 => n3046, A2 => n3047, A3 => n11282, ZN => 
                           n10653);
   U5683 : OR2_X1 port map( A1 => n11583, A2 => n10869, ZN => n6328);
   U5684 : NAND2_X1 port map( A1 => n11813, A2 => n11814, ZN => n12985);
   U5685 : NOR2_X1 port map( A1 => n11809, A2 => n11982, ZN => n4021);
   U5686 : OR2_X1 port map( A1 => n14426, A2 => n12534, ZN => n13871);
   U5687 : NOR2_X1 port map( A1 => n4046, A2 => n6482, ZN => n6481);
   U5688 : OR2_X1 port map( A1 => n11714, A2 => n11715, ZN => n3174);
   U5689 : XNOR2_X1 port map( A => n5122, B => n4041, ZN => n14440);
   U5690 : XNOR2_X1 port map( A => n12778, B => n12779, ZN => n14494);
   U5691 : XNOR2_X1 port map( A => n6895, B => n12584, ZN => n14309);
   U5692 : INV_X1 port map( A => n13257, ZN => n14312);
   U5693 : INV_X1 port map( A => n14106, ZN => n14231);
   U5694 : INV_X1 port map( A => n14440, ZN => n14432);
   U5695 : OR2_X1 port map( A1 => n14379, A2 => n4258, ZN => n14384);
   U5696 : INV_X1 port map( A => n15402, ZN => n14943);
   U5697 : OR2_X1 port map( A1 => n6699, A2 => n15503, ZN => n15267);
   U5698 : OR2_X1 port map( A1 => n15077, A2 => n15073, ZN => n14569);
   U5699 : AND2_X1 port map( A1 => n15511, A2 => n15275, ZN => n15279);
   U5701 : NAND2_X1 port map( A1 => n13601, A2 => n5024, ZN => n16477);
   U5702 : AND2_X1 port map( A1 => n4288, A2 => n4287, ZN => n6080);
   U5703 : AOI22_X1 port map( A1 => n3841, A2 => n3784, B1 => n426, B2 => n3840
                           , ZN => n4324);
   U5704 : INV_X1 port map( A => n4493, ZN => n15862);
   U5705 : XNOR2_X1 port map( A => n15212, B => n3792, ZN => n15745);
   U5706 : INV_X1 port map( A => n17710, ZN => n4156);
   U5707 : OR2_X1 port map( A1 => n15154, A2 => n15155, ZN => n5196);
   U5708 : OR2_X1 port map( A1 => n17190, A2 => n424, ZN => n4241);
   U5709 : INV_X1 port map( A => n4687, ZN => n17124);
   U5712 : AND2_X1 port map( A1 => n6337, A2 => n6336, ZN => n3529);
   U5713 : INV_X1 port map( A => n18106, ZN => n17903);
   U5715 : OAI21_X1 port map( B1 => n2707, B2 => n18537, A => n17699, ZN => 
                           n2704);
   U5717 : XNOR2_X1 port map( A => n19701, B => n18638, ZN => n2993);
   U5719 : INV_X1 port map( A => n20205, ZN => n4340);
   U5720 : XNOR2_X1 port map( A => n19465, B => n18653, ZN => n18815);
   U5721 : OR2_X1 port map( A1 => n17761, A2 => n525, ZN => n5417);
   U5722 : INV_X1 port map( A => n19480, ZN => n4976);
   U5723 : XNOR2_X1 port map( A => n19273, B => n19535, ZN => n19084);
   U5724 : AND2_X1 port map( A1 => n19938, A2 => n506, ZN => n2487);
   U5725 : XNOR2_X1 port map( A => n19483, B => n19085, ZN => n19634);
   U5727 : OAI21_X1 port map( B1 => n18406, B2 => n5021, A => n18706, ZN => 
                           n17778);
   U5728 : OR2_X1 port map( A1 => n17862, A2 => n18516, ZN => n17863);
   U5730 : INV_X1 port map( A => n4569, ZN => n4306);
   U5731 : AOI21_X1 port map( B1 => n20404, B2 => n20549, A => n3747, ZN => 
                           n19857);
   U5732 : AND2_X1 port map( A1 => n20551, A2 => n20405, ZN => n3747);
   U5733 : OR2_X1 port map( A1 => n20401, A2 => n5680, ZN => n20566);
   U5734 : XNOR2_X1 port map( A => n19479, B => n19478, ZN => n20133);
   U5735 : XNOR2_X1 port map( A => n4030, B => n19492, ZN => n19493);
   U5737 : INV_X1 port map( A => n23642, ZN => n2138);
   U5738 : XNOR2_X1 port map( A => n22231, B => n22230, ZN => n23177);
   U5739 : INV_X1 port map( A => n23102, ZN => n22686);
   U5744 : INV_X1 port map( A => n23227, ZN => n23399);
   U5745 : INV_X1 port map( A => n23289, ZN => n4950);
   U5746 : XNOR2_X1 port map( A => n6017, B => n21988, ZN => n21989);
   U5748 : INV_X1 port map( A => n23702, ZN => n6099);
   U5749 : XNOR2_X1 port map( A => n22588, B => n22587, ZN => n22592);
   U5750 : OR2_X1 port map( A1 => n23770, A2 => n23769, ZN => n6355);
   U5751 : OR2_X1 port map( A1 => n4561, A2 => n23611, ZN => n4560);
   U5752 : AOI21_X1 port map( B1 => n4336, B2 => n23803, A => n2004, ZN => 
                           n2835);
   U5753 : XNOR2_X1 port map( A => n25738, B => n25921, ZN => n25563);
   U5754 : INV_X1 port map( A => n7584, ZN => n7885);
   U5755 : OR2_X1 port map( A1 => n8141, A2 => n7560, ZN => n7565);
   U5756 : OR2_X1 port map( A1 => n7840, A2 => n7836, ZN => n7368);
   U5757 : OR2_X1 port map( A1 => n6209, A2 => n7506, ZN => n7133);
   U5758 : OR2_X1 port map( A1 => n7912, A2 => n7911, ZN => n8286);
   U5759 : OR2_X1 port map( A1 => n8018, A2 => n28161, ZN => n6807);
   U5762 : OR2_X1 port map( A1 => n8716, A2 => n8786, ZN => n7607);
   U5765 : INV_X1 port map( A => n8073, ZN => n9100);
   U5766 : OR2_X1 port map( A1 => n9026, A2 => n9228, ZN => n3675);
   U5767 : INV_X1 port map( A => n10087, ZN => n10009);
   U5768 : AND2_X1 port map( A1 => n8974, A2 => n8819, ZN => n6689);
   U5770 : OR2_X1 port map( A1 => n9398, A2 => n8983, ZN => n3139);
   U5771 : INV_X1 port map( A => n10251, ZN => n5995);
   U5772 : XNOR2_X1 port map( A => n9626, B => n9754, ZN => n9683);
   U5773 : INV_X1 port map( A => n11123, ZN => n11118);
   U5774 : INV_X1 port map( A => n9590, ZN => n4807);
   U5775 : NOR2_X1 port map( A1 => n9034, A2 => n8792, ZN => n6860);
   U5776 : AND2_X1 port map( A1 => n8330, A2 => n9144, ZN => n2335);
   U5777 : XNOR2_X1 port map( A => n10228, B => n10184, ZN => n10046);
   U5778 : INV_X1 port map( A => n8742, ZN => n2908);
   U5779 : INV_X1 port map( A => n11144, ZN => n10806);
   U5780 : XNOR2_X1 port map( A => n8063, B => n8062, ZN => n11149);
   U5781 : XNOR2_X1 port map( A => n10206, B => n10205, ZN => n11240);
   U5782 : OAI21_X1 port map( B1 => n12132, B2 => n12266, A => n12267, ZN => 
                           n5964);
   U5783 : INV_X1 port map( A => n12504, ZN => n12867);
   U5784 : OR2_X1 port map( A1 => n6282, A2 => n6281, ZN => n6280);
   U5785 : OR2_X1 port map( A1 => n12151, A2 => n11856, ZN => n3796);
   U5786 : OR2_X1 port map( A1 => n10771, A2 => n567, ZN => n2538);
   U5787 : OAI21_X1 port map( B1 => n11879, B2 => n11876, A => n11582, ZN => 
                           n6561);
   U5789 : NOR2_X1 port map( A1 => n11297, A2 => n3558, ZN => n3557);
   U5790 : OR2_X1 port map( A1 => n11837, A2 => n3653, ZN => n3646);
   U5791 : XNOR2_X1 port map( A => n12738, B => n12632, ZN => n13220);
   U5792 : OR2_X1 port map( A1 => n569, A2 => n10701, ZN => n2217);
   U5793 : INV_X1 port map( A => n14126, ZN => n4897);
   U5794 : OR2_X1 port map( A1 => n29089, A2 => n13589, ZN => n2144);
   U5795 : XNOR2_X1 port map( A => n6052, B => n13439, ZN => n14373);
   U5796 : XNOR2_X1 port map( A => n13438, B => n13437, ZN => n6052);
   U5799 : XNOR2_X1 port map( A => n12419, B => n12418, ZN => n14398);
   U5800 : XNOR2_X1 port map( A => n12757, B => n12756, ZN => n14464);
   U5801 : INV_X1 port map( A => n16090, ZN => n16282);
   U5802 : XNOR2_X1 port map( A => n11203, B => n11202, ZN => n14106);
   U5804 : OR2_X1 port map( A1 => n13871, A2 => n13706, ZN => n3435);
   U5805 : XNOR2_X1 port map( A => n12375, B => n12376, ZN => n14408);
   U5806 : INV_X1 port map( A => n13877, ZN => n4509);
   U5807 : XNOR2_X1 port map( A => n2172, B => n13462, ZN => n2171);
   U5808 : XNOR2_X1 port map( A => n6297, B => n6298, ZN => n2173);
   U5811 : XNOR2_X1 port map( A => n13273, B => n4501, ZN => n11543);
   U5812 : OR2_X1 port map( A1 => n5531, A2 => n13730, ZN => n3799);
   U5813 : OR2_X1 port map( A1 => n14321, A2 => n14320, ZN => n6794);
   U5814 : OR3_X1 port map( A1 => n29306, A2 => n14165, A3 => n14481, ZN => 
                           n3408);
   U5815 : INV_X1 port map( A => n16567, ZN => n15723);
   U5816 : INV_X1 port map( A => n15135, ZN => n15252);
   U5817 : OR2_X1 port map( A1 => n15025, A2 => n15444, ZN => n4491);
   U5818 : AND2_X1 port map( A1 => n14111, A2 => n2727, ZN => n2726);
   U5819 : AND2_X1 port map( A1 => n14484, A2 => n14166, ZN => n4074);
   U5820 : OR2_X1 port map( A1 => n14896, A2 => n5025, ZN => n6851);
   U5821 : XNOR2_X1 port map( A => n4765, B => n4766, ZN => n17315);
   U5822 : INV_X1 port map( A => n17492, ZN => n17496);
   U5823 : INV_X1 port map( A => n14846, ZN => n5614);
   U5824 : OR2_X1 port map( A1 => n15091, A2 => n15090, ZN => n3022);
   U5825 : INV_X1 port map( A => n16937, ZN => n17340);
   U5827 : XNOR2_X1 port map( A => n15817, B => n15790, ZN => n5621);
   U5829 : XNOR2_X1 port map( A => n16012, B => n15977, ZN => n16224);
   U5830 : XNOR2_X1 port map( A => n14561, B => n14562, ZN => n17269);
   U5832 : NOR2_X1 port map( A1 => n28768, A2 => n17012, ZN => n17423);
   U5833 : XNOR2_X1 port map( A => n15575, B => n6319, ZN => n15577);
   U5834 : OR2_X1 port map( A1 => n17469, A2 => n17516, ZN => n2610);
   U5835 : XNOR2_X1 port map( A => n16050, B => n259, ZN => n4588);
   U5836 : INV_X1 port map( A => n16918, ZN => n17314);
   U5837 : XNOR2_X1 port map( A => n15883, B => n15882, ZN => n17567);
   U5838 : INV_X1 port map( A => n17484, ZN => n4271);
   U5840 : XNOR2_X1 port map( A => n2671, B => n16610, ZN => n17110);
   U5841 : XNOR2_X1 port map( A => n1977, B => n16140, ZN => n2671);
   U5842 : XNOR2_X1 port map( A => n16090, B => n5892, ZN => n13926);
   U5843 : AND2_X1 port map( A1 => n29406, A2 => n17110, ZN => n17473);
   U5844 : OR2_X1 port map( A1 => n17570, A2 => n423, ZN => n4157);
   U5845 : XNOR2_X1 port map( A => n6870, B => n6869, ZN => n17143);
   U5846 : AND2_X1 port map( A1 => n17528, A2 => n16706, ZN => n6161);
   U5847 : XNOR2_X1 port map( A => n15860, B => n15861, ZN => n4316);
   U5848 : INV_X1 port map( A => n17355, ZN => n4283);
   U5850 : INV_X1 port map( A => n17553, ZN => n16913);
   U5851 : INV_X1 port map( A => n17524, ZN => n4979);
   U5853 : INV_X1 port map( A => n17361, ZN => n17046);
   U5854 : OR2_X1 port map( A1 => n17546, A2 => n211, ZN => n2375);
   U5855 : INV_X1 port map( A => n18035, ZN => n2500);
   U5856 : XNOR2_X1 port map( A => n19445, B => n3255, ZN => n4339);
   U5857 : XNOR2_X1 port map( A => n18691, B => n4029, ZN => n3255);
   U5858 : INV_X1 port map( A => n20221, ZN => n20168);
   U5859 : XNOR2_X1 port map( A => n17334, B => n17333, ZN => n20406);
   U5860 : INV_X1 port map( A => n20547, ZN => n6261);
   U5861 : INV_X1 port map( A => n21092, ZN => n20145);
   U5862 : XNOR2_X1 port map( A => n19648, B => n19649, ZN => n20282);
   U5863 : INV_X1 port map( A => n20475, ZN => n5408);
   U5864 : INV_X1 port map( A => n415, ZN => n5935);
   U5865 : XNOR2_X1 port map( A => n19633, B => n6535, ZN => n6534);
   U5866 : BUF_X1 port map( A => n20176, Z => n20171);
   U5868 : AND2_X1 port map( A1 => n28658, A2 => n29145, ZN => n20084);
   U5869 : NOR2_X1 port map( A1 => n20176, A2 => n6114, ZN => n19052);
   U5870 : OR2_X1 port map( A1 => n20099, A2 => n18887, ZN => n20042);
   U5871 : AND2_X1 port map( A1 => n5056, A2 => n20099, ZN => n2715);
   U5872 : INV_X1 port map( A => n29146, ZN => n18837);
   U5873 : INV_X1 port map( A => n20334, ZN => n20005);
   U5874 : INV_X1 port map( A => n20406, ZN => n20556);
   U5875 : XNOR2_X1 port map( A => n16869, B => n5062, ZN => n16870);
   U5876 : XNOR2_X1 port map( A => n5539, B => n5538, ZN => n20319);
   U5877 : AND2_X1 port map( A1 => n20388, A2 => n20539, ZN => n19958);
   U5878 : OR2_X1 port map( A1 => n19820, A2 => n20539, ZN => n19959);
   U5879 : AND2_X1 port map( A1 => n20293, A2 => n20125, ZN => n19973);
   U5880 : INV_X1 port map( A => n20039, ZN => n20087);
   U5881 : XNOR2_X1 port map( A => n18734, B => n18733, ZN => n2735);
   U5882 : XNOR2_X1 port map( A => n4838, B => n4030, ZN => n6701);
   U5884 : OAI21_X1 port map( B1 => n20444, B2 => n3247, A => n3246, ZN => 
                           n20448);
   U5885 : INV_X1 port map( A => n4567, ZN => n4570);
   U5886 : OR2_X1 port map( A1 => n20153, A2 => n28188, ZN => n5034);
   U5887 : INV_X1 port map( A => n22386, ZN => n21325);
   U5889 : INV_X1 port map( A => n3838, ZN => n20841);
   U5891 : XNOR2_X1 port map( A => n6837, B => n6836, ZN => n23637);
   U5892 : XNOR2_X1 port map( A => n22572, B => n22573, ZN => n23827);
   U5893 : XNOR2_X1 port map( A => n21386, B => n21385, ZN => n23338);
   U5894 : XNOR2_X1 port map( A => n21911, B => n21910, ZN => n23492);
   U5895 : OR2_X1 port map( A1 => n23149, A2 => n23461, ZN => n4892);
   U5896 : INV_X1 port map( A => n23493, ZN => n6608);
   U5898 : OR2_X1 port map( A1 => n23741, A2 => n22944, ZN => n3149);
   U5899 : INV_X1 port map( A => n23564, ZN => n22995);
   U5900 : INV_X1 port map( A => n4003, ZN => n23761);
   U5903 : INV_X1 port map( A => n23637, ZN => n23557);
   U5904 : INV_X1 port map( A => n2141, ZN => n23397);
   U5905 : OAI21_X1 port map( B1 => n4256, B2 => n4255, A => n22996, ZN => 
                           n4254);
   U5906 : OR2_X1 port map( A1 => n23646, A2 => n23645, ZN => n3723);
   U5907 : NOR2_X1 port map( A1 => n23529, A2 => n23531, ZN => n5482);
   U5908 : NAND2_X1 port map( A1 => n23677, A2 => n3901, ZN => n24808);
   U5909 : OR2_X1 port map( A1 => n23360, A2 => n23673, ZN => n2575);
   U5910 : AOI21_X1 port map( B1 => n6267, B2 => n24404, A => n24405, ZN => 
                           n23306);
   U5911 : INV_X1 port map( A => n3797, ZN => n6267);
   U5912 : INV_X1 port map( A => n6110, ZN => n25179);
   U5913 : XNOR2_X1 port map( A => n25398, B => n25249, ZN => n25069);
   U5915 : XNOR2_X1 port map( A => n25907, B => n25906, ZN => n26510);
   U5916 : XNOR2_X1 port map( A => n3837, B => n25191, ZN => n25915);
   U5917 : NAND2_X1 port map( A1 => n24150, A2 => n5922, ZN => n25546);
   U5918 : OAI22_X1 port map( A1 => n5137, A2 => n5138, B1 => n24612, B2 => 
                           n24611, ZN => n5136);
   U5919 : NAND2_X1 port map( A1 => n24614, A2 => n29109, ZN => n5138);
   U5920 : XNOR2_X1 port map( A => n23244, B => n23243, ZN => n23862);
   U5921 : INV_X1 port map( A => n25418, ZN => n26792);
   U5922 : INV_X1 port map( A => n26278, ZN => n26798);
   U5923 : XNOR2_X1 port map( A => n24923, B => n24925, ZN => n5754);
   U5924 : OR2_X1 port map( A1 => n26868, A2 => n27110, ZN => n26310);
   U5926 : AND2_X1 port map( A1 => n7162, A2 => n7320, ZN => n7279);
   U5927 : OR2_X1 port map( A1 => n7865, A2 => n7308, ZN => n3664);
   U5928 : OR2_X1 port map( A1 => n7787, A2 => n7330, ZN => n7293);
   U5929 : INV_X1 port map( A => n7591, ZN => n7957);
   U5931 : OAI21_X1 port map( B1 => n7303, B2 => n7305, A => n7237, ZN => n5173
                           );
   U5932 : OR2_X1 port map( A1 => n8525, A2 => n8687, ZN => n9223);
   U5933 : NAND2_X1 port map( A1 => n6316, A2 => n8898, ZN => n6318);
   U5934 : OAI21_X1 port map( B1 => n8840, B2 => n8839, A => n8961, ZN => n3182
                           );
   U5935 : OR2_X1 port map( A1 => n8842, A2 => n605, ZN => n3181);
   U5936 : INV_X1 port map( A => n10372, ZN => n10201);
   U5937 : OR2_X1 port map( A1 => n8762, A2 => n9566, ZN => n7273);
   U5938 : INV_X1 port map( A => n8472, ZN => n6662);
   U5940 : OAI21_X1 port map( B1 => n6344, B2 => n9042, A => n8110, ZN => n7159
                           );
   U5943 : XNOR2_X1 port map( A => n9786, B => n9785, ZN => n5984);
   U5944 : XNOR2_X1 port map( A => n8649, B => n10334, ZN => n11144);
   U5945 : XNOR2_X1 port map( A => n9639, B => n10426, ZN => n10189);
   U5946 : XNOR2_X1 port map( A => n10265, B => n10302, ZN => n9961);
   U5947 : AND2_X1 port map( A1 => n7413, A2 => n7411, ZN => n2676);
   U5948 : OR2_X1 port map( A1 => n8407, A2 => n3297, ZN => n3296);
   U5949 : XNOR2_X1 port map( A => n10007, B => n4714, ZN => n10424);
   U5950 : OR2_X1 port map( A1 => n9224, A2 => n8685, ZN => n5959);
   U5951 : OR2_X1 port map( A1 => n8802, A2 => n8801, ZN => n8803);
   U5952 : INV_X1 port map( A => n11335, ZN => n11341);
   U5954 : NOR2_X1 port map( A1 => n3804, A2 => n10989, ZN => n3803);
   U5955 : AND2_X1 port map( A1 => n10775, A2 => n6108, ZN => n5706);
   U5956 : XNOR2_X1 port map( A => n9683, B => n10027, ZN => n4589);
   U5957 : INV_X1 port map( A => n11056, ZN => n10851);
   U5958 : INV_X1 port map( A => n11350, ZN => n3161);
   U5959 : INV_X1 port map( A => n333, ZN => n6816);
   U5960 : OR2_X1 port map( A1 => n10911, A2 => n10913, ZN => n5904);
   U5961 : XNOR2_X1 port map( A => n9811, B => n9887, ZN => n2662);
   U5962 : INV_X1 port map( A => n11090, ZN => n5277);
   U5963 : XNOR2_X1 port map( A => n6133, B => n6135, ZN => n11022);
   U5964 : XNOR2_X1 port map( A => n5414, B => n5413, ZN => n10937);
   U5965 : XNOR2_X1 port map( A => n9683, B => n9416, ZN => n5413);
   U5966 : XNOR2_X1 port map( A => n5411, B => n5410, ZN => n5414);
   U5967 : INV_X1 port map( A => n10936, ZN => n11002);
   U5968 : INV_X1 port map( A => n10620, ZN => n11099);
   U5969 : OR2_X1 port map( A1 => n11056, A2 => n10855, ZN => n10856);
   U5970 : OR2_X1 port map( A1 => n591, A2 => n2211, ZN => n2210);
   U5972 : XNOR2_X1 port map( A => n9350, B => n10046, ZN => n5860);
   U5973 : INV_X1 port map( A => n6108, ZN => n5710);
   U5974 : AND2_X1 port map( A1 => n11933, A2 => n12070, ZN => n11595);
   U5975 : INV_X1 port map( A => n12559, ZN => n13034);
   U5976 : XNOR2_X1 port map( A => n12377, B => n4277, ZN => n12379);
   U5977 : INV_X1 port map( A => n12788, ZN => n4277);
   U5978 : OR2_X1 port map( A1 => n12080, A2 => n29499, ZN => n5715);
   U5979 : INV_X1 port map( A => n285, ZN => n12322);
   U5981 : INV_X1 port map( A => n12472, ZN => n13231);
   U5982 : INV_X1 port map( A => n12236, ZN => n11979);
   U5985 : AND2_X1 port map( A1 => n12330, A2 => n6431, ZN => n3281);
   U5986 : OR2_X1 port map( A1 => n12003, A2 => n12004, ZN => n2603);
   U5987 : INV_X1 port map( A => n13538, ZN => n12885);
   U5988 : XNOR2_X1 port map( A => n12542, B => n13493, ZN => n13315);
   U5989 : XNOR2_X1 port map( A => n13406, B => n13538, ZN => n13027);
   U5990 : INV_X1 port map( A => n13872, ZN => n14428);
   U5992 : INV_X1 port map( A => n11676, ZN => n11674);
   U5994 : XNOR2_X1 port map( A => n12658, B => n12723, ZN => n13243);
   U5998 : OR2_X1 port map( A1 => n6581, A2 => n28201, ZN => n6519);
   U5999 : INV_X1 port map( A => n12978, ZN => n4375);
   U6000 : INV_X1 port map( A => n28805, ZN => n4433);
   U6001 : NOR2_X1 port map( A1 => n14475, A2 => n13936, ZN => n14473);
   U6002 : OR2_X1 port map( A1 => n14480, A2 => n14157, ZN => n13847);
   U6003 : XNOR2_X1 port map( A => n4199, B => n4198, ZN => n14487);
   U6004 : XNOR2_X1 port map( A => n4200, B => n12065, ZN => n4199);
   U6005 : XNOR2_X1 port map( A => n12064, B => n2916, ZN => n4200);
   U6006 : INV_X1 port map( A => n14450, ZN => n2972);
   U6007 : XNOR2_X1 port map( A => n11669, B => n3870, ZN => n5805);
   U6008 : AOI21_X1 port map( B1 => n14232, B2 => n14102, A => n4054, ZN => 
                           n14104);
   U6009 : AND2_X1 port map( A1 => n4056, A2 => n14106, ZN => n2608);
   U6010 : INV_X1 port map( A => n15431, ZN => n15031);
   U6012 : XNOR2_X1 port map( A => n13338, B => n2570, ZN => n11838);
   U6013 : XNOR2_X1 port map( A => n4474, B => n13035, ZN => n2570);
   U6014 : OR2_X1 port map( A1 => n15494, A2 => n14702, ZN => n6246);
   U6015 : XNOR2_X1 port map( A => n12635, B => n12636, ZN => n14177);
   U6016 : OR2_X1 port map( A1 => n14498, A2 => n29036, ZN => n13973);
   U6017 : XNOR2_X1 port map( A => n12963, B => n12964, ZN => n14123);
   U6019 : AND2_X1 port map( A1 => n15053, A2 => n15261, ZN => n2161);
   U6020 : INV_X1 port map( A => n15310, ZN => n15315);
   U6021 : NOR2_X1 port map( A1 => n4088, A2 => n4897, ZN => n4896);
   U6022 : AND2_X1 port map( A1 => n14262, A2 => n14259, ZN => n13747);
   U6025 : INV_X1 port map( A => n15515, ZN => n6293);
   U6026 : OAI211_X1 port map( C1 => n15249, C2 => n15247, A => n13715, B => 
                           n13714, ZN => n16126);
   U6027 : OR2_X1 port map( A1 => n15053, A2 => n14761, ZN => n6391);
   U6028 : INV_X1 port map( A => n4811, ZN => n16384);
   U6029 : INV_X1 port map( A => n15073, ZN => n14571);
   U6031 : INV_X1 port map( A => n4992, ZN => n6674);
   U6032 : OR2_X1 port map( A1 => n15266, A2 => n14922, ZN => n5722);
   U6033 : INV_X1 port map( A => n3673, ZN => n4492);
   U6034 : OR2_X1 port map( A1 => n14598, A2 => n14762, ZN => n3550);
   U6035 : XNOR2_X1 port map( A => n3856, B => n16373, ZN => n16640);
   U6036 : XNOR2_X1 port map( A => n16084, B => n2117, ZN => n16643);
   U6039 : OR2_X1 port map( A1 => n14728, A2 => n15395, ZN => n3605);
   U6040 : OR2_X1 port map( A1 => n13519, A2 => n14884, ZN => n3487);
   U6041 : INV_X1 port map( A => n17298, ZN => n5430);
   U6042 : NOR2_X1 port map( A1 => n5471, A2 => n17143, ZN => n17087);
   U6043 : XNOR2_X1 port map( A => n15106, B => n16229, ZN => n16191);
   U6044 : BUF_X1 port map( A => n14871, Z => n17395);
   U6045 : BUF_X1 port map( A => n16679, Z => n17282);
   U6047 : AND2_X1 port map( A1 => n4414, A2 => n4413, ZN => n17828);
   U6048 : AOI21_X1 port map( B1 => n17074, B2 => n17505, A => n17829, ZN => 
                           n4414);
   U6049 : INV_X1 port map( A => n17556, ZN => n16916);
   U6050 : INV_X1 port map( A => n538, ZN => n4314);
   U6051 : OR2_X1 port map( A1 => n29547, A2 => n18028, ZN => n3932);
   U6052 : OR2_X1 port map( A1 => n18410, A2 => n18121, ZN => n18416);
   U6054 : XNOR2_X1 port map( A => n5859, B => n16658, ZN => n17438);
   U6055 : NAND2_X1 port map( A1 => n17081, A2 => n6067, ZN => n18589);
   U6056 : INV_X1 port map( A => n17151, ZN => n6067);
   U6057 : NOR2_X1 port map( A1 => n28194, A2 => n5891, ZN => n16973);
   U6059 : OR2_X1 port map( A1 => n2825, A2 => n5891, ZN => n2827);
   U6060 : AND2_X1 port map( A1 => n18305, A2 => n18306, ZN => n6576);
   U6062 : NAND2_X1 port map( A1 => n4830, A2 => n4829, ZN => n17834);
   U6064 : OAI211_X1 port map( C1 => n17518, C2 => n17470, A => n6889, B => 
                           n17516, ZN => n17084);
   U6065 : AND2_X1 port map( A1 => n17017, A2 => n17016, ZN => n4866);
   U6066 : AND3_X1 port map( A1 => n17844, A2 => n18241, A3 => n3848, ZN => 
                           n3847);
   U6067 : AND3_X1 port map( A1 => n524, A2 => n18018, A3 => n1888, ZN => n6429
                           );
   U6068 : OR2_X1 port map( A1 => n18251, A2 => n1888, ZN => n18254);
   U6069 : AND2_X1 port map( A1 => n18216, A2 => n18215, ZN => n4824);
   U6070 : OR2_X1 port map( A1 => n17596, A2 => n18227, ZN => n5747);
   U6071 : OR2_X1 port map( A1 => n18261, A2 => n18324, ZN => n17986);
   U6072 : OR2_X1 port map( A1 => n17815, A2 => n4762, ZN => n4761);
   U6073 : OR2_X1 port map( A1 => n17266, A2 => n29298, ZN => n16971);
   U6074 : OAI21_X1 port map( B1 => n18445, B2 => n4928, A => n4927, ZN => 
                           n19252);
   U6075 : AOI21_X1 port map( B1 => n18178, B2 => n4930, A => n4929, ZN => 
                           n4928);
   U6076 : XNOR2_X1 port map( A => n19389, B => n3385, ZN => n19048);
   U6077 : XNOR2_X1 port map( A => n6445, B => n4883, ZN => n19026);
   U6078 : INV_X1 port map( A => n19103, ZN => n6445);
   U6080 : OR2_X1 port map( A1 => n17693, A2 => n18078, ZN => n18079);
   U6081 : OAI22_X1 port map( A1 => n18311, A2 => n17918, B1 => n6225, B2 => 
                           n18355, ZN => n17922);
   U6082 : NOR2_X1 port map( A1 => n2776, A2 => n18123, ZN => n2775);
   U6083 : AND2_X1 port map( A1 => n2778, A2 => n17818, ZN => n2776);
   U6084 : AND2_X1 port map( A1 => n4210, A2 => n4212, ZN => n3402);
   U6085 : XNOR2_X1 port map( A => n19152, B => n4746, ZN => n4745);
   U6086 : AND2_X1 port map( A1 => n18376, A2 => n18380, ZN => n17166);
   U6087 : XNOR2_X1 port map( A => n19496, B => n28516, ZN => n19402);
   U6088 : XNOR2_X1 port map( A => n19553, B => n19552, ZN => n20451);
   U6090 : INV_X1 port map( A => n18691, ZN => n4030);
   U6092 : OR2_X1 port map( A1 => n17756, A2 => n18243, ZN => n2771);
   U6093 : INV_X1 port map( A => n18653, ZN => n19568);
   U6094 : AND2_X1 port map( A1 => n5000, A2 => n21425, ZN => n20896);
   U6095 : AND2_X1 port map( A1 => n21087, A2 => n5827, ZN => n20895);
   U6096 : XNOR2_X1 port map( A => n19543, B => n2993, ZN => n19544);
   U6097 : OAI22_X1 port map( A1 => n19174, A2 => n5491, B1 => n19692, B2 => 
                           n5490, ZN => n19176);
   U6098 : INV_X1 port map( A => n5225, ZN => n5303);
   U6099 : NOR2_X1 port map( A1 => n499, A2 => n6834, ZN => n2797);
   U6100 : AND2_X1 port map( A1 => n19752, A2 => n5937, ZN => n19781);
   U6101 : INV_X1 port map( A => n19761, ZN => n20069);
   U6102 : OR2_X1 port map( A1 => n20089, A2 => n29114, ZN => n6399);
   U6103 : OR2_X1 port map( A1 => n5684, A2 => n20713, ZN => n20714);
   U6104 : OR2_X1 port map( A1 => n20715, A2 => n5684, ZN => n5683);
   U6106 : AND2_X1 port map( A1 => n20451, A2 => n19554, ZN => n21063);
   U6107 : OR2_X1 port map( A1 => n28491, A2 => n21359, ZN => n4167);
   U6108 : OR2_X1 port map( A1 => n19935, A2 => n20607, ZN => n19936);
   U6109 : INV_X1 port map( A => n20647, ZN => n5783);
   U6110 : INV_X1 port map( A => n2081, ZN => n4096);
   U6111 : NAND2_X1 port map( A1 => n20229, A2 => n29426, ZN => n3852);
   U6112 : INV_X1 port map( A => n21642, ZN => n21402);
   U6113 : AND2_X1 port map( A1 => n5778, A2 => n20088, ZN => n18749);
   U6114 : INV_X1 port map( A => n3238, ZN => n5928);
   U6115 : AND2_X1 port map( A1 => n4242, A2 => n19974, ZN => n3243);
   U6116 : INV_X1 port map( A => n21253, ZN => n2125);
   U6117 : OR2_X1 port map( A1 => n21078, A2 => n495, ZN => n21076);
   U6118 : AND2_X1 port map( A1 => n21075, A2 => n21071, ZN => n2992);
   U6119 : INV_X1 port map( A => n21075, ZN => n2989);
   U6120 : OR2_X1 port map( A1 => n21052, A2 => n21051, ZN => n3039);
   U6122 : OR2_X1 port map( A1 => n19921, A2 => n28894, ZN => n20257);
   U6123 : OAI211_X1 port map( C1 => n21818, C2 => n20108, A => n5124, B => 
                           n5123, ZN => n22099);
   U6124 : OR2_X1 port map( A1 => n20043, A2 => n20151, ZN => n4409);
   U6126 : NOR2_X1 port map( A1 => n20152, A2 => n18887, ZN => n18831);
   U6127 : INV_X1 port map( A => n21875, ZN => n22093);
   U6128 : OR2_X1 port map( A1 => n20557, A2 => n20556, ZN => n3193);
   U6129 : INV_X1 port map( A => n19743, ZN => n4362);
   U6130 : AND2_X1 port map( A1 => n5443, A2 => n5442, ZN => n5441);
   U6131 : OR2_X1 port map( A1 => n29530, A2 => n21309, ZN => n5442);
   U6132 : INV_X1 port map( A => n21567, ZN => n6247);
   U6134 : XNOR2_X1 port map( A => n22337, B => n6504, ZN => n22852);
   U6135 : OR2_X1 port map( A1 => n21542, A2 => n20393, ZN => n2725);
   U6136 : XNOR2_X1 port map( A => n22811, B => n22363, ZN => n21454);
   U6137 : AND2_X1 port map( A1 => n23768, A2 => n23765, ZN => n5355);
   U6138 : XNOR2_X1 port map( A => n22710, B => n22320, ZN => n22545);
   U6139 : OAI21_X1 port map( B1 => n481, B2 => n29602, A => n22962, ZN => 
                           n2367);
   U6140 : INV_X1 port map( A => n22923, ZN => n4229);
   U6141 : XNOR2_X1 port map( A => n22882, B => n3321, ZN => n3091);
   U6142 : OAI21_X1 port map( B1 => n20955, B2 => n20802, A => n2296, ZN => 
                           n21102);
   U6143 : OAI21_X1 port map( B1 => n21449, B2 => n21673, A => n3132, ZN => 
                           n3131);
   U6144 : OAI21_X1 port map( B1 => n20830, B2 => n20831, A => n412, ZN => 
                           n20832);
   U6145 : INV_X1 port map( A => n21675, ZN => n3132);
   U6147 : OR2_X1 port map( A1 => n21572, A2 => n21571, ZN => n3562);
   U6148 : OR2_X1 port map( A1 => n20950, A2 => n21538, ZN => n5878);
   U6149 : XNOR2_X1 port map( A => n22896, B => n22692, ZN => n22502);
   U6150 : OR2_X1 port map( A1 => n21202, A2 => n21509, ZN => n3288);
   U6152 : NAND2_X1 port map( A1 => n21393, A2 => n21392, ZN => n2395);
   U6153 : AOI22_X1 port map( A1 => n4143, A2 => n20031, B1 => n3588, B2 => 
                           n21638, ZN => n20035);
   U6154 : NOR2_X1 port map( A1 => n21392, A2 => n21632, ZN => n3588);
   U6155 : XNOR2_X1 port map( A => n28449, B => n3451, ZN => n5840);
   U6156 : OR2_X1 port map( A1 => n21261, A2 => n21718, ZN => n3407);
   U6157 : OR2_X1 port map( A1 => n28789, A2 => n21497, ZN => n6750);
   U6158 : OR2_X1 port map( A1 => n20928, A2 => n21198, ZN => n4566);
   U6160 : INV_X1 port map( A => n5080, ZN => n24092);
   U6161 : INV_X1 port map( A => n23492, ZN => n23791);
   U6162 : XNOR2_X1 port map( A => n22466, B => n22465, ZN => n23392);
   U6163 : OR2_X1 port map( A1 => n23127, A2 => n23126, ZN => n23128);
   U6165 : NOR2_X1 port map( A1 => n24120, A2 => n29726, ZN => n23888);
   U6166 : INV_X1 port map( A => n24305, ZN => n24365);
   U6167 : OAI21_X1 port map( B1 => n24673, B2 => n23334, A => n2130, ZN => 
                           n25444);
   U6168 : AND2_X1 port map( A1 => n24323, A2 => n404, ZN => n4025);
   U6169 : AND2_X1 port map( A1 => n24547, A2 => n24160, ZN => n2820);
   U6170 : XNOR2_X1 port map( A => n24254, B => n24255, ZN => n25406);
   U6171 : XNOR2_X1 port map( A => n25191, B => n4861, ZN => n24784);
   U6172 : AND3_X1 port map( A1 => n5479, A2 => n5478, A3 => n220, ZN => n23698
                           );
   U6173 : OR2_X1 port map( A1 => n24817, A2 => n24809, ZN => n5479);
   U6174 : OR2_X1 port map( A1 => n24237, A2 => n24195, ZN => n24571);
   U6175 : OR2_X1 port map( A1 => n24551, A2 => n24552, ZN => n5509);
   U6176 : OR2_X1 port map( A1 => n5094, A2 => n24593, ZN => n4690);
   U6177 : INV_X1 port map( A => n24257, ZN => n2175);
   U6178 : XNOR2_X1 port map( A => n28465, B => n3493, ZN => n5431);
   U6179 : XNOR2_X1 port map( A => n5146, B => n26899, ZN => n25140);
   U6182 : OR2_X1 port map( A1 => n24972, A2 => n24256, ZN => n3121);
   U6183 : OAI21_X1 port map( B1 => n24716, B2 => n4136, A => n4135, ZN => 
                           n23869);
   U6184 : XNOR2_X1 port map( A => n25546, B => n26093, ZN => n26007);
   U6185 : NOR2_X1 port map( A1 => n5105, A2 => n24227, ZN => n5104);
   U6186 : NAND2_X1 port map( A1 => n2880, A2 => n2878, ZN => n4161);
   U6187 : INV_X1 port map( A => n24237, ZN => n6239);
   U6189 : AND2_X1 port map( A1 => n24711, A2 => n24713, ZN => n23070);
   U6190 : XNOR2_X1 port map( A => n26083, B => n26053, ZN => n25533);
   U6193 : XNOR2_X1 port map( A => n26101, B => n25411, ZN => n2812);
   U6194 : INV_X1 port map( A => n24797, ZN => n25786);
   U6195 : XNOR2_X1 port map( A => n25577, B => n25282, ZN => n25875);
   U6196 : XNOR2_X1 port map( A => n25430, B => n25369, ZN => n25898);
   U6197 : OR2_X1 port map( A1 => n26466, A2 => n26191, ZN => n26192);
   U6198 : AND2_X1 port map( A1 => n29028, A2 => n25406, ZN => n6685);
   U6199 : XNOR2_X1 port map( A => n1958, B => n25311, ZN => n4643);
   U6200 : AND2_X1 port map( A1 => n26581, A2 => n26927, ZN => n4401);
   U6201 : INV_X1 port map( A => n26927, ZN => n4402);
   U6202 : XNOR2_X1 port map( A => n24982, B => n24983, ZN => n26385);
   U6203 : OR2_X1 port map( A1 => n27055, A2 => n27902, ZN => n26851);
   U6205 : XNOR2_X1 port map( A => n3168, B => n25712, ZN => n27063);
   U6207 : AND2_X1 port map( A1 => n29524, A2 => n29058, ZN => n27001);
   U6208 : OR2_X1 port map( A1 => n26623, A2 => n27050, ZN => n26246);
   U6209 : NOR2_X1 port map( A1 => n28468, A2 => n27548, ZN => n2617);
   U6210 : INV_X1 port map( A => n27287, ZN => n27281);
   U6211 : OAI21_X1 port map( B1 => n29022, B2 => n27772, A => n6419, ZN => 
                           n6418);
   U6212 : AND2_X1 port map( A1 => n7584, A2 => n7303, ZN => n3004);
   U6213 : INV_X1 port map( A => n7257, ZN => n6209);
   U6214 : AND2_X1 port map( A1 => n29639, A2 => n7488, ZN => n7664);
   U6215 : INV_X1 port map( A => n7585, ZN => n2224);
   U6216 : NOR2_X1 port map( A1 => n7580, A2 => n7071, ZN => n2223);
   U6217 : INV_X1 port map( A => n8724, ZN => n10241);
   U6218 : OR2_X1 port map( A1 => n8720, A2 => n8787, ZN => n4322);
   U6219 : AND2_X1 port map( A1 => n8810, A2 => n8523, ZN => n3225);
   U6220 : NAND3_X1 port map( A1 => n3094, A2 => n8283, A3 => n3093, ZN => 
                           n8956);
   U6221 : OR2_X1 port map( A1 => n8285, A2 => n8284, ZN => n3093);
   U6222 : INV_X1 port map( A => n8658, ZN => n8501);
   U6223 : AND2_X1 port map( A1 => n2740, A2 => n2739, ZN => n7302);
   U6224 : OR2_X1 port map( A1 => n9004, A2 => n9184, ZN => n3755);
   U6226 : OR3_X1 port map( A1 => n9184, A2 => n8782, A3 => n9009, ZN => n7755)
                           ;
   U6227 : OR2_X1 port map( A1 => n8642, A2 => n8984, ZN => n9176);
   U6229 : OR2_X1 port map( A1 => n8752, A2 => n8751, ZN => n3050);
   U6232 : OR2_X1 port map( A1 => n6590, A2 => n5944, ZN => n4730);
   U6233 : NAND4_X1 port map( A1 => n8076, A2 => n2698, A3 => n8075, A4 => 
                           n8074, ZN => n10028);
   U6234 : INV_X1 port map( A => n9097, ZN => n2698);
   U6235 : AND2_X1 port map( A1 => n8666, A2 => n8490, ZN => n9097);
   U6237 : OAI211_X1 port map( C1 => n610, C2 => n8897, A => n3274, B => n2980,
                           ZN => n3273);
   U6239 : OR2_X1 port map( A1 => n8888, A2 => n8886, ZN => n8010);
   U6240 : XNOR2_X1 port map( A => n9794, B => n2677, ZN => n9658);
   U6241 : OR2_X1 port map( A1 => n9026, A2 => n597, ZN => n3780);
   U6242 : XNOR2_X1 port map( A => n10144, B => n1225, ZN => n4507);
   U6243 : OR2_X1 port map( A1 => n11166, A2 => n10820, ZN => n2103);
   U6244 : OR2_X1 port map( A1 => n8327, A2 => n606, ZN => n3609);
   U6245 : AND2_X1 port map( A1 => n9120, A2 => n9119, ZN => n4969);
   U6246 : MUX2_X1 port map( A => n9149, B => n11, S => n9146, Z => n9155);
   U6247 : AND2_X1 port map( A1 => n8338, A2 => n8337, ZN => n2712);
   U6248 : XNOR2_X1 port map( A => n9296, B => n9977, ZN => n5268);
   U6249 : XNOR2_X1 port map( A => n9931, B => n4713, ZN => n10303);
   U6250 : OR2_X1 port map( A1 => n8753, A2 => n9132, ZN => n8341);
   U6251 : OR2_X1 port map( A1 => n8631, A2 => n8490, ZN => n8494);
   U6252 : XNOR2_X1 port map( A => n10227, B => n9899, ZN => n9825);
   U6253 : OR2_X1 port map( A1 => n8852, A2 => n9079, ZN => n7493);
   U6254 : OR2_X1 port map( A1 => n8851, A2 => n8724, ZN => n7491);
   U6255 : OR2_X1 port map( A1 => n11351, A2 => n11350, ZN => n11190);
   U6256 : INV_X1 port map( A => n11165, ZN => n9686);
   U6257 : NOR2_X1 port map( A1 => n8422, A2 => n10821, ZN => n2127);
   U6258 : OR2_X1 port map( A1 => n10522, A2 => n279, ZN => n11276);
   U6259 : INV_X1 port map( A => n10051, ZN => n10730);
   U6260 : OR2_X1 port map( A1 => n5366, A2 => n28208, ZN => n4902);
   U6262 : AND2_X1 port map( A1 => n11435, A2 => n12266, ZN => n2466);
   U6264 : XNOR2_X1 port map( A => n1990, B => n8845, ZN => n11335);
   U6265 : INV_X1 port map( A => n12206, ZN => n4038);
   U6266 : OR2_X1 port map( A1 => n4037, A2 => n12109, ZN => n2683);
   U6267 : INV_X1 port map( A => n11671, ZN => n5079);
   U6268 : OR2_X1 port map( A1 => n11165, A2 => n11053, ZN => n11309);
   U6269 : AND2_X1 port map( A1 => n10833, A2 => n11033, ZN => n4801);
   U6270 : NOR2_X1 port map( A1 => n11047, A2 => n11261, ZN => n6515);
   U6272 : AND2_X1 port map( A1 => n11185, A2 => n11186, ZN => n3907);
   U6273 : OR2_X1 port map( A1 => n10431, A2 => n5279, ZN => n10577);
   U6274 : AND2_X1 port map( A1 => n10620, A2 => n11226, ZN => n10623);
   U6275 : NOR2_X1 port map( A1 => n11990, A2 => n10863, ZN => n11617);
   U6276 : INV_X1 port map( A => n12566, ZN => n13557);
   U6277 : AOI21_X1 port map( B1 => n12512, B2 => n10863, A => n6374, ZN => 
                           n5090);
   U6278 : NOR2_X1 port map( A1 => n12211, A2 => n12111, ZN => n4449);
   U6279 : INV_X1 port map( A => n10648, ZN => n12343);
   U6280 : INV_X1 port map( A => n12200, ZN => n11807);
   U6281 : AND2_X1 port map( A1 => n11007, A2 => n11006, ZN => n3013);
   U6282 : INV_X1 port map( A => n11990, ZN => n5637);
   U6283 : INV_X1 port map( A => n3653, ZN => n3108);
   U6284 : OR2_X1 port map( A1 => n10923, A2 => n10920, ZN => n3776);
   U6285 : AND2_X1 port map( A1 => n11195, A2 => n11194, ZN => n12261);
   U6286 : INV_X1 port map( A => n4341, ZN => n11954);
   U6288 : INV_X1 port map( A => n10905, ZN => n11927);
   U6289 : INV_X1 port map( A => n11921, ZN => n11549);
   U6291 : NOR2_X1 port map( A1 => n11022, A2 => n11315, ZN => n3882);
   U6292 : AND2_X1 port map( A1 => n3817, A2 => n11248, ZN => n3275);
   U6293 : OR2_X1 port map( A1 => n11540, A2 => n572, ZN => n6659);
   U6294 : INV_X1 port map( A => n4474, ZN => n12808);
   U6295 : OR2_X1 port map( A1 => n10685, A2 => n28405, ZN => n6780);
   U6296 : OR2_X1 port map( A1 => n10691, A2 => n4538, ZN => n4537);
   U6297 : AND2_X1 port map( A1 => n10957, A2 => n10962, ZN => n6775);
   U6299 : OR2_X1 port map( A1 => n11116, A2 => n11115, ZN => n3807);
   U6300 : AND2_X1 port map( A1 => n12042, A2 => n11962, ZN => n12043);
   U6301 : OR2_X1 port map( A1 => n11963, A2 => n11968, ZN => n2976);
   U6302 : OR2_X1 port map( A1 => n11514, A2 => n12244, ZN => n3021);
   U6303 : AOI21_X1 port map( B1 => n12155, B2 => n12991, A => n430, ZN => 
                           n11387);
   U6304 : OR2_X1 port map( A1 => n5964, A2 => n2008, ZN => n4997);
   U6305 : INV_X1 port map( A => n13457, ZN => n6298);
   U6306 : XNOR2_X1 port map( A => n13460, B => n13459, ZN => n2172);
   U6307 : OR2_X1 port map( A1 => n14593, A2 => n14101, ZN => n4150);
   U6308 : AND2_X1 port map( A1 => n2440, A2 => n11946, ZN => n11950);
   U6310 : AND2_X1 port map( A1 => n15503, A2 => n15506, ZN => n5575);
   U6311 : NOR2_X1 port map( A1 => n12146, A2 => n11715, ZN => n5169);
   U6312 : OR2_X1 port map( A1 => n11415, A2 => n11715, ZN => n3688);
   U6314 : INV_X1 port map( A => n12377, ZN => n13562);
   U6315 : XNOR2_X1 port map( A => n2975, B => n13209, ZN => n13402);
   U6316 : INV_X1 port map( A => n13025, ZN => n2975);
   U6317 : OR3_X1 port map( A1 => n15180, A2 => n28803, A3 => n15174, ZN => 
                           n13841);
   U6318 : OR2_X1 port map( A1 => n14407, A2 => n5584, ZN => n4974);
   U6319 : AND2_X1 port map( A1 => n14398, A2 => n13877, ZN => n4009);
   U6320 : INV_X1 port map( A => n28806, ZN => n2959);
   U6321 : INV_X1 port map( A => n14166, ZN => n13947);
   U6322 : AND2_X1 port map( A1 => n14241, A2 => n15194, ZN => n6571);
   U6323 : AND2_X1 port map( A1 => n14078, A2 => n14250, ZN => n5789);
   U6324 : AND2_X1 port map( A1 => n14165, A2 => n14487, ZN => n13948);
   U6325 : OAI211_X1 port map( C1 => n5693, C2 => n14181, A => n5451, B => 
                           n1320, ZN => n15345);
   U6326 : INV_X1 port map( A => n14480, ZN => n14161);
   U6328 : OR2_X1 port map( A1 => n14084, A2 => n14287, ZN => n14080);
   U6329 : NAND2_X1 port map( A1 => n1848, A2 => n15171, ZN => n13865);
   U6330 : OR2_X1 port map( A1 => n14262, A2 => n14259, ZN => n13761);
   U6331 : OR2_X1 port map( A1 => n15491, A2 => n15485, ZN => n14618);
   U6332 : OAI211_X1 port map( C1 => n14575, C2 => n2733, A => n2732, B => 
                           n2731, ZN => n16304);
   U6333 : OAI21_X1 port map( B1 => n14172, B2 => n14173, A => n15199, ZN => 
                           n3012);
   U6334 : INV_X1 port map( A => n16283, ZN => n16486);
   U6335 : INV_X1 port map( A => n14645, ZN => n2191);
   U6336 : OR2_X1 port map( A1 => n13847, A2 => n293, ZN => n6725);
   U6337 : NOR2_X1 port map( A1 => n4992, A2 => n15060, ZN => n15062);
   U6339 : AOI21_X1 port map( B1 => n14496, B2 => n14154, A => n6798, ZN => 
                           n14501);
   U6340 : AND2_X1 port map( A1 => n14495, A2 => n14494, ZN => n6798);
   U6341 : OR2_X1 port map( A1 => n14453, A2 => n1320, ZN => n5641);
   U6342 : OR2_X1 port map( A1 => n15164, A2 => n15464, ZN => n4677);
   U6343 : OR2_X1 port map( A1 => n15010, A2 => n15374, ZN => n6877);
   U6344 : OAI211_X1 port map( C1 => n15008, C2 => n426, A => n15369, B => 
                           n3783, ZN => n6880);
   U6345 : AOI22_X1 port map( A1 => n2608, A2 => n14230, B1 => n14108, B2 => 
                           n14107, ZN => n14109);
   U6346 : OAI22_X1 port map( A1 => n14390, A2 => n14601, B1 => n15288, B2 => 
                           n14391, ZN => n2208);
   U6347 : OR2_X1 port map( A1 => n15691, A2 => n13989, ZN => n4407);
   U6348 : AND2_X1 port map( A1 => n13932, A2 => n2493, ZN => n13930);
   U6349 : AND2_X1 port map( A1 => n14784, A2 => n15184, ZN => n14533);
   U6350 : AND2_X1 port map( A1 => n14677, A2 => n15098, ZN => n4660);
   U6351 : AND2_X1 port map( A1 => n15183, A2 => n15182, ZN => n13818);
   U6353 : AND2_X1 port map( A1 => n15015, A2 => n15014, ZN => n15320);
   U6354 : OR2_X1 port map( A1 => n14516, A2 => n15115, ZN => n5444);
   U6355 : INV_X1 port map( A => n14928, ZN => n14960);
   U6356 : INV_X1 port map( A => n14697, ZN => n15512);
   U6357 : INV_X1 port map( A => n13587, ZN => n14038);
   U6358 : OAI21_X1 port map( B1 => n15335, B2 => n15338, A => n28802, ZN => 
                           n15240);
   U6359 : OR2_X1 port map( A1 => n15104, A2 => n15420, ZN => n5379);
   U6360 : XNOR2_X1 port map( A => n15397, B => n1957, ZN => n17296);
   U6361 : OR2_X1 port map( A1 => n14187, A2 => n12743, ZN => n14189);
   U6362 : OR2_X1 port map( A1 => n14261, A2 => n3395, ZN => n3750);
   U6363 : OR2_X1 port map( A1 => n14098, A2 => n3396, ZN => n3749);
   U6364 : OAI21_X1 port map( B1 => n13758, B2 => n15152, A => n2448, ZN => 
                           n16318);
   U6365 : OAI21_X1 port map( B1 => n28222, B2 => n2028, A => n15056, ZN => 
                           n2162);
   U6366 : AND3_X1 port map( A1 => n15264, A2 => n4097, A3 => n2738, ZN => 
                           n14711);
   U6367 : OR2_X1 port map( A1 => n15260, A2 => n15054, ZN => n2738);
   U6368 : XNOR2_X1 port map( A => n6454, B => n16625, ZN => n6453);
   U6369 : AND2_X1 port map( A1 => n14021, A2 => n14024, ZN => n3782);
   U6370 : INV_X1 port map( A => n16878, ZN => n17388);
   U6371 : XNOR2_X1 port map( A => n16051, B => n1967, ZN => n16525);
   U6372 : OR2_X1 port map( A1 => n14706, A2 => n15506, ZN => n6216);
   U6373 : OR2_X1 port map( A1 => n14641, A2 => n15082, ZN => n2592);
   U6374 : AND2_X1 port map( A1 => n2744, A2 => n14982, ZN => n2743);
   U6375 : OR2_X1 port map( A1 => n14797, A2 => n14534, ZN => n2742);
   U6376 : XNOR2_X1 port map( A => n15545, B => n6295, ZN => n15874);
   U6377 : INV_X1 port map( A => n3856, ZN => n6295);
   U6378 : AND2_X1 port map( A1 => n17348, A2 => n29632, ZN => n16948);
   U6379 : XNOR2_X1 port map( A => n28406, B => n4852, ZN => n16203);
   U6380 : AND2_X1 port map( A1 => n16724, A2 => n4687, ZN => n6559);
   U6381 : XNOR2_X1 port map( A => n15909, B => n5406, ZN => n15682);
   U6382 : INV_X1 port map( A => n16377, ZN => n5406);
   U6383 : XNOR2_X1 port map( A => n15660, B => n15659, ZN => n16944);
   U6384 : INV_X1 port map( A => n15174, ZN => n3080);
   U6385 : OR2_X1 port map( A1 => n15326, A2 => n15014, ZN => n2699);
   U6386 : INV_X1 port map( A => n3565, ZN => n4978);
   U6388 : INV_X1 port map( A => n16467, ZN => n6296);
   U6389 : NOR2_X1 port map( A1 => n4218, A2 => n17548, ZN => n16946);
   U6390 : INV_X1 port map( A => n17338, ZN => n17201);
   U6392 : OR2_X1 port map( A1 => n17459, A2 => n16812, ZN => n16813);
   U6396 : AND2_X1 port map( A1 => n16860, A2 => n16814, ZN => n16687);
   U6397 : INV_X1 port map( A => n17137, ZN => n17502);
   U6398 : OR2_X1 port map( A1 => n17304, A2 => n6002, ZN => n6001);
   U6399 : AND2_X1 port map( A1 => n17304, A2 => n17421, ZN => n17616);
   U6400 : OR2_X1 port map( A1 => n4269, A2 => n17830, ZN => n2856);
   U6401 : INV_X1 port map( A => n4218, ZN => n2133);
   U6402 : NOR2_X1 port map( A1 => n5398, A2 => n17552, ZN => n2632);
   U6404 : AND2_X1 port map( A1 => n18197, A2 => n16718, ZN => n4174);
   U6405 : AOI21_X1 port map( B1 => n511, B2 => n18500, A => n18506, ZN => 
                           n5392);
   U6407 : AND2_X1 port map( A1 => n18325, A2 => n18262, ZN => n4058);
   U6408 : OR2_X1 port map( A1 => n337, A2 => n17437, ZN => n17308);
   U6409 : AND3_X1 port map( A1 => n18441, A2 => n4929, A3 => n18444, ZN => 
                           n4786);
   U6410 : OR2_X1 port map( A1 => n18012, A2 => n18480, ZN => n5179);
   U6412 : INV_X1 port map( A => n17336, ZN => n2664);
   U6413 : INV_X1 port map( A => n387, ZN => n6830);
   U6414 : OR2_X1 port map( A1 => n17441, A2 => n336, ZN => n5458);
   U6415 : NAND2_X1 port map( A1 => n3250, A2 => n17422, ZN => n18231);
   U6416 : AND2_X1 port map( A1 => n17695, A2 => n18276, ZN => n17804);
   U6417 : AND2_X1 port map( A1 => n18124, A2 => n17834, ZN => n17840);
   U6418 : AND2_X1 port map( A1 => n18596, A2 => n18595, ZN => n2341);
   U6419 : INV_X1 port map( A => n18332, ZN => n18372);
   U6420 : AND2_X1 port map( A1 => n18232, A2 => n18402, ZN => n3285);
   U6421 : OAI21_X1 port map( B1 => n17715, B2 => n17720, A => n6588, ZN => 
                           n18526);
   U6422 : OR2_X1 port map( A1 => n17990, A2 => n6927, ZN => n6713);
   U6423 : OR2_X1 port map( A1 => n15647, A2 => n28793, ZN => n5610);
   U6424 : OR2_X1 port map( A1 => n16714, A2 => n4283, ZN => n5609);
   U6425 : OR2_X1 port map( A1 => n518, A2 => n18356, ZN => n2317);
   U6426 : OR2_X1 port map( A1 => n6030, A2 => n16611, ZN => n2838);
   U6427 : OR2_X1 port map( A1 => n4059, A2 => n18268, ZN => n4119);
   U6429 : AND2_X1 port map( A1 => n6230, A2 => n6229, ZN => n6228);
   U6430 : AND2_X1 port map( A1 => n18285, A2 => n18081, ZN => n18083);
   U6431 : INV_X1 port map( A => n19706, ZN => n3284);
   U6432 : AOI22_X1 port map( A1 => n16980, A2 => n18523, B1 => n18524, B2 => 
                           n373, ZN => n16981);
   U6433 : INV_X1 port map( A => n19111, ZN => n18980);
   U6435 : INV_X1 port map( A => n5492, ZN => n5491);
   U6436 : AND2_X1 port map( A1 => n20193, A2 => n20414, ZN => n20578);
   U6437 : OR2_X1 port map( A1 => n17918, A2 => n18354, ZN => n5842);
   U6438 : INV_X1 port map( A => n20200, ZN => n20304);
   U6439 : XNOR2_X1 port map( A => n18857, B => n18856, ZN => n19269);
   U6440 : INV_X1 port map( A => n18877, ZN => n3403);
   U6441 : OR2_X1 port map( A1 => n17639, A2 => n29125, ZN => n17640);
   U6445 : OR2_X1 port map( A1 => n18458, A2 => n18459, ZN => n6670);
   U6446 : AND2_X1 port map( A1 => n18455, A2 => n18456, ZN => n6671);
   U6447 : INV_X1 port map( A => n20302, ZN => n5436);
   U6448 : INV_X1 port map( A => n18690, ZN => n18927);
   U6449 : XNOR2_X1 port map( A => n19139, B => n1179, ZN => n5746);
   U6450 : XNOR2_X1 port map( A => n18867, B => n19108, ZN => n19599);
   U6451 : XNOR2_X1 port map( A => n19247, B => n4030, ZN => n19248);
   U6452 : OR2_X1 port map( A1 => n18042, A2 => n18423, ZN => n4802);
   U6453 : OAI21_X1 port map( B1 => n18202, B2 => n18201, A => n18200, ZN => 
                           n6488);
   U6454 : XNOR2_X1 port map( A => n19252, B => n18948, ZN => n6276);
   U6455 : AND2_X1 port map( A1 => n20533, A2 => n20933, ZN => n5125);
   U6456 : OR2_X1 port map( A1 => n20144, A2 => n21091, ZN => n5854);
   U6457 : INV_X1 port map( A => n21087, ZN => n21426);
   U6458 : AND2_X1 port map( A1 => n20283, A2 => n20282, ZN => n19896);
   U6459 : NOR2_X1 port map( A1 => n20443, A2 => n20299, ZN => n20446);
   U6460 : OR2_X1 port map( A1 => n22145, A2 => n22139, ZN => n21030);
   U6461 : NOR2_X1 port map( A1 => n20406, A2 => n28501, ZN => n6315);
   U6462 : XNOR2_X1 port map( A => n5522, B => n5521, ZN => n5520);
   U6464 : AND2_X1 port map( A1 => n20474, A2 => n5408, ZN => n21275);
   U6465 : OR2_X1 port map( A1 => n20477, A2 => n20475, ZN => n20352);
   U6466 : OR2_X1 port map( A1 => n21143, A2 => n4395, ZN => n4394);
   U6467 : AND2_X1 port map( A1 => n20351, A2 => n21547, ZN => n20362);
   U6468 : OAI21_X1 port map( B1 => n18846, B2 => n18776, A => n19765, ZN => 
                           n5469);
   U6470 : OR2_X1 port map( A1 => n20450, A2 => n5375, ZN => n2747);
   U6471 : OR2_X1 port map( A1 => n20183, A2 => n499, ZN => n19185);
   U6472 : OR2_X1 port map( A1 => n20721, A2 => n21599, ZN => n5720);
   U6473 : INV_X1 port map( A => n22320, ZN => n22379);
   U6474 : OR2_X1 port map( A1 => n20466, A2 => n21932, ZN => n20184);
   U6475 : AND2_X1 port map( A1 => n21119, A2 => n21144, ZN => n21122);
   U6476 : NAND3_X1 port map( A1 => n21412, A2 => n4937, A3 => n28184, ZN => 
                           n2653);
   U6478 : INV_X1 port map( A => n5684, ZN => n5983);
   U6479 : OAI21_X1 port map( B1 => n21447, B2 => n21080, A => n20213, ZN => 
                           n21959);
   U6480 : NOR2_X1 port map( A1 => n21674, A2 => n21679, ZN => n21080);
   U6481 : INV_X1 port map( A => n22633, ZN => n22691);
   U6482 : OR2_X1 port map( A1 => n21625, A2 => n22145, ZN => n21028);
   U6483 : OR2_X1 port map( A1 => n22149, A2 => n22148, ZN => n2097);
   U6485 : AND2_X1 port map( A1 => n20276, A2 => n6016, ZN => n2666);
   U6486 : AND2_X1 port map( A1 => n20269, A2 => n2669, ZN => n2668);
   U6487 : OR2_X1 port map( A1 => n21645, A2 => n21642, ZN => n4071);
   U6488 : OR2_X1 port map( A1 => n22288, A2 => n21208, ZN => n3858);
   U6489 : AOI21_X1 port map( B1 => n6240, B2 => n20781, A => n20780, ZN => 
                           n20885);
   U6490 : INV_X1 port map( A => n5782, ZN => n5780);
   U6491 : OR2_X1 port map( A1 => n20441, A2 => n20440, ZN => n3547);
   U6492 : XNOR2_X1 port map( A => n22822, B => n22132, ZN => n22571);
   U6493 : XNOR2_X1 port map( A => n22132, B => n21959, ZN => n22800);
   U6494 : INV_X1 port map( A => n20885, ZN => n22787);
   U6495 : XNOR2_X1 port map( A => n5395, B => n22903, ZN => n6364);
   U6496 : XNOR2_X1 port map( A => n22337, B => n634, ZN => n5395);
   U6497 : OR2_X1 port map( A1 => n20888, A2 => n20889, ZN => n6039);
   U6498 : AND2_X1 port map( A1 => n21237, A2 => n21399, ZN => n21751);
   U6499 : XNOR2_X1 port map( A => n6141, B => n22791, ZN => n22164);
   U6500 : NAND2_X1 port map( A1 => n4638, A2 => n4634, ZN => n22594);
   U6502 : OR2_X1 port map( A1 => n21382, A2 => n4266, ZN => n4265);
   U6503 : OR2_X1 port map( A1 => n29488, A2 => n21269, ZN => n6427);
   U6504 : INV_X1 port map( A => n20989, ZN => n6116);
   U6505 : XNOR2_X1 port map( A => n21903, B => n22488, ZN => n22727);
   U6506 : OR2_X1 port map( A1 => n21257, A2 => n5772, ZN => n3319);
   U6507 : XNOR2_X1 port map( A => n22417, B => n22416, ZN => n23651);
   U6508 : OR2_X1 port map( A1 => n23733, A2 => n2141, ZN => n2951);
   U6510 : OR2_X1 port map( A1 => n23790, A2 => n23492, ZN => n23319);
   U6511 : OR2_X1 port map( A1 => n21445, A2 => n20833, ZN => n6349);
   U6512 : XNOR2_X1 port map( A => n20682, B => n20681, ZN => n3887);
   U6513 : NOR2_X1 port map( A1 => n2138, A2 => n1838, ZN => n4255);
   U6514 : NOR2_X1 port map( A1 => n28390, A2 => n29074, ZN => n4256);
   U6515 : INV_X1 port map( A => n23177, ZN => n23645);
   U6517 : OR2_X1 port map( A1 => n23501, A2 => n28554, ZN => n5354);
   U6518 : INV_X1 port map( A => n4726, ZN => n23537);
   U6519 : OR2_X1 port map( A1 => n23800, A2 => n28444, ZN => n23536);
   U6520 : AND2_X1 port map( A1 => n22284, A2 => n29061, ZN => n23554);
   U6521 : AOI22_X1 port map( A1 => n5541, A2 => n23835, B1 => n23833, B2 => 
                           n23834, ZN => n4532);
   U6522 : AND2_X1 port map( A1 => n23662, A2 => n23163, ZN => n23524);
   U6523 : INV_X1 port map( A => n23769, ZN => n23499);
   U6525 : OR2_X1 port map( A1 => n23765, A2 => n23764, ZN => n23501);
   U6527 : OR2_X1 port map( A1 => n23586, A2 => n23262, ZN => n4234);
   U6528 : NOR2_X1 port map( A1 => n23455, A2 => n23456, ZN => n23357);
   U6529 : XNOR2_X1 port map( A => n22922, B => n4229, ZN => n4228);
   U6530 : AND2_X1 port map( A1 => n29120, A2 => n28523, ZN => n6596);
   U6531 : NOR2_X1 port map( A1 => n24581, A2 => n24468, ZN => n3295);
   U6532 : OR2_X1 port map( A1 => n23789, A2 => n23790, ZN => n6609);
   U6533 : OR2_X1 port map( A1 => n23809, A2 => n22742, ZN => n2202);
   U6534 : OR2_X1 port map( A1 => n24709, A2 => n24341, ZN => n24705);
   U6535 : INV_X1 port map( A => n23606, ZN => n5347);
   U6537 : XNOR2_X1 port map( A => n22137, B => n22138, ZN => n23712);
   U6538 : OR2_X1 port map( A1 => n23228, A2 => n23227, ZN => n23229);
   U6539 : AND2_X1 port map( A1 => n2823, A2 => n23126, ZN => n2822);
   U6540 : OR2_X1 port map( A1 => n4664, A2 => n24376, ZN => n3205);
   U6541 : INV_X1 port map( A => n24613, ZN => n24057);
   U6542 : OR2_X1 port map( A1 => n24593, A2 => n24141, ZN => n3481);
   U6543 : INV_X1 port map( A => n23467, ZN => n6787);
   U6544 : NAND4_X1 port map( A1 => n6109, A2 => n23409, A3 => n23410, A4 => 
                           n23507, ZN => n6110);
   U6545 : NOR2_X1 port map( A1 => n24614, A2 => n29109, ZN => n5217);
   U6546 : NAND2_X1 port map( A1 => n24339, A2 => n24334, ZN => n24709);
   U6547 : AND2_X1 port map( A1 => n24706, A2 => n24708, ZN => n5751);
   U6548 : OR2_X1 port map( A1 => n23042, A2 => n23632, ZN => n23043);
   U6549 : INV_X1 port map( A => n2153, ZN => n2154);
   U6551 : INV_X1 port map( A => n22747, ZN => n23979);
   U6552 : AND2_X1 port map( A1 => n5210, A2 => n25007, ZN => n24065);
   U6553 : AOI22_X1 port map( A1 => n23303, A2 => n5699, B1 => n5530, B2 => 
                           n4019, ZN => n4177);
   U6554 : INV_X1 port map( A => n24582, ZN => n24054);
   U6555 : OAI211_X1 port map( C1 => n22998, C2 => n23563, A => n2623, B => 
                           n2622, ZN => n24437);
   U6557 : INV_X1 port map( A => n24188, ZN => n2240);
   U6558 : BUF_X1 port map( A => n24984, Z => n25781);
   U6560 : XNOR2_X1 port map( A => n24958, B => n24957, ZN => n26384);
   U6562 : INV_X1 port map( A => n5263, ZN => n25750);
   U6563 : AND2_X1 port map( A1 => n29622, A2 => n5263, ZN => n27079);
   U6564 : INV_X1 port map( A => n25815, ZN => n27086);
   U6565 : AND2_X1 port map( A1 => n26614, A2 => n27067, ZN => n27065);
   U6566 : AND2_X1 port map( A1 => n24501, A2 => n24500, ZN => n3206);
   U6567 : XNOR2_X1 port map( A => n26118, B => n25849, ZN => n25311);
   U6569 : INV_X1 port map( A => n27038, ZN => n5314);
   U6570 : BUF_X1 port map( A => n25633, Z => n26960);
   U6571 : NOR2_X1 port map( A1 => n23862, A2 => n25418, ZN => n23863);
   U6572 : NAND2_X1 port map( A1 => n24575, A2 => n26560, ZN => n5504);
   U6573 : NOR2_X1 port map( A1 => n377, A2 => n4913, ZN => n24575);
   U6574 : NOR2_X1 port map( A1 => n26435, A2 => n26935, ZN => n26558);
   U6575 : OR2_X1 port map( A1 => n28471, A2 => n28423, ZN => n2323);
   U6576 : OR2_X1 port map( A1 => n26801, A2 => n26800, ZN => n6322);
   U6577 : AND2_X1 port map( A1 => n26132, A2 => n28642, ZN => n26260);
   U6581 : INV_X1 port map( A => n2145, ZN => n27123);
   U6582 : INV_X1 port map( A => n26851, ZN => n27838);
   U6583 : INV_X1 port map( A => n26310, ZN => n26866);
   U6584 : NOR2_X1 port map( A1 => n26125, A2 => n27140, ZN => n26519);
   U6585 : INV_X1 port map( A => n26507, ZN => n27087);
   U6586 : OR2_X1 port map( A1 => n26251, A2 => n26733, ZN => n5390);
   U6587 : OR2_X1 port map( A1 => n5388, A2 => n26995, ZN => n5391);
   U6588 : OR2_X1 port map( A1 => n27043, A2 => n29058, ZN => n4497);
   U6589 : AND2_X1 port map( A1 => n27052, A2 => n25983, ZN => n27017);
   U6591 : XNOR2_X1 port map( A => n2153, B => n1928, ZN => n25257);
   U6592 : OR2_X1 port map( A1 => n26222, A2 => n29159, ZN => n28101);
   U6593 : INV_X1 port map( A => n26652, ZN => n27537);
   U6594 : INV_X1 port map( A => n27038, ZN => n27209);
   U6595 : NOR2_X1 port map( A1 => n26197, A2 => n26196, ZN => n5373);
   U6597 : AND2_X1 port map( A1 => n342, A2 => n26960, ZN => n4921);
   U6598 : AND2_X1 port map( A1 => n27465, A2 => n29468, ZN => n6712);
   U6599 : INV_X1 port map( A => n27525, ZN => n4809);
   U6600 : NOR3_X1 port map( A1 => n27505, A2 => n27527, A3 => n27523, ZN => 
                           n27513);
   U6601 : OR2_X1 port map( A1 => n26804, A2 => n26280, ZN => n3075);
   U6602 : OR2_X1 port map( A1 => n26785, A2 => n6070, ZN => n3703);
   U6603 : NOR2_X1 port map( A1 => n26787, A2 => n26788, ZN => n3702);
   U6605 : AND2_X1 port map( A1 => n26880, A2 => n27301, ZN => n27259);
   U6606 : OAI21_X1 port map( B1 => n26918, B2 => n26782, A => n26920, ZN => 
                           n6633);
   U6607 : NOR2_X1 port map( A1 => n27547, A2 => n27203, ZN => n27546);
   U6608 : AND2_X1 port map( A1 => n27567, A2 => n3087, ZN => n2268);
   U6609 : AOI21_X1 port map( B1 => n28421, B2 => n6724, A => n26935, ZN => 
                           n6723);
   U6610 : NOR2_X1 port map( A1 => n27591, A2 => n27596, ZN => n27592);
   U6612 : INV_X1 port map( A => n27672, ZN => n5877);
   U6614 : NOR2_X1 port map( A1 => n27780, A2 => n29070, ZN => n27769);
   U6616 : NAND2_X1 port map( A1 => n6025, A2 => n6024, ZN => n27772);
   U6617 : OR2_X1 port map( A1 => n6008, A2 => n26297, ZN => n6024);
   U6618 : INV_X1 port map( A => n27826, ZN => n2378);
   U6619 : AND2_X1 port map( A1 => n27827, A2 => n27841, ZN => n2767);
   U6620 : OAI211_X1 port map( C1 => n27056, C2 => n27902, A => n5301, B => 
                           n26849, ZN => n5300);
   U6621 : AND3_X1 port map( A1 => n26624, A2 => n28446, A3 => n26246, ZN => 
                           n26626);
   U6622 : OAI22_X1 port map( A1 => n4411, A2 => n27041, B1 => n28783, B2 => 
                           n28130, ZN => n25555);
   U6623 : AOI21_X1 port map( B1 => n25506, B2 => n25505, A => n25504, ZN => 
                           n6857);
   U6624 : OR2_X1 port map( A1 => n7828, A2 => n7635, ZN => n8203);
   U6625 : INV_X1 port map( A => n8207, ZN => n3447);
   U6626 : INV_X1 port map( A => n7318, ZN => n6384);
   U6627 : OR2_X1 port map( A1 => n7349, A2 => n8158, ZN => n2944);
   U6628 : AND2_X1 port map( A1 => n7288, A2 => n4856, ZN => n2624);
   U6629 : AND2_X1 port map( A1 => n7499, A2 => n7500, ZN => n8589);
   U6630 : AND2_X1 port map( A1 => n7986, A2 => n631, ZN => n7662);
   U6632 : NAND2_X1 port map( A1 => n5160, A2 => n9045, ZN => n5159);
   U6633 : OR2_X1 port map( A1 => n9041, A2 => n9243, ZN => n9244);
   U6634 : INV_X1 port map( A => n8941, ZN => n9566);
   U6635 : OR2_X1 port map( A1 => n8141, A2 => n7336, ZN => n7723);
   U6636 : INV_X1 port map( A => n8465, ZN => n8463);
   U6637 : INV_X1 port map( A => n7279, ZN => n2115);
   U6638 : INV_X1 port map( A => n7320, ZN => n5242);
   U6639 : INV_X1 port map( A => n8610, ZN => n8609);
   U6640 : INV_X1 port map( A => n8762, ZN => n9561);
   U6641 : OR2_X1 port map( A1 => n7550, A2 => n7330, ZN => n7789);
   U6642 : AND2_X1 port map( A1 => n7330, A2 => n7782, ZN => n2670);
   U6645 : INV_X1 port map( A => n7914, ZN => n3329);
   U6647 : NOR2_X1 port map( A1 => n6908, A2 => n29304, ZN => n6316);
   U6649 : AND2_X1 port map( A1 => n7585, A2 => n7303, ZN => n5558);
   U6650 : INV_X1 port map( A => n7664, ZN => n2099);
   U6651 : OR2_X1 port map( A1 => n7485, A2 => n7665, ZN => n7486);
   U6652 : OR2_X1 port map( A1 => n8873, A2 => n8877, ZN => n8532);
   U6653 : OR2_X1 port map( A1 => n7313, A2 => n7898, ZN => n6545);
   U6654 : AOI22_X1 port map( A1 => n8245, A2 => n8246, B1 => n8243, B2 => 
                           n8244, ZN => n5911);
   U6655 : OR2_X1 port map( A1 => n7924, A2 => n7626, ZN => n8218);
   U6656 : OR2_X1 port map( A1 => n7520, A2 => n29321, ZN => n5072);
   U6657 : INV_X1 port map( A => n8035, ZN => n7510);
   U6658 : OR2_X1 port map( A1 => n7376, A2 => n7692, ZN => n8242);
   U6659 : OR2_X1 port map( A1 => n8560, A2 => n8562, ZN => n8568);
   U6660 : AND2_X1 port map( A1 => n8490, A2 => n9095, ZN => n2977);
   U6661 : AND2_X1 port map( A1 => n8955, A2 => n8801, ZN => n8472);
   U6662 : OR2_X1 port map( A1 => n6908, A2 => n284, ZN => n2980);
   U6663 : INV_X1 port map( A => n9531, ZN => n6892);
   U6664 : AND2_X1 port map( A1 => n7258, A2 => n29629, ZN => n2170);
   U6665 : AND2_X1 port map( A1 => n8685, A2 => n8687, ZN => n4729);
   U6667 : INV_X1 port map( A => n8872, ZN => n9061);
   U6668 : AND2_X1 port map( A1 => n7216, A2 => n3301, ZN => n3300);
   U6669 : OR2_X1 port map( A1 => n8685, A2 => n8687, ZN => n9026);
   U6670 : INV_X1 port map( A => n8717, ZN => n4321);
   U6671 : OR2_X1 port map( A1 => n7594, A2 => n7870, ZN => n6801);
   U6672 : OR2_X1 port map( A1 => n7604, A2 => n7864, ZN => n3034);
   U6674 : OR2_X1 port map( A1 => n9227, A2 => n597, ZN => n8102);
   U6675 : OAI22_X1 port map( A1 => n8234, A2 => n7619, B1 => n6973, B2 => 
                           n7919, ZN => n6976);
   U6677 : INV_X1 port map( A => n7114, ZN => n8829);
   U6678 : OR2_X1 port map( A1 => n8827, A2 => n8192, ZN => n8464);
   U6679 : INV_X1 port map( A => n8327, ZN => n5594);
   U6680 : AND3_X1 port map( A1 => n8498, A2 => n8497, A3 => n8651, ZN => n3128
                           );
   U6681 : INV_X1 port map( A => n9029, ZN => n9027);
   U6682 : INV_X1 port map( A => n9034, ZN => n7714);
   U6685 : OR2_X1 port map( A1 => n7748, A2 => n7749, ZN => n2358);
   U6686 : OAI21_X1 port map( B1 => n8873, B2 => n8403, A => n8404, ZN => n3297
                           );
   U6687 : OR2_X1 port map( A1 => n7736, A2 => n7268, ZN => n3115);
   U6688 : AND2_X1 port map( A1 => n7792, A2 => n28149, ZN => n2546);
   U6690 : OR3_X1 port map( A1 => n8958, A2 => n8802, A3 => n8955, ZN => n8316)
                           ;
   U6691 : OR2_X1 port map( A1 => n8154, A2 => n7550, ZN => n3282);
   U6692 : INV_X1 port map( A => n8886, ZN => n8334);
   U6693 : INV_X1 port map( A => n8605, ZN => n2320);
   U6694 : OR2_X1 port map( A1 => n8914, A2 => n8669, ZN => n8512);
   U6695 : BUF_X1 port map( A => n8499, Z => n8652);
   U6696 : INV_X1 port map( A => n8499, ZN => n8656);
   U6697 : AOI21_X1 port map( B1 => n7383, B2 => n617, A => n3639, ZN => n6748)
                           ;
   U6698 : INV_X1 port map( A => n6718, ZN => n8753);
   U6699 : INV_X1 port map( A => n8320, ZN => n9533);
   U6700 : OAI211_X1 port map( C1 => n7989, C2 => n7990, A => n7988, B => n7987
                           , ZN => n8664);
   U6701 : OR2_X1 port map( A1 => n8211, A2 => n439, ZN => n3117);
   U6702 : OR2_X1 port map( A1 => n8811, A2 => n2238, ZN => n8679);
   U6703 : OR2_X1 port map( A1 => n8292, A2 => n8287, ZN => n2568);
   U6705 : AND2_X1 port map( A1 => n9196, A2 => n329, ZN => n9199);
   U6706 : INV_X1 port map( A => n8726, ZN => n8603);
   U6707 : INV_X1 port map( A => n8984, ZN => n8982);
   U6708 : OR2_X1 port map( A1 => n8157, A2 => n8156, ZN => n6874);
   U6709 : INV_X1 port map( A => n8966, ZN => n8837);
   U6710 : OAI21_X1 port map( B1 => n3225, B2 => n29241, A => n3224, ZN => 
                           n8255);
   U6711 : AOI22_X1 port map( A1 => n9168, A2 => n9167, B1 => n9165, B2 => 
                           n9166, ZN => n9312);
   U6712 : NOR2_X1 port map( A1 => n28638, A2 => n11197, ZN => n5916);
   U6713 : INV_X1 port map( A => n9684, ZN => n10146);
   U6714 : OR2_X1 port map( A1 => n10497, A2 => n10502, ZN => n11133);
   U6715 : XNOR2_X1 port map( A => n301, B => n9991, ZN => n5410);
   U6716 : AND2_X1 port map( A1 => n8734, A2 => n8733, ZN => n2983);
   U6717 : AND2_X1 port map( A1 => n9221, A2 => n9220, ZN => n2352);
   U6719 : OR2_X1 port map( A1 => n8855, A2 => n9070, ZN => n8862);
   U6720 : OAI211_X1 port map( C1 => n9012, C2 => n8910, A => n9015, B => n6147
                           , ZN => n8085);
   U6721 : INV_X1 port map( A => n11163, ZN => n3904);
   U6723 : XNOR2_X1 port map( A => n9312, B => n9991, ZN => n10373);
   U6724 : OR2_X1 port map( A1 => n10740, A2 => n582, ZN => n6703);
   U6725 : AND2_X1 port map( A1 => n28876, A2 => n11149, ZN => n10512);
   U6726 : OR2_X1 port map( A1 => n10806, A2 => n28627, ZN => n6360);
   U6727 : INV_X1 port map( A => n11778, ZN => n11553);
   U6728 : AND2_X1 port map( A1 => n10966, A2 => n10965, ZN => n4715);
   U6729 : OR2_X1 port map( A1 => n10872, A2 => n435, ZN => n2283);
   U6730 : OR2_X1 port map( A1 => n4908, A2 => n11094, ZN => n2464);
   U6731 : OAI21_X1 port map( B1 => n10505, B2 => n4383, A => n11121, ZN => 
                           n9914);
   U6732 : OR2_X1 port map( A1 => n10504, A2 => n10507, ZN => n3460);
   U6733 : INV_X1 port map( A => n29149, ZN => n3816);
   U6734 : INV_X1 port map( A => n12158, ZN => n12157);
   U6735 : AND2_X1 port map( A1 => n10713, A2 => n1834, ZN => n4553);
   U6736 : OR2_X1 port map( A1 => n4844, A2 => n11599, ZN => n4843);
   U6739 : OR2_X1 port map( A1 => n12058, A2 => n11795, ZN => n12060);
   U6740 : AND2_X1 port map( A1 => n28174, A2 => n29122, ZN => n6386);
   U6741 : AND2_X1 port map( A1 => n12236, A2 => n375, ZN => n5008);
   U6742 : INV_X1 port map( A => n11491, ZN => n12302);
   U6743 : OR2_X1 port map( A1 => n10713, A2 => n5672, ZN => n11131);
   U6744 : AND2_X1 port map( A1 => n11114, A2 => n11113, ZN => n5109);
   U6745 : OR2_X1 port map( A1 => n12109, A2 => n12110, ZN => n6282);
   U6746 : OR2_X1 port map( A1 => n10819, A2 => n10820, ZN => n3536);
   U6747 : OR2_X1 port map( A1 => n11152, A2 => n5150, ZN => n10802);
   U6748 : XNOR2_X1 port map( A => n10086, B => n10089, ZN => n6183);
   U6749 : XNOR2_X1 port map( A => n10085, B => n10090, ZN => n6184);
   U6750 : INV_X1 port map( A => n29078, ZN => n9348);
   U6751 : AND2_X1 port map( A1 => n4296, A2 => n2690, ZN => n2688);
   U6752 : INV_X1 port map( A => n11332, ZN => n4463);
   U6753 : INV_X1 port map( A => n11956, ZN => n5603);
   U6754 : OR2_X1 port map( A1 => n10972, A2 => n10970, ZN => n6368);
   U6755 : OR2_X1 port map( A1 => n11551, A2 => n11778, ZN => n5170);
   U6756 : INV_X1 port map( A => n11206, ZN => n5258);
   U6757 : AND2_X1 port map( A1 => n11754, A2 => n11536, ZN => n11756);
   U6758 : AND2_X1 port map( A1 => n10603, A2 => n10966, ZN => n3322);
   U6759 : INV_X1 port map( A => n12156, ZN => n12159);
   U6760 : INV_X1 port map( A => n12507, ZN => n6374);
   U6761 : AND2_X1 port map( A1 => n11955, A2 => n12257, ZN => n4018);
   U6762 : OAI21_X1 port map( B1 => n10637, B2 => n5281, A => n11093, ZN => 
                           n5280);
   U6763 : NOR2_X1 port map( A1 => n10431, A2 => n11207, ZN => n5281);
   U6764 : INV_X1 port map( A => n11640, ZN => n11401);
   U6765 : AND2_X1 port map( A1 => n12151, A2 => n12150, ZN => n3603);
   U6767 : AND2_X1 port map( A1 => n5533, A2 => n11193, ZN => n4903);
   U6768 : INV_X1 port map( A => n11458, ZN => n11874);
   U6769 : INV_X1 port map( A => n11980, ZN => n11809);
   U6770 : AND2_X1 port map( A1 => n6482, A2 => n10717, ZN => n11489);
   U6771 : OR2_X1 port map( A1 => n6411, A2 => n10851, ZN => n3934);
   U6772 : INV_X1 port map( A => n574, ZN => n3201);
   U6774 : INV_X1 port map( A => n13444, ZN => n12600);
   U6775 : OR2_X1 port map( A1 => n12156, A2 => n12158, ZN => n11512);
   U6776 : OR2_X1 port map( A1 => n10894, A2 => n11290, ZN => n6430);
   U6777 : OR2_X1 port map( A1 => n12177, A2 => n12181, ZN => n3604);
   U6778 : AND2_X1 port map( A1 => n12516, A2 => n12517, ZN => n11941);
   U6779 : OR2_X1 port map( A1 => n12270, A2 => n28202, ZN => n12075);
   U6781 : OAI21_X1 port map( B1 => n10883, B2 => n11086, A => n11212, ZN => 
                           n2143);
   U6782 : OR2_X1 port map( A1 => n10918, A2 => n2968, ZN => n10105);
   U6783 : INV_X1 port map( A => n13086, ZN => n11810);
   U6784 : INV_X1 port map( A => n3871, ZN => n4297);
   U6785 : OR2_X1 port map( A1 => n10113, A2 => n10946, ZN => n6373);
   U6786 : OR2_X1 port map( A1 => n10927, A2 => n10930, ZN => n2948);
   U6787 : OR2_X1 port map( A1 => n11487, A2 => n11787, ZN => n6480);
   U6788 : INV_X1 port map( A => n12077, ZN => n5947);
   U6789 : AND2_X1 port map( A1 => n12339, A2 => n12338, ZN => n12028);
   U6790 : OR2_X1 port map( A1 => n10648, A2 => n12338, ZN => n12030);
   U6791 : OR2_X1 port map( A1 => n11340, A2 => n11335, ZN => n11342);
   U6792 : OR2_X1 port map( A1 => n11344, A2 => n11345, ZN => n2580);
   U6793 : NOR2_X1 port map( A1 => n4105, A2 => n11505, ZN => n6132);
   U6794 : AND2_X1 port map( A1 => n12303, A2 => n11491, ZN => n11608);
   U6797 : OR2_X1 port map( A1 => n28568, A2 => n333, ZN => n4101);
   U6798 : OR2_X1 port map( A1 => n12155, A2 => n12150, ZN => n12099);
   U6799 : AND3_X1 port map( A1 => n7813, A2 => n28206, A3 => n10808, ZN => 
                           n4389);
   U6800 : INV_X1 port map( A => n12145, ZN => n11708);
   U6801 : AND2_X1 port map( A1 => n11417, A2 => n11648, ZN => n12142);
   U6802 : INV_X1 port map( A => n11599, ZN => n12204);
   U6803 : OR2_X1 port map( A1 => n10859, A2 => n11181, ZN => n9055);
   U6804 : OR2_X1 port map( A1 => n11043, A2 => n11260, ZN => n11051);
   U6805 : INV_X1 port map( A => n12284, ZN => n12279);
   U6806 : AND2_X1 port map( A1 => n11859, A2 => n11944, ZN => n11860);
   U6807 : INV_X1 port map( A => n12332, ZN => n12018);
   U6810 : INV_X1 port map( A => n12273, ZN => n4869);
   U6811 : OR2_X1 port map( A1 => n12346, A2 => n12338, ZN => n3592);
   U6812 : AND2_X1 port map( A1 => n12206, A2 => n12109, ZN => n11373);
   U6813 : AND2_X1 port map( A1 => n3113, A2 => n11316, ZN => n9502);
   U6814 : OR2_X1 port map( A1 => n10993, A2 => n10992, ZN => n2165);
   U6815 : OAI211_X1 port map( C1 => n10628, C2 => n3441, A => n2413, B => 
                           n6108, ZN => n2847);
   U6816 : INV_X1 port map( A => n11962, ZN => n12221);
   U6817 : OR2_X1 port map( A1 => n10569, A2 => n10795, ZN => n3103);
   U6818 : OR2_X1 port map( A1 => n6604, A2 => n10572, ZN => n10574);
   U6819 : INV_X1 port map( A => n12453, ZN => n13080);
   U6820 : XNOR2_X1 port map( A => n13445, B => n3374, ZN => n12262);
   U6821 : INV_X1 port map( A => n2981, ZN => n4502);
   U6822 : INV_X1 port map( A => n4298, ZN => n12064);
   U6823 : INV_X1 port map( A => n14600, ZN => n6048);
   U6824 : INV_X1 port map( A => n13523, ZN => n12816);
   U6825 : AOI21_X1 port map( B1 => n12315, B2 => n5464, A => n11615, ZN => 
                           n5463);
   U6826 : OR2_X1 port map( A1 => n14146, A2 => n3860, ZN => n3859);
   U6827 : INV_X1 port map( A => n12799, ZN => n12568);
   U6828 : INV_X1 port map( A => n12632, ZN => n12603);
   U6829 : INV_X1 port map( A => n13521, ZN => n13520);
   U6831 : INV_X1 port map( A => n14262, ZN => n3071);
   U6832 : OR2_X1 port map( A1 => n11682, A2 => n12236, ZN => n10676);
   U6833 : OR2_X1 port map( A1 => n5578, A2 => n12232, ZN => n10674);
   U6834 : INV_X1 port map( A => n12813, ZN => n13144);
   U6835 : AND2_X1 port map( A1 => n5058, A2 => n14376, ZN => n5057);
   U6836 : OR2_X1 port map( A1 => n14434, A2 => n14433, ZN => n12887);
   U6837 : OR2_X1 port map( A1 => n14842, A2 => n15285, ZN => n5931);
   U6838 : OR2_X1 port map( A1 => n14695, A2 => n15285, ZN => n2893);
   U6839 : INV_X1 port map( A => n14047, ZN => n6011);
   U6840 : OAI211_X1 port map( C1 => n2112, C2 => n28804, A => n2111, B => 
                           n2110, ZN => n14621);
   U6841 : OR2_X1 port map( A1 => n13868, A2 => n28805, ZN => n3228);
   U6842 : OR2_X1 port map( A1 => n14195, A2 => n14193, ZN => n4500);
   U6843 : OR2_X1 port map( A1 => n14451, A2 => n14178, ZN => n13932);
   U6844 : NOR2_X1 port map( A1 => n14294, A2 => n14295, ZN => n13808);
   U6845 : INV_X1 port map( A => n13306, ZN => n14291);
   U6846 : AND2_X1 port map( A1 => n13893, A2 => n13892, ZN => n4836);
   U6847 : INV_X1 port map( A => n15388, ZN => n6517);
   U6848 : AND2_X1 port map( A1 => n14142, A2 => n2000, ZN => n13410);
   U6850 : AND2_X1 port map( A1 => n14773, A2 => n14807, ZN => n14555);
   U6851 : AND2_X1 port map( A1 => n15103, A2 => n15420, ZN => n5381);
   U6853 : INV_X1 port map( A => n13639, ZN => n13637);
   U6854 : INV_X1 port map( A => n2974, ZN => n2874);
   U6857 : INV_X1 port map( A => n14373, ZN => n13726);
   U6858 : INV_X1 port map( A => n14763, ZN => n4162);
   U6859 : OR2_X1 port map( A1 => n15208, A2 => n14928, ZN => n13785);
   U6860 : AOI21_X1 port map( B1 => n28195, B2 => n6854, A => n28196, ZN => 
                           n6853);
   U6861 : INV_X1 port map( A => n14944, ZN => n6854);
   U6862 : INV_X1 port map( A => n15046, ZN => n15226);
   U6863 : OR2_X1 port map( A1 => n2974, A2 => n29589, ZN => n3379);
   U6866 : OR2_X1 port map( A1 => n4436, A2 => n28805, ZN => n4431);
   U6867 : AND2_X1 port map( A1 => n29320, A2 => n293, ZN => n3868);
   U6868 : AND3_X1 port map( A1 => n3843, A2 => n13854, A3 => n4840, ZN => 
                           n5598);
   U6869 : OR2_X1 port map( A1 => n14839, A2 => n4359, ZN => n4358);
   U6870 : INV_X1 port map( A => n14969, ZN => n14793);
   U6871 : INV_X1 port map( A => n5378, ZN => n14397);
   U6873 : INV_X1 port map( A => n14534, ZN => n15460);
   U6874 : INV_X1 port map( A => n15503, ZN => n15497);
   U6875 : INV_X1 port map( A => n14922, ZN => n15500);
   U6876 : INV_X1 port map( A => n13785, ZN => n14796);
   U6877 : INV_X1 port map( A => n16388, ZN => n16471);
   U6878 : OAI21_X1 port map( B1 => n2800, B2 => n15209, A => n15201, ZN => 
                           n2691);
   U6880 : AND3_X1 port map( A1 => n14746, A2 => n14747, A3 => n14998, ZN => 
                           n4720);
   U6881 : INV_X1 port map( A => n13796, ZN => n6640);
   U6882 : OR2_X1 port map( A1 => n15238, A2 => n15239, ZN => n14220);
   U6883 : AND2_X1 port map( A1 => n14415, A2 => n6232, ZN => n6231);
   U6884 : INV_X1 port map( A => n14826, ZN => n15430);
   U6885 : OR2_X1 port map( A1 => n4893, A2 => n14354, ZN => n14013);
   U6886 : OR2_X1 port map( A1 => n13815, A2 => n14408, ZN => n4284);
   U6887 : AND2_X1 port map( A1 => n14969, A2 => n14972, ZN => n14792);
   U6888 : OR2_X1 port map( A1 => n15361, A2 => n4992, ZN => n15363);
   U6889 : AND2_X1 port map( A1 => n15486, A2 => n15491, ZN => n6245);
   U6890 : INV_X1 port map( A => n15071, ZN => n5229);
   U6891 : AND2_X1 port map( A1 => n15182, A2 => n15190, ZN => n14645);
   U6892 : AOI22_X1 port map( A1 => n13799, A2 => n14063, B1 => n14064, B2 => 
                           n13798, ZN => n3564);
   U6893 : OR2_X1 port map( A1 => n13817, A2 => n14303, ZN => n5283);
   U6894 : INV_X1 port map( A => n14533, ZN => n14649);
   U6896 : AND2_X1 port map( A1 => n3348, A2 => n14346, ZN => n4121);
   U6897 : MUX2_X1 port map( A => n15108, B => n15410, S => n14937, Z => n5788)
                           ;
   U6898 : OR2_X1 port map( A1 => n15109, A2 => n15406, ZN => n5785);
   U6900 : OR2_X1 port map( A1 => n15310, A2 => n15306, ZN => n5189);
   U6902 : INV_X1 port map( A => n15155, ZN => n2203);
   U6903 : NAND2_X1 port map( A1 => n14733, A2 => n15248, ZN => n4622);
   U6904 : OR2_X1 port map( A1 => n14730, A2 => n15246, ZN => n4619);
   U6905 : INV_X1 port map( A => n17232, ZN => n4478);
   U6906 : AND2_X1 port map( A1 => n3926, A2 => n15224, ZN => n3925);
   U6907 : OR2_X1 port map( A1 => n13840, A2 => n14007, ZN => n2561);
   U6908 : OR2_X1 port map( A1 => n14134, A2 => n14342, ZN => n6235);
   U6909 : OR2_X1 port map( A1 => n3799, A2 => n3798, ZN => n13732);
   U6910 : OR2_X1 port map( A1 => n15369, A2 => n14737, ZN => n4458);
   U6911 : NOR2_X1 port map( A1 => n14761, A2 => n14248, ZN => n2729);
   U6912 : AOI21_X1 port map( B1 => n14917, B2 => n15489, A => n14916, ZN => 
                           n5643);
   U6913 : AND2_X1 port map( A1 => n6457, A2 => n15316, ZN => n6456);
   U6914 : OR2_X1 port map( A1 => n16888, A2 => n17139, ZN => n2185);
   U6915 : XNOR2_X1 port map( A => n15281, B => n15280, ZN => n5714);
   U6916 : OAI211_X1 port map( C1 => n15243, C2 => n15355, A => n6675, B => 
                           n6674, ZN => n6673);
   U6917 : AOI21_X1 port map( B1 => n14149, B2 => n15361, A => n14751, ZN => 
                           n6672);
   U6918 : XNOR2_X1 port map( A => n2700, B => n16176, ZN => n16591);
   U6920 : AND2_X1 port map( A1 => n15420, A2 => n15101, ZN => n14935);
   U6921 : XNOR2_X1 port map( A => n16556, B => n27422, ZN => n15568);
   U6922 : XNOR2_X1 port map( A => n16084, B => n27730, ZN => n15630);
   U6923 : INV_X1 port map( A => n15781, ZN => n15654);
   U6924 : INV_X1 port map( A => n17555, ZN => n17220);
   U6925 : OAI21_X1 port map( B1 => n15084, B2 => n4407, A => n13305, ZN => 
                           n13313);
   U6926 : INV_X1 port map( A => n3374, ZN => n3138);
   U6927 : XNOR2_X1 port map( A => n16606, B => n5513, ZN => n6159);
   U6928 : OR2_X1 port map( A1 => n15326, A2 => n15327, ZN => n3626);
   U6929 : OR2_X1 port map( A1 => n14540, A2 => n15202, ZN => n14541);
   U6930 : OAI21_X1 port map( B1 => n14964, B2 => n14539, A => n14963, ZN => 
                           n14542);
   U6931 : AND2_X1 port map( A1 => n17556, A2 => n17553, ZN => n4099);
   U6932 : OR2_X1 port map( A1 => n17455, A2 => n16797, ZN => n5987);
   U6933 : OR2_X1 port map( A1 => n17155, A2 => n28564, ZN => n5226);
   U6934 : INV_X1 port map( A => n18467, ZN => n17915);
   U6935 : INV_X1 port map( A => n17138, ZN => n6727);
   U6936 : AND3_X1 port map( A1 => n16612, A2 => n17497, A3 => n17498, ZN => 
                           n18222);
   U6937 : OAI21_X1 port map( B1 => n17530, B2 => n17531, A => n17529, ZN => 
                           n18224);
   U6938 : AND2_X1 port map( A1 => n17830, A2 => n4270, ZN => n5808);
   U6939 : AND2_X1 port map( A1 => n17412, A2 => n16831, ZN => n2485);
   U6940 : INV_X1 port map( A => n17745, ZN => n2499);
   U6941 : AND2_X1 port map( A1 => n17864, A2 => n18527, ZN => n18541);
   U6943 : AOI21_X1 port map( B1 => n18215, B2 => n18216, A => n520, ZN => 
                           n17868);
   U6945 : INV_X1 port map( A => n18526, ZN => n5909);
   U6947 : OR2_X1 port map( A1 => n18506, A2 => n18215, ZN => n5157);
   U6948 : NOR2_X1 port map( A1 => n18215, A2 => n520, ZN => n18214);
   U6949 : AND2_X1 port map( A1 => n18018, A2 => n18251, ZN => n2316);
   U6950 : AND2_X1 port map( A1 => n1888, A2 => n18020, ZN => n2814);
   U6951 : OR2_X1 port map( A1 => n18471, A2 => n18469, ZN => n17659);
   U6952 : INV_X1 port map( A => n2819, ZN => n17709);
   U6953 : NOR2_X1 port map( A1 => n18539, A2 => n18260, ZN => n2707);
   U6955 : OR2_X1 port map( A1 => n5695, A2 => n17540, ZN => n5694);
   U6956 : INV_X1 port map( A => n17261, ZN => n16779);
   U6957 : OR2_X1 port map( A1 => n3880, A2 => n17269, ZN => n2985);
   U6958 : OAI211_X1 port map( C1 => n16802, C2 => n534, A => n16727, B => 
                           n5585, ZN => n17695);
   U6960 : INV_X1 port map( A => n17347, ZN => n17345);
   U6961 : OR2_X1 port map( A1 => n17439, A2 => n17437, ZN => n5639);
   U6962 : XNOR2_X1 port map( A => n16464, B => n4977, ZN => n16428);
   U6963 : AND2_X1 port map( A1 => n16762, A2 => n5398, ZN => n4787);
   U6964 : INV_X1 port map( A => n17046, ZN => n6180);
   U6965 : MUX2_X1 port map( A => n16678, B => n16677, S => n17456, Z => n16932
                           );
   U6966 : OR2_X1 port map( A1 => n18595, A2 => n17834, ZN => n3450);
   U6967 : INV_X1 port map( A => n17695, ZN => n17803);
   U6968 : INV_X1 port map( A => n17719, ZN => n18524);
   U6969 : INV_X1 port map( A => n18529, ZN => n18539);
   U6970 : AND2_X1 port map( A1 => n18538, A2 => n18537, ZN => n18054);
   U6971 : AND2_X1 port map( A1 => n17942, A2 => n17872, ZN => n17940);
   U6972 : AND2_X1 port map( A1 => n5383, A2 => n18379, ZN => n17997);
   U6973 : OR2_X1 port map( A1 => n2985, A2 => n16996, ZN => n3343);
   U6974 : INV_X1 port map( A => n17402, ZN => n4571);
   U6975 : OR2_X1 port map( A1 => n14915, A2 => n17402, ZN => n4112);
   U6977 : NOR2_X1 port map( A1 => n20147, A2 => n4877, ZN => n19010);
   U6978 : OAI21_X1 port map( B1 => n17390, B2 => n424, A => n3090, ZN => n4040
                           );
   U6980 : AND2_X1 port map( A1 => n17562, A2 => n17314, ZN => n4763);
   U6981 : OR2_X1 port map( A1 => n17551, A2 => n17548, ZN => n17245);
   U6982 : AND3_X1 port map( A1 => n17569, A2 => n17229, A3 => n29098, ZN => 
                           n17230);
   U6983 : AND2_X1 port map( A1 => n16547, A2 => n16548, ZN => n16552);
   U6984 : OR2_X1 port map( A1 => n16550, A2 => n17508, ZN => n16551);
   U6985 : INV_X1 port map( A => n3812, ZN => n16661);
   U6986 : AND2_X1 port map( A1 => n18380, A2 => n18379, ZN => n17165);
   U6987 : INV_X1 port map( A => n17969, ZN => n18238);
   U6989 : INV_X1 port map( A => n6526, ZN => n18600);
   U6990 : OR2_X1 port map( A1 => n18354, A2 => n18353, ZN => n5084);
   U6991 : OR2_X1 port map( A1 => n18355, A2 => n18353, ZN => n5589);
   U6992 : INV_X1 port map( A => n17126, ZN => n3471);
   U6993 : AND2_X1 port map( A1 => n18449, A2 => n18195, ZN => n18454);
   U6994 : OAI21_X1 port map( B1 => n16833, B2 => n16834, A => n16916, ZN => 
                           n16835);
   U6995 : OR2_X1 port map( A1 => n17518, A2 => n17516, ZN => n17108);
   U6996 : INV_X1 port map( A => n18260, ZN => n2151);
   U6997 : OR2_X1 port map( A1 => n4706, A2 => n17451, ZN => n4702);
   U6998 : INV_X1 port map( A => n5759, ZN => n19585);
   U6999 : AND2_X1 port map( A1 => n17978, A2 => n17979, ZN => n3439);
   U7000 : AOI21_X1 port map( B1 => n18500, B2 => n18213, A => n18216, ZN => 
                           n5692);
   U7001 : INV_X1 port map( A => n3597, ZN => n2758);
   U7002 : OR2_X1 port map( A1 => n18122, A2 => n18416, ZN => n3933);
   U7003 : OAI211_X1 port map( C1 => n2242, C2 => n17209, A => n2243, B => 
                           n2241, ZN => n18690);
   U7004 : AND2_X1 port map( A1 => n17837, A2 => n18591, ZN => n2242);
   U7005 : INV_X1 port map( A => n2855, ZN => n2123);
   U7006 : OR2_X1 port map( A1 => n18109, A2 => n17798, ZN => n18458);
   U7007 : OR2_X1 port map( A1 => n18456, A2 => n18107, ZN => n6038);
   U7008 : AND2_X1 port map( A1 => n6912, A2 => n17584, ZN => n17585);
   U7009 : OR2_X1 port map( A1 => n16907, A2 => n17037, ZN => n5999);
   U7010 : INV_X1 port map( A => n18180, ZN => n18444);
   U7011 : OR2_X1 port map( A1 => n17254, A2 => n17251, ZN => n5081);
   U7012 : INV_X1 port map( A => n18589, ZN => n18128);
   U7013 : OR2_X1 port map( A1 => n17802, A2 => n18422, ZN => n17823);
   U7014 : NOR2_X1 port map( A1 => n4707, A2 => n18215, ZN => n4450);
   U7015 : INV_X1 port map( A => n18248, ZN => n18406);
   U7016 : INV_X1 port map( A => n17858, ZN => n2694);
   U7017 : INV_X1 port map( A => n18081, ZN => n18523);
   U7018 : AND2_X1 port map( A1 => n18242, A2 => n18236, ZN => n17967);
   U7019 : INV_X1 port map( A => n18268, ZN => n18329);
   U7020 : AND2_X1 port map( A1 => n18261, A2 => n18268, ZN => n16930);
   U7021 : INV_X1 port map( A => n16718, ZN => n18451);
   U7023 : AND2_X1 port map( A1 => n18528, A2 => n17701, ZN => n17703);
   U7024 : AND3_X1 port map( A1 => n21066, A2 => n21065, A3 => n21064, ZN => 
                           n21663);
   U7026 : OAI211_X1 port map( C1 => n18239, C2 => n29034, A => n2785, B => 
                           n2784, ZN => n19354);
   U7027 : OR2_X1 port map( A1 => n18230, A2 => n1887, ZN => n2723);
   U7028 : AND2_X1 port map( A1 => n21091, A2 => n29134, ZN => n20149);
   U7029 : AND3_X1 port map( A1 => n4412, A2 => n18371, A3 => n18337, ZN => 
                           n5164);
   U7030 : XNOR2_X1 port map( A => n18735, B => n6653, ZN => n18569);
   U7031 : INV_X1 port map( A => n20032, ZN => n3717);
   U7032 : OR2_X1 port map( A1 => n16867, A2 => n5059, ZN => n5060);
   U7033 : INV_X1 port map( A => n20109, ZN => n20320);
   U7034 : INV_X1 port map( A => n19669, ZN => n18726);
   U7035 : INV_X1 port map( A => n3232, ZN => n4881);
   U7036 : OR2_X1 port map( A1 => n17212, A2 => n17211, ZN => n3719);
   U7037 : INV_X1 port map( A => n19491, ZN => n6489);
   U7038 : AOI21_X1 port map( B1 => n18525, B2 => n18526, A => n5325, ZN => 
                           n5324);
   U7039 : INV_X1 port map( A => n16990, ZN => n19525);
   U7040 : INV_X1 port map( A => n19687, ZN => n5952);
   U7041 : OR2_X1 port map( A1 => n20088, A2 => n20090, ZN => n4006);
   U7042 : INV_X1 port map( A => n20563, ZN => n20395);
   U7043 : AND2_X1 port map( A1 => n20064, A2 => n413, ZN => n20068);
   U7044 : OR2_X1 port map( A1 => n20374, A2 => n19841, ZN => n20070);
   U7045 : AND2_X1 port map( A1 => n19814, A2 => n19815, ZN => n4657);
   U7046 : NOR2_X1 port map( A1 => n2641, A2 => n21442, ZN => n2640);
   U7047 : INV_X1 port map( A => n2735, ZN => n20093);
   U7048 : OR2_X1 port map( A1 => n20875, A2 => n20814, ZN => n21265);
   U7049 : INV_X1 port map( A => n20155, ZN => n19773);
   U7050 : OAI21_X1 port map( B1 => n28186, B2 => n20334, A => n3186, ZN => 
                           n20007);
   U7051 : AND2_X1 port map( A1 => n20966, A2 => n21218, ZN => n20999);
   U7052 : OR2_X1 port map( A1 => n20200, A2 => n20205, ZN => n4338);
   U7053 : AND2_X1 port map( A1 => n20121, A2 => n20120, ZN => n20891);
   U7054 : AND2_X1 port map( A1 => n20205, A2 => n20201, ZN => n2978);
   U7055 : OR2_X1 port map( A1 => n20148, A2 => n20146, ZN => n5794);
   U7056 : OR2_X1 port map( A1 => n5334, A2 => n20580, ZN => n5333);
   U7057 : INV_X1 port map( A => n20404, ZN => n20554);
   U7059 : INV_X1 port map( A => n21156, ZN => n3401);
   U7060 : AOI22_X1 port map( A1 => n5935, A2 => n20446, B1 => n5934, B2 => 
                           n5933, ZN => n6771);
   U7061 : AND3_X1 port map( A1 => n21587, A2 => n20591, A3 => n3789, ZN => 
                           n20594);
   U7062 : OR2_X1 port map( A1 => n20404, A2 => n20549, ZN => n20408);
   U7063 : OR2_X1 port map( A1 => n20401, A2 => n20208, ZN => n19743);
   U7064 : NOR2_X1 port map( A1 => n20498, A2 => n1624, ZN => n20008);
   U7065 : AND2_X1 port map( A1 => n4148, A2 => n21334, ZN => n2307);
   U7066 : OR2_X1 port map( A1 => n20226, A2 => n1624, ZN => n5385);
   U7067 : OR2_X1 port map( A1 => n21664, A2 => n21665, ZN => n3692);
   U7068 : INV_X1 port map( A => n5151, ZN => n21662);
   U7069 : OR2_X1 port map( A1 => n4312, A2 => n4309, ZN => n4308);
   U7070 : OR2_X1 port map( A1 => n20513, A2 => n20509, ZN => n4909);
   U7071 : AND2_X1 port map( A1 => n20623, A2 => n20626, ZN => n6059);
   U7072 : AOI21_X1 port map( B1 => n20500, B2 => n20504, A => n3761, ZN => 
                           n6635);
   U7074 : INV_X1 port map( A => n5106, ZN => n19860);
   U7075 : NOR2_X1 port map( A1 => n21541, A2 => n21539, ZN => n21499);
   U7076 : OR2_X1 port map( A1 => n21500, A2 => n28611, ZN => n20779);
   U7078 : AND2_X1 port map( A1 => n20645, A2 => n21063, ZN => n5782);
   U7079 : NAND2_X1 port map( A1 => n4874, A2 => n4878, ZN => n20954);
   U7080 : AND2_X1 port map( A1 => n21389, A2 => n21387, ZN => n2572);
   U7081 : AND2_X1 port map( A1 => n19993, A2 => n20165, ZN => n19991);
   U7083 : INV_X1 port map( A => n6314, ZN => n6311);
   U7084 : OR2_X1 port map( A1 => n21265, A2 => n21269, ZN => n6396);
   U7085 : OR2_X1 port map( A1 => n21481, A2 => n21577, ZN => n6698);
   U7086 : INV_X1 port map( A => n19505, ZN => n6842);
   U7088 : OR2_X1 port map( A1 => n20107, A2 => n20106, ZN => n3126);
   U7089 : OR2_X1 port map( A1 => n20183, A2 => n20182, ZN => n3076);
   U7090 : NOR2_X1 port map( A1 => n21615, A2 => n2339, ZN => n2338);
   U7091 : INV_X1 port map( A => n21610, ZN => n2339);
   U7092 : INV_X1 port map( A => n21163, ZN => n21619);
   U7093 : OR2_X1 port map( A1 => n21601, A2 => n21596, ZN => n21597);
   U7094 : OR2_X1 port map( A1 => n19417, A2 => n20688, ZN => n19418);
   U7096 : OR2_X1 port map( A1 => n20746, A2 => n20858, ZN => n4959);
   U7097 : OR2_X1 port map( A1 => n20644, A2 => n5783, ZN => n4267);
   U7098 : INV_X1 port map( A => n20833, ZN => n21654);
   U7099 : OR2_X1 port map( A1 => n20217, A2 => n5303, ZN => n2799);
   U7101 : INV_X1 port map( A => n21140, ZN => n20851);
   U7102 : AOI21_X1 port map( B1 => n19779, B2 => n29146, A => n20084, ZN => 
                           n19780);
   U7103 : OR2_X1 port map( A1 => n21311, A2 => n21306, ZN => n20768);
   U7104 : OR2_X1 port map( A1 => n21265, A2 => n29553, ZN => n6425);
   U7105 : OR2_X1 port map( A1 => n19058, A2 => n20174, ZN => n19009);
   U7107 : AND2_X1 port map( A1 => n19966, A2 => n21032, ZN => n2091);
   U7108 : INV_X1 port map( A => n5194, ZN => n19965);
   U7109 : INV_X1 port map( A => n5827, ZN => n21421);
   U7111 : NOR2_X1 port map( A1 => n20954, A2 => n20953, ZN => n21934);
   U7112 : AND2_X1 port map( A1 => n3560, A2 => n3559, ZN => n21936);
   U7113 : OR2_X1 port map( A1 => n18787, A2 => n2804, ZN => n2803);
   U7114 : OR2_X1 port map( A1 => n22026, A2 => n22290, ZN => n3548);
   U7115 : INV_X1 port map( A => n22618, ZN => n6863);
   U7116 : BUF_X1 port map( A => n21625, Z => n5339);
   U7117 : OR2_X1 port map( A1 => n20600, A2 => n386, ZN => n4933);
   U7118 : INV_X1 port map( A => n20362, ZN => n2830);
   U7119 : AOI21_X1 port map( B1 => n6533, B2 => n6532, A => n21106, ZN => 
                           n6531);
   U7120 : INV_X1 port map( A => n21029, ZN => n6533);
   U7121 : OR2_X1 port map( A1 => n20239, A2 => n6512, ZN => n20003);
   U7122 : INV_X1 port map( A => n21461, ZN => n5176);
   U7123 : INV_X1 port map( A => n21638, ZN => n21631);
   U7125 : OR2_X1 port map( A1 => n20865, A2 => n20864, ZN => n21494);
   U7127 : OR2_X1 port map( A1 => n5560, A2 => n4877, ZN => n6894);
   U7128 : OR2_X1 port map( A1 => n21113, A2 => n5953, ZN => n5544);
   U7129 : INV_X1 port map( A => n21464, ZN => n21560);
   U7130 : OAI21_X1 port map( B1 => n5782, B2 => n20646, A => n5781, ZN => 
                           n20721);
   U7132 : INV_X1 port map( A => n5273, ZN => n21439);
   U7133 : AOI22_X1 port map( A1 => n20232, A2 => n383, B1 => n20231, B2 => 
                           n19032, ZN => n5273);
   U7134 : NOR2_X1 port map( A1 => n21655, A2 => n21657, ZN => n21443);
   U7135 : INV_X1 port map( A => n3954, ZN => n3952);
   U7136 : INV_X1 port map( A => n21534, ZN => n21198);
   U7137 : INV_X1 port map( A => n21519, ZN => n21180);
   U7138 : XNOR2_X1 port map( A => n21825, B => n3380, ZN => n3222);
   U7139 : INV_X1 port map( A => n22464, ZN => n4862);
   U7140 : INV_X1 port map( A => n22337, ZN => n21889);
   U7141 : INV_X1 port map( A => n22800, ZN => n20214);
   U7142 : XNOR2_X1 port map( A => n29549, B => n5797, ZN => n22706);
   U7143 : INV_X1 port map( A => n3643, ZN => n5797);
   U7144 : AND2_X1 port map( A1 => n339, A2 => n23772, ZN => n23488);
   U7145 : INV_X1 port map( A => n21872, ZN => n2752);
   U7146 : XNOR2_X1 port map( A => n22204, B => n4565, ZN => n22206);
   U7147 : INV_X1 port map( A => n21789, ZN => n4565);
   U7148 : OR2_X1 port map( A1 => n23741, A2 => n29564, ZN => n6472);
   U7149 : OR2_X1 port map( A1 => n21462, A2 => n20841, ZN => n3620);
   U7150 : OAI21_X1 port map( B1 => n21568, B2 => n21460, A => n6247, ZN => 
                           n3621);
   U7151 : OR2_X1 port map( A1 => n20276, A2 => n6016, ZN => n6015);
   U7152 : AOI21_X1 port map( B1 => n1974, B2 => n20271, A => n2668, ZN => 
                           n2667);
   U7153 : OR2_X1 port map( A1 => n4071, A2 => n21749, ZN => n6528);
   U7154 : AND2_X1 port map( A1 => n23303, A2 => n4178, ZN => n5697);
   U7155 : INV_X1 port map( A => n4178, ZN => n5699);
   U7156 : INV_X1 port map( A => n2637, ZN => n21894);
   U7157 : OR2_X1 port map( A1 => n23738, A2 => n23827, ZN => n3940);
   U7158 : AND2_X1 port map( A1 => n23769, A2 => n28554, ZN => n5237);
   U7159 : NOR2_X1 port map( A1 => n23250, A2 => n23406, ZN => n5042);
   U7160 : INV_X1 port map( A => n23777, ZN => n23514);
   U7161 : BUF_X1 port map( A => n23167, Z => n23169);
   U7163 : INV_X1 port map( A => n23656, ZN => n4772);
   U7164 : INV_X1 port map( A => n24269, ZN => n2937);
   U7165 : NOR2_X1 port map( A1 => n24726, A2 => n24596, ZN => n5767);
   U7166 : OR2_X1 port map( A1 => n5741, A2 => n5448, ZN => n23191);
   U7167 : INV_X1 port map( A => n407, ZN => n2281);
   U7168 : INV_X1 port map( A => n4086, ZN => n4429);
   U7169 : INV_X1 port map( A => n24503, ZN => n6600);
   U7170 : OR2_X1 port map( A1 => n23221, A2 => n6099, ZN => n5552);
   U7171 : OR2_X1 port map( A1 => n24437, A2 => n24436, ZN => n24121);
   U7172 : AND2_X1 port map( A1 => n22977, A2 => n23250, ZN => n23746);
   U7173 : NOR2_X1 port map( A1 => n24288, A2 => n24596, ZN => n24598);
   U7174 : NOR2_X1 port map( A1 => n4020, A2 => n29018, ZN => n4019);
   U7175 : AND2_X1 port map( A1 => n23768, A2 => n23767, ZN => n6358);
   U7176 : OR2_X1 port map( A1 => n2779, A2 => n23651, ZN => n3135);
   U7177 : AOI21_X1 port map( B1 => n22949, B2 => n23398, A => n23736, ZN => 
                           n22010);
   U7179 : NOR2_X1 port map( A1 => n23005, A2 => n23787, ZN => n6081);
   U7180 : INV_X1 port map( A => n23408, ZN => n2239);
   U7181 : INV_X1 port map( A => n24447, ZN => n24761);
   U7182 : INV_X1 port map( A => n23772, ZN => n23778);
   U7183 : INV_X1 port map( A => n24735, ZN => n3310);
   U7185 : OR2_X1 port map( A1 => n23735, A2 => n2141, ZN => n3502);
   U7186 : INV_X1 port map( A => n23790, ZN => n23320);
   U7187 : OR2_X1 port map( A1 => n24097, A2 => n24098, ZN => n3599);
   U7188 : INV_X1 port map( A => n24676, ZN => n6406);
   U7189 : OR2_X1 port map( A1 => n23344, A2 => n23339, ZN => n6195);
   U7190 : OAI211_X1 port map( C1 => n23146, C2 => n4872, A => n4892, B => 
                           n4891, ZN => n24295);
   U7191 : NAND2_X1 port map( A1 => n24610, A2 => n24614, ZN => n6746);
   U7192 : OR2_X1 port map( A1 => n23441, A2 => n2842, ZN => n23092);
   U7193 : NAND2_X1 port map( A1 => n24655, A2 => n2810, ZN => n24656);
   U7194 : OR2_X1 port map( A1 => n23205, A2 => n24555, ZN => n22747);
   U7196 : OAI21_X1 port map( B1 => n3519, B2 => n407, A => n3518, ZN => n4175)
                           ;
   U7197 : INV_X1 port map( A => n5591, ZN => n3519);
   U7198 : INV_X1 port map( A => n4917, ZN => n22869);
   U7199 : OR2_X1 port map( A1 => n23457, A2 => n23460, ZN => n23464);
   U7200 : OR2_X1 port map( A1 => n23099, A2 => n23418, ZN => n23100);
   U7202 : AND2_X1 port map( A1 => n24666, A2 => n24383, ZN => n24315);
   U7203 : NOR2_X1 port map( A1 => n4851, A2 => n4232, ZN => n4602);
   U7204 : NOR2_X1 port map( A1 => n24592, A2 => n24591, ZN => n24279);
   U7205 : AND2_X1 port map( A1 => n3612, A2 => n23096, ZN => n22929);
   U7206 : INV_X1 port map( A => n24589, ZN => n2997);
   U7207 : AND2_X1 port map( A1 => n24728, A2 => n24595, ZN => n5768);
   U7208 : INV_X1 port map( A => n24726, ZN => n24291);
   U7209 : INV_X1 port map( A => n24479, ZN => n24210);
   U7210 : INV_X1 port map( A => n23867, ZN => n24714);
   U7211 : NOR2_X1 port map( A1 => n24700, A2 => n24428, ZN => n24429);
   U7212 : INV_X1 port map( A => n23435, ZN => n3986);
   U7213 : AND2_X1 port map( A1 => n28524, A2 => n24716, ZN => n24106);
   U7214 : INV_X1 port map( A => n24713, ZN => n24412);
   U7215 : AND2_X1 port map( A1 => n24331, A2 => n2134, ZN => n3630);
   U7216 : NOR2_X1 port map( A1 => n24631, A2 => n24532, ZN => n24227);
   U7217 : NOR2_X1 port map( A1 => n24383, A2 => n24666, ZN => n24075);
   U7218 : INV_X1 port map( A => n24800, ZN => n24802);
   U7219 : AND2_X1 port map( A1 => n23798, A2 => n23799, ZN => n6599);
   U7220 : AND2_X1 port map( A1 => n4125, A2 => n4124, ZN => n20656);
   U7221 : NOR2_X1 port map( A1 => n24637, A2 => n24636, ZN => n25797);
   U7222 : INV_X1 port map( A => n23599, ZN => n23597);
   U7223 : AND2_X1 port map( A1 => n24817, A2 => n24809, ZN => n24496);
   U7225 : INV_X1 port map( A => n2649, ZN => n24683);
   U7226 : OR2_X1 port map( A1 => n405, A2 => n2697, ZN => n3743);
   U7227 : INV_X1 port map( A => n4596, ZN => n4595);
   U7228 : NOR2_X1 port map( A1 => n24645, A2 => n24638, ZN => n2107);
   U7229 : INV_X1 port map( A => n24665, ZN => n4605);
   U7230 : INV_X1 port map( A => n23994, ZN => n24376);
   U7231 : OAI21_X1 port map( B1 => n6211, B2 => n23829, A => n2188, ZN => 
                           n22947);
   U7232 : NAND2_X1 port map( A1 => n23721, A2 => n23394, ZN => n4473);
   U7233 : OR2_X1 port map( A1 => n23287, A2 => n2202, ZN => n2612);
   U7234 : AND2_X1 port map( A1 => n6741, A2 => n24584, ZN => n22130);
   U7235 : INV_X1 port map( A => n24133, ZN => n23389);
   U7236 : INV_X1 port map( A => n24081, ZN => n24386);
   U7237 : INV_X1 port map( A => n24138, ZN => n25006);
   U7238 : INV_X1 port map( A => n25008, ZN => n24304);
   U7239 : AND2_X1 port map( A1 => n24757, A2 => n24756, ZN => n2865);
   U7240 : AND2_X1 port map( A1 => n24757, A2 => n24447, ZN => n2866);
   U7241 : AND2_X1 port map( A1 => n24800, A2 => n24502, ZN => n4335);
   U7242 : NOR2_X1 port map( A1 => n24789, A2 => n4576, ZN => n4575);
   U7246 : INV_X1 port map( A => n23004, ZN => n5350);
   U7247 : AND2_X1 port map( A1 => n3199, A2 => n23840, ZN => n5309);
   U7248 : OR2_X1 port map( A1 => n24758, A2 => n24447, ZN => n24448);
   U7249 : INV_X1 port map( A => n5168, ZN => n5137);
   U7250 : OR2_X1 port map( A1 => n23281, A2 => n23392, ZN => n5292);
   U7252 : NOR2_X1 port map( A1 => n29467, A2 => n26447, ZN => n26160);
   U7253 : OR2_X1 port map( A1 => n6422, A2 => n5633, ZN => n5632);
   U7255 : OR2_X1 port map( A1 => n26386, A2 => n27165, ZN => n3190);
   U7256 : OR2_X1 port map( A1 => n24708, A2 => n24707, ZN => n5750);
   U7257 : INV_X1 port map( A => n24963, ZN => n26120);
   U7258 : AND3_X1 port map( A1 => n24138, A2 => n24369, A3 => n25008, ZN => 
                           n24139);
   U7259 : OAI21_X1 port map( B1 => n26739, B2 => n25655, A => n26737, ZN => 
                           n5422);
   U7260 : NOR2_X1 port map( A1 => n25618, A2 => n280, ZN => n27392);
   U7261 : NOR2_X1 port map( A1 => n25404, A2 => n27395, ZN => n26463);
   U7262 : INV_X1 port map( A => n26447, ZN => n3498);
   U7263 : OR2_X1 port map( A1 => n26447, A2 => n26448, ZN => n3497);
   U7264 : OR2_X1 port map( A1 => n26920, A2 => n4820, ZN => n3066);
   U7265 : INV_X1 port map( A => n4820, ZN => n26173);
   U7266 : AND2_X1 port map( A1 => n26172, A2 => n26919, ZN => n26918);
   U7267 : OR2_X1 port map( A1 => n26366, A2 => n29293, ZN => n2139);
   U7268 : OR2_X1 port map( A1 => n27181, A2 => n25034, ZN => n26270);
   U7269 : XNOR2_X1 port map( A => n24918, B => n24919, ZN => n2145);
   U7270 : OAI211_X1 port map( C1 => n26858, C2 => n28487, A => n27138, B => 
                           n29633, ZN => n27688);
   U7271 : NOR2_X1 port map( A1 => n28536, A2 => n27131, ZN => n4080);
   U7272 : INV_X1 port map( A => n27175, ZN => n27173);
   U7273 : OAI211_X1 port map( C1 => n27073, C2 => n27072, A => n3786, B => 
                           n3785, ZN => n27080);
   U7274 : AOI21_X1 port map( B1 => n28101, B2 => n5036, A => n26747, ZN => 
                           n26635);
   U7275 : AND2_X1 port map( A1 => n5144, A2 => n26251, ZN => n26253);
   U7276 : OR2_X1 port map( A1 => n29482, A2 => n26995, ZN => n5144);
   U7277 : AND2_X1 port map( A1 => n26757, A2 => n29479, ZN => n6625);
   U7278 : NOR2_X1 port map( A1 => n28107, A2 => n28794, ZN => n28110);
   U7279 : OR2_X1 port map( A1 => n25665, A2 => n26723, ZN => n6288);
   U7281 : AND2_X1 port map( A1 => n29541, A2 => n623, ZN => n6621);
   U7282 : NOR2_X1 port map( A1 => n27362, A2 => n25358, ZN => n25360);
   U7283 : OR2_X1 port map( A1 => n27377, A2 => n27213, ZN => n4091);
   U7284 : OR2_X1 port map( A1 => n27213, A2 => n28393, ZN => n5374);
   U7285 : OR2_X1 port map( A1 => n5581, A2 => n27382, ZN => n4033);
   U7286 : OR2_X1 port map( A1 => n27394, A2 => n6685, ZN => n27396);
   U7287 : INV_X1 port map( A => n27425, ZN => n6738);
   U7288 : AOI21_X1 port map( B1 => n26171, B2 => n26782, A => n26917, ZN => 
                           n4816);
   U7289 : AND2_X1 port map( A1 => n29468, A2 => n449, ZN => n27446);
   U7290 : OAI211_X1 port map( C1 => n26926, C2 => n4400, A => n2050, B => 
                           n4399, ZN => n4823);
   U7291 : AOI21_X1 port map( B1 => n5505, B2 => n4402, A => n4401, ZN => n4400
                           );
   U7292 : OR2_X1 port map( A1 => n27498, A2 => n27493, ZN => n5605);
   U7293 : AOI21_X1 port map( B1 => n6768, B2 => n26935, A => n456, ZN => n6766
                           );
   U7294 : OAI21_X1 port map( B1 => n26562, B2 => n26561, A => n26457, ZN => 
                           n2966);
   U7295 : BUF_X1 port map( A => n27526, Z => n27505);
   U7296 : NOR2_X1 port map( A1 => n27524, A2 => n3067, ZN => n4164);
   U7297 : INV_X1 port map( A => n26151, ZN => n26921);
   U7298 : AND2_X1 port map( A1 => n6095, A2 => n27527, ZN => n27524);
   U7299 : OR2_X1 port map( A1 => n27286, A2 => n2438, ZN => n2437);
   U7300 : NOR2_X1 port map( A1 => n27304, A2 => n27306, ZN => n6226);
   U7301 : MUX2_X1 port map( A => n26261, B => n26260, S => n27168, Z => n26262
                           );
   U7302 : OAI21_X1 port map( B1 => n26381, B2 => n26426, A => n4944, ZN => 
                           n26277);
   U7303 : INV_X1 port map( A => n27628, ZN => n27617);
   U7304 : INV_X1 port map( A => n27614, ZN => n27627);
   U7305 : INV_X1 port map( A => n27650, ZN => n27636);
   U7306 : OR2_X1 port map( A1 => n28655, A2 => n27663, ZN => n5874);
   U7307 : AND2_X1 port map( A1 => n27165, A2 => n27166, ZN => n6185);
   U7308 : INV_X1 port map( A => n27662, ZN => n27676);
   U7309 : INV_X1 port map( A => n29117, ZN => n4250);
   U7310 : AND2_X1 port map( A1 => n26311, A2 => n26310, ZN => n6669);
   U7311 : OR2_X1 port map( A1 => n26867, A2 => n29048, ZN => n3220);
   U7312 : OR2_X1 port map( A1 => n29118, A2 => n27772, ZN => n4248);
   U7313 : INV_X1 port map( A => n27777, ZN => n27780);
   U7314 : NOR2_X1 port map( A1 => n27795, A2 => n27807, ZN => n27791);
   U7315 : OR3_X1 port map( A1 => n29232, A2 => n27790, A3 => n27817, ZN => 
                           n6902);
   U7316 : OR2_X1 port map( A1 => n27109, A2 => n26332, ZN => n3589);
   U7317 : AND2_X1 port map( A1 => n3791, A2 => n27859, ZN => n5294);
   U7318 : INV_X1 port map( A => n27855, ZN => n3791);
   U7319 : NOR2_X1 port map( A1 => n27855, A2 => n27859, ZN => n4536);
   U7320 : OR2_X1 port map( A1 => n27051, A2 => n28446, ZN => n3351);
   U7321 : AND2_X1 port map( A1 => n27925, A2 => n27244, ZN => n27934);
   U7322 : OR2_X1 port map( A1 => n28456, A2 => n27982, ZN => n3271);
   U7323 : NOR2_X1 port map( A1 => n4499, A2 => n398, ZN => n4498);
   U7324 : AOI21_X1 port map( B1 => n4411, B2 => n25968, A => n27003, ZN => 
                           n25970);
   U7325 : AND2_X1 port map( A1 => n29161, A2 => n376, ZN => n5017);
   U7326 : AND2_X1 port map( A1 => n28063, A2 => n28067, ZN => n28047);
   U7327 : OR2_X1 port map( A1 => n26761, A2 => n26754, ZN => n26238);
   U7328 : AND2_X1 port map( A1 => n28065, A2 => n28066, ZN => n28052);
   U7329 : INV_X1 port map( A => n28101, ZN => n5037);
   U7330 : NOR2_X1 port map( A1 => n28591, A2 => n28107, ZN => n3691);
   U7331 : INV_X1 port map( A => n2541, ZN => n3897);
   U7332 : INV_X1 port map( A => n3554, ZN => n5649);
   U7333 : INV_X1 port map( A => n3660, ZN => n4923);
   U7334 : INV_X1 port map( A => n3493, ZN => n3610);
   U7335 : INV_X1 port map( A => n27286, ZN => n27280);
   U7336 : INV_X1 port map( A => n27259, ZN => n5426);
   U7337 : AND3_X1 port map( A1 => n2267, A2 => n27570, A3 => n27569, ZN => 
                           Ciphertext(79));
   U7338 : OR2_X1 port map( A1 => n27227, A2 => n27732, ZN => n2792);
   U7339 : OR2_X1 port map( A1 => n26872, A2 => n27101, ZN => n2376);
   U7341 : OR2_X1 port map( A1 => n26544, A2 => n3378, ZN => n26550);
   U7342 : OAI21_X1 port map( B1 => n28438, B2 => n4998, A => n3571, ZN => 
                           n27246);
   U7343 : OR2_X1 port map( A1 => n28037, A2 => n26602, ZN => n5850);
   U7344 : OR3_X1 port map( A1 => n22140, A2 => n21627, A3 => n21624, ZN => 
                           n1940);
   U7345 : INV_X1 port map( A => n7867, ZN => n5149);
   U7347 : XNOR2_X1 port map( A => n13281, B => n13282, ZN => n14304);
   U7348 : INV_X1 port map( A => n29610, ZN => n4751);
   U7350 : INV_X1 port map( A => n20444, ZN => n5933);
   U7351 : INV_X1 port map( A => n26510, ZN => n5299);
   U7352 : INV_X1 port map( A => n27854, ZN => n5295);
   U7354 : INV_X1 port map( A => n20323, ZN => n2181);
   U7355 : XNOR2_X1 port map( A => n9389, B => n4716, ZN => n10687);
   U7356 : OR2_X1 port map( A1 => n21601, A2 => n21314, ZN => n1941);
   U7357 : OR2_X1 port map( A1 => n29594, A2 => n18421, ZN => n1942);
   U7359 : INV_X1 port map( A => n14399, ZN => n2549);
   U7360 : NAND3_X1 port map( A1 => n6899, A2 => n3839, A3 => n4873, ZN => 
                           n17772);
   U7361 : INV_X1 port map( A => n11022, ZN => n11314);
   U7362 : OR2_X1 port map( A1 => n18229, A2 => n29023, ZN => n1943);
   U7363 : XNOR2_X1 port map( A => n13094, B => n13093, ZN => n14132);
   U7364 : XNOR2_X1 port map( A => n12425, B => n12424, ZN => n14401);
   U7365 : OR3_X1 port map( A1 => n26195, A2 => n29617, A3 => n26469, ZN => 
                           n1944);
   U7366 : OR2_X1 port map( A1 => n333, A2 => n6815, ZN => n1945);
   U7367 : OR2_X1 port map( A1 => n20306, A2 => n19947, ZN => n1946);
   U7368 : OR2_X1 port map( A1 => n11361, A2 => n15576, ZN => n1947);
   U7369 : OR2_X1 port map( A1 => n21626, A2 => n22139, ZN => n1948);
   U7370 : OR2_X1 port map( A1 => n19939, A2 => n28657, ZN => n1949);
   U7371 : AND2_X1 port map( A1 => n28536, A2 => n28480, ZN => n1950);
   U7373 : OR2_X1 port map( A1 => n498, A2 => n20636, ZN => n1951);
   U7374 : AND2_X1 port map( A1 => n2735, A2 => n20088, ZN => n1952);
   U7375 : OR2_X1 port map( A1 => n17502, A2 => n17140, ZN => n1953);
   U7376 : OR2_X1 port map( A1 => n17764, A2 => n28073, ZN => n1954);
   U7377 : INV_X1 port map( A => n1928, ZN => n4359);
   U7378 : INV_X1 port map( A => n24141, ZN => n24277);
   U7379 : INV_X1 port map( A => n12264, ZN => n12134);
   U7380 : NAND2_X1 port map( A1 => n9865, A2 => n12194, ZN => n11816);
   U7381 : INV_X1 port map( A => n6114, ZN => n20174);
   U7382 : INV_X1 port map( A => n7362, ZN => n3431);
   U7383 : INV_X1 port map( A => n12231, ZN => n13087);
   U7384 : XOR2_X1 port map( A => n13040, B => n13510, Z => n1956);
   U7385 : INV_X1 port map( A => n27701, ZN => n6008);
   U7386 : INV_X1 port map( A => n17829, ZN => n4273);
   U7387 : XOR2_X1 port map( A => n15396, B => n16468, Z => n1957);
   U7388 : XOR2_X1 port map( A => n25249, B => n3607, Z => n1958);
   U7392 : OAI211_X1 port map( C1 => n11952, C2 => n11951, A => n11950, B => 
                           n11949, ZN => n13008);
   U7393 : INV_X1 port map( A => n20443, ZN => n3247);
   U7394 : INV_X1 port map( A => n23305, ZN => n4020);
   U7395 : INV_X1 port map( A => n4037, ZN => n12207);
   U7396 : INV_X1 port map( A => n23764, ZN => n4759);
   U7397 : XNOR2_X1 port map( A => n26078, B => n26079, ZN => n27136);
   U7399 : AND2_X1 port map( A1 => n14193, A2 => n14192, ZN => n1959);
   U7401 : INV_X1 port map( A => n10453, ZN => n11875);
   U7402 : INV_X1 port map( A => n18233, ZN => n18399);
   U7403 : INV_X1 port map( A => n21481, ZN => n21580);
   U7404 : INV_X1 port map( A => n17359, ZN => n2449);
   U7406 : OR2_X1 port map( A1 => n14366, A2 => n14123, ZN => n1960);
   U7407 : OR2_X1 port map( A1 => n13907, A2 => n14051, ZN => n1961);
   U7408 : INV_X1 port map( A => n23529, ZN => n23697);
   U7410 : INV_X1 port map( A => n18179, ZN => n4929);
   U7411 : OR2_X1 port map( A1 => n21369, A2 => n21716, ZN => n1962);
   U7412 : AND2_X1 port map( A1 => n5919, A2 => n5921, ZN => n1963);
   U7413 : OR2_X1 port map( A1 => n15395, A2 => n15394, ZN => n1964);
   U7414 : OR2_X1 port map( A1 => n28506, A2 => n5193, ZN => n1965);
   U7415 : INV_X1 port map( A => n2846, ZN => n12224);
   U7416 : AND2_X1 port map( A1 => n6704, A2 => n6703, ZN => n1966);
   U7417 : INV_X1 port map( A => n9312, ZN => n5412);
   U7418 : INV_X1 port map( A => n24751, ZN => n2879);
   U7419 : NOR2_X1 port map( A1 => n26260, A2 => n6087, ZN => n1968);
   U7420 : INV_X1 port map( A => n22143, ZN => n6532);
   U7421 : AOI21_X1 port map( B1 => n27021, B2 => n27020, A => n27019, ZN => 
                           n27938);
   U7422 : INV_X1 port map( A => n18595, ZN => n5476);
   U7425 : INV_X1 port map( A => n15415, ZN => n3922);
   U7426 : AND2_X1 port map( A1 => n14101, A2 => n14231, ZN => n1969);
   U7427 : AND3_X1 port map( A1 => n20294, A2 => n19814, A3 => n19818, ZN => 
                           n1970);
   U7428 : NAND2_X1 port map( A1 => n27010, A2 => n27013, ZN => n1971);
   U7429 : OR2_X1 port map( A1 => n19829, A2 => n20588, ZN => n1972);
   U7430 : INV_X1 port map( A => n21346, ZN => n3260);
   U7431 : XNOR2_X1 port map( A => n25941, B => n5186, ZN => n26299);
   U7432 : INV_X1 port map( A => n17552, ZN => n4624);
   U7434 : INV_X1 port map( A => n18171, ZN => n4884);
   U7435 : AND2_X1 port map( A1 => n20270, A2 => n3666, ZN => n1974);
   U7436 : INV_X1 port map( A => n22013, ZN => n4828);
   U7437 : INV_X1 port map( A => n18527, ZN => n18535);
   U7438 : XNOR2_X1 port map( A => n9405, B => n9404, ZN => n11003);
   U7439 : INV_X1 port map( A => n23768, ZN => n6462);
   U7440 : INV_X1 port map( A => n10786, ZN => n4538);
   U7441 : INV_X1 port map( A => n23827, ZN => n2187);
   U7442 : AOI22_X1 port map( A1 => n22745, A2 => n23285, B1 => n22638, B2 => 
                           n28594, ZN => n23922);
   U7443 : INV_X1 port map( A => n23922, ZN => n5168);
   U7446 : OR3_X1 port map( A1 => n24502, A2 => n24800, A3 => n24804, ZN => 
                           n1976);
   U7447 : XNOR2_X1 port map( A => n6890, B => n16537, ZN => n17065);
   U7448 : XNOR2_X1 port map( A => n7229, B => n7230, ZN => n10544);
   U7449 : XNOR2_X1 port map( A => n19600, B => n19601, ZN => n20322);
   U7450 : INV_X1 port map( A => n20322, ZN => n2180);
   U7451 : XNOR2_X1 port map( A => n19142, B => n19143, ZN => n20339);
   U7452 : INV_X1 port map( A => n20451, ZN => n5377);
   U7453 : XNOR2_X1 port map( A => n21799, B => n21798, ZN => n23763);
   U7454 : XNOR2_X1 port map( A => n15587, B => n15586, ZN => n17335);
   U7455 : XNOR2_X1 port map( A => n25395, B => n25394, ZN => n26911);
   U7457 : XNOR2_X1 port map( A => Plaintext(84), B => Key(84), ZN => n7839);
   U7459 : XNOR2_X1 port map( A => n21992, B => n21993, ZN => n23736);
   U7460 : XOR2_X1 port map( A => n16605, B => n16604, Z => n1977);
   U7461 : AND3_X1 port map( A1 => n26927, A2 => n26489, A3 => n26933, ZN => 
                           n1978);
   U7462 : INV_X1 port map( A => n18203, ZN => n3995);
   U7463 : XNOR2_X1 port map( A => n24488, B => n25529, ZN => n26459);
   U7464 : INV_X1 port map( A => n18033, ZN => n18155);
   U7465 : XOR2_X1 port map( A => n16339, B => n16405, Z => n1979);
   U7466 : INV_X1 port map( A => n27410, ZN => n4922);
   U7467 : XNOR2_X1 port map( A => n25258, B => n25259, ZN => n26761);
   U7469 : NAND2_X1 port map( A1 => n25159, A2 => n25158, ZN => n27202);
   U7471 : XNOR2_X1 port map( A => n18822, B => n18823, ZN => n20099);
   U7473 : XOR2_X1 port map( A => n15801, B => n2995, Z => n1980);
   U7474 : XOR2_X1 port map( A => n18778, B => n19225, Z => n1981);
   U7475 : XNOR2_X1 port map( A => n18555, B => n18554, ZN => n19843);
   U7476 : XNOR2_X1 port map( A => n22559, B => n22560, ZN => n23738);
   U7477 : XOR2_X1 port map( A => n19110, B => n1927, Z => n1982);
   U7478 : XOR2_X1 port map( A => n10363, B => n3244, Z => n1983);
   U7479 : XNOR2_X1 port map( A => n20839, B => n20838, ZN => n23658);
   U7480 : XOR2_X1 port map( A => n22633, B => n28294, Z => n1984);
   U7481 : XOR2_X1 port map( A => n9575, B => n9512, Z => n1985);
   U7482 : XNOR2_X1 port map( A => n8455, B => n8454, ZN => n10748);
   U7483 : XOR2_X1 port map( A => n13445, B => n13446, Z => n1987);
   U7484 : XOR2_X1 port map( A => n9466, B => n9465, Z => n1988);
   U7485 : XOR2_X1 port map( A => n19704, B => n2995, Z => n1989);
   U7486 : XNOR2_X1 port map( A => n22804, B => n22803, ZN => n23418);
   U7487 : XNOR2_X1 port map( A => n22335, B => n22336, ZN => n23760);
   U7488 : INV_X1 port map( A => n18251, ZN => n2834);
   U7489 : INV_X1 port map( A => n6504, ZN => n22427);
   U7490 : XOR2_X1 port map( A => n8844, B => n8843, Z => n1990);
   U7493 : AND2_X1 port map( A1 => n8014, A2 => n7141, ZN => n1991);
   U7494 : INV_X1 port map( A => n21145, ZN => n21120);
   U7495 : OR2_X1 port map( A1 => n18451, A2 => n18198, ZN => n1992);
   U7496 : OR3_X1 port map( A1 => n11979, A2 => n1986, A3 => n375, ZN => n1993)
                           ;
   U7497 : INV_X1 port map( A => n22991, ZN => n22996);
   U7498 : AND2_X1 port map( A1 => n27191, A2 => n28513, ZN => n1994);
   U7499 : OR3_X1 port map( A1 => n27175, A2 => n27177, A3 => n27178, ZN => 
                           n1995);
   U7500 : OR3_X1 port map( A1 => n26920, A2 => n26782, A3 => n26919, ZN => 
                           n1996);
   U7501 : INV_X1 port map( A => n21095, ZN => n20147);
   U7502 : INV_X1 port map( A => n20137, ZN => n2152);
   U7503 : XOR2_X1 port map( A => n16052, B => n16476, Z => n1998);
   U7504 : AND2_X1 port map( A1 => n11235, A2 => n3441, ZN => n1999);
   U7505 : OR2_X1 port map( A1 => n13716, A2 => n13902, ZN => n2000);
   U7506 : XNOR2_X1 port map( A => n15579, B => n15580, ZN => n17204);
   U7507 : NAND2_X1 port map( A1 => n4640, A2 => n20169, ZN => n21089);
   U7508 : XNOR2_X1 port map( A => n16209, B => n16210, ZN => n16887);
   U7510 : AND2_X1 port map( A1 => n15382, A2 => n15383, ZN => n2001);
   U7511 : INV_X1 port map( A => n19995, ZN => n19997);
   U7512 : INV_X1 port map( A => n18500, ZN => n18217);
   U7513 : AND2_X1 port map( A1 => n15420, A2 => n15102, ZN => n2002);
   U7514 : XOR2_X1 port map( A => n13552, B => n27225, Z => n2003);
   U7515 : AND2_X1 port map( A1 => n23801, A2 => n23802, ZN => n2004);
   U7516 : INV_X1 port map( A => n20858, ZN => n4960);
   U7517 : INV_X1 port map( A => n2108, ZN => n4109);
   U7519 : XNOR2_X1 port map( A => Key(0), B => Plaintext(0), ZN => n7889);
   U7522 : AND2_X1 port map( A1 => n9062, A2 => n8872, ZN => n2006);
   U7523 : AND2_X1 port map( A1 => n20064, A2 => n20069, ZN => n2007);
   U7524 : INV_X1 port map( A => n18261, ZN => n3833);
   U7525 : AND2_X1 port map( A1 => n11574, A2 => n12132, ZN => n2008);
   U7526 : OR2_X1 port map( A1 => n14948, A2 => n15073, ZN => n2009);
   U7527 : INV_X1 port map( A => n7830, ZN => n8205);
   U7529 : AND2_X1 port map( A1 => n27851, A2 => n27854, ZN => n2010);
   U7530 : OR2_X1 port map( A1 => n27704, A2 => n27161, ZN => n2011);
   U7531 : OR3_X1 port map( A1 => n12578, A2 => n12272, A3 => n12270, ZN => 
                           n2012);
   U7532 : OR3_X1 port map( A1 => n24794, A2 => n2937, A3 => n24791, ZN => 
                           n2013);
   U7533 : OR3_X1 port map( A1 => n26362, A2 => n26799, A3 => n29573, ZN => 
                           n2014);
   U7534 : AND2_X1 port map( A1 => n25239, A2 => n27395, ZN => n2015);
   U7535 : AND2_X1 port map( A1 => n23663, A2 => n23662, ZN => n2016);
   U7536 : INV_X1 port map( A => n22141, ZN => n21627);
   U7537 : AND2_X1 port map( A1 => n14302, A2 => n29611, ZN => n2017);
   U7538 : OR2_X1 port map( A1 => n14373, A2 => n3860, ZN => n2018);
   U7539 : OR2_X1 port map( A1 => n17686, A2 => n28779, ZN => n2019);
   U7540 : AND2_X1 port map( A1 => n14131, A2 => n13842, ZN => n2020);
   U7541 : INV_X1 port map( A => n16977, ZN => n16774);
   U7542 : INV_X1 port map( A => n13602, ZN => n15404);
   U7543 : AND2_X1 port map( A1 => n28090, A2 => n4359, ZN => n2021);
   U7544 : OR2_X1 port map( A1 => n21634, A2 => n21638, ZN => n2022);
   U7545 : OR2_X1 port map( A1 => n20283, A2 => n28657, ZN => n2023);
   U7547 : AND2_X1 port map( A1 => n8593, A2 => n8817, ZN => n2024);
   U7548 : XOR2_X1 port map( A => n12883, B => n623, Z => n2025);
   U7549 : AND2_X1 port map( A1 => n21603, A2 => n28442, ZN => n2026);
   U7550 : INV_X1 port map( A => n6741, ZN => n24578);
   U7551 : AND2_X1 port map( A1 => n12266, A2 => n12267, ZN => n2027);
   U7552 : AND2_X1 port map( A1 => n15054, A2 => n14763, ZN => n2028);
   U7553 : AND2_X1 port map( A1 => n8955, A2 => n8956, ZN => n2029);
   U7554 : AND2_X1 port map( A1 => n17004, A2 => n17003, ZN => n2030);
   U7555 : OR2_X1 port map( A1 => n18588, A2 => n17206, ZN => n2031);
   U7556 : AND2_X1 port map( A1 => n4900, A2 => n4901, ZN => n2032);
   U7557 : XOR2_X1 port map( A => n10250, B => n3003, Z => n2034);
   U7558 : XOR2_X1 port map( A => n10137, B => n2912, Z => n2035);
   U7559 : INV_X1 port map( A => n24403, ZN => n2762);
   U7560 : INV_X1 port map( A => n23648, ZN => n23654);
   U7561 : OR2_X1 port map( A1 => n23612, A2 => n28582, ZN => n2036);
   U7562 : AND2_X1 port map( A1 => n5435, A2 => n5437, ZN => n2037);
   U7563 : INV_X1 port map( A => n27827, ZN => n27825);
   U7565 : OR2_X1 port map( A1 => n27134, A2 => n27129, ZN => n2038);
   U7566 : INV_X1 port map( A => n5383, ZN => n18380);
   U7567 : INV_X1 port map( A => n24709, ZN => n5752);
   U7568 : AND2_X1 port map( A1 => n5399, A2 => n4795, ZN => n2039);
   U7570 : AND2_X1 port map( A1 => n15382, A2 => n15151, ZN => n2040);
   U7571 : OR2_X1 port map( A1 => n22142, A2 => n19760, ZN => n2041);
   U7572 : AND2_X1 port map( A1 => n24515, A2 => n24514, ZN => n3671);
   U7573 : AND2_X1 port map( A1 => n8077, A2 => n8428, ZN => n2042);
   U7574 : OR2_X1 port map( A1 => n26455, A2 => n26454, ZN => n2043);
   U7575 : OR2_X1 port map( A1 => n18129, A2 => n17839, ZN => n2044);
   U7576 : NOR2_X1 port map( A1 => n13684, A2 => n3580, ZN => n14989);
   U7577 : INV_X1 port map( A => n14989, ZN => n3210);
   U7580 : OR2_X1 port map( A1 => n23469, A2 => n3135, ZN => n2046);
   U7581 : INV_X1 port map( A => n12201, ZN => n5825);
   U7582 : OR2_X1 port map( A1 => n5777, A2 => n15235, ZN => n2047);
   U7583 : NAND2_X1 port map( A1 => n17527, A2 => n6161, ZN => n2048);
   U7584 : INV_X1 port map( A => n10558, ZN => n11345);
   U7585 : INV_X1 port map( A => n27843, ZN => n27828);
   U7586 : AND2_X1 port map( A1 => n2259, A2 => n2258, ZN => n2049);
   U7587 : NAND2_X1 port map( A1 => n26929, A2 => n26489, ZN => n2050);
   U7588 : OR2_X1 port map( A1 => n26234, A2 => n26235, ZN => n2051);
   U7589 : XNOR2_X1 port map( A => n9489, B => n9490, ZN => n11253);
   U7590 : OR2_X1 port map( A1 => n17156, A2 => n17336, ZN => n2052);
   U7591 : NAND3_X1 port map( A1 => n29161, A2 => n29032, A3 => n29031, ZN => 
                           n2053);
   U7592 : OR2_X1 port map( A1 => n23724, A2 => n22455, ZN => n2054);
   U7594 : AND2_X1 port map( A1 => n3811, A2 => n5620, ZN => n2055);
   U7595 : AND2_X1 port map( A1 => n29572, A2 => n17395, ZN => n2056);
   U7596 : INV_X1 port map( A => n15828, ZN => n15007);
   U7597 : OR2_X1 port map( A1 => n17386, A2 => n17385, ZN => n2057);
   U7598 : NAND2_X1 port map( A1 => n23141, A2 => n5773, ZN => n2058);
   U7599 : OR2_X1 port map( A1 => n7651, A2 => n29081, ZN => n2059);
   U7600 : INV_X1 port map( A => n21586, ZN => n3789);
   U7601 : INV_X1 port map( A => n11550, ZN => n3900);
   U7602 : AND2_X1 port map( A1 => n27938, A2 => n28439, ZN => n2060);
   U7603 : OR2_X1 port map( A1 => n17313, A2 => n17315, ZN => n2061);
   U7606 : AND2_X1 port map( A1 => n20476, A2 => n20475, ZN => n2062);
   U7607 : INV_X1 port map( A => n11194, ZN => n5838);
   U7608 : INV_X1 port map( A => n21575, ZN => n21577);
   U7609 : OAI211_X1 port map( C1 => n20070, C2 => n20379, A => n20071, B => 
                           n19842, ZN => n21575);
   U7610 : INV_X1 port map( A => n24155, ZN => n24523);
   U7611 : NAND2_X1 port map( A1 => n28206, A2 => n11144, ZN => n2063);
   U7612 : NAND2_X1 port map( A1 => n25750, A2 => n27076, ZN => n2064);
   U7613 : OR2_X1 port map( A1 => n24609, A2 => n29109, ZN => n2065);
   U7614 : OR2_X1 port map( A1 => n23637, A2 => n29061, ZN => n2066);
   U7615 : AND2_X1 port map( A1 => n20783, A2 => n21177, ZN => n2067);
   U7616 : OR2_X1 port map( A1 => n3830, A2 => n13910, ZN => n2068);
   U7617 : OR2_X1 port map( A1 => n17342, A2 => n16711, ZN => n2069);
   U7618 : AND2_X1 port map( A1 => n23839, A2 => n23392, ZN => n2070);
   U7619 : OR2_X1 port map( A1 => n7534, A2 => n7749, ZN => n2071);
   U7621 : INV_X1 port map( A => n11430, ZN => n2748);
   U7622 : OR2_X1 port map( A1 => n4097, A2 => n15261, ZN => n2073);
   U7623 : OR2_X1 port map( A1 => n11927, A2 => n11852, ZN => n2074);
   U7624 : OR2_X1 port map( A1 => n14142, A2 => n13900, ZN => n2075);
   U7625 : INV_X1 port map( A => n28035, ZN => n6859);
   U7626 : INV_X1 port map( A => n20580, ZN => n20416);
   U7627 : AND2_X1 port map( A1 => n28506, A2 => n5192, ZN => n2076);
   U7628 : OAI21_X1 port map( B1 => n3986, B2 => n23434, A => n3985, ZN => 
                           n24509);
   U7629 : INV_X1 port map( A => n12257, ZN => n6687);
   U7630 : INV_X1 port map( A => n24794, ZN => n4576);
   U7632 : INV_X1 port map( A => n10497, ZN => n2646);
   U7633 : INV_X1 port map( A => n17977, ZN => n18234);
   U7634 : BUF_X1 port map( A => n10622, Z => n11896);
   U7636 : INV_X1 port map( A => n21656, ZN => n21440);
   U7638 : NAND3_X1 port map( A1 => n27076, A2 => n28521, A3 => n29622, ZN => 
                           n2078);
   U7639 : INV_X1 port map( A => n18383, ZN => n3283);
   U7640 : INV_X1 port map( A => n8929, ZN => n5958);
   U7641 : OR2_X1 port map( A1 => n23576, A2 => n23956, ZN => n2079);
   U7642 : OR2_X1 port map( A1 => n7633, A2 => n7915, ZN => n2080);
   U7643 : AND2_X1 port map( A1 => n4581, A2 => n20282, ZN => n2081);
   U7644 : OR2_X1 port map( A1 => n20321, A2 => n2180, ZN => n2082);
   U7646 : INV_X1 port map( A => n17088, ZN => n17504);
   U7647 : INV_X1 port map( A => n3501, ZN => n5513);
   U7648 : INV_X1 port map( A => n900, ZN => n4501);
   U7649 : INV_X1 port map( A => n3666, ZN => n6016);
   U7650 : INV_X1 port map( A => n1172, ZN => n4607);
   U7651 : INV_X1 port map( A => n72, ZN => n4070);
   U7652 : INV_X1 port map( A => n1923, ZN => n4222);
   U7653 : INV_X1 port map( A => n3036, ZN => n2116);
   U7654 : INV_X1 port map( A => n3062, ZN => n6653);
   U7655 : INV_X1 port map( A => n26032, ZN => n2117);
   U7656 : INV_X1 port map( A => n1215, ZN => n5892);
   U7657 : INV_X1 port map( A => n3003, ZN => n6174);
   U7658 : INV_X1 port map( A => n3710, ZN => n5802);
   U7659 : INV_X1 port map( A => n15576, ZN => n6319);
   U7660 : NAND2_X1 port map( A1 => n2083, A2 => n21032, ZN => n21389);
   U7661 : NAND3_X1 port map( A1 => n2091, A2 => n19965, A3 => n2083, ZN => 
                           n21731);
   U7662 : OAI21_X1 port map( B1 => n19963, B2 => n20548, A => n20556, ZN => 
                           n2083);
   U7663 : NAND2_X1 port map( A1 => n10640, A2 => n11242, ZN => n2085);
   U7664 : NAND2_X1 port map( A1 => n10639, A2 => n1900, ZN => n2086);
   U7665 : NAND2_X1 port map( A1 => n10629, A2 => n11235, ZN => n2087);
   U7666 : OAI22_X1 port map( A1 => n2090, A2 => n7619, B1 => n2088, B2 => 
                           n5946, ZN => n6060);
   U7667 : NAND2_X1 port map( A1 => n8236, A2 => n2089, ZN => n2088);
   U7668 : INV_X1 port map( A => n6973, ZN => n2089);
   U7669 : NAND2_X1 port map( A1 => n7919, A2 => n5946, ZN => n2090);
   U7670 : INV_X1 port map( A => n8231, ZN => n5946);
   U7671 : INV_X1 port map( A => n6973, ZN => n8234);
   U7672 : XNOR2_X2 port map( A => n6970, B => Key(107), ZN => n6973);
   U7673 : OAI21_X1 port map( B1 => n28114, B2 => n29480, A => n2092, ZN => 
                           n2093);
   U7674 : OAI21_X1 port map( B1 => n28109, B2 => n28110, A => n28075, ZN => 
                           n2092);
   U7675 : XNOR2_X1 port map( A => n2093, B => n28116, ZN => Ciphertext(191));
   U7676 : NAND2_X1 port map( A1 => n26996, A2 => n28532, ZN => n2094);
   U7677 : NAND2_X1 port map( A1 => n2096, A2 => n20222, ZN => n6577);
   U7680 : XNOR2_X1 port map( A => n2098, B => n22697, ZN => n22151);
   U7681 : NAND2_X1 port map( A1 => n22147, A2 => n2097, ZN => n2098);
   U7682 : XNOR2_X1 port map( A => n2098, B => n22525, ZN => n22470);
   U7685 : NAND2_X1 port map( A1 => n6260, A2 => n6259, ZN => n2101);
   U7687 : NOR2_X1 port map( A1 => n20829, A2 => n2101, ZN => n20831);
   U7688 : OR2_X1 port map( A1 => n2103, A2 => n10821, ZN => n4945);
   U7689 : NOR2_X1 port map( A1 => n4463, A2 => n2102, ZN => n4462);
   U7690 : AND2_X1 port map( A1 => n2103, A2 => n11331, ZN => n2102);
   U7691 : NAND2_X1 port map( A1 => n2104, A2 => n8941, ZN => n3595);
   U7692 : INV_X1 port map( A => n8553, ZN => n2104);
   U7693 : NAND2_X1 port map( A1 => n24641, A2 => n2107, ZN => n2105);
   U7694 : NAND2_X1 port map( A1 => n23176, A2 => n24195, ZN => n2106);
   U7696 : NAND2_X1 port map( A1 => n27193, A2 => n29585, ZN => n26140);
   U7697 : OAI211_X1 port map( C1 => n4243, C2 => n29585, A => n27123, B => 
                           n28595, ZN => n26292);
   U7698 : NAND2_X1 port map( A1 => n1994, A2 => n29585, ZN => n4110);
   U7699 : MUX2_X1 port map( A => n27193, B => n26291, S => n4109, Z => n26294)
                           ;
   U7700 : XNOR2_X2 port map( A => n12434, B => n4510, ZN => n13877);
   U7701 : NAND3_X1 port map( A1 => n28804, A2 => n13877, A3 => n14402, ZN => 
                           n2110);
   U7703 : NAND2_X1 port map( A1 => n14403, A2 => n4509, ZN => n2111);
   U7704 : XNOR2_X1 port map( A => n29140, B => n12450, ZN => n2113);
   U7705 : NAND2_X1 port map( A1 => n2114, A2 => n17497, ZN => n5587);
   U7706 : NOR2_X1 port map( A1 => n17496, A2 => n2114, ZN => n18223);
   U7707 : NAND2_X1 port map( A1 => n538, A2 => n17062, ZN => n2114);
   U7708 : NAND2_X1 port map( A1 => n4052, A2 => n2115, ZN => n4051);
   U7710 : NAND2_X1 port map( A1 => n2119, A2 => n23446, ZN => n2118);
   U7712 : NAND2_X1 port map( A1 => n2118, A2 => n2120, ZN => n22740);
   U7713 : NAND2_X1 port map( A1 => n2119, A2 => n23449, ZN => n4916);
   U7714 : NAND2_X1 port map( A1 => n23109, A2 => n23442, ZN => n2120);
   U7715 : NAND2_X1 port map( A1 => n2121, A2 => n5397, ZN => n4795);
   U7716 : NOR2_X1 port map( A1 => n16946, A2 => n2122, ZN => n2121);
   U7717 : INV_X1 port map( A => n17242, ZN => n2122);
   U7718 : NAND2_X1 port map( A1 => n18149, A2 => n2855, ZN => n17814);
   U7719 : NOR2_X1 port map( A1 => n18148, A2 => n2123, ZN => n18151);
   U7720 : NOR2_X1 port map( A1 => n3467, A2 => n2855, ZN => n18049);
   U7721 : NAND3_X1 port map( A1 => n420, A2 => n2123, A3 => n3467, ZN => 
                           n18434);
   U7723 : XNOR2_X1 port map( A => n18763, B => n18764, ZN => n2124);
   U7724 : XNOR2_X2 port map( A => n2124, B => n3912, ZN => n20049);
   U7725 : AND2_X1 port map( A1 => n20066, A2 => n413, ZN => n6477);
   U7726 : NAND2_X1 port map( A1 => n2125, A2 => n21811, ZN => n21382);
   U7727 : NOR2_X1 port map( A1 => n19732, A2 => n2125, ZN => n20983);
   U7728 : NOR2_X1 port map( A1 => n21809, A2 => n2125, ZN => n20980);
   U7729 : NAND3_X1 port map( A1 => n21809, A2 => n21806, A3 => n2125, ZN => 
                           n21255);
   U7730 : NAND3_X1 port map( A1 => n21809, A2 => n19732, A3 => n2125, ZN => 
                           n19734);
   U7731 : NAND2_X1 port map( A1 => n2127, A2 => n28208, ZN => n10745);
   U7733 : NAND2_X1 port map( A1 => n10467, A2 => n2127, ZN => n8423);
   U7734 : NOR2_X1 port map( A1 => n29310, A2 => n2128, ZN => n10233);
   U7735 : INV_X1 port map( A => n8605, ZN => n2128);
   U7736 : NAND2_X1 port map( A1 => n2129, A2 => n9087, ZN => n9088);
   U7737 : INV_X1 port map( A => n9081, ZN => n2129);
   U7738 : INV_X1 port map( A => n2131, ZN => n2130);
   U7739 : NAND2_X1 port map( A1 => n24676, A2 => n29555, ZN => n2132);
   U7740 : MUX2_X1 port map( A => n29483, B => n17548, S => n4218, Z => n17054)
                           ;
   U7741 : NAND2_X1 port map( A1 => n4787, A2 => n2133, ZN => n16763);
   U7742 : OAI22_X1 port map( A1 => n2134, A2 => n24426, B1 => n28531, B2 => 
                           n24772, ZN => n24430);
   U7743 : NAND2_X1 port map( A1 => n5248, A2 => n24769, ZN => n2134);
   U7746 : NAND2_X1 port map( A1 => n2137, A2 => n13718, ZN => n13723);
   U7749 : NAND2_X1 port map( A1 => n27134, A2 => n29293, ZN => n2140);
   U7750 : NAND2_X1 port map( A1 => n23256, A2 => n2141, ZN => n23732);
   U7751 : NOR2_X1 port map( A1 => n23398, A2 => n2141, ZN => n22950);
   U7752 : MUX2_X1 port map( A => n3432, B => n22949, S => n23397, Z => n23232)
                           ;
   U7753 : NAND2_X1 port map( A1 => n11377, A2 => n12102, ZN => n11655);
   U7754 : XNOR2_X2 port map( A => Key(11), B => Plaintext(11), ZN => n7770);
   U7755 : INV_X1 port map( A => n12104, ZN => n11662);
   U7757 : NAND2_X1 port map( A1 => n11659, A2 => n29116, ZN => n2142);
   U7758 : AOI21_X1 port map( B1 => n2144, B2 => n14037, A => n14036, ZN => 
                           n14042);
   U7759 : NAND2_X1 port map( A1 => n28513, A2 => n27190, ZN => n24920);
   U7760 : MUX2_X1 port map( A => n27190, B => n28513, S => n27191, Z => n27192
                           );
   U7761 : MUX2_X1 port map( A => n28595, B => n4227, S => n27123, Z => n27126)
                           ;
   U7762 : NAND2_X1 port map( A1 => n6177, A2 => n2146, ZN => n16957);
   U7763 : NAND2_X1 port map( A1 => n18537, A2 => n18527, ZN => n2146);
   U7764 : NAND2_X1 port map( A1 => n2148, A2 => n18536, ZN => n2147);
   U7765 : NAND2_X1 port map( A1 => n18537, A2 => n2149, ZN => n2148);
   U7766 : NAND2_X1 port map( A1 => n18538, A2 => n18527, ZN => n2149);
   U7767 : NAND2_X1 port map( A1 => n16957, A2 => n2151, ZN => n2150);
   U7768 : XNOR2_X1 port map( A => n2154, B => n2509, ZN => n24671);
   U7769 : XNOR2_X1 port map( A => n25773, B => n2154, ZN => n25099);
   U7770 : XNOR2_X1 port map( A => n25391, B => n2154, ZN => n25735);
   U7773 : NAND3_X1 port map( A1 => n17496, A2 => n4314, A3 => n17062, ZN => 
                           n2157);
   U7774 : NAND2_X1 port map( A1 => n2159, A2 => n17492, ZN => n2158);
   U7775 : XNOR2_X2 port map( A => n16308, B => n16307, ZN => n17492);
   U7776 : NAND2_X1 port map( A1 => n17497, A2 => n17491, ZN => n2159);
   U7777 : NAND2_X1 port map( A1 => n2161, A2 => n6207, ZN => n2160);
   U7778 : INV_X1 port map( A => n14761, ZN => n15261);
   U7780 : NAND2_X1 port map( A1 => n2164, A2 => n10991, ZN => n11694);
   U7781 : NAND2_X1 port map( A1 => n10635, A2 => n2165, ZN => n2164);
   U7783 : NAND2_X1 port map( A1 => n12286, A2 => n2166, ZN => n11625);
   U7784 : INV_X1 port map( A => n12281, ZN => n2166);
   U7785 : INV_X1 port map( A => n12407, ZN => n2167);
   U7786 : INV_X1 port map( A => n2168, ZN => n9567);
   U7788 : NAND2_X1 port map( A1 => n23110, A2 => n4794, ZN => n2169);
   U7790 : NAND2_X1 port map( A1 => n6209, A2 => n7506, ZN => n4129);
   U7791 : XNOR2_X2 port map( A => n7022, B => Key(56), ZN => n7257);
   U7792 : NAND2_X1 port map( A1 => n2174, A2 => n23468, ZN => n25282);
   U7793 : NAND3_X1 port map( A1 => n2176, A2 => n6786, A3 => n2175, ZN => 
                           n2174);
   U7794 : NAND2_X1 port map( A1 => n6788, A2 => n6787, ZN => n2176);
   U7795 : NAND2_X1 port map( A1 => n20325, A2 => n502, ZN => n2177);
   U7797 : NAND3_X1 port map( A1 => n20324, A2 => n2181, A3 => n2180, ZN => 
                           n2179);
   U7798 : NAND2_X1 port map( A1 => n2884, A2 => n20320, ZN => n2182);
   U7799 : OAI21_X1 port map( B1 => n2183, B2 => n17088, A => n1953, ZN => 
                           n17207);
   U7800 : NAND2_X1 port map( A1 => n2186, A2 => n2184, ZN => n2183);
   U7801 : NAND2_X1 port map( A1 => n17501, A2 => n2185, ZN => n2184);
   U7802 : NAND2_X1 port map( A1 => n29127, A2 => n16888, ZN => n17501);
   U7803 : INV_X1 port map( A => n17087, ZN => n2186);
   U7804 : NAND2_X1 port map( A1 => n23385, A2 => n23825, ZN => n2189);
   U7805 : NAND3_X1 port map( A1 => n23385, A2 => n23825, A3 => n2187, ZN => 
                           n2188);
   U7806 : AND2_X1 port map( A1 => n2189, A2 => n3940, ZN => n23743);
   U7807 : AND2_X1 port map( A1 => n4483, A2 => n2189, ZN => n24090);
   U7808 : NAND2_X1 port map( A1 => n20841, A2 => n21459, ZN => n21571);
   U7810 : NAND2_X1 port map( A1 => n2192, A2 => n2191, ZN => n2190);
   U7811 : NAND2_X1 port map( A1 => n14799, A2 => n547, ZN => n2192);
   U7812 : NAND2_X1 port map( A1 => n15185, A2 => n14784, ZN => n14799);
   U7813 : NAND2_X1 port map( A1 => n11487, A2 => n28436, ZN => n2360);
   U7814 : OAI211_X1 port map( C1 => n11430, C2 => n11487, A => n10717, B => 
                           n2193, ZN => n2303);
   U7816 : INV_X1 port map( A => n11787, ZN => n2194);
   U7818 : NAND2_X1 port map( A1 => n2200, A2 => n2199, ZN => n4954);
   U7819 : NAND2_X1 port map( A1 => n523, A2 => n18441, ZN => n2199);
   U7820 : NAND2_X1 port map( A1 => n18444, A2 => n18178, ZN => n2200);
   U7821 : NAND2_X1 port map( A1 => n18090, A2 => n18093, ZN => n18180);
   U7822 : NAND2_X1 port map( A1 => n16755, A2 => n16756, ZN => n18178);
   U7823 : AND2_X1 port map( A1 => n22745, A2 => n2202, ZN => n2201);
   U7824 : NAND2_X1 port map( A1 => n2203, A2 => n15379, ZN => n15380);
   U7825 : NAND2_X1 port map( A1 => n2040, A2 => n15155, ZN => n5815);
   U7826 : OAI21_X1 port map( B1 => n15384, B2 => n2203, A => n2001, ZN => 
                           n15385);
   U7827 : INV_X1 port map( A => n24240, ZN => n2205);
   U7829 : INV_X1 port map( A => n15565, ZN => n15452);
   U7830 : XNOR2_X1 port map( A => n15565, B => n2206, ZN => n15852);
   U7831 : INV_X1 port map( A => n15940, ZN => n2206);
   U7832 : OAI211_X1 port map( C1 => n28555, C2 => n20614, A => n20611, B => 
                           n19935, ZN => n4587);
   U7833 : OR2_X1 port map( A1 => n29646, A2 => n8131, ZN => n8050);
   U7834 : INV_X1 port map( A => n7129, ZN => n8049);
   U7835 : OR2_X1 port map( A1 => n6000, A2 => n14091, ZN => n4721);
   U7836 : INV_X1 port map( A => n24520, ZN => n3618);
   U7838 : XNOR2_X1 port map( A => n25948, B => n1172, ZN => n24529);
   U7839 : NOR2_X1 port map( A1 => n17487, A2 => n17489, ZN => n17151);
   U7840 : OR2_X1 port map( A1 => n4884, A2 => n28649, ZN => n3349);
   U7841 : OR2_X1 port map( A1 => n10995, A2 => n10786, ZN => n10597);
   U7842 : NOR2_X1 port map( A1 => n4231, A2 => n5773, ZN => n4769);
   U7843 : AND3_X1 port map( A1 => n5774, A2 => n23011, A3 => n4231, ZN => 
                           n4848);
   U7844 : INV_X1 port map( A => n19025, ZN => n4883);
   U7845 : OAI21_X1 port map( B1 => n8670, B2 => n9107, A => n8914, ZN => n8920
                           );
   U7846 : INV_X1 port map( A => n8670, ZN => n8511);
   U7847 : XNOR2_X1 port map( A => n22526, B => n21980, ZN => n22880);
   U7848 : AND2_X1 port map( A1 => n7488, A2 => n341, ZN => n3298);
   U7849 : XNOR2_X1 port map( A => n19685, B => n3686, ZN => n4043);
   U7850 : XNOR2_X1 port map( A => n19685, B => n27811, ZN => n4746);
   U7851 : XNOR2_X1 port map( A => n15971, B => n3661, ZN => n16140);
   U7853 : MUX2_X1 port map( A => n6608, B => n23792, S => n23790, Z => n23498)
                           ;
   U7854 : NOR2_X1 port map( A1 => n5764, A2 => n2640, ZN => n2639);
   U7855 : OR2_X1 port map( A1 => n4734, A2 => n29153, ZN => n14805);
   U7856 : OR2_X1 port map( A1 => n13257, A2 => n14314, ZN => n6307);
   U7857 : OR2_X1 port map( A1 => n11237, A2 => n11236, ZN => n2413);
   U7858 : OR2_X1 port map( A1 => n7898, A2 => n7900, ZN => n7596);
   U7859 : AND2_X1 port map( A1 => n20319, A2 => n20323, ZN => n2884);
   U7860 : AOI21_X1 port map( B1 => n6376, B2 => n18344, A => n18343, ZN => 
                           n18345);
   U7861 : OR2_X1 port map( A1 => n2717, A2 => n7340, ZN => n2716);
   U7862 : INV_X1 port map( A => n2452, ZN => n23415);
   U7863 : OR2_X1 port map( A1 => n23416, A2 => n2452, ZN => n2435);
   U7864 : OR2_X1 port map( A1 => n15447, A2 => n15323, ZN => n6521);
   U7865 : OR2_X1 port map( A1 => n23535, A2 => n23531, ZN => n4125);
   U7866 : XNOR2_X1 port map( A => n22698, B => n22594, ZN => n3092);
   U7867 : NOR2_X1 port map( A1 => n17719, A2 => n18286, ZN => n18525);
   U7868 : AND3_X1 port map( A1 => n17858, A2 => n17719, A3 => n18081, ZN => 
                           n5325);
   U7869 : AND2_X1 port map( A1 => n17719, A2 => n17859, ZN => n16980);
   U7870 : AND2_X1 port map( A1 => n4046, A2 => n11430, ZN => n11302);
   U7872 : NOR2_X1 port map( A1 => n24484, A2 => n23968, ZN => n24212);
   U7873 : OR2_X1 port map( A1 => n20488, A2 => n20485, ZN => n3532);
   U7874 : INV_X1 port map( A => n28620, ZN => n20240);
   U7875 : OR2_X1 port map( A1 => n28620, A2 => n20483, ZN => n19092);
   U7876 : OR2_X1 port map( A1 => n9530, A2 => n9531, ZN => n3156);
   U7877 : NAND2_X1 port map( A1 => n6892, A2 => n9530, ZN => n7419);
   U7879 : INV_X1 port map( A => n27724, ZN => n27714);
   U7880 : OR2_X1 port map( A1 => n11135, A2 => n3829, ZN => n3828);
   U7881 : XOR2_X1 port map( A => n10177, B => n8863, Z => n8885);
   U7882 : XNOR2_X1 port map( A => n19213, B => n19214, ZN => n20343);
   U7883 : OR2_X1 port map( A1 => n20725, A2 => n21598, ZN => n3530);
   U7884 : INV_X1 port map( A => n27773, ZN => n6419);
   U7885 : OR2_X1 port map( A1 => n29537, A2 => n27762, ZN => n5776);
   U7886 : AND2_X1 port map( A1 => n27904, A2 => n29536, ZN => n27839);
   U7887 : INV_X1 port map( A => n26299, ZN => n27060);
   U7888 : XNOR2_X1 port map( A => n25942, B => n25940, ZN => n5186);
   U7889 : XNOR2_X1 port map( A => n22302, B => n2752, ZN => n22235);
   U7890 : INV_X1 port map( A => n14304, ZN => n5956);
   U7891 : AND2_X1 port map( A1 => n11877, A2 => n10868, ZN => n11879);
   U7892 : AND2_X1 port map( A1 => n20636, A2 => n20639, ZN => n2528);
   U7893 : XNOR2_X1 port map( A => n18900, B => n28571, ZN => n6468);
   U7894 : INV_X1 port map( A => n18900, ZN => n19162);
   U7895 : OAI21_X1 port map( B1 => n4667, B2 => n14278, A => n14363, ZN => 
                           n4666);
   U7897 : OAI21_X1 port map( B1 => n27087, B2 => n26841, A => n2877, ZN => 
                           n27021);
   U7899 : OR2_X1 port map( A1 => n17282, A2 => n17283, ZN => n6380);
   U7900 : INV_X1 port map( A => n13725, ZN => n5404);
   U7901 : MUX2_X1 port map( A => n8351, B => n261, S => n8353, Z => n8356);
   U7902 : OR2_X1 port map( A1 => n23235, A2 => n23716, ZN => n23265);
   U7903 : NAND2_X1 port map( A1 => n23537, A2 => n23541, ZN => n2636);
   U7904 : AND2_X1 port map( A1 => n29508, A2 => n20614, ZN => n4684);
   U7905 : INV_X1 port map( A => n15727, ZN => n16427);
   U7906 : OR2_X1 port map( A1 => n8785, A2 => n8717, ZN => n4320);
   U7907 : OR2_X1 port map( A1 => n8047, A2 => n7127, ZN => n7716);
   U7908 : INV_X1 port map( A => n16846, ZN => n17009);
   U7909 : OR2_X1 port map( A1 => n21322, A2 => n5983, ZN => n21137);
   U7910 : NOR2_X1 port map( A1 => n29569, A2 => n21322, ZN => n20887);
   U7911 : XNOR2_X1 port map( A => n19272, B => n19534, ZN => n19598);
   U7912 : INV_X1 port map( A => n2728, ZN => n5978);
   U7913 : INV_X1 port map( A => n12022, ZN => n12353);
   U7914 : AND2_X1 port map( A1 => n12022, A2 => n11901, ZN => n10587);
   U7915 : INV_X1 port map( A => n7175, ZN => n8730);
   U7917 : INV_X1 port map( A => n14008, ZN => n4586);
   U7918 : NOR2_X1 port map( A1 => n10114, A2 => n11120, ZN => n4383);
   U7919 : OR2_X1 port map( A1 => n13932, A2 => n14452, ZN => n2327);
   U7921 : AND2_X1 port map( A1 => n14451, A2 => n14452, ZN => n3526);
   U7922 : OR2_X1 port map( A1 => n12234, A2 => n375, ZN => n6581);
   U7923 : OR2_X1 port map( A1 => n11176, A2 => n434, ZN => n11340);
   U7924 : AOI21_X1 port map( B1 => n7273, B2 => n2104, A => n9562, ZN => n7274
                           );
   U7925 : OR2_X1 port map( A1 => n10853, A2 => n11163, ZN => n11057);
   U7926 : INV_X1 port map( A => n15009, ZN => n3784);
   U7927 : AND2_X1 port map( A1 => n15371, A2 => n15009, ZN => n3840);
   U7928 : XNOR2_X1 port map( A => n19251, B => n5246, ZN => n19473);
   U7929 : INV_X1 port map( A => n18799, ZN => n5246);
   U7930 : OR2_X1 port map( A1 => n29152, A2 => n6002, ZN => n16964);
   U7931 : XNOR2_X1 port map( A => n12787, B => n13159, ZN => n12421);
   U7932 : AND2_X1 port map( A1 => n29058, A2 => n25676, ZN => n27003);
   U7933 : INV_X1 port map( A => n25676, ZN => n27045);
   U7934 : XNOR2_X1 port map( A => n25545, B => n25544, ZN => n25676);
   U7935 : OR2_X1 port map( A1 => n19761, A2 => n20066, ZN => n3436);
   U7936 : NOR2_X1 port map( A1 => n23233, A2 => n22174, ZN => n6728);
   U7937 : OR2_X1 port map( A1 => n21432, A2 => n21431, ZN => n4312);
   U7938 : OAI21_X1 port map( B1 => n1916, B2 => n20601, A => n20599, ZN => 
                           n5357);
   U7940 : AOI21_X1 port map( B1 => n7362, B2 => n7363, A => n8205, ZN => n3429
                           );
   U7941 : OR2_X1 port map( A1 => n7886, A2 => n7071, ZN => n2882);
   U7942 : NOR2_X1 port map( A1 => n7585, A2 => n7886, ZN => n2226);
   U7943 : OR2_X1 port map( A1 => n6617, A2 => n27363, ZN => n6616);
   U7944 : NOR2_X1 port map( A1 => n27908, A2 => n27913, ZN => n27889);
   U7945 : OR3_X1 port map( A1 => n27010, A2 => n27013, A3 => n27052, ZN => 
                           n5686);
   U7946 : INV_X1 port map( A => n7967, ZN => n4697);
   U7947 : AND3_X1 port map( A1 => n7965, A2 => n29302, A3 => n7967, ZN => 
                           n5255);
   U7948 : OR2_X1 port map( A1 => n7966, A2 => n7967, ZN => n3226);
   U7949 : AOI21_X1 port map( B1 => n27357, B2 => n27356, A => n6287, ZN => 
                           n2426);
   U7950 : OR2_X1 port map( A1 => n20383, A2 => n19836, ZN => n6237);
   U7951 : OR2_X1 port map( A1 => n526, A2 => n18136, ZN => n18143);
   U7952 : OR2_X1 port map( A1 => n14192, A2 => n13953, ZN => n5378);
   U7953 : NAND2_X1 port map( A1 => n10532, A2 => n11294, ZN => n5563);
   U7954 : OR2_X1 port map( A1 => n10891, A2 => n11294, ZN => n10892);
   U7955 : OR2_X1 port map( A1 => n23800, A2 => n4726, ZN => n5193);
   U7956 : OR2_X1 port map( A1 => n4193, A2 => n21459, ZN => n20754);
   U7957 : NAND3_X1 port map( A1 => n2210, A2 => n10951, A3 => n10950, ZN => 
                           n11859);
   U7958 : NAND2_X1 port map( A1 => n2211, A2 => n10972, ZN => n10949);
   U7959 : NAND2_X1 port map( A1 => n10971, A2 => n10970, ZN => n2211);
   U7960 : OAI211_X1 port map( C1 => n18599, C2 => n28142, A => n2213, B => 
                           n6526, ZN => n2212);
   U7961 : NAND2_X1 port map( A1 => n17989, A2 => n28142, ZN => n2213);
   U7962 : NAND2_X1 port map( A1 => n28142, A2 => n6927, ZN => n2215);
   U7964 : NAND2_X1 port map( A1 => n2218, A2 => n2217, ZN => n13036);
   U7965 : NAND3_X1 port map( A1 => n2219, A2 => n10700, A3 => n11363, ZN => 
                           n2218);
   U7966 : NAND2_X1 port map( A1 => n2220, A2 => n4712, ZN => n10515);
   U7967 : NAND2_X1 port map( A1 => n6075, A2 => n11870, ZN => n2220);
   U7968 : AND2_X1 port map( A1 => n8658, A2 => n8502, ZN => n8634);
   U7969 : NAND2_X1 port map( A1 => n2226, A2 => n2225, ZN => n2221);
   U7970 : NAND2_X1 port map( A1 => n2224, A2 => n2223, ZN => n2222);
   U7971 : INV_X1 port map( A => n7885, ZN => n2225);
   U7972 : NAND3_X1 port map( A1 => n591, A2 => n10972, A3 => n28608, ZN => 
                           n4045);
   U7974 : INV_X1 port map( A => n2232, ZN => n12015);
   U7975 : NAND3_X1 port map( A1 => n11887, A2 => n11886, A3 => n12332, ZN => 
                           n2232);
   U7976 : NAND2_X1 port map( A1 => n10535, A2 => n10878, ZN => n2227);
   U7977 : AOI21_X1 port map( B1 => n11222, B2 => n435, A => n11219, ZN => 
                           n2228);
   U7978 : AOI21_X1 port map( B1 => n7410, B2 => n9340, A => n2230, ZN => n2229
                           );
   U7979 : OAI21_X1 port map( B1 => n9132, B2 => n9340, A => n8342, ZN => n2230
                           );
   U7980 : OAI21_X1 port map( B1 => n601, B2 => n9131, A => n2231, ZN => n9341)
                           ;
   U7981 : NAND3_X1 port map( A1 => n7410, A2 => n8753, A3 => n600, ZN => n2231
                           );
   U7984 : NAND3_X1 port map( A1 => n1166, A2 => n17229, A3 => n17038, ZN => 
                           n2234);
   U7986 : NAND3_X1 port map( A1 => n7585, A2 => n7886, A3 => n7071, ZN => 
                           n2236);
   U7987 : INV_X2 port map( A => n7887, ZN => n7585);
   U7988 : NAND3_X1 port map( A1 => n7580, A2 => n7885, A3 => n7583, ZN => 
                           n2237);
   U7989 : NAND2_X1 port map( A1 => n2238, A2 => n8521, ZN => n8524);
   U7990 : NAND2_X1 port map( A1 => n2238, A2 => n8811, ZN => n8813);
   U7991 : NAND3_X1 port map( A1 => n2238, A2 => n8521, A3 => n8809, ZN => 
                           n8252);
   U7992 : AOI21_X1 port map( B1 => n8460, B2 => n8681, A => n2238, ZN => n8461
                           );
   U7993 : MUX2_X1 port map( A => n20444, B => n20443, S => n6843, Z => n19926)
                           ;
   U7994 : OAI22_X1 port map( A1 => n23747, A2 => n2239, B1 => n22978, B2 => 
                           n409, ZN => n22983);
   U7995 : OAI21_X1 port map( B1 => n23404, B2 => n23746, A => n2239, ZN => 
                           n5971);
   U7996 : NAND2_X1 port map( A1 => n2240, A2 => n24435, ZN => n24348);
   U7997 : NAND2_X1 port map( A1 => n403, A2 => n2240, ZN => n5348);
   U7998 : NAND2_X1 port map( A1 => n24433, A2 => n24434, ZN => n24188);
   U7999 : NAND2_X1 port map( A1 => n18588, A2 => n18595, ZN => n17837);
   U8000 : NAND2_X1 port map( A1 => n17840, A2 => n17835, ZN => n2241);
   U8001 : NAND2_X1 port map( A1 => n17208, A2 => n18129, ZN => n2243);
   U8003 : OAI21_X1 port map( B1 => n14958, B2 => n13865, A => n2244, ZN => 
                           n13866);
   U8004 : NAND2_X1 port map( A1 => n13861, A2 => n14958, ZN => n2244);
   U8006 : NAND2_X1 port map( A1 => n2246, A2 => n24810, ZN => n3001);
   U8007 : NOR2_X1 port map( A1 => n2251, A2 => n9009, ZN => n2248);
   U8009 : INV_X1 port map( A => n9009, ZN => n9191);
   U8010 : INV_X1 port map( A => n9184, ZN => n2251);
   U8012 : OR2_X1 port map( A1 => n7362, A2 => n7363, ZN => n8200);
   U8013 : NAND2_X1 port map( A1 => n10110, A2 => n10592, ZN => n2255);
   U8014 : NAND2_X1 port map( A1 => n9281, A2 => n10705, ZN => n2256);
   U8015 : NAND2_X1 port map( A1 => n2688, A2 => n2689, ZN => n11024);
   U8017 : XNOR2_X1 port map( A => n4042, B => n4043, ZN => n2257);
   U8020 : NAND2_X1 port map( A1 => n20980, A2 => n21811, ZN => n2258);
   U8022 : MUX2_X1 port map( A => n24736, B => n24735, S => n24734, Z => n24743
                           );
   U8023 : NAND2_X1 port map( A1 => n6118, A2 => n2260, ZN => n6117);
   U8024 : NAND2_X1 port map( A1 => n20726, A2 => n20986, ZN => n2260);
   U8025 : NAND2_X1 port map( A1 => n20177, A2 => n20173, ZN => n19058);
   U8026 : XNOR2_X1 port map( A => n19606, B => n19103, ZN => n18746);
   U8028 : NAND3_X1 port map( A1 => n18524, A2 => n18523, A3 => n17858, ZN => 
                           n17722);
   U8030 : XNOR2_X1 port map( A => n15007, B => n15452, ZN => n4990);
   U8031 : AND3_X2 port map( A1 => n2796, A2 => n2799, A3 => n2798, ZN => 
                           n21655);
   U8032 : INV_X1 port map( A => n7525, ZN => n7531);
   U8033 : NAND2_X1 port map( A1 => n8014, A2 => n7533, ZN => n7525);
   U8035 : NAND2_X1 port map( A1 => n14776, A2 => n14777, ZN => n16012);
   U8036 : NAND2_X1 port map( A1 => n18488, A2 => n18489, ZN => n15734);
   U8037 : NAND2_X1 port map( A1 => n17146, A2 => n17076, ZN => n16734);
   U8038 : NAND2_X1 port map( A1 => n1831, A2 => n11755, ZN => n11760);
   U8039 : OR2_X1 port map( A1 => n29114, A2 => n28820, ZN => n18790);
   U8040 : INV_X1 port map( A => n17235, ZN => n2701);
   U8043 : NAND3_X1 port map( A1 => n28068, A2 => n28067, A3 => n28069, ZN => 
                           n3262);
   U8044 : NAND2_X1 port map( A1 => n2263, A2 => n2262, ZN => n26725);
   U8045 : NAND2_X1 port map( A1 => n26720, A2 => n26215, ZN => n2262);
   U8046 : NAND2_X1 port map( A1 => n26719, A2 => n26718, ZN => n2263);
   U8049 : NAND2_X1 port map( A1 => n23894, A2 => n24322, ZN => n2265);
   U8050 : OR2_X1 port map( A1 => n23896, A2 => n24678, ZN => n2266);
   U8051 : NAND2_X1 port map( A1 => n27568, A2 => n2268, ZN => n2267);
   U8053 : MUX2_X1 port map( A => n25833, B => n25832, S => n26842, Z => n25834
                           );
   U8054 : NAND3_X1 port map( A1 => n2332, A2 => n2333, A3 => n811, ZN => 
                           n24080);
   U8056 : NAND2_X1 port map( A1 => n26333, A2 => n26836, ZN => n2269);
   U8057 : NAND2_X1 port map( A1 => n9197, A2 => n9206, ZN => n9000);
   U8058 : NAND2_X1 port map( A1 => n7637, A2 => n3428, ZN => n9197);
   U8059 : NAND2_X1 port map( A1 => n7362, A2 => n7634, ZN => n7636);
   U8061 : NAND2_X1 port map( A1 => n6685, A2 => n28908, ZN => n24362);
   U8062 : NAND2_X1 port map( A1 => n24827, A2 => n24828, ZN => n24829);
   U8063 : NAND2_X1 port map( A1 => n20027, A2 => n20273, ZN => n20030);
   U8065 : NAND2_X1 port map( A1 => n10447, A2 => n10446, ZN => n2271);
   U8067 : NAND2_X1 port map( A1 => n7813, A2 => n28627, ZN => n2273);
   U8069 : NAND2_X1 port map( A1 => n27827, A2 => n2275, ZN => n5336);
   U8070 : NAND2_X1 port map( A1 => n27841, A2 => n27101, ZN => n2275);
   U8071 : NAND3_X1 port map( A1 => n2276, A2 => n27765, A3 => n27764, ZN => 
                           n27767);
   U8072 : NAND2_X1 port map( A1 => n27785, A2 => n6419, ZN => n2276);
   U8075 : OAI21_X1 port map( B1 => n15055, B2 => n15259, A => n2278, ZN => 
                           n4418);
   U8076 : NAND2_X1 port map( A1 => n15259, A2 => n14761, ZN => n2278);
   U8077 : NAND2_X1 port map( A1 => n5684, A2 => n21322, ZN => n21588);
   U8078 : NAND3_X2 port map( A1 => n3194, A2 => n3193, A3 => n20555, ZN => 
                           n21322);
   U8081 : NAND2_X1 port map( A1 => n19561, A2 => n19562, ZN => n17797);
   U8083 : NAND2_X1 port map( A1 => n3552, A2 => n12255, ZN => n2709);
   U8084 : NAND3_X1 port map( A1 => n7769, A2 => n7768, A3 => n7767, ZN => 
                           n3183);
   U8086 : XOR2_X1 port map( A => n9619, B => n629, Z => n5896);
   U8087 : AOI21_X2 port map( B1 => n2281, B2 => n2282, A => n22862, ZN => 
                           n4917);
   U8088 : INV_X1 port map( A => n22861, ZN => n2282);
   U8089 : INV_X1 port map( A => n10657, ZN => n11222);
   U8090 : XNOR2_X1 port map( A => n4493, B => n16283, ZN => n15965);
   U8091 : INV_X1 port map( A => n7496, ZN => n3594);
   U8092 : AND2_X1 port map( A1 => n4320, A2 => n8367, ZN => n2340);
   U8093 : XNOR2_X1 port map( A => n10063, B => n10062, ZN => n5150);
   U8097 : NAND2_X1 port map( A1 => n8993, A2 => n9434, ZN => n3056);
   U8098 : XNOR2_X1 port map( A => n2285, B => n25054, ZN => n25058);
   U8099 : XNOR2_X1 port map( A => n25053, B => n26108, ZN => n2285);
   U8100 : NAND2_X1 port map( A1 => n26781, A2 => n26919, ZN => n3390);
   U8102 : NAND2_X1 port map( A1 => n4672, A2 => n22863, ZN => n6338);
   U8105 : NOR2_X1 port map( A1 => n23067, A2 => n28164, ZN => n2286);
   U8107 : INV_X1 port map( A => n23137, ZN => n23136);
   U8108 : NAND2_X1 port map( A1 => n23067, A2 => n28164, ZN => n23137);
   U8109 : NAND2_X1 port map( A1 => n2289, A2 => n9169, ZN => n9172);
   U8113 : OR2_X1 port map( A1 => n7654, A2 => n7653, ZN => n7679);
   U8114 : AND2_X1 port map( A1 => n10856, A2 => n5835, ZN => n11313);
   U8115 : XNOR2_X1 port map( A => n2291, B => n9770, ZN => n9343);
   U8116 : XNOR2_X1 port map( A => n9339, B => n10385, ZN => n2291);
   U8117 : INV_X1 port map( A => n18273, ZN => n2292);
   U8118 : NOR2_X1 port map( A1 => n4211, A2 => n18516, ZN => n18273);
   U8119 : NAND2_X1 port map( A1 => n8178, A2 => n8179, ZN => n8180);
   U8120 : NAND2_X1 port map( A1 => n29631, A2 => n26950, ZN => n26442);
   U8121 : AND2_X1 port map( A1 => n2748, A2 => n6482, ZN => n11789);
   U8122 : OR2_X1 port map( A1 => n20333, A2 => n20630, ZN => n19328);
   U8124 : INV_X1 port map( A => n14807, ZN => n14715);
   U8125 : INV_X1 port map( A => n4105, ZN => n12408);
   U8126 : XNOR2_X1 port map( A => n19183, B => n18649, ZN => n20563);
   U8127 : XNOR2_X1 port map( A => n12831, B => n12828, ZN => n2293);
   U8128 : OR2_X1 port map( A1 => n10318, A2 => n11287, ZN => n10664);
   U8129 : OR2_X1 port map( A1 => n9364, A2 => n3274, ZN => n3272);
   U8130 : INV_X1 port map( A => n21714, ZN => n20976);
   U8132 : NAND2_X1 port map( A1 => n17004, A2 => n15981, ZN => n4614);
   U8133 : NAND2_X1 port map( A1 => n15423, A2 => n15102, ZN => n15421);
   U8135 : NAND2_X1 port map( A1 => n12888, A2 => n14438, ZN => n2294);
   U8136 : OAI22_X1 port map( A1 => n24674, A2 => n29555, B1 => n24322, B2 => 
                           n24397, ZN => n2379);
   U8137 : OR2_X1 port map( A1 => n4854, A2 => n18159, ZN => n17326);
   U8138 : NAND2_X1 port map( A1 => n20955, A2 => n21090, ZN => n2296);
   U8139 : XNOR2_X2 port map( A => n2297, B => Key(15), ZN => n8177);
   U8140 : INV_X1 port map( A => Plaintext(15), ZN => n2297);
   U8142 : NOR2_X2 port map( A1 => n23491, A2 => n23490, ZN => n23946);
   U8145 : XNOR2_X1 port map( A => n25772, B => n2300, ZN => n25259);
   U8146 : XNOR2_X1 port map( A => n25257, B => n25546, ZN => n2300);
   U8147 : OAI21_X1 port map( B1 => n21515, B2 => n21516, A => n2301, ZN => 
                           n21517);
   U8148 : NAND3_X1 port map( A1 => n21532, A2 => n21514, A3 => n21513, ZN => 
                           n2301);
   U8150 : NAND3_X1 port map( A1 => n3740, A2 => n2832, A3 => n7590, ZN => 
                           n6802);
   U8152 : NAND2_X1 port map( A1 => n2335, A2 => n8560, ZN => n2334);
   U8153 : AND2_X1 port map( A1 => n11473, A2 => n12337, ZN => n5466);
   U8154 : NAND2_X1 port map( A1 => n13850, A2 => n14176, ZN => n2304);
   U8155 : OAI211_X1 port map( C1 => n20157, C2 => n20160, A => n19985, B => 
                           n2305, ZN => n4235);
   U8156 : NAND2_X1 port map( A1 => n20157, A2 => n29066, ZN => n2305);
   U8157 : NAND2_X1 port map( A1 => n21608, A2 => n2307, ZN => n21335);
   U8158 : NAND3_X2 port map( A1 => n2308, A2 => n8450, A3 => n8449, ZN => 
                           n10038);
   U8159 : OAI211_X1 port map( C1 => n9195, C2 => n9201, A => n2309, B => n8779
                           , ZN => n2308);
   U8160 : INV_X1 port map( A => n8451, ZN => n2309);
   U8161 : INV_X1 port map( A => n2311, ZN => n2310);
   U8162 : OAI21_X1 port map( B1 => n7347, B2 => n7759, A => n7763, ZN => n2311
                           );
   U8163 : NAND2_X1 port map( A1 => n21367, A2 => n21366, ZN => n2312);
   U8165 : XOR2_X1 port map( A => n9678, B => n9619, Z => n6796);
   U8166 : AOI22_X2 port map( A1 => n4176, A2 => n24408, B1 => n24407, B2 => 
                           n24406, ZN => n25345);
   U8167 : NOR2_X1 port map( A1 => n17249, A2 => n16977, ZN => n4863);
   U8168 : NAND2_X1 port map( A1 => n2313, A2 => n6699, ZN => n5577);
   U8169 : NAND4_X1 port map( A1 => n14705, A2 => n14447, A3 => n14448, A4 => 
                           n14449, ZN => n2313);
   U8170 : XNOR2_X1 port map( A => n15914, B => n16296, ZN => n16103);
   U8171 : AOI21_X2 port map( B1 => n6262, B2 => n15405, A => n15404, ZN => 
                           n15914);
   U8172 : AOI22_X1 port map( A1 => n421, A2 => n17119, B1 => n17121, B2 => 
                           n17120, ZN => n2314);
   U8173 : NAND2_X1 port map( A1 => n15462, A2 => n15464, ZN => n4513);
   U8174 : AND3_X2 port map( A1 => n13883, A2 => n13882, A3 => n13881, ZN => 
                           n15462);
   U8175 : NAND2_X1 port map( A1 => n16925, A2 => n16926, ZN => n16927);
   U8176 : NAND2_X1 port map( A1 => n24046, A2 => n24484, ZN => n24047);
   U8178 : NAND3_X1 port map( A1 => n11999, A2 => n11998, A3 => n11997, ZN => 
                           n2604);
   U8179 : AOI21_X1 port map( B1 => n21625, B2 => n22145, A => n22143, ZN => 
                           n21109);
   U8181 : OAI21_X1 port map( B1 => n8501, B2 => n8502, A => n8115, ZN => n8118
                           );
   U8182 : OR2_X2 port map( A1 => n2315, A2 => n9476, ZN => n13081);
   U8183 : AOI21_X1 port map( B1 => n9467, B2 => n10108, A => n588, ZN => n2315
                           );
   U8184 : NAND2_X1 port map( A1 => n524, A2 => n2316, ZN => n17578);
   U8185 : NAND2_X1 port map( A1 => n2837, A2 => n2836, ZN => n2318);
   U8186 : INV_X1 port map( A => n10834, ZN => n3820);
   U8189 : INV_X1 port map( A => n9793, ZN => n9515);
   U8190 : XNOR2_X1 port map( A => n5818, B => n9514, ZN => n9793);
   U8191 : XNOR2_X2 port map( A => n7087, B => Key(5), ZN => n7775);
   U8192 : AOI22_X1 port map( A1 => n4433, A2 => n1959, B1 => n13951, B2 => 
                           n4049, ZN => n4050);
   U8194 : NAND2_X1 port map( A1 => n8767, A2 => n604, ZN => n8580);
   U8195 : NAND2_X1 port map( A1 => n2496, A2 => n15098, ZN => n2495);
   U8197 : NAND2_X1 port map( A1 => n6069, A2 => n29610, ZN => n6068);
   U8199 : NAND2_X1 port map( A1 => n10682, A2 => n5265, ZN => n11493);
   U8200 : OR2_X1 port map( A1 => n20916, A2 => n18934, ZN => n18933);
   U8201 : INV_X1 port map( A => n7770, ZN => n7767);
   U8202 : AND2_X1 port map( A1 => n14958, A2 => n15476, ZN => n15169);
   U8205 : OR2_X1 port map( A1 => n12228, A2 => n13081, ZN => n11688);
   U8206 : INV_X1 port map( A => n18193, ZN => n6663);
   U8207 : INV_X1 port map( A => n23433, ZN => n5530);
   U8208 : INV_X1 port map( A => n1938, ZN => n7964);
   U8209 : NOR2_X1 port map( A1 => n14158, A2 => n14475, ZN => n3867);
   U8210 : OAI211_X1 port map( C1 => n27508, C2 => n27520, A => n4165, B => 
                           n4164, ZN => n27519);
   U8211 : XNOR2_X1 port map( A => n10070, B => n10069, ZN => n10752);
   U8212 : AND2_X1 port map( A1 => n28776, A2 => n17379, ZN => n6501);
   U8213 : XNOR2_X1 port map( A => n4298, B => n12559, ZN => n12775);
   U8214 : XNOR2_X1 port map( A => n19500, B => n1923, ZN => n4221);
   U8215 : NAND2_X1 port map( A1 => n11846, A2 => n11515, ZN => n2319);
   U8216 : NAND2_X1 port map( A1 => n8155, A2 => n7785, ZN => n7171);
   U8217 : NAND2_X1 port map( A1 => n7168, A2 => n7167, ZN => n8155);
   U8218 : AND3_X2 port map( A1 => n4398, A2 => n14011, A3 => n14012, ZN => 
                           n14821);
   U8219 : NOR2_X1 port map( A1 => n18261, A2 => n18326, ZN => n17713);
   U8220 : INV_X1 port map( A => n2779, ZN => n23470);
   U8221 : NOR2_X1 port map( A1 => n2735, A2 => n20088, ZN => n20040);
   U8222 : NAND2_X1 port map( A1 => n2128, A2 => n8726, ZN => n8852);
   U8224 : NAND2_X1 port map( A1 => n28210, A2 => n9029, ZN => n8795);
   U8226 : NAND2_X1 port map( A1 => n2324, A2 => n2323, ZN => n27304);
   U8227 : NAND2_X1 port map( A1 => n26421, A2 => n28471, ZN => n2324);
   U8228 : NAND3_X1 port map( A1 => n11856, A2 => n12155, A3 => n12088, ZN => 
                           n3008);
   U8230 : NAND2_X1 port map( A1 => n29241, A2 => n8251, ZN => n3224);
   U8231 : OR2_X1 port map( A1 => n7890, A2 => n7891, ZN => n7275);
   U8232 : NAND2_X1 port map( A1 => n25406, A2 => n26191, ZN => n25618);
   U8233 : OR2_X2 port map( A1 => n11200, A2 => n5660, ZN => n13118);
   U8234 : INV_X1 port map( A => Plaintext(156), ZN => n7046);
   U8235 : NAND3_X1 port map( A1 => n23538, A2 => n23536, A3 => n23689, ZN => 
                           n2326);
   U8236 : NAND2_X1 port map( A1 => n5567, A2 => n9232, ZN => n9049);
   U8237 : NAND2_X1 port map( A1 => n15022, A2 => n15303, ZN => n15025);
   U8238 : NAND2_X1 port map( A1 => n13931, A2 => n2327, ZN => n15303);
   U8240 : NAND2_X1 port map( A1 => n18172, A2 => n18170, ZN => n2329);
   U8241 : NAND2_X1 port map( A1 => n17783, A2 => n18173, ZN => n2330);
   U8242 : NAND2_X1 port map( A1 => n5272, A2 => n5728, ZN => n2332);
   U8243 : NAND2_X1 port map( A1 => n5272, A2 => n24079, ZN => n2333);
   U8244 : NAND2_X1 port map( A1 => n4193, A2 => n21457, ZN => n6803);
   U8245 : OR2_X1 port map( A1 => n13646, A2 => n13816, ZN => n5180);
   U8246 : XNOR2_X1 port map( A => n12069, B => n12699, ZN => n13438);
   U8247 : OR2_X1 port map( A1 => n3936, A2 => n28580, ZN => n3619);
   U8248 : NOR2_X1 port map( A1 => n11449, A2 => n12328, ZN => n12014);
   U8249 : INV_X1 port map( A => n13646, ZN => n14299);
   U8250 : INV_X1 port map( A => n9913, ZN => n11127);
   U8251 : XNOR2_X1 port map( A => n19520, B => n18691, ZN => n19066);
   U8252 : NAND3_X1 port map( A1 => n10586, A2 => n12354, A3 => n11467, ZN => 
                           n11469);
   U8253 : NAND2_X1 port map( A1 => n5001, A2 => n17018, ZN => n17254);
   U8254 : NAND2_X1 port map( A1 => n7980, A2 => n7641, ZN => n7193);
   U8255 : NAND2_X1 port map( A1 => n29077, A2 => n10912, ZN => n10688);
   U8256 : NAND3_X1 port map( A1 => n21614, A2 => n28791, A3 => n2337, ZN => 
                           n21616);
   U8257 : NAND2_X1 port map( A1 => n21609, A2 => n2338, ZN => n2337);
   U8258 : NAND3_X1 port map( A1 => n6293, A2 => n15512, A3 => n15514, ZN => 
                           n15517);
   U8259 : NAND2_X1 port map( A1 => n4318, A2 => n2340, ZN => n9823);
   U8260 : OAI21_X1 port map( B1 => n10476, B2 => n11347, A => n2342, ZN => 
                           n11356);
   U8261 : NAND2_X1 port map( A1 => n11347, A2 => n11350, ZN => n2342);
   U8263 : NAND2_X1 port map( A1 => n6210, A2 => n7507, ZN => n2789);
   U8265 : NAND2_X1 port map( A1 => n2345, A2 => n14400, ZN => n2344);
   U8266 : INV_X1 port map( A => n13877, ZN => n2345);
   U8267 : OR2_X1 port map( A1 => n14398, A2 => n14400, ZN => n2346);
   U8268 : NAND2_X1 port map( A1 => n15514, A2 => n14697, ZN => n2347);
   U8270 : XNOR2_X1 port map( A => n15642, B => n16421, ZN => n15644);
   U8271 : NAND2_X2 port map( A1 => n4708, A2 => n14699, ZN => n16421);
   U8272 : NAND2_X1 port map( A1 => n11880, A2 => n11881, ZN => n2348);
   U8273 : NAND2_X1 port map( A1 => n11879, A2 => n287, ZN => n2349);
   U8274 : NAND2_X1 port map( A1 => n21661, A2 => n20833, ZN => n21073);
   U8275 : NAND2_X1 port map( A1 => n7746, A2 => n7533, ZN => n7143);
   U8277 : NAND2_X1 port map( A1 => n2614, A2 => n10712, ZN => n11774);
   U8278 : NAND3_X1 port map( A1 => n6738, A2 => n27427, A3 => n29542, ZN => 
                           n26968);
   U8279 : NAND2_X1 port map( A1 => n17116, A2 => n29539, ZN => n3100);
   U8280 : OAI211_X2 port map( C1 => n24045, C2 => n24044, A => n2828, B => 
                           n2829, ZN => n26053);
   U8281 : NAND2_X1 port map( A1 => n5888, A2 => n2352, ZN => n9226);
   U8283 : NAND3_X1 port map( A1 => n2794, A2 => n27746, A3 => n2795, ZN => 
                           n2793);
   U8287 : NAND2_X1 port map( A1 => n15315, A2 => n15319, ZN => n15316);
   U8288 : MUX2_X1 port map( A => n18337, B => n18331, S => n18332, Z => n17651
                           );
   U8292 : NAND3_X1 port map( A1 => n11196, A2 => n10751, A3 => n28207, ZN => 
                           n2431);
   U8294 : AOI21_X1 port map( B1 => n14924, B2 => n14923, A => n15497, ZN => 
                           n14925);
   U8296 : NAND2_X1 port map( A1 => n10646, A2 => n12027, ZN => n10647);
   U8299 : NAND3_X1 port map( A1 => n1931, A2 => n12162, A3 => n2357, ZN => 
                           n11380);
   U8300 : INV_X1 port map( A => n12103, ZN => n2357);
   U8301 : XOR2_X1 port map( A => n19699, B => n19698, Z => n5006);
   U8302 : OR2_X1 port map( A1 => n17269, A2 => n29299, ZN => n3038);
   U8303 : OAI22_X1 port map( A1 => n6034, A2 => n23686, B1 => n23168, B2 => 
                           n23679, ZN => n23134);
   U8304 : NAND3_X2 port map( A1 => n2359, A2 => n2780, A3 => n2358, ZN => 
                           n9184);
   U8305 : NAND2_X1 port map( A1 => n2781, A2 => n7141, ZN => n2359);
   U8306 : NAND3_X1 port map( A1 => n11790, A2 => n11791, A3 => n2360, ZN => 
                           n11792);
   U8307 : NAND2_X1 port map( A1 => n2361, A2 => n26729, ZN => n25628);
   U8308 : OAI21_X1 port map( B1 => n2361, B2 => n26729, A => n26728, ZN => 
                           n26730);
   U8309 : INV_X1 port map( A => n26481, ZN => n2361);
   U8310 : MUX2_X1 port map( A => n10912, B => n29078, S => n10911, Z => n10917
                           );
   U8311 : OAI21_X1 port map( B1 => n10689, B2 => n10911, A => n29078, ZN => 
                           n10690);
   U8312 : AOI21_X1 port map( B1 => n10914, B2 => n10605, A => n29077, ZN => 
                           n10452);
   U8313 : NAND2_X1 port map( A1 => n10915, A2 => n29077, ZN => n10606);
   U8315 : AND2_X1 port map( A1 => n2363, A2 => n18215, ZN => n18502);
   U8316 : INV_X1 port map( A => n18216, ZN => n2363);
   U8317 : NAND2_X1 port map( A1 => n5692, A2 => n2364, ZN => n5691);
   U8318 : INV_X1 port map( A => n18215, ZN => n2364);
   U8319 : NAND2_X1 port map( A1 => n5154, A2 => n2365, ZN => n17727);
   U8320 : NAND2_X1 port map( A1 => n5690, A2 => n18215, ZN => n2365);
   U8321 : NAND2_X1 port map( A1 => n14634, A2 => n14635, ZN => n16567);
   U8322 : OR2_X2 port map( A1 => n13845, A2 => n13846, ZN => n15738);
   U8324 : INV_X1 port map( A => n10985, ZN => n3802);
   U8325 : AOI22_X2 port map( A1 => n23933, A2 => n24291, B1 => n23934, B2 => 
                           n24730, ZN => n25808);
   U8327 : XNOR2_X1 port map( A => n12753, B => n13136, ZN => n13328);
   U8328 : NAND3_X1 port map( A1 => n5659, A2 => n514, A3 => n17906, ZN => 
                           n4076);
   U8329 : NAND2_X1 port map( A1 => n2366, A2 => n23830, ZN => n24095);
   U8330 : NAND2_X1 port map( A1 => n481, A2 => n23833, ZN => n23830);
   U8331 : INV_X1 port map( A => n2367, ZN => n2366);
   U8332 : NAND3_X1 port map( A1 => n2368, A2 => n8977, A3 => n8818, ZN => 
                           n8822);
   U8333 : NAND2_X1 port map( A1 => n8974, A2 => n8817, ZN => n2368);
   U8334 : XNOR2_X1 port map( A => n9977, B => n2034, ZN => n6916);
   U8335 : NAND2_X1 port map( A1 => n2369, A2 => n4554, ZN => n10102);
   U8336 : NAND2_X1 port map( A1 => n4553, A2 => n4555, ZN => n2369);
   U8337 : NAND2_X1 port map( A1 => n20579, A2 => n20417, ZN => n2371);
   U8338 : NAND2_X1 port map( A1 => n20578, A2 => n20577, ZN => n2372);
   U8340 : OAI22_X1 port map( A1 => n5064, A2 => n6011, B1 => n13909, B2 => 
                           n14043, ZN => n2373);
   U8341 : XNOR2_X2 port map( A => n2374, B => Key(108), ZN => n8217);
   U8342 : INV_X1 port map( A => Plaintext(108), ZN => n2374);
   U8344 : NAND2_X1 port map( A1 => n2377, A2 => n2376, ZN => n26873);
   U8345 : OAI21_X1 port map( B1 => n3236, B2 => n26902, A => n2378, ZN => 
                           n2377);
   U8346 : NOR2_X2 port map( A1 => n24069, A2 => n2379, ZN => n25809);
   U8347 : OAI211_X1 port map( C1 => n27478, C2 => n27492, A => n2380, B => 
                           n5606, ZN => n26704);
   U8348 : NAND2_X1 port map( A1 => n2882, A2 => n2883, ZN => n2382);
   U8352 : NAND2_X1 port map( A1 => n3005, A2 => n20481, ZN => n2383);
   U8354 : NAND2_X1 port map( A1 => n5147, A2 => n7604, ZN => n8735);
   U8355 : XNOR2_X1 port map( A => n2384, B => n9932, ZN => n4600);
   U8356 : XNOR2_X1 port map( A => n9928, B => n9929, ZN => n2384);
   U8357 : AND2_X1 port map( A1 => n14336, A2 => n14408, ZN => n13813);
   U8358 : OR2_X1 port map( A1 => n17304, A2 => n5714, ZN => n16788);
   U8359 : OR2_X1 port map( A1 => n18456, A2 => n4230, ZN => n16793);
   U8360 : INV_X1 port map( A => n20090, ZN => n20091);
   U8361 : NAND2_X1 port map( A1 => n2386, A2 => n1568, ZN => n4695);
   U8362 : OAI21_X1 port map( B1 => n4696, B2 => n29301, A => n3642, ZN => 
                           n2386);
   U8363 : OAI21_X1 port map( B1 => n12232, B2 => n776, A => n2412, ZN => 
                           n12039);
   U8365 : INV_X1 port map( A => Plaintext(164), ZN => n2387);
   U8366 : NAND2_X1 port map( A1 => n2917, A2 => n3331, ZN => n2388);
   U8368 : NAND2_X1 port map( A1 => n6843, A2 => n20133, ZN => n2390);
   U8369 : NAND2_X1 port map( A1 => n2391, A2 => n8168, ZN => n2942);
   U8370 : NAND2_X1 port map( A1 => n7536, A2 => n7352, ZN => n2391);
   U8372 : XNOR2_X1 port map( A => n2392, B => n3633, ZN => Ciphertext(76));
   U8373 : NOR2_X1 port map( A1 => n27206, A2 => n27207, ZN => n2392);
   U8374 : OR2_X1 port map( A1 => n14197, A2 => n28199, ZN => n14198);
   U8377 : XNOR2_X1 port map( A => n22275, B => n22485, ZN => n2393);
   U8378 : XNOR2_X1 port map( A => n2394, B => n22170, ZN => n22173);
   U8379 : XNOR2_X1 port map( A => n22171, B => n28387, ZN => n2394);
   U8380 : NAND2_X1 port map( A1 => n21394, A2 => n2395, ZN => n2409);
   U8382 : NAND2_X1 port map( A1 => n2918, A2 => n20863, ZN => n2396);
   U8384 : NAND3_X2 port map( A1 => n2397, A2 => n3487, A3 => n13518, ZN => 
                           n16312);
   U8385 : NAND2_X1 port map( A1 => n6668, A2 => n14884, ZN => n2397);
   U8386 : NAND3_X1 port map( A1 => n15717, A2 => n17366, A3 => n15731, ZN => 
                           n15733);
   U8387 : NOR2_X1 port map( A1 => n8301, A2 => n7400, ZN => n3203);
   U8388 : NAND2_X1 port map( A1 => n11908, A2 => n12363, ZN => n11446);
   U8389 : NAND2_X1 port map( A1 => n14231, A2 => n14230, ZN => n3645);
   U8390 : OR2_X1 port map( A1 => n17374, A2 => n17379, ZN => n4651);
   U8391 : NAND2_X1 port map( A1 => n21328, A2 => n21330, ZN => n21163);
   U8392 : NOR2_X1 port map( A1 => n29526, A2 => n21373, ZN => n21273);
   U8393 : NAND2_X1 port map( A1 => n2399, A2 => n2398, ZN => n3058);
   U8394 : AOI21_X1 port map( B1 => n349, B2 => n12072, A => n12251, ZN => 
                           n2398);
   U8395 : NAND2_X1 port map( A1 => n11933, A2 => n12249, ZN => n2399);
   U8396 : OAI21_X1 port map( B1 => n23417, B2 => n485, A => n2400, ZN => 
                           n23420);
   U8397 : XNOR2_X1 port map( A => n9811, B => n2401, ZN => n9813);
   U8398 : XNOR2_X1 port map( A => n9810, B => n10071, ZN => n2401);
   U8400 : INV_X1 port map( A => Plaintext(168), ZN => n6208);
   U8401 : INV_X1 port map( A => n18762, ZN => n3913);
   U8402 : NAND3_X1 port map( A1 => n9436, A2 => n9211, A3 => n9209, ZN => 
                           n7682);
   U8406 : AOI21_X1 port map( B1 => n2898, B2 => n8291, A => n8287, ZN => n2406
                           );
   U8407 : OAI21_X1 port map( B1 => n27791, B2 => n2407, A => n27800, ZN => 
                           n27792);
   U8408 : NOR2_X1 port map( A1 => n27790, A2 => n27819, ZN => n2407);
   U8409 : NAND2_X1 port map( A1 => n17763, A2 => n17873, ZN => n17764);
   U8410 : NAND2_X1 port map( A1 => n19833, A2 => n20382, ZN => n5943);
   U8412 : NAND2_X1 port map( A1 => n11235, A2 => n11013, ZN => n11016);
   U8413 : AOI21_X1 port map( B1 => n3464, B2 => n7238, A => n7885, ZN => n5174
                           );
   U8414 : INV_X1 port map( A => n8801, ZN => n9160);
   U8415 : OAI21_X1 port map( B1 => n2945, B2 => n13747, A => n13763, ZN => 
                           n2408);
   U8416 : OR2_X1 port map( A1 => n9124, A2 => n284, ZN => n4060);
   U8417 : NOR2_X1 port map( A1 => n10706, A2 => n10942, ZN => n10447);
   U8418 : INV_X1 port map( A => n8136, ZN => n7127);
   U8419 : INV_X1 port map( A => n23448, ZN => n4794);
   U8420 : INV_X1 port map( A => n14259, ZN => n2681);
   U8421 : INV_X1 port map( A => n14981, ZN => n5635);
   U8422 : NAND2_X1 port map( A1 => n21398, A2 => n2409, ZN => n22158);
   U8423 : XNOR2_X2 port map( A => n7108, B => Key(188), ZN => n7900);
   U8424 : NAND2_X1 port map( A1 => n7800, A2 => n7801, ZN => n7802);
   U8425 : NAND2_X1 port map( A1 => n7127, A2 => n29646, ZN => n8052);
   U8426 : NAND2_X1 port map( A1 => n14262, A2 => n14260, ZN => n14098);
   U8428 : NAND2_X1 port map( A1 => n23376, A2 => n23377, ZN => n23381);
   U8430 : NAND2_X1 port map( A1 => n23497, A2 => n23493, ZN => n23796);
   U8432 : NAND3_X1 port map( A1 => n8830, A2 => n1839, A3 => n8829, ZN => 
                           n2410);
   U8433 : NOR2_X1 port map( A1 => n18286, A2 => n18524, ZN => n18082);
   U8434 : AND2_X2 port map( A1 => n4427, A2 => n4428, ZN => n17719);
   U8435 : INV_X1 port map( A => n2413, ZN => n10629);
   U8436 : NAND2_X1 port map( A1 => n12232, A2 => n12234, ZN => n2412);
   U8437 : NAND2_X1 port map( A1 => n14702, A2 => n14916, ZN => n15495);
   U8438 : NAND2_X1 port map( A1 => n27631, A2 => n27630, ZN => n2415);
   U8439 : INV_X1 port map( A => n17415, ZN => n15811);
   U8440 : NAND2_X1 port map( A1 => n2417, A2 => n17415, ZN => n2416);
   U8441 : INV_X1 port map( A => n17413, ZN => n2417);
   U8442 : NAND2_X1 port map( A1 => n2419, A2 => n9188, ZN => n2418);
   U8443 : NAND2_X1 port map( A1 => n9187, A2 => n9186, ZN => n2419);
   U8444 : NAND2_X1 port map( A1 => n9189, A2 => n8445, ZN => n2420);
   U8447 : NAND2_X1 port map( A1 => n10697, A2 => n10989, ZN => n2423);
   U8449 : NAND2_X1 port map( A1 => n4577, A2 => n7579, ZN => n2424);
   U8450 : NAND2_X1 port map( A1 => n3379, A2 => n14141, ZN => n13717);
   U8452 : NOR2_X1 port map( A1 => n8956, A2 => n8954, ZN => n2425);
   U8453 : INV_X1 port map( A => n21364, ZN => n5772);
   U8454 : XOR2_X1 port map( A => n13398, B => n13397, Z => n2875);
   U8455 : OAI21_X1 port map( B1 => n27359, B2 => n27360, A => n2426, ZN => 
                           n27361);
   U8456 : NAND2_X1 port map( A1 => n6766, A2 => n6767, ZN => n6769);
   U8457 : NAND2_X1 port map( A1 => n20853, A2 => n2427, ZN => n20855);
   U8460 : NAND3_X1 port map( A1 => n4560, A2 => n4562, A3 => n2036, ZN => 
                           n24138);
   U8461 : NOR2_X1 port map( A1 => n27230, A2 => n2428, ZN => n27232);
   U8462 : OAI22_X1 port map( A1 => n27229, A2 => n27757, B1 => n27228, B2 => 
                           n29049, ZN => n2428);
   U8463 : OAI211_X2 port map( C1 => n9194, C2 => n7639, A => n7638, B => n2429
                           , ZN => n9772);
   U8464 : NAND2_X1 port map( A1 => n6897, A2 => n9202, ZN => n2429);
   U8466 : NAND2_X1 port map( A1 => n10869, A2 => n11453, ZN => n2430);
   U8467 : NAND2_X1 port map( A1 => n11595, A2 => n12251, ZN => n2710);
   U8468 : XNOR2_X2 port map( A => n9432, B => n5895, ZN => n10936);
   U8469 : OR2_X1 port map( A1 => n8762, A2 => n8553, ZN => n8557);
   U8472 : NAND3_X1 port map( A1 => n8488, A2 => n8899, A3 => n1793, ZN => 
                           n6317);
   U8474 : NAND2_X1 port map( A1 => n4941, A2 => n3148, ZN => n8132);
   U8476 : NAND2_X1 port map( A1 => n27217, A2 => n2433, ZN => n2432);
   U8477 : INV_X1 port map( A => n27562, ZN => n2433);
   U8478 : NAND2_X1 port map( A1 => n27216, A2 => n27562, ZN => n2434);
   U8483 : INV_X1 port map( A => n27277, ZN => n2438);
   U8484 : NAND2_X1 port map( A1 => n27290, A2 => n27286, ZN => n2439);
   U8485 : INV_X1 port map( A => n21292, ZN => n20985);
   U8486 : OR2_X1 port map( A1 => n28626, A2 => n23099, ZN => n2451);
   U8489 : NAND2_X1 port map( A1 => n2442, A2 => n464, ZN => n3713);
   U8490 : INV_X1 port map( A => n9116, ZN => n8071);
   U8492 : NAND2_X1 port map( A1 => n17796, A2 => n2445, ZN => n2444);
   U8493 : INV_X1 port map( A => n18087, ZN => n2445);
   U8494 : NAND2_X1 port map( A1 => n13678, A2 => n12743, ZN => n14182);
   U8495 : NAND2_X1 port map( A1 => n4261, A2 => n1993, ZN => n13133);
   U8496 : NAND2_X1 port map( A1 => n13852, A2 => n13933, ZN => n14187);
   U8499 : NAND2_X1 port map( A1 => n15381, A2 => n15384, ZN => n2448);
   U8500 : NAND2_X1 port map( A1 => n4283, A2 => n17357, ZN => n2450);
   U8502 : XOR2_X1 port map( A => n13482, B => n27515, Z => n6652);
   U8503 : NAND2_X1 port map( A1 => n11072, A2 => n11075, ZN => n10891);
   U8504 : NAND2_X1 port map( A1 => n5352, A2 => n13827, ZN => n5351);
   U8505 : OAI211_X1 port map( C1 => n25954, C2 => n27317, A => n2454, B => 
                           n2453, ZN => n25955);
   U8506 : NAND2_X1 port map( A1 => n26594, A2 => n27317, ZN => n2453);
   U8507 : NAND2_X1 port map( A1 => n25897, A2 => n27873, ZN => n2454);
   U8508 : INV_X1 port map( A => n10008, ZN => n3073);
   U8509 : OR2_X1 port map( A1 => n5775, A2 => n22284, ZN => n23040);
   U8510 : XNOR2_X1 port map( A => n10138, B => n9735, ZN => n9918);
   U8511 : NAND2_X1 port map( A1 => n15294, A2 => n2455, ZN => n14836);
   U8512 : XNOR2_X1 port map( A => n6665, B => n6666, ZN => n10875);
   U8515 : XNOR2_X1 port map( A => n22439, B => n22440, ZN => n2779);
   U8517 : NAND2_X1 port map( A1 => n2458, A2 => n3831, ZN => n19277);
   U8518 : NAND3_X1 port map( A1 => n17714, A2 => n3832, A3 => n18323, ZN => 
                           n2458);
   U8520 : NAND2_X1 port map( A1 => n11414, A2 => n11415, ZN => n11418);
   U8521 : NAND3_X1 port map( A1 => n7952, A2 => n28614, A3 => n2461, ZN => 
                           n7951);
   U8522 : NAND2_X1 port map( A1 => n7946, A2 => n7947, ZN => n2461);
   U8524 : OAI21_X1 port map( B1 => n14281, B2 => n14285, A => n2462, ZN => 
                           n13621);
   U8525 : NAND2_X1 port map( A1 => n14285, A2 => n14287, ZN => n2462);
   U8526 : NAND4_X2 port map( A1 => n11624, A2 => n11625, A3 => n11627, A4 => 
                           n11626, ZN => n13567);
   U8527 : OAI21_X1 port map( B1 => n6386, B2 => n6385, A => n10888, ZN => 
                           n10889);
   U8530 : AND2_X2 port map( A1 => n3304, A2 => n3305, ZN => n22139);
   U8531 : XNOR2_X2 port map( A => n7166, B => Key(20), ZN => n7291);
   U8532 : NAND3_X1 port map( A1 => n5659, A2 => n17906, A3 => n17663, ZN => 
                           n5701);
   U8533 : NAND2_X1 port map( A1 => n28105, A2 => n29056, ZN => n2463);
   U8534 : OAI21_X2 port map( B1 => n17495, B2 => n16733, A => n16732, ZN => 
                           n18203);
   U8535 : OAI21_X1 port map( B1 => n7954, B2 => n8670, A => n7953, ZN => n7955
                           );
   U8536 : XOR2_X1 port map( A => n9672, B => n9671, Z => n4601);
   U8537 : NAND2_X1 port map( A1 => n12265, A2 => n2466, ZN => n11060);
   U8539 : OAI22_X1 port map( A1 => n14119, A2 => n14369, B1 => n14093, B2 => 
                           n564, ZN => n13835);
   U8540 : NAND2_X1 port map( A1 => n559, A2 => n14366, ZN => n14119);
   U8542 : NAND2_X1 port map( A1 => n11688, A2 => n11689, ZN => n11691);
   U8543 : OAI21_X1 port map( B1 => n612, B2 => n7981, A => n7642, ZN => n7454)
                           ;
   U8545 : NAND2_X1 port map( A1 => n8724, A2 => n8605, ZN => n2890);
   U8546 : XNOR2_X1 port map( A => n19412, B => n18857, ZN => n19097);
   U8547 : NAND2_X1 port map( A1 => n17167, A2 => n2468, ZN => n19412);
   U8548 : NAND2_X1 port map( A1 => n9221, A2 => n8525, ZN => n9224);
   U8549 : NAND4_X2 port map( A1 => n6330, A2 => n6329, A3 => n6328, A4 => 
                           n10465, ZN => n13097);
   U8551 : AOI21_X1 port map( B1 => n8893, B2 => n8892, A => n8891, ZN => n8894
                           );
   U8552 : NAND2_X1 port map( A1 => n8504, A2 => n8009, ZN => n8892);
   U8553 : NOR2_X1 port map( A1 => n2469, A2 => n2016, ZN => n23008);
   U8554 : OAI21_X1 port map( B1 => n21896, B2 => n23663, A => n23522, ZN => 
                           n2469);
   U8555 : NAND3_X1 port map( A1 => n3157, A2 => n3156, A3 => n9529, ZN => 
                           n9536);
   U8557 : NAND3_X1 port map( A1 => n7990, A2 => n2472, A3 => n2471, ZN => 
                           n2470);
   U8558 : NAND2_X1 port map( A1 => n29639, A2 => n341, ZN => n2471);
   U8559 : NAND3_X1 port map( A1 => n4647, A2 => n4646, A3 => n6206, ZN => 
                           n22227);
   U8560 : NAND2_X1 port map( A1 => n6526, A2 => n6927, ZN => n2935);
   U8562 : OAI21_X1 port map( B1 => n24496, B2 => n24497, A => n24810, ZN => 
                           n2473);
   U8563 : OR2_X1 port map( A1 => n14491, A2 => n14498, ZN => n2964);
   U8564 : NAND2_X1 port map( A1 => n28651, A2 => n28467, ZN => n25035);
   U8565 : INV_X1 port map( A => n20597, ZN => n20603);
   U8566 : XNOR2_X1 port map( A => n12872, B => n4375, ZN => n12652);
   U8567 : OR2_X2 port map( A1 => n5031, A2 => n3405, ZN => n4364);
   U8568 : OR2_X1 port map( A1 => n26679, A2 => n27821, ZN => n3561);
   U8569 : OR2_X1 port map( A1 => n14451, A2 => n13753, ZN => n2970);
   U8570 : AND2_X1 port map( A1 => n23599, A2 => n23467, ZN => n24257);
   U8571 : NOR2_X1 port map( A1 => n24257, A2 => n5548, ZN => n2806);
   U8572 : INV_X1 port map( A => n15290, ZN => n15294);
   U8573 : INV_X1 port map( A => n6080, ZN => n6449);
   U8574 : AND2_X1 port map( A1 => n3227, A2 => n21626, ZN => n5338);
   U8576 : OR2_X1 port map( A1 => n15027, A2 => n15431, ZN => n15029);
   U8577 : INV_X1 port map( A => n18646, ZN => n19668);
   U8579 : OR2_X1 port map( A1 => n7786, A2 => n7787, ZN => n7167);
   U8580 : INV_X1 port map( A => n18231, ZN => n18400);
   U8581 : AND2_X1 port map( A1 => n21625, A2 => n22141, ZN => n2911);
   U8582 : OAI22_X1 port map( A1 => n3992, A2 => n10031, B1 => n10718, B2 => 
                           n11137, ZN => n3991);
   U8583 : XNOR2_X1 port map( A => n25836, B => n25903, ZN => n25207);
   U8584 : XNOR2_X1 port map( A => n25207, B => n26038, ZN => n25502);
   U8585 : OR2_X1 port map( A1 => n15101, A2 => n15103, ZN => n2576);
   U8586 : INV_X1 port map( A => n14893, ZN => n15107);
   U8588 : INV_X1 port map( A => n22992, ZN => n23643);
   U8589 : OAI21_X1 port map( B1 => n2020, B2 => n14344, A => n14341, ZN => 
                           n6234);
   U8590 : NAND3_X2 port map( A1 => n17329, A2 => n17330, A3 => n2720, ZN => 
                           n19136);
   U8591 : NAND2_X1 port map( A1 => n2475, A2 => n2474, ZN => n27639);
   U8592 : OR2_X1 port map( A1 => n26357, A2 => n28651, ZN => n2474);
   U8593 : NAND3_X1 port map( A1 => n25043, A2 => n26270, A3 => n25042, ZN => 
                           n2475);
   U8594 : INV_X1 port map( A => n29565, ZN => n14486);
   U8595 : INV_X1 port map( A => n17570, ZN => n17573);
   U8596 : XNOR2_X1 port map( A => n429, B => n13414, ZN => n12087);
   U8599 : AOI22_X1 port map( A1 => n28422, A2 => n27537, B1 => n28468, B2 => 
                           n27547, ZN => n27543);
   U8600 : NOR2_X1 port map( A1 => n24420, A2 => n24517, ZN => n24513);
   U8601 : XNOR2_X1 port map( A => n19634, B => n19599, ZN => n6487);
   U8602 : NAND3_X1 port map( A1 => n4332, A2 => n17560, A3 => n2061, ZN => 
                           n5428);
   U8607 : NAND2_X1 port map( A1 => n4774, A2 => n17980, ZN => n17981);
   U8611 : NAND2_X1 port map( A1 => n7421, A2 => n7420, ZN => n2480);
   U8612 : NAND2_X1 port map( A1 => n2482, A2 => n2481, ZN => n23745);
   U8614 : NAND2_X1 port map( A1 => n23737, A2 => n23228, ZN => n2482);
   U8615 : OAI21_X1 port map( B1 => n13410, B2 => n2874, A => n2873, ZN => 
                           n13411);
   U8618 : NAND2_X1 port map( A1 => n20458, A2 => n4569, ZN => n20600);
   U8620 : OAI211_X1 port map( C1 => n14498, C2 => n14493, A => n2488, B => 
                           n13672, ZN => n12804);
   U8621 : NAND2_X1 port map( A1 => n2489, A2 => n17089, ZN => n18695);
   U8622 : OAI21_X1 port map( B1 => n17082, B2 => n18596, A => n5476, ZN => 
                           n2489);
   U8623 : XNOR2_X1 port map( A => n19101, B => n2490, ZN => n19006);
   U8624 : XNOR2_X1 port map( A => n19004, B => n19003, ZN => n2490);
   U8625 : AOI21_X1 port map( B1 => n7407, B2 => n7408, A => n7480, ZN => n2491
                           );
   U8627 : NAND2_X1 port map( A1 => n5693, A2 => n14178, ZN => n2493);
   U8629 : NOR2_X1 port map( A1 => n14006, A2 => n14386, ZN => n13573);
   U8630 : NAND2_X1 port map( A1 => n13572, A2 => n14380, ZN => n14006);
   U8633 : XNOR2_X1 port map( A => n15966, B => n15989, ZN => n15042);
   U8634 : OAI211_X1 port map( C1 => n23636, C2 => n23557, A => n2494, B => 
                           n23556, ZN => n23561);
   U8635 : NOR2_X1 port map( A1 => n23555, A2 => n23554, ZN => n2494);
   U8636 : NAND2_X1 port map( A1 => n184, A2 => n15094, ZN => n2496);
   U8638 : NAND2_X1 port map( A1 => n2500, A2 => n2499, ZN => n2498);
   U8639 : OR2_X1 port map( A1 => n5837, A2 => n11955, ZN => n12258);
   U8641 : NAND2_X1 port map( A1 => n7619, A2 => n8232, ZN => n7620);
   U8644 : NAND2_X1 port map( A1 => n2504, A2 => n2503, ZN => n11900);
   U8645 : NAND2_X1 port map( A1 => n11898, A2 => n29461, ZN => n2503);
   U8646 : NAND2_X1 port map( A1 => n11897, A2 => n11896, ZN => n2504);
   U8650 : OR2_X1 port map( A1 => n18215, A2 => n5155, ZN => n5154);
   U8651 : INV_X1 port map( A => n7554, ZN => n8133);
   U8652 : INV_X1 port map( A => n10937, ZN => n10999);
   U8653 : XNOR2_X1 port map( A => n5412, B => n10392, ZN => n5411);
   U8654 : AND3_X2 port map( A1 => n2071, A2 => n2564, A3 => n2565, ZN => n9062
                           );
   U8655 : OR2_X1 port map( A1 => n7079, A2 => n7092, ZN => n2507);
   U8656 : XNOR2_X1 port map( A => n15536, B => n16201, ZN => n15540);
   U8659 : NAND2_X1 port map( A1 => n23529, A2 => n23531, ZN => n23135);
   U8660 : NAND2_X1 port map( A1 => n18235, A2 => n17977, ZN => n2508);
   U8662 : NAND2_X1 port map( A1 => n7634, A2 => n7828, ZN => n7832);
   U8664 : XNOR2_X1 port map( A => n15761, B => n4767, ZN => n4766);
   U8666 : NAND2_X1 port map( A1 => n16946, A2 => n16945, ZN => n6176);
   U8667 : OR2_X1 port map( A1 => n11449, A2 => n11747, ZN => n11450);
   U8670 : NOR2_X1 port map( A1 => n18053, A2 => n18054, ZN => n18055);
   U8671 : NAND2_X1 port map( A1 => n4680, A2 => n16667, ZN => n16685);
   U8672 : BUF_X1 port map( A => n16764, Z => n17002);
   U8673 : NAND2_X1 port map( A1 => n7194, A2 => n7985, ZN => n2514);
   U8674 : NAND2_X1 port map( A1 => n7193, A2 => n7644, ZN => n2516);
   U8676 : NAND3_X1 port map( A1 => n20710, A2 => n20816, A3 => n21268, ZN => 
                           n6426);
   U8677 : NAND2_X1 port map( A1 => n11492, A2 => n4404, ZN => n11497);
   U8680 : NOR2_X1 port map( A1 => n11086, A2 => n28624, ZN => n2518);
   U8681 : INV_X1 port map( A => n19891, ZN => n3421);
   U8682 : NAND2_X1 port map( A1 => n8133, A2 => n8047, ZN => n7718);
   U8683 : NAND2_X1 port map( A1 => n2519, A2 => n20718, ZN => n22759);
   U8684 : NAND2_X1 port map( A1 => n5206, A2 => n5205, ZN => n2519);
   U8685 : NAND2_X1 port map( A1 => n20514, A2 => n20513, ZN => n19241);
   U8686 : NAND2_X1 port map( A1 => n20343, A2 => n20342, ZN => n20514);
   U8687 : NAND2_X1 port map( A1 => n2521, A2 => n2520, ZN => n11632);
   U8688 : NAND2_X1 port map( A1 => n10757, A2 => n11345, ZN => n2520);
   U8689 : NAND2_X1 port map( A1 => n1926, A2 => n15320, ZN => n3627);
   U8690 : INV_X1 port map( A => n27248, ZN => n5335);
   U8691 : OAI211_X2 port map( C1 => n27167, C2 => n26369, A => n2525, B => 
                           n2524, ZN => n27625);
   U8692 : NAND2_X1 port map( A1 => n27171, A2 => n27169, ZN => n2524);
   U8693 : NAND2_X1 port map( A1 => n26368, A2 => n29487, ZN => n2525);
   U8694 : INV_X1 port map( A => n13260, ZN => n13485);
   U8695 : OR2_X1 port map( A1 => n26819, A2 => n6568, ZN => n4926);
   U8696 : NOR2_X1 port map( A1 => n26447, A2 => n26449, ZN => n4832);
   U8698 : OAI22_X1 port map( A1 => n2526, A2 => n24220, B1 => n24219, B2 => 
                           n23956, ZN => n24221);
   U8699 : NAND2_X1 port map( A1 => n28509, A2 => n24760, ZN => n2526);
   U8700 : NOR2_X1 port map( A1 => n7708, A2 => n7382, ZN => n2897);
   U8701 : XNOR2_X1 port map( A => n6569, B => n19387, ZN => n20248);
   U8702 : AOI21_X1 port map( B1 => n3504, B2 => n3503, A => n20636, ZN => 
                           n2529);
   U8703 : NAND2_X1 port map( A1 => n15119, A2 => n14743, ZN => n13660);
   U8704 : NAND2_X1 port map( A1 => n4179, A2 => n7497, ZN => n7499);
   U8705 : NAND2_X1 port map( A1 => n2718, A2 => n18405, ZN => n5022);
   U8706 : NAND4_X2 port map( A1 => n24763, A2 => n24762, A3 => n2531, A4 => 
                           n2530, ZN => n25810);
   U8707 : NAND2_X1 port map( A1 => n2866, A2 => n378, ZN => n2530);
   U8708 : NAND2_X1 port map( A1 => n2865, A2 => n23588, ZN => n2531);
   U8709 : XNOR2_X1 port map( A => n22388, B => n22523, ZN => n2532);
   U8711 : OAI211_X1 port map( C1 => n27199, C2 => n27198, A => n3899, B => 
                           n2618, ZN => n3898);
   U8712 : NAND2_X1 port map( A1 => n18009, A2 => n2533, ZN => n18762);
   U8713 : OR2_X1 port map( A1 => n18010, A2 => n6079, ZN => n2533);
   U8715 : XNOR2_X2 port map( A => n13529, B => n13528, ZN => n14007);
   U8718 : OAI22_X1 port map( A1 => n19752, A2 => n20083, B1 => n5126, B2 => 
                           n18837, ZN => n2534);
   U8721 : NAND2_X1 port map( A1 => n12180, A2 => n12181, ZN => n11411);
   U8722 : NAND2_X1 port map( A1 => n24416, A2 => n24709, ZN => n6513);
   U8723 : OAI21_X1 port map( B1 => n24707, B2 => n24417, A => n5795, ZN => 
                           n24416);
   U8724 : NAND3_X1 port map( A1 => n27825, A2 => n27101, A3 => n26901, ZN => 
                           n26875);
   U8725 : XNOR2_X1 port map( A => n10328, B => n10184, ZN => n10185);
   U8727 : AOI21_X1 port map( B1 => n8180, B2 => n8181, A => n4856, ZN => n8182
                           );
   U8728 : OAI21_X2 port map( B1 => n7647, B2 => n7648, A => n7646, ZN => n9211
                           );
   U8729 : NAND2_X1 port map( A1 => n11584, A2 => n567, ZN => n11587);
   U8730 : NAND2_X1 port map( A1 => n8028, A2 => n8032, ZN => n7736);
   U8734 : OAI211_X1 port map( C1 => n10499, C2 => n1834, A => n10715, B => 
                           n2539, ZN => n10455);
   U8735 : NAND2_X1 port map( A1 => n5672, A2 => n10498, ZN => n2539);
   U8736 : INV_X1 port map( A => n10022, ZN => n3452);
   U8737 : AOI21_X1 port map( B1 => n11456, B2 => n11455, A => n2542, ZN => 
                           n13017);
   U8738 : OAI21_X1 port map( B1 => n8829, B2 => n8826, A => n8462, ZN => n3706
                           );
   U8739 : NAND2_X1 port map( A1 => n8192, A2 => n4675, ZN => n8462);
   U8745 : XNOR2_X1 port map( A => n18166, B => n18167, ZN => n19820);
   U8746 : OR2_X1 port map( A1 => n13639, A2 => n14944, ZN => n13586);
   U8747 : XNOR2_X1 port map( A => n3403, B => n18913, ZN => n19604);
   U8748 : NOR2_X1 port map( A1 => n18214, A2 => n4824, ZN => n18218);
   U8750 : OAI21_X1 port map( B1 => n2546, B2 => n8147, A => n2545, ZN => n7151
                           );
   U8751 : OR2_X1 port map( A1 => n17439, A2 => n336, ZN => n16926);
   U8752 : NAND3_X2 port map( A1 => n3140, A2 => n8184, A3 => n3139, ZN => 
                           n10321);
   U8753 : XNOR2_X2 port map( A => n8318, B => n8319, ZN => n11168);
   U8754 : NAND2_X1 port map( A1 => n7928, A2 => n7927, ZN => n2547);
   U8755 : OAI21_X1 port map( B1 => n14064, B2 => n14065, A => n3393, ZN => 
                           n13164);
   U8756 : XOR2_X1 port map( A => n16444, B => n16519, Z => n5858);
   U8757 : AOI21_X2 port map( B1 => n18419, B2 => n18418, A => n18417, ZN => 
                           n19206);
   U8759 : XNOR2_X1 port map( A => n2551, B => n21766, ZN => n21768);
   U8760 : XNOR2_X1 port map( A => n21765, B => n22757, ZN => n2551);
   U8761 : NAND2_X1 port map( A1 => n27021, A2 => n27018, ZN => n2552);
   U8763 : NAND3_X1 port map( A1 => n29718, A2 => n17202, A3 => n17203, ZN => 
                           n6335);
   U8764 : XOR2_X1 port map( A => n25188, B => n28496, Z => n6789);
   U8766 : NAND2_X1 port map( A1 => n2839, A2 => n2840, ZN => n6718);
   U8767 : INV_X1 port map( A => n14419, ZN => n14420);
   U8768 : NAND3_X1 port map( A1 => n13924, A2 => n14775, A3 => n13923, ZN => 
                           n5893);
   U8769 : INV_X1 port map( A => n11330, ZN => n8422);
   U8770 : XNOR2_X1 port map( A => n10145, B => n2403, ZN => n9935);
   U8774 : NAND3_X1 port map( A1 => n23144, A2 => n24630, A3 => n24629, ZN => 
                           n4365);
   U8776 : NAND3_X1 port map( A1 => n8218, A2 => n7624, A3 => n7625, ZN => 
                           n2556);
   U8777 : INV_X1 port map( A => n28195, ZN => n5025);
   U8779 : NAND2_X1 port map( A1 => n7896, A2 => n7897, ZN => n7899);
   U8780 : INV_X1 port map( A => Plaintext(47), ZN => n2638);
   U8781 : OR3_X2 port map( A1 => n21701, A2 => n21700, A3 => n21699, ZN => 
                           n21872);
   U8782 : OAI21_X1 port map( B1 => n499, B2 => n20180, A => n20217, ZN => 
                           n3078);
   U8783 : XNOR2_X2 port map( A => n21840, B => n21839, ZN => n23772);
   U8785 : NAND2_X1 port map( A1 => n4849, A2 => n2557, ZN => n24769);
   U8786 : NOR2_X1 port map( A1 => n4847, A2 => n4848, ZN => n2557);
   U8787 : NAND2_X1 port map( A1 => n3429, A2 => n3430, ZN => n3428);
   U8788 : NAND2_X1 port map( A1 => n18020, A2 => n18018, ZN => n2558);
   U8789 : NAND3_X1 port map( A1 => n18603, A2 => n6714, A3 => n6713, ZN => 
                           n18812);
   U8790 : NOR2_X1 port map( A1 => n17475, A2 => n17478, ZN => n2559);
   U8791 : INV_X1 port map( A => n17480, ZN => n2560);
   U8792 : AND2_X1 port map( A1 => n10810, A2 => n10473, ZN => n11324);
   U8794 : NAND2_X1 port map( A1 => n13839, A2 => n13838, ZN => n2562);
   U8795 : INV_X1 port map( A => n11795, ZN => n3558);
   U8796 : NAND2_X1 port map( A1 => n3124, A2 => n24793, ZN => n3714);
   U8797 : INV_X1 port map( A => n18330, ZN => n6403);
   U8798 : NAND2_X1 port map( A1 => n2563, A2 => n2663, ZN => n10728);
   U8799 : NAND2_X1 port map( A1 => n2661, A2 => n10927, ZN => n2563);
   U8800 : NAND2_X1 port map( A1 => n7531, A2 => n7141, ZN => n2564);
   U8801 : NAND2_X1 port map( A1 => n7532, A2 => n7523, ZN => n2565);
   U8802 : OAI211_X1 port map( C1 => n18591, C2 => n17837, A => n17836, B => 
                           n2044, ZN => n2566);
   U8803 : INV_X1 port map( A => n20437, ZN => n20611);
   U8805 : INV_X1 port map( A => n5945, ZN => n6590);
   U8807 : XNOR2_X1 port map( A => n2567, B => n15641, ZN => n17030);
   U8808 : XNOR2_X1 port map( A => n15645, B => n15640, ZN => n2567);
   U8809 : NOR2_X1 port map( A1 => n5164, A2 => n17888, ZN => n5162);
   U8810 : NAND2_X1 port map( A1 => n14084, A2 => n14286, ZN => n13770);
   U8811 : XNOR2_X2 port map( A => n16225, B => n16226, ZN => n17138);
   U8812 : NAND3_X1 port map( A1 => n21496, A2 => n28789, A3 => n21495, ZN => 
                           n6749);
   U8813 : NAND2_X1 port map( A1 => n11549, A2 => n11851, ZN => n11548);
   U8814 : NAND3_X1 port map( A1 => n7917, A2 => n7915, A3 => n7916, ZN => 
                           n2569);
   U8815 : NOR2_X2 port map( A1 => n3197, A2 => n18152, ZN => n19376);
   U8816 : OAI211_X1 port map( C1 => n18016, C2 => n18493, A => n1997, B => 
                           n3768, ZN => n2571);
   U8817 : AOI21_X1 port map( B1 => n21478, B2 => n1930, A => n2572, ZN => 
                           n21391);
   U8818 : OR2_X1 port map( A1 => n15248, A2 => n15137, ZN => n14116);
   U8819 : NAND2_X1 port map( A1 => n2573, A2 => n14970, ZN => n14977);
   U8820 : NAND2_X1 port map( A1 => n5813, A2 => n14969, ZN => n2573);
   U8823 : XNOR2_X1 port map( A => n2574, B => n13522, ZN => n12683);
   U8824 : XNOR2_X1 port map( A => n12680, B => n13171, ZN => n2574);
   U8825 : NAND2_X1 port map( A1 => n6022, A2 => n6286, ZN => n15583);
   U8827 : NAND3_X1 port map( A1 => n2575, A2 => n23363, A3 => n3902, ZN => 
                           n3901);
   U8828 : NAND2_X1 port map( A1 => n16728, A2 => n17484, ZN => n2578);
   U8829 : NAND2_X1 port map( A1 => n17830, A2 => n17829, ZN => n2579);
   U8830 : OR2_X1 port map( A1 => n9220, A2 => n9221, ZN => n9024);
   U8831 : OAI21_X1 port map( B1 => n14843, B2 => n14844, A => n15284, ZN => 
                           n14848);
   U8832 : INV_X1 port map( A => n20551, ZN => n6086);
   U8834 : NAND2_X1 port map( A1 => n2581, A2 => n11816, ZN => n11433);
   U8835 : OAI21_X1 port map( B1 => n11724, B2 => n11819, A => n11818, ZN => 
                           n2581);
   U8836 : NAND2_X1 port map( A1 => n2583, A2 => n2582, ZN => n13863);
   U8837 : NAND2_X1 port map( A1 => n13862, A2 => n14460, ZN => n2582);
   U8838 : NAND2_X1 port map( A1 => n2584, A2 => n3580, ZN => n2583);
   U8839 : NAND2_X1 port map( A1 => n14204, A2 => n14200, ZN => n2584);
   U8841 : NOR2_X1 port map( A1 => n14194, A2 => n29604, ZN => n4434);
   U8842 : NAND2_X1 port map( A1 => n2634, A2 => n526, ZN => n2633);
   U8843 : OAI21_X1 port map( B1 => n8532, B2 => n8709, A => n2585, ZN => n7035
                           );
   U8844 : NAND2_X1 port map( A1 => n8407, A2 => n8876, ZN => n2585);
   U8845 : NOR2_X1 port map( A1 => n8699, A2 => n8881, ZN => n8407);
   U8846 : XNOR2_X1 port map( A => n19167, B => n1989, ZN => n19168);
   U8847 : NAND3_X1 port map( A1 => n2586, A2 => n24593, A3 => n4692, ZN => 
                           n4691);
   U8848 : NAND2_X1 port map( A1 => n404, A2 => n24397, ZN => n24674);
   U8850 : NAND2_X1 port map( A1 => n2589, A2 => n29735, ZN => n2587);
   U8852 : NAND2_X1 port map( A1 => n7004, A2 => n2590, ZN => n7005);
   U8853 : NOR2_X1 port map( A1 => n2591, A2 => n17689, ZN => n5201);
   U8854 : NAND3_X2 port map( A1 => n2593, A2 => n2592, A3 => n2009, ZN => 
                           n16272);
   U8855 : NAND2_X1 port map( A1 => n14640, A2 => n15082, ZN => n2593);
   U8857 : NAND2_X1 port map( A1 => n20006, A2 => n20258, ZN => n2594);
   U8859 : XNOR2_X1 port map( A => n9601, B => n10228, ZN => n10285);
   U8860 : NAND2_X1 port map( A1 => n8597, A2 => n8819, ZN => n2596);
   U8861 : INV_X1 port map( A => n8596, ZN => n2597);
   U8863 : NAND2_X1 port map( A1 => n2599, A2 => n16799, ZN => n3017);
   U8864 : NAND3_X1 port map( A1 => n3672, A2 => n17129, A3 => n2600, ZN => 
                           n2599);
   U8865 : INV_X1 port map( A => n17990, ZN => n18598);
   U8866 : NAND2_X1 port map( A1 => n2601, A2 => n6152, ZN => n6151);
   U8867 : NAND2_X1 port map( A1 => n11133, A2 => n10457, ZN => n2601);
   U8868 : OR2_X2 port map( A1 => n6044, A2 => n13835, ZN => n15180);
   U8869 : NAND2_X1 port map( A1 => n8303, A2 => n8296, ZN => n8299);
   U8870 : NAND2_X1 port map( A1 => n17834, A2 => n18595, ZN => n18130);
   U8871 : MUX2_X1 port map( A => n2610, B => n17110, S => n17106, Z => n2609);
   U8872 : AOI21_X1 port map( B1 => n10401, B2 => n8763, A => n2104, ZN => 
                           n8646);
   U8873 : NAND2_X1 port map( A1 => n2611, A2 => n22742, ZN => n2613);
   U8874 : NAND2_X1 port map( A1 => n3043, A2 => n23286, ZN => n2611);
   U8875 : MUX2_X1 port map( A => n24405, B => n24404, S => n24403, Z => n23506
                           );
   U8876 : AND3_X2 port map( A1 => n2613, A2 => n3042, A3 => n2612, ZN => 
                           n24403);
   U8877 : OAI22_X1 port map( A1 => n11131, A2 => n2646, B1 => n4555, B2 => 
                           n2614, ZN => n2655);
   U8878 : NAND2_X1 port map( A1 => n10713, A2 => n10502, ZN => n2614);
   U8879 : NAND2_X1 port map( A1 => n27130, A2 => n29293, ZN => n2615);
   U8880 : NOR2_X1 port map( A1 => n27548, A2 => n27202, ZN => n27545);
   U8881 : NAND2_X1 port map( A1 => n2617, A2 => n28422, ZN => n2618);
   U8882 : INV_X1 port map( A => n24437, ZN => n23886);
   U8883 : INV_X1 port map( A => n24347, ZN => n2619);
   U8884 : INV_X1 port map( A => n2621, ZN => n2620);
   U8886 : OAI21_X1 port map( B1 => n22994, B2 => n22995, A => n22993, ZN => 
                           n2623);
   U8887 : NAND2_X1 port map( A1 => n2624, A2 => n7766, ZN => n2629);
   U8888 : NAND2_X1 port map( A1 => n2630, A2 => n2631, ZN => n2625);
   U8889 : NAND2_X1 port map( A1 => n8177, A2 => n2630, ZN => n2626);
   U8890 : NAND3_X1 port map( A1 => n2628, A2 => n2627, A3 => n2629, ZN => 
                           n8335);
   U8891 : NAND2_X1 port map( A1 => n2630, A2 => n2631, ZN => n2627);
   U8892 : NAND2_X1 port map( A1 => n8177, A2 => n2630, ZN => n2628);
   U8893 : NAND2_X1 port map( A1 => n8179, A2 => n8176, ZN => n7766);
   U8895 : INV_X1 port map( A => n7289, ZN => n2631);
   U8896 : NAND2_X1 port map( A1 => n2632, A2 => n2122, ZN => n5399);
   U8897 : NOR2_X1 port map( A1 => n2632, A2 => n29483, ZN => n15688);
   U8898 : NAND3_X1 port map( A1 => n14376, A2 => n29059, A3 => n2849, ZN => 
                           n6613);
   U8899 : NOR2_X1 port map( A1 => n17847, A2 => n17846, ZN => n2634);
   U8900 : NAND3_X1 port map( A1 => n23024, A2 => n23539, A3 => n2637, ZN => 
                           n6764);
   U8901 : NAND2_X1 port map( A1 => n23687, A2 => n23801, ZN => n2637);
   U8902 : NAND2_X1 port map( A1 => n2637, A2 => n4337, ZN => n4336);
   U8903 : AND2_X1 port map( A1 => n21894, A2 => n2636, ZN => n21895);
   U8904 : NAND2_X1 port map( A1 => n7129, A2 => n29119, ZN => n3148);
   U8908 : NAND3_X1 port map( A1 => n14851, A2 => n2644, A3 => n2643, ZN => 
                           n2642);
   U8909 : NAND2_X1 port map( A1 => n15312, A2 => n15310, ZN => n2643);
   U8910 : NAND3_X2 port map( A1 => n5949, A2 => n6794, A3 => n14316, ZN => 
                           n15310);
   U8911 : NAND2_X1 port map( A1 => n15309, A2 => n15306, ZN => n2644);
   U8912 : NAND2_X1 port map( A1 => n14854, A2 => n14852, ZN => n2645);
   U8913 : XNOR2_X2 port map( A => n9975, B => n9974, ZN => n10713);
   U8914 : NAND2_X1 port map( A1 => n2648, A2 => n2647, ZN => n24314);
   U8915 : NAND2_X1 port map( A1 => n2649, A2 => n24391, ZN => n2647);
   U8917 : NAND3_X1 port map( A1 => n490, A2 => n21410, A3 => n20663, ZN => 
                           n2650);
   U8918 : NAND2_X1 port map( A1 => n21047, A2 => n2652, ZN => n2651);
   U8919 : NOR2_X1 port map( A1 => n21410, A2 => n21171, ZN => n2652);
   U8923 : INV_X1 port map( A => n17889, ZN => n2656);
   U8924 : NAND2_X1 port map( A1 => n2659, A2 => n2657, ZN => n7114);
   U8925 : OAI21_X1 port map( B1 => n2658, B2 => n2631, A => n8179, ZN => n2657
                           );
   U8926 : INV_X1 port map( A => n7290, ZN => n2658);
   U8929 : NAND2_X1 port map( A1 => n7289, A2 => n8173, ZN => n7347);
   U8930 : NAND2_X1 port map( A1 => n10930, A2 => n10932, ZN => n2661);
   U8931 : NAND2_X1 port map( A1 => n10727, A2 => n10929, ZN => n2663);
   U8933 : NAND2_X1 port map( A1 => n2741, A2 => n2664, ZN => n16938);
   U8935 : AND2_X1 port map( A1 => n21665, A2 => n3666, ZN => n2669);
   U8936 : NAND3_X1 port map( A1 => n9142, A2 => n8564, A3 => n599, ZN => n8565
                           );
   U8937 : NAND2_X1 port map( A1 => n2670, A2 => n7331, ZN => n7335);
   U8942 : AND2_X1 port map( A1 => n13827, A2 => n14278, ZN => n4369);
   U8943 : OAI21_X1 port map( B1 => n28507, B2 => n4166, A => n29691, ZN => 
                           n13618);
   U8945 : XNOR2_X2 port map( A => n2675, B => Key(23), ZN => n7330);
   U8946 : INV_X1 port map( A => Plaintext(23), ZN => n2675);
   U8947 : XNOR2_X1 port map( A => n2677, B => n27952, ZN => n7415);
   U8948 : XNOR2_X1 port map( A => n2677, B => n3114, ZN => n9740);
   U8949 : XNOR2_X1 port map( A => n9639, B => n2677, ZN => n9403);
   U8950 : XNOR2_X1 port map( A => n9702, B => n2677, ZN => n10368);
   U8951 : INV_X1 port map( A => n11310, ZN => n2680);
   U8952 : NAND2_X1 port map( A1 => n11163, A2 => n29637, ZN => n11310);
   U8953 : NOR2_X1 port map( A1 => n2681, A2 => n14260, ZN => n2945);
   U8954 : NAND2_X1 port map( A1 => n13614, A2 => n2681, ZN => n12369);
   U8957 : NAND2_X1 port map( A1 => n28203, A2 => n12109, ZN => n2684);
   U8958 : NAND2_X1 port map( A1 => n9655, A2 => n12109, ZN => n2685);
   U8960 : AND2_X1 port map( A1 => n11258, A2 => n2690, ZN => n4326);
   U8961 : NAND2_X1 port map( A1 => n2689, A2 => n2687, ZN => n11023);
   U8962 : AND2_X1 port map( A1 => n2690, A2 => n11318, ZN => n2687);
   U8963 : MUX2_X1 port map( A => n2690, B => n11254, S => n594, Z => n9503);
   U8964 : NAND2_X1 port map( A1 => n14929, A2 => n2691, ZN => n15781);
   U8965 : NAND2_X1 port map( A1 => n7163, A2 => n7164, ZN => n7771);
   U8966 : AOI21_X1 port map( B1 => n2694, B2 => n17719, A => n18081, ZN => 
                           n6229);
   U8967 : OAI22_X1 port map( A1 => n2694, A2 => n18285, B1 => n373, B2 => 
                           n17719, ZN => n3753);
   U8968 : OAI21_X1 port map( B1 => n18525, B2 => n18523, A => n2694, ZN => 
                           n18287);
   U8970 : NAND2_X1 port map( A1 => n2696, A2 => n7985, ZN => n2695);
   U8971 : NAND2_X1 port map( A1 => n7983, A2 => n7984, ZN => n2696);
   U8973 : NAND2_X1 port map( A1 => n23656, A2 => n4232, ZN => n2697);
   U8974 : NOR2_X1 port map( A1 => n11666, A2 => n3946, ZN => n11667);
   U8975 : XNOR2_X1 port map( A => n2700, B => n2996, ZN => n14675);
   U8976 : XNOR2_X1 port map( A => n2700, B => n1046, ZN => n16034);
   U8977 : XNOR2_X1 port map( A => n2700, B => n3323, ZN => n16511);
   U8978 : XNOR2_X1 port map( A => n16470, B => n2700, ZN => n16375);
   U8979 : NAND2_X1 port map( A1 => n535, A2 => n17368, ZN => n17233);
   U8980 : NAND2_X1 port map( A1 => n2701, A2 => n17046, ZN => n15732);
   U8981 : NAND2_X1 port map( A1 => n535, A2 => n17234, ZN => n17235);
   U8982 : NAND2_X1 port map( A1 => n17043, A2 => n535, ZN => n3549);
   U8985 : NOR2_X1 port map( A1 => n18530, A2 => n29476, ZN => n2702);
   U8988 : NAND2_X1 port map( A1 => n509, A2 => n18529, ZN => n18259);
   U8989 : NAND2_X1 port map( A1 => n22084, A2 => n2708, ZN => n6220);
   U8990 : AOI21_X1 port map( B1 => n28431, B2 => n2708, A => n28622, ZN => 
                           n22085);
   U8991 : INV_X1 port map( A => n23706, ZN => n2708);
   U8992 : XNOR2_X1 port map( A => n10344, B => n3067, ZN => n2711);
   U8993 : XNOR2_X1 port map( A => n2711, B => n9698, ZN => n9301);
   U8994 : INV_X1 port map( A => n8506, ZN => n2713);
   U8995 : NAND2_X1 port map( A1 => n563, A2 => n2714, ZN => n13767);
   U8996 : NAND2_X1 port map( A1 => n2715, A2 => n20155, ZN => n4410);
   U8997 : OAI22_X1 port map( A1 => n2815, A2 => n2715, B1 => n20100, B2 => 
                           n20101, ZN => n20533);
   U8998 : NAND2_X1 port map( A1 => n2717, A2 => n614, ZN => n7165);
   U8999 : NAND2_X1 port map( A1 => n7321, A2 => n7770, ZN => n2717);
   U9000 : AND2_X1 port map( A1 => n2718, A2 => n4756, ZN => n6264);
   U9001 : NAND2_X1 port map( A1 => n5021, A2 => n5023, ZN => n2718);
   U9002 : NOR2_X1 port map( A1 => n5439, A2 => n18230, ZN => n19024);
   U9003 : OAI211_X1 port map( C1 => n5439, C2 => n2723, A => n2722, B => n2721
                           , ZN => n18767);
   U9004 : NAND2_X1 port map( A1 => n18230, A2 => n1887, ZN => n2721);
   U9005 : NAND2_X1 port map( A1 => n5439, A2 => n1887, ZN => n2722);
   U9008 : INV_X1 port map( A => n14744, ZN => n2727);
   U9009 : NAND2_X1 port map( A1 => n29604, A2 => n14393, ZN => n4436);
   U9010 : NAND2_X1 port map( A1 => n2728, A2 => n14194, ZN => n14394);
   U9011 : NAND2_X1 port map( A1 => n14395, A2 => n29604, ZN => n4047);
   U9012 : NAND2_X1 port map( A1 => n13951, A2 => n29604, ZN => n13870);
   U9013 : OAI22_X1 port map( A1 => n5745, A2 => n14393, B1 => n28805, B2 => 
                           n29604, ZN => n6283);
   U9014 : NAND4_X1 port map( A1 => n14597, A2 => n6921, A3 => n2729, A4 => 
                           n14258, ZN => n2730);
   U9016 : NAND2_X1 port map( A1 => n15105, A2 => n15423, ZN => n14934);
   U9017 : NAND2_X1 port map( A1 => n2002, A2 => n15105, ZN => n2732);
   U9018 : NAND2_X1 port map( A1 => n15423, A2 => n549, ZN => n2733);
   U9019 : NAND2_X1 port map( A1 => n29104, A2 => n2735, ZN => n6409);
   U9020 : OAI21_X1 port map( B1 => n20093, B2 => n20041, A => n2734, ZN => 
                           n18789);
   U9021 : NAND2_X1 port map( A1 => n20041, A2 => n20088, ZN => n2734);
   U9022 : OAI22_X1 port map( A1 => n20087, A2 => n19757, B1 => n20092, B2 => 
                           n2735, ZN => n19758);
   U9023 : NAND2_X1 port map( A1 => n24705, A2 => n2736, ZN => n24710);
   U9024 : NAND2_X1 port map( A1 => n24709, A2 => n29043, ZN => n2736);
   U9025 : NAND2_X1 port map( A1 => n2737, A2 => n14761, ZN => n15264);
   U9026 : NAND3_X2 port map( A1 => n14245, A2 => n14247, A3 => n14246, ZN => 
                           n14761);
   U9027 : INV_X1 port map( A => n14762, ZN => n2737);
   U9028 : NAND2_X1 port map( A1 => n4162, A2 => n15260, ZN => n4097);
   U9029 : NAND2_X1 port map( A1 => n8504, A2 => n8886, ZN => n2739);
   U9031 : NAND3_X1 port map( A1 => n8504, A2 => n8336, A3 => n8889, ZN => 
                           n2740);
   U9033 : NAND2_X1 port map( A1 => n17335, A2 => n28564, ZN => n17203);
   U9034 : NAND3_X1 port map( A1 => n15180, A2 => n28803, A3 => n14534, ZN => 
                           n2744);
   U9036 : OR2_X1 port map( A1 => n3954, A2 => n1908, ZN => n2746);
   U9037 : NAND3_X1 port map( A1 => n20455, A2 => n20454, A3 => n20632, ZN => 
                           n20456);
   U9038 : NAND2_X1 port map( A1 => n20033, A2 => n20634, ZN => n20455);
   U9040 : NAND2_X1 port map( A1 => n5172, A2 => n5171, ZN => n2749);
   U9041 : AND2_X1 port map( A1 => n23363, A2 => n23360, ZN => n21302);
   U9042 : OAI211_X2 port map( C1 => n486, C2 => n23069, A => n2751, B => n2750
                           , ZN => n24711);
   U9043 : NAND2_X1 port map( A1 => n23674, A2 => n23363, ZN => n2750);
   U9044 : NAND2_X1 port map( A1 => n23068, A2 => n486, ZN => n2751);
   U9045 : NAND3_X1 port map( A1 => n29122, A2 => n11047, A3 => n2753, ZN => 
                           n9653);
   U9046 : NAND3_X1 port map( A1 => n11260, A2 => n11266, A3 => n2753, ZN => 
                           n10669);
   U9047 : INV_X1 port map( A => n11267, ZN => n2753);
   U9050 : NAND2_X1 port map( A1 => n11260, A2 => n11045, ZN => n2755);
   U9051 : NAND3_X1 port map( A1 => n1954, A2 => n2757, A3 => n2756, ZN => 
                           n17770);
   U9052 : NAND3_X1 port map( A1 => n17764, A2 => n3597, A3 => n28073, ZN => 
                           n2756);
   U9053 : NAND2_X1 port map( A1 => n2758, A2 => n1133, ZN => n2757);
   U9054 : XNOR2_X1 port map( A => n2759, B => n3321, ZN => n19341);
   U9055 : XNOR2_X1 port map( A => n2759, B => n3643, ZN => n19633);
   U9056 : XNOR2_X1 port map( A => n2759, B => n2986, ZN => n18662);
   U9057 : XNOR2_X1 port map( A => n19688, B => n2759, ZN => n18868);
   U9058 : XNOR2_X1 port map( A => n19111, B => n2759, ZN => n19112);
   U9059 : NAND2_X1 port map( A1 => n2761, A2 => n2760, ZN => n23909);
   U9060 : NAND3_X1 port map( A1 => n24405, A2 => n24083, A3 => n24403, ZN => 
                           n2760);
   U9061 : NAND3_X1 port map( A1 => n24408, A2 => n24404, A3 => n2762, ZN => 
                           n2761);
   U9062 : INV_X1 port map( A => n27846, ZN => n2765);
   U9063 : NAND3_X1 port map( A1 => n27843, A2 => n27826, A3 => n27825, ZN => 
                           n2763);
   U9064 : NAND2_X1 port map( A1 => n2767, A2 => n3542, ZN => n2764);
   U9066 : INV_X1 port map( A => n17567, ZN => n2769);
   U9067 : NAND2_X1 port map( A1 => n17759, A2 => n17758, ZN => n2770);
   U9068 : NAND2_X1 port map( A1 => n17969, A2 => n18236, ZN => n17756);
   U9069 : NAND2_X1 port map( A1 => n2773, A2 => n1354, ZN => n2772);
   U9070 : NAND2_X1 port map( A1 => n7888, A2 => n7777, ZN => n2773);
   U9071 : NAND2_X1 port map( A1 => n7778, A2 => n7315, ZN => n7888);
   U9072 : INV_X1 port map( A => n17818, ZN => n18413);
   U9073 : INV_X1 port map( A => n18120, ZN => n2777);
   U9074 : NOR2_X1 port map( A1 => n18414, A2 => n18410, ZN => n2778);
   U9075 : NOR2_X1 port map( A1 => n18411, A2 => n17818, ZN => n18120);
   U9077 : NAND2_X1 port map( A1 => n23651, A2 => n2779, ZN => n23194);
   U9078 : NAND2_X1 port map( A1 => n23046, A2 => n23654, ZN => n23652);
   U9079 : MUX2_X1 port map( A => n23649, B => n23650, S => n23470, Z => n23653
                           );
   U9080 : NAND2_X1 port map( A1 => n8019, A2 => n7747, ZN => n2780);
   U9081 : OAI22_X1 port map( A1 => n7746, A2 => n7745, B1 => n7743, B2 => 
                           n7744, ZN => n2781);
   U9082 : NAND2_X1 port map( A1 => n2783, A2 => n13703, ZN => n14424);
   U9083 : NAND2_X1 port map( A1 => n2783, A2 => n14426, ZN => n14305);
   U9084 : NAND2_X1 port map( A1 => n4522, A2 => n2783, ZN => n12532);
   U9086 : AND2_X1 port map( A1 => n2783, A2 => n29558, ZN => n2782);
   U9087 : INV_X1 port map( A => n12534, ZN => n2783);
   U9089 : MUX2_X1 port map( A => n23657, B => n23351, S => n29583, Z => n23143
                           );
   U9090 : INV_X1 port map( A => n19354, ZN => n19655);
   U9091 : NAND3_X1 port map( A1 => n2786, A2 => n17844, A3 => n18243, ZN => 
                           n2784);
   U9092 : NAND2_X1 port map( A1 => n2787, A2 => n17843, ZN => n2785);
   U9093 : INV_X1 port map( A => n7506, ZN => n6210);
   U9094 : XNOR2_X2 port map( A => Key(57), B => Plaintext(57), ZN => n7506);
   U9095 : NAND2_X1 port map( A1 => n7514, A2 => n7506, ZN => n2788);
   U9096 : XNOR2_X1 port map( A => n15853, B => n15852, ZN => n2790);
   U9097 : NAND2_X1 port map( A1 => n18062, A2 => n2791, ZN => n4348);
   U9099 : OAI22_X1 port map( A1 => n17929, A2 => n2791, B1 => n18061, B2 => 
                           n17928, ZN => n17930);
   U9100 : NAND2_X1 port map( A1 => n397, A2 => n27744, ZN => n2795);
   U9102 : NAND2_X1 port map( A1 => n2797, A2 => n5303, ZN => n2796);
   U9103 : NAND2_X1 port map( A1 => n15208, A2 => n14928, ZN => n15206);
   U9104 : INV_X1 port map( A => n15206, ZN => n2800);
   U9105 : OAI211_X1 port map( C1 => n2803, C2 => n18788, A => n2802, B => 
                           n2801, ZN => n22312);
   U9106 : NAND2_X1 port map( A1 => n18788, A2 => n2804, ZN => n2801);
   U9107 : NAND2_X1 port map( A1 => n18787, A2 => n2804, ZN => n2802);
   U9108 : INV_X1 port map( A => Key(15), ZN => n2804);
   U9109 : XNOR2_X1 port map( A => n2805, B => n22295, ZN => n21850);
   U9110 : XNOR2_X1 port map( A => n2805, B => n22073, ZN => n20680);
   U9111 : NOR2_X1 port map( A1 => n2806, A2 => n24976, ZN => n24512);
   U9112 : OAI21_X1 port map( B1 => n24975, B2 => n2806, A => n24259, ZN => 
                           n25059);
   U9113 : OAI211_X2 port map( C1 => n23804, C2 => n28919, A => n1976, B => 
                           n2807, ZN => n26054);
   U9114 : NAND2_X1 port map( A1 => n2808, A2 => n24653, ZN => n24028);
   U9115 : INV_X1 port map( A => n24651, ZN => n2808);
   U9116 : NAND2_X1 port map( A1 => n24029, A2 => n2809, ZN => n24031);
   U9117 : NOR2_X1 port map( A1 => n28481, A2 => n24523, ZN => n2809);
   U9118 : NOR2_X1 port map( A1 => n24651, A2 => n629, ZN => n2810);
   U9119 : INV_X1 port map( A => n17846, ZN => n2811);
   U9120 : XNOR2_X1 port map( A => n25343, B => n25340, ZN => n2813);
   U9121 : NAND3_X1 port map( A1 => n1888, A2 => n18020, A3 => n18251, ZN => 
                           n3069);
   U9122 : NAND2_X1 port map( A1 => n2814, A2 => n2834, ZN => n3084);
   U9123 : INV_X1 port map( A => n20156, ZN => n2815);
   U9124 : NAND2_X1 port map( A1 => n24513, A2 => n24421, ZN => n2816);
   U9126 : NAND2_X1 port map( A1 => n23748, A2 => n23749, ZN => n2817);
   U9127 : XNOR2_X2 port map( A => n15931, B => n15930, ZN => n17570);
   U9128 : AOI21_X2 port map( B1 => n2821, B2 => n6868, A => n2820, ZN => 
                           n25903);
   U9129 : NOR2_X1 port map( A1 => n23126, A2 => n24020, ZN => n24160);
   U9130 : INV_X1 port map( A => n24538, ZN => n2823);
   U9131 : NAND2_X1 port map( A1 => n24159, A2 => n24542, ZN => n2824);
   U9132 : NAND2_X1 port map( A1 => n23126, A2 => n24001, ZN => n24159);
   U9133 : INV_X1 port map( A => n17424, ZN => n2826);
   U9134 : INV_X1 port map( A => n17424, ZN => n2825);
   U9135 : NAND2_X1 port map( A1 => n2825, A2 => n17425, ZN => n17008);
   U9137 : NAND2_X1 port map( A1 => n24450, A2 => n24757, ZN => n2828);
   U9138 : NAND3_X1 port map( A1 => n24761, A2 => n28509, A3 => n24758, ZN => 
                           n2829);
   U9139 : OAI211_X2 port map( C1 => n21522, C2 => n21550, A => n21521, B => 
                           n2830, ZN => n22567);
   U9140 : AND2_X1 port map( A1 => n17393, A2 => n17293, ZN => n16958);
   U9141 : NAND2_X1 port map( A1 => n5487, A2 => n533, ZN => n17000);
   U9142 : NAND2_X1 port map( A1 => n16961, A2 => n533, ZN => n5326);
   U9143 : AOI22_X1 port map( A1 => n2831, A2 => n15268, B1 => n14703, B2 => 
                           n15269, ZN => n14704);
   U9144 : INV_X1 port map( A => n14618, ZN => n2831);
   U9145 : OAI21_X1 port map( B1 => n15269, B2 => n3748, A => n2831, ZN => 
                           n15270);
   U9146 : INV_X1 port map( A => n7233, ZN => n2832);
   U9148 : INV_X1 port map( A => n7589, ZN => n2833);
   U9149 : NOR3_X1 port map( A1 => n18017, A2 => n2834, A3 => n18020, ZN => 
                           n17960);
   U9150 : NAND2_X1 port map( A1 => n18022, A2 => n2834, ZN => n3068);
   U9151 : NOR2_X1 port map( A1 => n18353, A2 => n18354, ZN => n2836);
   U9152 : NAND2_X1 port map( A1 => n18311, A2 => n518, ZN => n2837);
   U9153 : NAND3_X1 port map( A1 => n6719, A2 => n6905, A3 => n7926, ZN => 
                           n2839);
   U9154 : NAND3_X1 port map( A1 => n7398, A2 => n6719, A3 => n7625, ZN => 
                           n2840);
   U9156 : NAND3_X1 port map( A1 => n7514, A2 => n7506, A3 => n29629, ZN => 
                           n2841);
   U9157 : NAND2_X1 port map( A1 => n28182, A2 => n23289, ZN => n2842);
   U9158 : NAND2_X1 port map( A1 => n2842, A2 => n23816, ZN => n4415);
   U9159 : NAND2_X1 port map( A1 => n2027, A2 => n12132, ZN => n5039);
   U9160 : MUX2_X1 port map( A => n29149, B => n3820, S => n11033, Z => n2843);
   U9161 : NAND2_X1 port map( A1 => n8898, A2 => n8900, ZN => n2844);
   U9162 : NOR2_X1 port map( A1 => n81, A2 => n9124, ZN => n8900);
   U9163 : XNOR2_X1 port map( A => n10251, B => n2845, ZN => n9907);
   U9164 : XNOR2_X1 port map( A => n10151, B => n2845, ZN => n10152);
   U9165 : XNOR2_X1 port map( A => n2845, B => n15576, ZN => n9621);
   U9167 : NAND3_X1 port map( A1 => n6163, A2 => n10638, A3 => n6165, ZN => 
                           n2846);
   U9168 : NOR2_X1 port map( A1 => n2846, A2 => n12042, ZN => n12044);
   U9170 : INV_X1 port map( A => n14372, ZN => n2849);
   U9171 : NAND2_X1 port map( A1 => n16985, A2 => n19560, ZN => n17639);
   U9172 : XNOR2_X1 port map( A => n2850, B => n24906, ZN => Ciphertext(13));
   U9173 : OAI21_X1 port map( B1 => n4090, B2 => n2852, A => n2851, ZN => n2850
                           );
   U9174 : INV_X1 port map( A => n27376, ZN => n2851);
   U9175 : NAND2_X1 port map( A1 => n5372, A2 => n5374, ZN => n2852);
   U9176 : INV_X1 port map( A => n2853, ZN => n18045);
   U9177 : NAND2_X1 port map( A1 => n17225, A2 => n17224, ZN => n2853);
   U9178 : NAND2_X1 port map( A1 => n2853, A2 => n18430, ZN => n17610);
   U9179 : NAND2_X1 port map( A1 => n1894, A2 => n2853, ZN => n18146);
   U9181 : NAND2_X1 port map( A1 => n18432, A2 => n2854, ZN => n18435);
   U9182 : NOR2_X1 port map( A1 => n2855, A2 => n18045, ZN => n2854);
   U9183 : NAND2_X1 port map( A1 => n17482, A2 => n4271, ZN => n2857);
   U9186 : NAND2_X1 port map( A1 => n2864, A2 => n9070, ZN => n2859);
   U9187 : NAND2_X1 port map( A1 => n602, A2 => n8819, ZN => n8475);
   U9188 : NAND2_X1 port map( A1 => n2024, A2 => n8594, ZN => n2860);
   U9189 : NAND2_X1 port map( A1 => n2862, A2 => n8977, ZN => n2861);
   U9190 : NAND2_X1 port map( A1 => n5962, A2 => n8593, ZN => n2862);
   U9191 : NAND3_X1 port map( A1 => n602, A2 => n8819, A3 => n8594, ZN => n2863
                           );
   U9192 : NAND2_X1 port map( A1 => n9072, A2 => n8741, ZN => n2864);
   U9193 : NAND2_X1 port map( A1 => n378, A2 => n24447, ZN => n5991);
   U9196 : AND2_X1 port map( A1 => n28996, A2 => n14695, ZN => n14846);
   U9197 : INV_X1 port map( A => n20152, ZN => n20097);
   U9198 : NAND2_X1 port map( A1 => n2871, A2 => n2870, ZN => n18890);
   U9199 : NAND3_X1 port map( A1 => n5053, A2 => n20096, A3 => n20152, ZN => 
                           n2870);
   U9200 : XNOR2_X2 port map( A => n18819, B => n18818, ZN => n20152);
   U9201 : NAND3_X1 port map( A1 => n28188, A2 => n20098, A3 => n20155, ZN => 
                           n2871);
   U9203 : INV_X1 port map( A => n2872, ZN => n20052);
   U9204 : NAND2_X1 port map( A1 => n20066, A2 => n20064, ZN => n2872);
   U9205 : NAND2_X1 port map( A1 => n3436, A2 => n2872, ZN => n20051);
   U9206 : NAND2_X1 port map( A1 => n6924, A2 => n2874, ZN => n2873);
   U9207 : NAND2_X1 port map( A1 => n2876, A2 => n26840, ZN => n2877);
   U9208 : INV_X1 port map( A => n25815, ZN => n2876);
   U9209 : XNOR2_X1 port map( A => n25813, B => n25812, ZN => n26507);
   U9210 : NAND3_X1 port map( A1 => n24747, A2 => n24745, A3 => n2879, ZN => 
                           n2878);
   U9211 : NAND2_X1 port map( A1 => n29545, A2 => n28550, ZN => n4980);
   U9212 : AND2_X1 port map( A1 => n21303, A2 => n24745, ZN => n24746);
   U9213 : INV_X1 port map( A => n4675, ZN => n8827);
   U9214 : NAND2_X1 port map( A1 => n3004, A2 => n7886, ZN => n2883);
   U9215 : NAND3_X1 port map( A1 => n15008, A2 => n15369, A3 => n426, ZN => 
                           n5093);
   U9217 : NAND2_X1 port map( A1 => n15236, A2 => n15235, ZN => n2885);
   U9219 : NAND2_X1 port map( A1 => n26385, A2 => n26384, ZN => n27166);
   U9220 : NAND2_X1 port map( A1 => n2888, A2 => n2887, ZN => n23132);
   U9221 : NAND2_X1 port map( A1 => n23360, A2 => n23673, ZN => n2887);
   U9222 : NAND2_X1 port map( A1 => n18521, A2 => n17724, ZN => n3544);
   U9223 : NAND2_X1 port map( A1 => n18286, A2 => n17719, ZN => n17724);
   U9224 : NAND2_X1 port map( A1 => n1925, A2 => n21425, ZN => n3238);
   U9226 : NAND2_X1 port map( A1 => n3266, A2 => n6543, ZN => n23491);
   U9228 : NAND2_X1 port map( A1 => n10403, A2 => n10402, ZN => n2892);
   U9229 : NAND3_X1 port map( A1 => n432, A2 => n5258, A3 => n11094, ZN => 
                           n11095);
   U9230 : NAND3_X1 port map( A1 => n19837, A2 => n20381, A3 => n20383, ZN => 
                           n4361);
   U9231 : OR2_X1 port map( A1 => n10003, A2 => n10002, ZN => n10004);
   U9232 : OAI21_X1 port map( B1 => n19960, B2 => n19819, A => n20545, ZN => 
                           n3473);
   U9233 : NOR2_X1 port map( A1 => n27551, A2 => n29578, ZN => n27217);
   U9234 : MUX2_X1 port map( A => n12371, B => n12370, S => n3362, Z => n2895);
   U9235 : NAND3_X2 port map( A1 => n4160, A2 => n4159, A3 => n2896, ZN => 
                           n9037);
   U9236 : NAND2_X1 port map( A1 => n7853, A2 => n2897, ZN => n2896);
   U9239 : OAI211_X2 port map( C1 => n21319, C2 => n21320, A => n21318, B => 
                           n21317, ZN => n22152);
   U9240 : NAND2_X1 port map( A1 => n21674, A2 => n21448, ZN => n4460);
   U9242 : NAND2_X1 port map( A1 => n5779, A2 => n5780, ZN => n21596);
   U9243 : INV_X1 port map( A => n10884, ZN => n11284);
   U9245 : NAND2_X1 port map( A1 => n18592, A2 => n3450, ZN => n2901);
   U9248 : INV_X1 port map( A => n4504, ZN => n16085);
   U9249 : AND2_X1 port map( A1 => n12234, A2 => n375, ZN => n6871);
   U9250 : XNOR2_X1 port map( A => n2902, B => n26113, ZN => n26125);
   U9251 : XNOR2_X1 port map( A => n2903, B => n22545, ZN => n22017);
   U9252 : XNOR2_X1 port map( A => n22016, B => n6141, ZN => n2903);
   U9253 : NOR2_X1 port map( A1 => n2904, A2 => n10920, ZN => n10921);
   U9254 : NAND2_X1 port map( A1 => n10919, A2 => n11135, ZN => n2904);
   U9256 : NAND2_X1 port map( A1 => n24377, A2 => n24376, ZN => n2905);
   U9257 : NAND2_X1 port map( A1 => n24379, A2 => n24378, ZN => n2906);
   U9259 : NAND2_X1 port map( A1 => n2908, A2 => n9071, ZN => n2907);
   U9260 : NOR2_X1 port map( A1 => n18223, A2 => n18222, ZN => n17499);
   U9262 : NAND2_X1 port map( A1 => n11294, A2 => n10318, ZN => n10309);
   U9263 : NAND2_X1 port map( A1 => n7750, A2 => n7349, ZN => n7751);
   U9264 : NAND2_X1 port map( A1 => n5694, A2 => n17215, ZN => n16751);
   U9266 : INV_X1 port map( A => n27065, ZN => n3178);
   U9267 : NAND2_X1 port map( A1 => n5016, A2 => n14652, ZN => n4642);
   U9268 : NOR2_X1 port map( A1 => n24244, A2 => n2913, ZN => n25065);
   U9269 : AND2_X1 port map( A1 => n24238, A2 => n24559, ZN => n2913);
   U9270 : INV_X1 port map( A => n11819, ZN => n12190);
   U9271 : INV_X1 port map( A => n24717, ZN => n4136);
   U9272 : AND2_X1 port map( A1 => n23474, A2 => n23761, ZN => n23190);
   U9273 : OAI21_X1 port map( B1 => n9868, B2 => n12186, A => n9867, ZN => 
                           n13396);
   U9275 : NAND2_X1 port map( A1 => n435, A2 => n10534, ZN => n11104);
   U9276 : INV_X1 port map( A => n24404, ZN => n24085);
   U9277 : OR3_X1 port map( A1 => n29602, A2 => n22531, A3 => n29020, ZN => 
                           n5713);
   U9278 : MUX2_X1 port map( A => n20051, B => n20050, S => n20063, Z => n21210
                           );
   U9280 : INV_X1 port map( A => n24316, ZN => n24667);
   U9281 : XNOR2_X1 port map( A => n13097, B => n12377, ZN => n13229);
   U9282 : OR2_X1 port map( A1 => n14195, A2 => n5978, ZN => n4435);
   U9283 : AND2_X1 port map( A1 => n18410, A2 => n17818, ZN => n4240);
   U9284 : INV_X1 port map( A => n13922, ZN => n14775);
   U9285 : XNOR2_X1 port map( A => n22316, B => n22317, ZN => n4003);
   U9286 : INV_X1 port map( A => n17620, ZN => n18159);
   U9287 : INV_X1 port map( A => n3315, ZN => n15099);
   U9288 : XNOR2_X1 port map( A => n9763, B => n10074, ZN => n10277);
   U9289 : INV_X1 port map( A => n12110, ZN => n12208);
   U9290 : INV_X1 port map( A => n6000, ZN => n12976);
   U9292 : OAI21_X1 port map( B1 => n14175, B2 => n14239, A => n14174, ZN => 
                           n3011);
   U9293 : XNOR2_X1 port map( A => n12490, B => n11389, ZN => n3687);
   U9295 : NAND2_X1 port map( A1 => n8448, A2 => n8451, ZN => n8449);
   U9296 : NAND2_X1 port map( A1 => n3330, A2 => n3329, ZN => n2917);
   U9297 : NAND2_X1 port map( A1 => n6718, A2 => n9132, ZN => n8550);
   U9298 : NOR2_X1 port map( A1 => n24892, A2 => n24227, ZN => n24229);
   U9299 : NAND2_X1 port map( A1 => n23134, A2 => n6035, ZN => n5884);
   U9300 : NAND2_X1 port map( A1 => n7438, A2 => n7626, ZN => n6719);
   U9301 : NAND2_X1 port map( A1 => n24245, A2 => n24246, ZN => n24247);
   U9302 : OR2_X1 port map( A1 => n11168, A2 => n10820, ZN => n10746);
   U9303 : NAND2_X1 port map( A1 => n2920, A2 => n2919, ZN => n23069);
   U9304 : NAND2_X1 port map( A1 => n23366, A2 => n23131, ZN => n2919);
   U9305 : NAND2_X1 port map( A1 => n23364, A2 => n2921, ZN => n2920);
   U9306 : INV_X1 port map( A => n23131, ZN => n2921);
   U9308 : NAND2_X1 port map( A1 => n20429, A2 => n20619, ZN => n2922);
   U9310 : NAND2_X1 port map( A1 => n2927, A2 => n2924, ZN => n9392);
   U9311 : NAND2_X1 port map( A1 => n2925, A2 => n8077, ZN => n2924);
   U9312 : OAI21_X1 port map( B1 => n8430, B2 => n8119, A => n2926, ZN => n2925
                           );
   U9313 : NAND2_X1 port map( A1 => n261, A2 => n8426, ZN => n2926);
   U9314 : NAND2_X1 port map( A1 => n8432, A2 => n8431, ZN => n2927);
   U9315 : NAND2_X1 port map( A1 => n8936, A2 => n2928, ZN => n8938);
   U9316 : NAND2_X1 port map( A1 => n3032, A2 => n377, ZN => n2929);
   U9317 : NAND2_X1 port map( A1 => n20574, A2 => n20568, ZN => n2930);
   U9318 : NAND2_X1 port map( A1 => n19836, A2 => n20573, ZN => n2931);
   U9325 : OAI21_X1 port map( B1 => n3072, B2 => n14261, A => n2934, ZN => 
                           n14270);
   U9326 : NAND2_X1 port map( A1 => n3071, A2 => n14263, ZN => n2934);
   U9330 : NAND2_X1 port map( A1 => n24792, A2 => n24269, ZN => n2938);
   U9331 : NAND2_X1 port map( A1 => n466, A2 => n29567, ZN => n2939);
   U9332 : NAND2_X1 port map( A1 => n29471, A2 => n24310, ZN => n2940);
   U9333 : NAND2_X1 port map( A1 => n7350, A2 => n7351, ZN => n2941);
   U9334 : NAND2_X1 port map( A1 => n11101, A2 => n11896, ZN => n2943);
   U9335 : XNOR2_X2 port map( A => n5066, B => n22901, ZN => n23456);
   U9337 : NOR2_X1 port map( A1 => n5403, A2 => n14376, ZN => n14377);
   U9338 : NOR2_X1 port map( A1 => n1991, A2 => n3031, ZN => n3030);
   U9339 : OAI211_X1 port map( C1 => n20240, C2 => n20239, A => n3532, B => 
                           n29527, ZN => n20361);
   U9340 : OAI21_X1 port map( B1 => n15098, B2 => n14901, A => n15099, ZN => 
                           n3316);
   U9342 : NAND2_X1 port map( A1 => n11982, A2 => n11980, ZN => n12227);
   U9343 : OR2_X1 port map( A1 => n13703, A2 => n12534, ZN => n4665);
   U9344 : NAND2_X1 port map( A1 => n7744, A2 => n8013, ZN => n8016);
   U9346 : OR2_X1 port map( A1 => n27119, A2 => n29016, ZN => n3456);
   U9347 : NAND3_X1 port map( A1 => n5771, A2 => n2950, A3 => n2949, ZN => 
                           n18646);
   U9348 : NAND2_X1 port map( A1 => n17907, A2 => n18343, ZN => n2949);
   U9349 : NAND2_X1 port map( A1 => n17909, A2 => n17908, ZN => n2950);
   U9350 : AND2_X1 port map( A1 => n19949, A2 => n20196, ZN => n20590);
   U9351 : NAND2_X1 port map( A1 => n21322, A2 => n20886, ZN => n6042);
   U9352 : NAND2_X1 port map( A1 => n23732, A2 => n2951, ZN => n23737);
   U9353 : NAND2_X1 port map( A1 => n2963, A2 => n2952, ZN => n7385);
   U9354 : NAND3_X1 port map( A1 => n7384, A2 => n7853, A3 => n7496, ZN => 
                           n2952);
   U9355 : NAND3_X2 port map( A1 => n6856, A2 => n6851, A3 => n6852, ZN => 
                           n16365);
   U9358 : AOI21_X1 port map( B1 => n7451, B2 => n7452, A => n8297, ZN => n3445
                           );
   U9360 : OR2_X1 port map( A1 => n10726, A2 => n10924, ZN => n10459);
   U9361 : OR2_X1 port map( A1 => n1899, A2 => n7291, ZN => n7332);
   U9364 : NAND2_X1 port map( A1 => n6729, A2 => n20324, ZN => n2956);
   U9365 : XOR2_X1 port map( A => n12432, B => n12433, Z => n4510);
   U9366 : XNOR2_X1 port map( A => n4360, B => n16480, ZN => n15779);
   U9368 : OAI21_X2 port map( B1 => n23582, B2 => n23583, A => n23581, ZN => 
                           n24757);
   U9369 : NAND2_X1 port map( A1 => n2958, A2 => n2957, ZN => n14990);
   U9370 : NAND2_X1 port map( A1 => n13682, A2 => n28806, ZN => n2957);
   U9371 : NAND2_X1 port map( A1 => n13683, A2 => n2959, ZN => n2958);
   U9372 : NOR2_X1 port map( A1 => n6565, A2 => n20433, ZN => n6564);
   U9373 : NAND2_X1 port map( A1 => n23799, A2 => n23793, ZN => n23495);
   U9374 : NOR2_X1 port map( A1 => n1938, A2 => n7675, ZN => n5256);
   U9375 : XNOR2_X1 port map( A => n22771, B => n22297, ZN => n6837);
   U9376 : NAND2_X1 port map( A1 => n1926, A2 => n15012, ZN => n6333);
   U9377 : NAND4_X2 port map( A1 => n4234, A2 => n4233, A3 => n6154, A4 => 
                           n6153, ZN => n24756);
   U9379 : XNOR2_X1 port map( A => n15796, B => n3813, ZN => n3937);
   U9380 : XNOR2_X1 port map( A => n13248, B => n12850, ZN => n2962);
   U9381 : NAND3_X1 port map( A1 => n7384, A2 => n7708, A3 => n7382, ZN => 
                           n2963);
   U9382 : NAND2_X1 port map( A1 => n12049, A2 => n12053, ZN => n12057);
   U9383 : OR3_X1 port map( A1 => n11951, A2 => n11943, A3 => n3946, ZN => 
                           n10952);
   U9385 : OR2_X1 port map( A1 => n13677, A2 => n12743, ZN => n14471);
   U9386 : NAND2_X1 port map( A1 => n2965, A2 => n2964, ZN => n14496);
   U9387 : NAND2_X1 port map( A1 => n2967, A2 => n9531, ZN => n6405);
   U9388 : OAI21_X1 port map( B1 => n5396, B2 => n8320, A => n8749, ZN => n2967
                           );
   U9389 : OAI21_X1 port map( B1 => n14101, B2 => n14230, A => n3645, ZN => 
                           n14595);
   U9391 : INV_X1 port map( A => n11136, ZN => n2968);
   U9392 : NAND2_X1 port map( A1 => n11135, A2 => n11140, ZN => n10918);
   U9393 : NAND3_X1 port map( A1 => n18018, A2 => n17564, A3 => n18017, ZN => 
                           n17773);
   U9395 : NAND2_X1 port map( A1 => n7309, A2 => n7306, ZN => n7307);
   U9396 : NAND2_X1 port map( A1 => n18150, A2 => n1894, ZN => n3468);
   U9397 : NAND2_X1 port map( A1 => n11708, A2 => n11417, ZN => n11415);
   U9399 : OAI211_X1 port map( C1 => n14181, C2 => n2972, A => n190, B => n2970
                           , ZN => n2969);
   U9400 : INV_X1 port map( A => n10809, ZN => n6347);
   U9403 : NOR2_X1 port map( A1 => n7982, A2 => n7981, ZN => n7648);
   U9404 : XNOR2_X1 port map( A => n9003, B => n9094, ZN => n5924);
   U9406 : NAND2_X1 port map( A1 => n8492, A2 => n2977, ZN => n8004);
   U9407 : NAND2_X1 port map( A1 => n20304, A2 => n2978, ZN => n20120);
   U9408 : OAI21_X2 port map( B1 => n11388, B2 => n11387, A => n11386, ZN => 
                           n4253);
   U9409 : NOR2_X1 port map( A1 => n20894, A2 => n20895, ZN => n5830);
   U9410 : NAND2_X1 port map( A1 => n8735, A2 => n2983, ZN => n8736);
   U9411 : NAND2_X1 port map( A1 => n8741, A2 => n9073, ZN => n8617);
   U9412 : NAND2_X1 port map( A1 => n3149, A2 => n3150, ZN => n22948);
   U9413 : NAND4_X2 port map( A1 => n11993, A2 => n11994, A3 => n11992, A4 => 
                           n11991, ZN => n13028);
   U9414 : NAND3_X1 port map( A1 => n24520, A2 => n24516, A3 => n24421, ZN => 
                           n3359);
   U9415 : OAI21_X1 port map( B1 => n5625, B2 => n28471, A => n4751, ZN => 
                           n4750);
   U9416 : OAI211_X1 port map( C1 => n17265, C2 => n16992, A => n16996, B => 
                           n2985, ZN => n16998);
   U9417 : XNOR2_X1 port map( A => n9952, B => n9951, ZN => n5316);
   U9418 : OR2_X1 port map( A1 => n20612, A2 => n29508, ZN => n4682);
   U9419 : INV_X1 port map( A => n11877, ZN => n11453);
   U9421 : NAND2_X1 port map( A1 => n7939, A2 => n7400, ZN => n8298);
   U9422 : NAND2_X1 port map( A1 => n21655, A2 => n2989, ZN => n2988);
   U9423 : NAND3_X1 port map( A1 => n21072, A2 => n21073, A3 => n2992, ZN => 
                           n2991);
   U9424 : INV_X1 port map( A => n18242, ZN => n4725);
   U9425 : OR2_X1 port map( A1 => n22991, A2 => n23640, ZN => n22256);
   U9426 : OAI21_X1 port map( B1 => n29315, B2 => n29146, A => n2994, ZN => 
                           n18574);
   U9427 : NAND2_X1 port map( A1 => n29146, A2 => n20081, ZN => n2994);
   U9428 : XNOR2_X2 port map( A => n7037, B => Key(150), ZN => n7456);
   U9429 : INV_X1 port map( A => n20658, ZN => n21750);
   U9430 : INV_X1 port map( A => n24809, ZN => n24499);
   U9431 : OAI211_X2 port map( C1 => n19731, C2 => n20117, A => n4682, B => 
                           n4683, ZN => n21811);
   U9432 : OR2_X1 port map( A1 => n17565, A2 => n4316, ZN => n17040);
   U9433 : INV_X1 port map( A => n21374, ZN => n21375);
   U9434 : XNOR2_X1 port map( A => n28433, B => n1119, ZN => n24847);
   U9436 : NAND2_X1 port map( A1 => n3001, A2 => n2999, ZN => n24208);
   U9437 : NAND2_X1 port map( A1 => n220, A2 => n24817, ZN => n2999);
   U9438 : XNOR2_X1 port map( A => n6100, B => n22056, ZN => n23702);
   U9439 : NOR2_X1 port map( A1 => n5706, A2 => n10777, ZN => n5705);
   U9440 : OR2_X1 port map( A1 => n7508, A2 => n7514, ZN => n7132);
   U9441 : NOR2_X2 port map( A1 => n17343, A2 => n3002, ZN => n18707);
   U9442 : NAND2_X1 port map( A1 => n2069, A2 => n17341, ZN => n3002);
   U9443 : NAND2_X1 port map( A1 => n21085, A2 => n20804, ZN => n20805);
   U9444 : NAND2_X1 port map( A1 => n24242, A2 => n24635, ZN => n24192);
   U9445 : NAND3_X1 port map( A1 => n23808, A2 => n22742, A3 => n28653, ZN => 
                           n3337);
   U9446 : NOR2_X1 port map( A1 => n384, A2 => n20239, ZN => n3005);
   U9448 : OAI21_X1 port map( B1 => n18539, B2 => n18535, A => n3006, ZN => 
                           n17700);
   U9449 : NAND2_X1 port map( A1 => n18539, A2 => n17864, ZN => n3006);
   U9450 : NAND2_X1 port map( A1 => n5616, A2 => n14349, ZN => n14015);
   U9451 : NOR2_X1 port map( A1 => n19895, A2 => n19896, ZN => n3009);
   U9452 : XNOR2_X1 port map( A => n4764, B => n29154, ZN => n24877);
   U9454 : INV_X1 port map( A => n14952, ZN => n14949);
   U9455 : NAND2_X1 port map( A1 => n15077, A2 => n14948, ZN => n14952);
   U9456 : NAND3_X1 port map( A1 => n3461, A2 => n3460, A3 => n9914, ZN => 
                           n11390);
   U9457 : INV_X1 port map( A => n3011, ZN => n3010);
   U9458 : MUX2_X1 port map( A => n11927, B => n11392, S => n11391, Z => n11393
                           );
   U9459 : NAND2_X1 port map( A1 => n11921, A2 => n11853, ZN => n11391);
   U9460 : NAND2_X1 port map( A1 => n10726, A2 => n10924, ZN => n10051);
   U9461 : NOR2_X2 port map( A1 => n3014, A2 => n11089, ZN => n12578);
   U9462 : AOI21_X1 port map( B1 => n11081, B2 => n11082, A => n433, ZN => 
                           n3014);
   U9463 : OR2_X1 port map( A1 => n8741, A2 => n9073, ZN => n8859);
   U9464 : INV_X1 port map( A => n14863, ZN => n15369);
   U9465 : XNOR2_X1 port map( A => n25508, B => n25322, ZN => n26107);
   U9466 : INV_X1 port map( A => n4166, ZN => n13827);
   U9468 : XNOR2_X1 port map( A => n9779, B => n9446, ZN => n10148);
   U9469 : NAND2_X1 port map( A1 => n3017, A2 => n4706, ZN => n18171);
   U9470 : XNOR2_X1 port map( A => n4669, B => n13260, ZN => n12966);
   U9472 : NAND2_X1 port map( A1 => n3019, A2 => n21599, ZN => n21319);
   U9473 : NAND2_X1 port map( A1 => n28442, A2 => n21601, ZN => n3019);
   U9474 : NAND3_X1 port map( A1 => n4443, A2 => n11512, A3 => n12035, ZN => 
                           n3020);
   U9475 : OAI22_X1 port map( A1 => n10933, A2 => n1879, B1 => n10932, B2 => 
                           n10931, ZN => n5905);
   U9476 : NAND3_X1 port map( A1 => n8187, A2 => n8186, A3 => n8562, ZN => 
                           n8190);
   U9477 : NAND2_X1 port map( A1 => n15089, A2 => n3022, ZN => n15092);
   U9478 : NAND2_X1 port map( A1 => n10725, A2 => n10724, ZN => n3023);
   U9479 : OAI211_X2 port map( C1 => n21415, C2 => n21414, A => n3025, B => 
                           n3024, ZN => n22473);
   U9480 : NAND2_X1 port map( A1 => n21413, A2 => n4937, ZN => n3024);
   U9481 : NAND2_X1 port map( A1 => n21411, A2 => n21412, ZN => n3025);
   U9483 : NAND2_X1 port map( A1 => n23159, A2 => n23512, ZN => n3026);
   U9484 : NOR2_X1 port map( A1 => n11108, A2 => n3027, ZN => n11109);
   U9485 : INV_X1 port map( A => n11942, ZN => n3027);
   U9486 : NAND2_X1 port map( A1 => n12271, A2 => n28202, ZN => n11942);
   U9488 : NAND2_X1 port map( A1 => n3205, A2 => n4662, ZN => n3028);
   U9489 : OAI21_X1 port map( B1 => n13612, B2 => n13611, A => n14261, ZN => 
                           n3346);
   U9493 : OAI211_X2 port map( C1 => n8352, C2 => n8431, A => n8060, B => n8059
                           , ZN => n10071);
   U9494 : NOR2_X1 port map( A1 => n26560, A2 => n28578, ZN => n3032);
   U9495 : NAND2_X1 port map( A1 => n26460, A2 => n28578, ZN => n3033);
   U9496 : NAND3_X1 port map( A1 => n8018, A2 => n7744, A3 => n7745, ZN => 
                           n7247);
   U9498 : NOR2_X1 port map( A1 => n15462, A2 => n15464, ZN => n13889);
   U9500 : NAND2_X1 port map( A1 => n10745, A2 => n4945, ZN => n11636);
   U9501 : XNOR2_X1 port map( A => n3037, B => n22471, ZN => n23391);
   U9502 : XNOR2_X1 port map( A => n22469, B => n22470, ZN => n3037);
   U9503 : NAND2_X1 port map( A1 => n17508, A2 => n17505, ZN => n16728);
   U9505 : BUF_X1 port map( A => n25268, Z => n25513);
   U9506 : AND2_X1 port map( A1 => n26682, A2 => n27433, ZN => n26833);
   U9507 : OR2_X1 port map( A1 => n24117, A2 => n24433, ZN => n24118);
   U9508 : OR2_X1 port map( A1 => n23261, A2 => n23712, ZN => n22972);
   U9509 : INV_X1 port map( A => n17872, ZN => n17937);
   U9510 : OR2_X1 port map( A1 => n21412, A2 => n20663, ZN => n21415);
   U9511 : NAND3_X1 port map( A1 => n16970, A2 => n16969, A3 => n3038, ZN => 
                           n16972);
   U9512 : NOR2_X1 port map( A1 => n13693, A2 => n29607, ZN => n4610);
   U9513 : INV_X1 port map( A => n23290, ZN => n23441);
   U9515 : AND2_X1 port map( A1 => n24583, A2 => n29026, ZN => n6056);
   U9517 : INV_X1 port map( A => n17438, ZN => n17434);
   U9518 : INV_X1 port map( A => n16980, ZN => n4002);
   U9519 : XNOR2_X1 port map( A => n3092, B => n3091, ZN => n22598);
   U9520 : OAI211_X1 port map( C1 => n20493, C2 => n20496, A => n3040, B => 
                           n5225, ZN => n5305);
   U9521 : NAND2_X1 port map( A1 => n3041, A2 => n29616, ZN => n3040);
   U9522 : INV_X1 port map( A => n20494, ZN => n3041);
   U9523 : INV_X1 port map( A => n13060, ZN => n14127);
   U9524 : INV_X1 port map( A => n18285, ZN => n17859);
   U9525 : NAND2_X1 port map( A1 => n28653, A2 => n23284, ZN => n3042);
   U9526 : OR2_X1 port map( A1 => n23809, A2 => n23806, ZN => n3043);
   U9529 : XNOR2_X1 port map( A => n3044, B => n13441, ZN => n12048);
   U9530 : XNOR2_X1 port map( A => n12034, B => n13167, ZN => n3044);
   U9531 : NAND2_X1 port map( A1 => n7565, A2 => n7562, ZN => n7124);
   U9532 : INV_X1 port map( A => n14414, ZN => n14216);
   U9534 : NAND2_X1 port map( A1 => n555, A2 => n14414, ZN => n3045);
   U9536 : NAND2_X1 port map( A1 => n585, A2 => n11284, ZN => n3046);
   U9537 : NAND2_X1 port map( A1 => n11029, A2 => n10884, ZN => n3047);
   U9538 : OAI211_X2 port map( C1 => n18002, C2 => n18337, A => n1973, B => 
                           n3048, ZN => n19427);
   U9539 : NAND2_X1 port map( A1 => n18001, A2 => n18337, ZN => n3048);
   U9540 : OAI21_X1 port map( B1 => n5870, B2 => n8523, A => n8524, ZN => n3679
                           );
   U9544 : NAND2_X1 port map( A1 => n8748, A2 => n8751, ZN => n3051);
   U9545 : NAND2_X1 port map( A1 => n3052, A2 => n23713, ZN => n23237);
   U9546 : NAND2_X1 port map( A1 => n23261, A2 => n23587, ZN => n3052);
   U9547 : NAND2_X1 port map( A1 => n3053, A2 => n23057, ZN => n6439);
   U9548 : OAI22_X1 port map( A1 => n23426, A2 => n28122, B1 => n23428, B2 => 
                           n29108, ZN => n3053);
   U9550 : NOR2_X2 port map( A1 => n4114, A2 => n11603, ZN => n6683);
   U9551 : OAI22_X1 port map( A1 => n11340, A2 => n11338, B1 => n11175, B2 => 
                           n11345, ZN => n6289);
   U9552 : NAND2_X1 port map( A1 => n3055, A2 => n29470, ZN => n23509);
   U9553 : INV_X1 port map( A => n23507, ZN => n3055);
   U9554 : NAND2_X1 port map( A1 => n24388, A2 => n24387, ZN => n23507);
   U9555 : INV_X1 port map( A => n12244, ZN => n5839);
   U9556 : NAND3_X1 port map( A1 => n10570, A2 => n11068, A3 => n10571, ZN => 
                           n11901);
   U9558 : XNOR2_X1 port map( A => n12529, B => n13563, ZN => n10538);
   U9559 : INV_X1 port map( A => n5593, ZN => n5592);
   U9560 : XNOR2_X1 port map( A => n19438, B => n18988, ZN => n3912);
   U9561 : NAND3_X1 port map( A1 => n12360, A2 => n12358, A3 => n6552, ZN => 
                           n6551);
   U9562 : NOR2_X2 port map( A1 => n17112, A2 => n17111, ZN => n17847);
   U9563 : NAND2_X1 port map( A1 => n11021, A2 => n3058, ZN => n13371);
   U9564 : NAND3_X1 port map( A1 => n14221, A2 => n5777, A3 => n14222, ZN => 
                           n16510);
   U9565 : NAND2_X1 port map( A1 => n3061, A2 => n3060, ZN => n3059);
   U9566 : INV_X1 port map( A => n24030, ZN => n3060);
   U9567 : NAND2_X1 port map( A1 => n6501, A2 => n4295, ZN => n6500);
   U9568 : NAND2_X1 port map( A1 => n13852, A2 => n14184, ZN => n14470);
   U9569 : NAND3_X1 port map( A1 => n8536, A2 => n8384, A3 => n8730, ZN => 
                           n7187);
   U9570 : NAND2_X1 port map( A1 => n6466, A2 => n14217, ZN => n14417);
   U9571 : NAND2_X1 port map( A1 => n26637, A2 => n29092, ZN => n3063);
   U9572 : NAND2_X1 port map( A1 => n27970, A2 => n26636, ZN => n3064);
   U9573 : NAND2_X1 port map( A1 => n7851, A2 => n7708, ZN => n7856);
   U9575 : INV_X1 port map( A => n10717, ZN => n6479);
   U9576 : INV_X1 port map( A => n21536, ZN => n20793);
   U9577 : NAND2_X1 port map( A1 => n21514, A2 => n21199, ZN => n21536);
   U9578 : NAND2_X1 port map( A1 => n3065, A2 => n27514, ZN => n27518);
   U9579 : NOR2_X1 port map( A1 => n27513, A2 => n27516, ZN => n3065);
   U9580 : NAND3_X1 port map( A1 => n6435, A2 => n26917, A3 => n3066, ZN => 
                           n6437);
   U9581 : INV_X1 port map( A => n27520, ZN => n27523);
   U9582 : XNOR2_X1 port map( A => n25521, B => n25069, ZN => n4810);
   U9583 : NAND2_X1 port map( A1 => n21210, A2 => n21209, ZN => n22026);
   U9584 : NAND2_X1 port map( A1 => n11922, A2 => n11852, ZN => n3410);
   U9587 : NAND2_X1 port map( A1 => n14268, A2 => n14262, ZN => n3072);
   U9588 : INV_X1 port map( A => n9577, ZN => n10192);
   U9589 : XNOR2_X1 port map( A => n9577, B => n3073, ZN => n9818);
   U9590 : OR2_X1 port map( A1 => n11819, A2 => n12198, ZN => n12127);
   U9591 : NAND2_X1 port map( A1 => n12041, A2 => n12042, ZN => n10643);
   U9593 : NAND2_X1 port map( A1 => n5498, A2 => n24364, ZN => n5501);
   U9594 : OAI211_X1 port map( C1 => n17902, C2 => n18111, A => n18110, B => 
                           n17798, ZN => n3074);
   U9595 : OAI21_X1 port map( B1 => n7321, B2 => n7116, A => n7768, ZN => n5244
                           );
   U9596 : NAND3_X1 port map( A1 => n27288, A2 => n27275, A3 => n27287, ZN => 
                           n3146);
   U9598 : INV_X1 port map( A => n3078, ZN => n3077);
   U9599 : OAI21_X1 port map( B1 => n5635, B2 => n3080, A => n3079, ZN => 
                           n15181);
   U9600 : AOI21_X2 port map( B1 => n11561, B2 => n11562, A => n11560, ZN => 
                           n13190);
   U9601 : XNOR2_X2 port map( A => n12903, B => n12902, ZN => n14084);
   U9602 : NAND3_X1 port map( A1 => n2014, A2 => n6322, A3 => n6323, ZN => 
                           n26652);
   U9603 : AOI22_X1 port map( A1 => n26653, A2 => n27548, B1 => n27541, B2 => 
                           n27547, ZN => n26654);
   U9604 : OAI22_X1 port map( A1 => n19032, A2 => n20232, B1 => n383, B2 => 
                           n20231, ZN => n5274);
   U9605 : NOR2_X1 port map( A1 => n20956, A2 => n20957, ZN => n3280);
   U9606 : NAND2_X1 port map( A1 => n5207, A2 => n14243, ZN => n3082);
   U9608 : NAND2_X1 port map( A1 => n17577, A2 => n18251, ZN => n3085);
   U9610 : INV_X1 port map( A => n4515, ZN => n14802);
   U9611 : NAND3_X2 port map( A1 => n13875, A2 => n13876, A3 => n5015, ZN => 
                           n4515);
   U9612 : NAND2_X1 port map( A1 => n25994, A2 => n27371, ZN => n25995);
   U9613 : NAND2_X1 port map( A1 => n14167, A2 => n14169, ZN => n6744);
   U9614 : NAND2_X1 port map( A1 => n8081, A2 => n8336, ZN => n8506);
   U9615 : INV_X1 port map( A => n21645, ZN => n4659);
   U9616 : NAND2_X1 port map( A1 => n2057, A2 => n424, ZN => n3090);
   U9617 : NAND3_X1 port map( A1 => n8277, A2 => n8279, A3 => n8278, ZN => 
                           n3094);
   U9619 : NAND2_X1 port map( A1 => n21216, A2 => n21000, ZN => n20998);
   U9620 : NAND2_X1 port map( A1 => n3095, A2 => n7967, ZN => n4698);
   U9621 : OAI21_X1 port map( B1 => n7963, B2 => n1938, A => n7236, ZN => n3095
                           );
   U9622 : AND3_X1 port map( A1 => n3541, A2 => n3481, A3 => n24588, ZN => 
                           n5863);
   U9623 : OR2_X1 port map( A1 => n10093, A2 => n11152, ZN => n3165);
   U9624 : NAND2_X1 port map( A1 => n5332, A2 => n2205, ZN => n24637);
   U9625 : NAND2_X1 port map( A1 => n5576, A2 => n3583, ZN => n15535);
   U9626 : NAND2_X1 port map( A1 => n18034, A2 => n18154, ZN => n4854);
   U9627 : XNOR2_X1 port map( A => n13505, B => n13134, ZN => n3097);
   U9628 : NAND3_X2 port map( A1 => n3668, A2 => n5371, A3 => n3667, ZN => 
                           n13451);
   U9630 : NOR2_X1 port map( A1 => n6374, A2 => n10863, ZN => n6372);
   U9631 : NAND2_X1 port map( A1 => n3100, A2 => n3099, ZN => n17122);
   U9633 : AOI21_X1 port map( B1 => n10686, B2 => n9362, A => n6775, ZN => 
                           n6774);
   U9634 : INV_X1 port map( A => n4852, ZN => n16654);
   U9635 : NOR2_X2 port map( A1 => n17257, A2 => n17256, ZN => n18240);
   U9636 : OR2_X2 port map( A1 => n12091, A2 => n12092, ZN => n11856);
   U9637 : NAND2_X1 port map( A1 => n14310, A2 => n14309, ZN => n13888);
   U9639 : NAND2_X1 port map( A1 => n3106, A2 => n3105, ZN => n10818);
   U9640 : NAND2_X1 port map( A1 => n10815, A2 => n28207, ZN => n3105);
   U9641 : NAND2_X1 port map( A1 => n3107, A2 => n28157, ZN => n3106);
   U9642 : OAI21_X1 port map( B1 => n28638, B2 => n3585, A => n3584, ZN => 
                           n3107);
   U9643 : NOR2_X1 port map( A1 => n24368, A2 => n24367, ZN => n24303);
   U9645 : INV_X1 port map( A => n15175, ZN => n15459);
   U9646 : OR2_X1 port map( A1 => n572, A2 => n11754, ZN => n11477);
   U9647 : OR2_X1 port map( A1 => n21936, A2 => n21935, ZN => n21937);
   U9648 : INV_X1 port map( A => n21424, ZN => n5000);
   U9649 : AND2_X1 port map( A1 => n3922, A2 => n14893, ZN => n12011);
   U9650 : XNOR2_X1 port map( A => n12849, B => n12554, ZN => n13332);
   U9651 : INV_X1 port map( A => n6482, ZN => n4744);
   U9653 : OAI21_X1 port map( B1 => n15169, B2 => n6925, A => n1850, ZN => 
                           n14553);
   U9654 : INV_X1 port map( A => n23765, ZN => n23766);
   U9655 : XNOR2_X1 port map( A => n6416, B => n6415, ZN => n17272);
   U9656 : INV_X1 port map( A => n24397, ZN => n24323);
   U9657 : INV_X1 port map( A => n23655, ZN => n24793);
   U9658 : XNOR2_X1 port map( A => n3913, B => n19584, ZN => n18988);
   U9659 : INV_X1 port map( A => n22735, ZN => n6119);
   U9660 : AOI21_X1 port map( B1 => n28916, B2 => n21089, A => n21930, ZN => 
                           n3560);
   U9661 : XNOR2_X1 port map( A => n29035, B => n19323, ZN => n19693);
   U9662 : NOR2_X1 port map( A1 => n8521, A2 => n8811, ZN => n5869);
   U9663 : AOI21_X1 port map( B1 => n28638, B2 => n10563, A => n11196, ZN => 
                           n6272);
   U9664 : NAND3_X1 port map( A1 => n12508, A2 => n3108, A3 => n10863, ZN => 
                           n11835);
   U9666 : INV_X1 port map( A => n26769, ZN => n6768);
   U9667 : NAND2_X1 port map( A1 => n296, A2 => n18972, ZN => n5106);
   U9668 : INV_X1 port map( A => n15642, ZN => n16425);
   U9669 : NAND3_X1 port map( A1 => n7673, A2 => n7481, A3 => n8281, ZN => 
                           n7482);
   U9670 : OR2_X1 port map( A1 => n7851, A2 => n7384, ZN => n7383);
   U9671 : AND2_X1 port map( A1 => n14435, A2 => n14207, ZN => n13957);
   U9672 : XNOR2_X1 port map( A => n12847, B => n12848, ZN => n3110);
   U9674 : XNOR2_X1 port map( A => n19263, B => n19639, ZN => n3111);
   U9675 : XNOR2_X1 port map( A => n9491, B => n9492, ZN => n6135);
   U9676 : NAND2_X1 port map( A1 => n11255, A2 => n11315, ZN => n3113);
   U9679 : NAND2_X1 port map( A1 => n3895, A2 => n3896, ZN => n5682);
   U9680 : XNOR2_X2 port map( A => n19107, B => n19106, ZN => n20488);
   U9681 : NAND3_X1 port map( A1 => n8890, A2 => n8507, A3 => n8886, ZN => 
                           n8508);
   U9683 : NAND3_X1 port map( A1 => n3118, A2 => n8210, A3 => n3117, ZN => 
                           n8838);
   U9684 : NAND2_X1 port map( A1 => n3159, A2 => n8209, ZN => n3118);
   U9689 : INV_X1 port map( A => n9431, ZN => n9678);
   U9690 : AND2_X1 port map( A1 => n20786, A2 => n21097, ZN => n20799);
   U9691 : AOI21_X1 port map( B1 => n3123, B2 => n7829, A => n8205, ZN => n7435
                           );
   U9692 : NAND2_X1 port map( A1 => n8201, A2 => n7828, ZN => n3123);
   U9693 : AND2_X1 port map( A1 => n24794, A2 => n28512, ZN => n3124);
   U9694 : NAND2_X1 port map( A1 => n16806, A2 => n17259, ZN => n16669);
   U9695 : INV_X1 port map( A => n26746, ZN => n5760);
   U9697 : NAND2_X1 port map( A1 => n3125, A2 => n14322, ZN => n14066);
   U9698 : NAND3_X1 port map( A1 => n15294, A2 => n15293, A3 => n15291, ZN => 
                           n14838);
   U9699 : OR2_X1 port map( A1 => n13909, A2 => n14047, ZN => n5730);
   U9700 : NAND2_X1 port map( A1 => n6661, A2 => n12004, ZN => n11686);
   U9701 : NOR2_X2 port map( A1 => n10567, A2 => n10566, ZN => n12004);
   U9702 : XNOR2_X1 port map( A => n6453, B => n15978, ZN => n6455);
   U9703 : OR2_X1 port map( A1 => n21736, A2 => n29314, ZN => n21477);
   U9704 : NAND2_X1 port map( A1 => n3375, A2 => n14359, ZN => n13032);
   U9705 : NAND3_X1 port map( A1 => n8286, A2 => n7913, A3 => n7914, ZN => 
                           n7918);
   U9706 : INV_X1 port map( A => n23658, ZN => n5773);
   U9707 : INV_X1 port map( A => n13902, ZN => n4425);
   U9708 : AND2_X1 port map( A1 => n15361, A2 => n4992, ZN => n14753);
   U9709 : NAND3_X1 port map( A1 => n9234, A2 => n9235, A3 => n9233, ZN => 
                           n9236);
   U9710 : NAND2_X1 port map( A1 => n20105, A2 => n3126, ZN => n20933);
   U9711 : INV_X1 port map( A => n7426, ZN => n6993);
   U9712 : INV_X1 port map( A => n17864, ZN => n18536);
   U9713 : OR2_X1 port map( A1 => n27056, A2 => n26850, ZN => n27055);
   U9714 : OR2_X1 port map( A1 => n14771, A2 => n14770, ZN => n3638);
   U9715 : OR2_X1 port map( A1 => n23010, A2 => n6227, ZN => n23140);
   U9716 : INV_X1 port map( A => n17957, ZN => n4905);
   U9717 : OAI21_X1 port map( B1 => n8658, B2 => n8654, A => n8503, ZN => n3127
                           );
   U9718 : INV_X1 port map( A => n581, ZN => n5914);
   U9720 : NAND2_X1 port map( A1 => n10750, A2 => n11198, ZN => n3130);
   U9721 : NAND2_X1 port map( A1 => n20832, A2 => n3131, ZN => n22718);
   U9722 : OR2_X1 port map( A1 => n7308, A2 => n7093, ZN => n7863);
   U9723 : AND2_X1 port map( A1 => n28197, A2 => n15361, ZN => n14750);
   U9724 : INV_X1 port map( A => n14922, ZN => n6699);
   U9725 : AND2_X1 port map( A1 => n10797, A2 => n11225, ZN => n10621);
   U9726 : INV_X1 port map( A => n19554, ZN => n19927);
   U9727 : AND2_X1 port map( A1 => n28207, A2 => n10814, ZN => n6677);
   U9728 : NAND3_X1 port map( A1 => n349, A2 => n12252, A3 => n12253, ZN => 
                           n3553);
   U9730 : INV_X1 port map( A => n20148, ZN => n20102);
   U9733 : INV_X1 port map( A => n18011, ZN => n18477);
   U9735 : NAND3_X1 port map( A1 => n3137, A2 => n5854, A3 => n4877, ZN => 
                           n3136);
   U9736 : INV_X1 port map( A => n20038, ZN => n3137);
   U9738 : NOR2_X1 port map( A1 => n4044, A2 => n17780, ZN => n17783);
   U9739 : XNOR2_X1 port map( A => n22173, B => n22483, ZN => n23261);
   U9741 : INV_X1 port map( A => n3441, ZN => n5709);
   U9742 : INV_X1 port map( A => n15265, ZN => n15499);
   U9744 : NOR2_X1 port map( A1 => n5584, A2 => n14331, ZN => n14410);
   U9745 : OAI21_X1 port map( B1 => n14410, B2 => n14409, A => n14408, ZN => 
                           n4001);
   U9746 : NOR2_X1 port map( A1 => n24293, A2 => n24533, ZN => n24892);
   U9747 : XNOR2_X1 port map( A => n25711, B => n25713, ZN => n3168);
   U9748 : OAI21_X1 port map( B1 => n12075, B2 => n5974, A => n5973, ZN => 
                           n5972);
   U9749 : XNOR2_X1 port map( A => n18779, B => n18991, ZN => n18499);
   U9750 : XNOR2_X1 port map( A => n16279, B => n3138, ZN => n16370);
   U9751 : NAND2_X1 port map( A1 => n17547, A2 => n4624, ZN => n4623);
   U9752 : NAND2_X1 port map( A1 => n4626, A2 => n4625, ZN => n17547);
   U9753 : NAND3_X1 port map( A1 => n6875, A2 => n9176, A3 => n8983, ZN => 
                           n3140);
   U9755 : OAI21_X2 port map( B1 => n8917, B2 => n8674, A => n8673, ZN => 
                           n10257);
   U9757 : XNOR2_X1 port map( A => n9272, B => n10148, ZN => n3141);
   U9758 : INV_X1 port map( A => n28523, ZN => n24027);
   U9759 : OAI211_X2 port map( C1 => n11408, C2 => n11645, A => n3143, B => 
                           n3142, ZN => n13405);
   U9760 : NAND2_X1 port map( A1 => n12142, A2 => n11715, ZN => n3142);
   U9762 : AOI21_X1 port map( B1 => n20336, B2 => n20625, A => n20623, ZN => 
                           n3144);
   U9763 : INV_X1 port map( A => n20889, ZN => n5205);
   U9764 : OAI22_X1 port map( A1 => n20643, A2 => n20905, B1 => n21605, B2 => 
                           n21599, ZN => n3145);
   U9765 : XNOR2_X2 port map( A => n16502, B => n16501, ZN => n16797);
   U9766 : NAND3_X1 port map( A1 => n3998, A2 => n3999, A3 => n11750, ZN => 
                           n4000);
   U9767 : OAI21_X1 port map( B1 => n27285, B2 => n27291, A => n3146, ZN => 
                           n27252);
   U9768 : NOR2_X1 port map( A1 => n23513, A2 => n339, ZN => n3147);
   U9770 : NAND2_X1 port map( A1 => n12037, A2 => n12158, ZN => n4443);
   U9771 : NOR2_X1 port map( A1 => n17927, A2 => n18301, ZN => n17929);
   U9772 : NAND2_X1 port map( A1 => n19764, A2 => n5424, ZN => n18847);
   U9773 : OAI22_X1 port map( A1 => n20048, A2 => n19761, B1 => n18892, B2 => 
                           n20049, ZN => n5424);
   U9775 : NOR2_X1 port map( A1 => n21291, A2 => n21290, ZN => n20913);
   U9776 : NAND2_X1 port map( A1 => n29564, A2 => n23827, ZN => n22944);
   U9777 : NAND2_X1 port map( A1 => n22945, A2 => n23741, ZN => n3150);
   U9778 : XNOR2_X1 port map( A => n9685, B => n6440, ZN => n4590);
   U9779 : XNOR2_X1 port map( A => n3151, B => n624, ZN => Ciphertext(111));
   U9780 : OAI211_X1 port map( C1 => n26893, C2 => n26894, A => n26891, B => 
                           n26892, ZN => n3151);
   U9782 : NAND2_X1 port map( A1 => n14518, A2 => n15217, ZN => n14837);
   U9783 : XNOR2_X2 port map( A => n16268, B => n16267, ZN => n17487);
   U9785 : NAND2_X1 port map( A1 => n803, A2 => n24803, ZN => n24261);
   U9786 : NAND2_X1 port map( A1 => n14767, A2 => n14810, ZN => n13924);
   U9788 : NAND4_X2 port map( A1 => n8833, A2 => n8834, A3 => n8832, A4 => 
                           n8831, ZN => n9941);
   U9789 : OAI21_X2 port map( B1 => n29119, B2 => n8137, A => n4940, ZN => 
                           n8981);
   U9790 : NAND2_X1 port map( A1 => n1834, A2 => n10713, ZN => n6152);
   U9791 : OR3_X1 port map( A1 => n29083, A2 => n16541, A3 => n17456, ZN => 
                           n16542);
   U9792 : NOR2_X1 port map( A1 => n30, A2 => n14400, ZN => n4010);
   U9795 : NAND2_X1 port map( A1 => n5724, A2 => n5726, ZN => n5721);
   U9796 : INV_X1 port map( A => n18301, ZN => n3153);
   U9797 : NAND2_X1 port map( A1 => n17278, A2 => n17277, ZN => n16767);
   U9798 : NAND2_X1 port map( A1 => n10528, A2 => n11047, ZN => n11264);
   U9800 : AOI21_X1 port map( B1 => n7210, B2 => n7211, A => n8264, ZN => n3155
                           );
   U9801 : NAND2_X1 port map( A1 => n29395, A2 => n9530, ZN => n3157);
   U9802 : OR2_X1 port map( A1 => n18919, A2 => n21091, ZN => n4876);
   U9803 : OR2_X1 port map( A1 => n14398, A2 => n14401, ZN => n14210);
   U9804 : NAND2_X1 port map( A1 => n11112, A2 => n11111, ZN => n3509);
   U9805 : NAND2_X1 port map( A1 => n29546, A2 => n17355, ZN => n17358);
   U9806 : OR2_X2 port map( A1 => n11663, A2 => n11664, ZN => n13444);
   U9807 : AOI21_X2 port map( B1 => n23195, B2 => n23470, A => n3158, ZN => 
                           n24559);
   U9808 : NAND2_X1 port map( A1 => n370, A2 => n8208, ZN => n3159);
   U9809 : INV_X1 port map( A => n5316, ZN => n11111);
   U9810 : INV_X1 port map( A => n22026, ZN => n22288);
   U9811 : OR2_X1 port map( A1 => n14045, A2 => n14046, ZN => n5064);
   U9812 : NAND2_X1 port map( A1 => n3162, A2 => n3160, ZN => n11473);
   U9813 : NAND3_X1 port map( A1 => n3636, A2 => n10477, A3 => n3161, ZN => 
                           n3160);
   U9814 : NAND2_X1 port map( A1 => n10479, A2 => n11350, ZN => n3162);
   U9816 : INV_X1 port map( A => n23228, ZN => n3432);
   U9817 : NOR2_X1 port map( A1 => n14842, A2 => n14695, ZN => n14060);
   U9818 : OAI22_X1 port map( A1 => n1076, A2 => n26426, B1 => n26431, B2 => 
                           n26425, ZN => n26276);
   U9819 : NAND2_X1 port map( A1 => n10696, A2 => n10989, ZN => n3801);
   U9820 : OAI21_X1 port map( B1 => n27121, B2 => n27122, A => n3456, ZN => 
                           n27128);
   U9821 : NAND3_X1 port map( A1 => n7706, A2 => n3163, A3 => n371, ZN => n4159
                           );
   U9822 : NAND2_X1 port map( A1 => n7705, A2 => n7852, ZN => n3163);
   U9823 : INV_X1 port map( A => n29647, ZN => n18509);
   U9824 : NOR2_X1 port map( A1 => n5265, A2 => n28608, ZN => n5264);
   U9825 : NAND3_X2 port map( A1 => n5082, A2 => n4629, A3 => n17668, ZN => 
                           n19232);
   U9826 : NAND2_X1 port map( A1 => n28188, A2 => n20152, ZN => n20043);
   U9827 : NAND2_X1 port map( A1 => n3166, A2 => n6027, ZN => n4733);
   U9830 : NAND2_X1 port map( A1 => n3171, A2 => n3170, ZN => n3169);
   U9831 : NAND2_X1 port map( A1 => n17124, A2 => n16723, ZN => n3170);
   U9832 : INV_X1 port map( A => n16725, ZN => n3172);
   U9834 : NAND2_X1 port map( A1 => n6407, A2 => n23331, ZN => n24397);
   U9836 : OAI21_X1 port map( B1 => n11742, B2 => n11740, A => n3176, ZN => 
                           n11448);
   U9837 : NAND2_X1 port map( A1 => n11742, A2 => n11907, ZN => n3176);
   U9838 : NAND3_X1 port map( A1 => n27066, A2 => n26616, A3 => n3178, ZN => 
                           n3177);
   U9839 : XNOR2_X1 port map( A => n16204, B => n16242, ZN => n16206);
   U9841 : INV_X1 port map( A => n14178, ZN => n14450);
   U9843 : NAND3_X1 port map( A1 => n8439, A2 => n8785, A3 => n8719, ZN => 
                           n8367);
   U9844 : NAND2_X1 port map( A1 => n3806, A2 => n4290, ZN => n14463);
   U9845 : NAND2_X1 port map( A1 => n19927, A2 => n20266, ZN => n19931);
   U9846 : OAI21_X1 port map( B1 => n10876, B2 => n11220, A => n11104, ZN => 
                           n10535);
   U9847 : INV_X1 port map( A => n6779, ZN => n5573);
   U9849 : NAND2_X1 port map( A1 => n18590, A2 => n18591, ZN => n18593);
   U9850 : NAND2_X1 port map( A1 => n17065, A2 => n17450, ZN => n17128);
   U9852 : AND3_X2 port map( A1 => n24165, A2 => n6946, A3 => n24164, ZN => 
                           n26039);
   U9853 : NAND2_X1 port map( A1 => n587, A2 => n11204, ZN => n11205);
   U9854 : NAND2_X1 port map( A1 => n7612, A2 => n7611, ZN => n3179);
   U9855 : NAND3_X1 port map( A1 => n17542, A2 => n17217, A3 => n28454, ZN => 
                           n6642);
   U9856 : OAI21_X1 port map( B1 => n11653, B2 => n3603, A => n12155, ZN => 
                           n3795);
   U9859 : XNOR2_X2 port map( A => n16364, B => n16363, ZN => n17374);
   U9860 : NAND3_X1 port map( A1 => n3184, A2 => n1840, A3 => n22401, ZN => 
                           n21069);
   U9861 : NAND2_X1 port map( A1 => n21068, A2 => n21664, ZN => n3184);
   U9862 : NAND3_X1 port map( A1 => n7883, A2 => n7585, A3 => n7882, ZN => 
                           n3185);
   U9863 : NAND2_X1 port map( A1 => n20334, A2 => n20625, ZN => n3186);
   U9864 : NAND3_X1 port map( A1 => n14370, A2 => n14120, A3 => n14366, ZN => 
                           n12977);
   U9866 : NAND2_X1 port map( A1 => n23679, A2 => n29544, ZN => n3189);
   U9867 : NOR2_X1 port map( A1 => n28535, A2 => n3190, ZN => n26133);
   U9868 : NAND2_X1 port map( A1 => n7521, A2 => n7266, ZN => n7710);
   U9869 : NAND2_X1 port map( A1 => n5611, A2 => n23761, ZN => n3192);
   U9870 : NAND3_X1 port map( A1 => n20550, A2 => n5982, A3 => n20551, ZN => 
                           n3194);
   U9871 : NAND2_X1 port map( A1 => n21321, A2 => n28584, ZN => n4342);
   U9872 : NAND2_X1 port map( A1 => n3797, A2 => n24403, ZN => n4081);
   U9873 : OAI21_X1 port map( B1 => n471, B2 => n24256, A => n24012, ZN => 
                           n6788);
   U9875 : NAND2_X1 port map( A1 => n3716, A2 => n4053, ZN => n21227);
   U9876 : NAND2_X1 port map( A1 => n4540, A2 => n4541, ZN => n9684);
   U9877 : INV_X1 port map( A => n24639, ZN => n24196);
   U9879 : NOR2_X1 port map( A1 => n20611, A2 => n3547, ZN => n20442);
   U9880 : XNOR2_X1 port map( A => n16196, B => n6159, ZN => n6158);
   U9881 : NAND3_X1 port map( A1 => n14446, A2 => n14421, A3 => n13954, ZN => 
                           n13956);
   U9882 : NAND2_X1 port map( A1 => n20119, A2 => n19947, ZN => n20307);
   U9885 : NAND2_X1 port map( A1 => n28721, A2 => n7821, ZN => n6987);
   U9886 : NAND2_X1 port map( A1 => n17880, A2 => n19828, ZN => n17958);
   U9887 : NAND2_X1 port map( A1 => n7669, A2 => n7670, ZN => n7672);
   U9889 : OR2_X1 port map( A1 => n12057, A2 => n12313, ZN => n11772);
   U9890 : INV_X1 port map( A => n15583, ZN => n16328);
   U9891 : NOR2_X1 port map( A1 => n9018, A2 => n9016, ZN => n8481);
   U9892 : OR2_X1 port map( A1 => n14534, A2 => n15456, ZN => n15177);
   U9893 : INV_X1 port map( A => n5150, ZN => n10804);
   U9894 : AOI22_X1 port map( A1 => n20691, A2 => n20690, B1 => n21366, B2 => 
                           n21713, ZN => n21718);
   U9895 : INV_X1 port map( A => n26222, ZN => n5035);
   U9896 : XNOR2_X1 port map( A => n6212, B => n21728, ZN => n22777);
   U9897 : NAND2_X1 port map( A1 => n3466, A2 => n3468, ZN => n3197);
   U9898 : NAND2_X1 port map( A1 => n3198, A2 => n10993, ZN => n3455);
   U9899 : NAND2_X1 port map( A1 => n10991, A2 => n10992, ZN => n3198);
   U9900 : NAND3_X1 port map( A1 => n23391, A2 => n23392, A3 => n23839, ZN => 
                           n3199);
   U9901 : NAND2_X1 port map( A1 => n11926, A2 => n3201, ZN => n3200);
   U9902 : NAND2_X1 port map( A1 => n11925, A2 => n574, ZN => n3202);
   U9903 : NAND2_X1 port map( A1 => n3203, A2 => n8303, ZN => n8306);
   U9904 : NAND2_X1 port map( A1 => n23304, A2 => n4178, ZN => n3204);
   U9905 : NOR2_X1 port map( A1 => n11347, A2 => n10476, ZN => n10849);
   U9906 : NAND2_X1 port map( A1 => n15409, A2 => n14893, ZN => n14940);
   U9908 : NAND2_X1 port map( A1 => n14994, A2 => n14992, ZN => n14993);
   U9910 : NAND2_X1 port map( A1 => n14916, A2 => n15490, ZN => n5645);
   U9911 : XNOR2_X1 port map( A => n25889, B => n25927, ZN => n24932);
   U9913 : AOI21_X1 port map( B1 => n19870, B2 => n3213, A => n20106, ZN => 
                           n20736);
   U9914 : NAND2_X1 port map( A1 => n20147, A2 => n20148, ZN => n3213);
   U9915 : NAND2_X1 port map( A1 => n3216, A2 => n3214, ZN => n23671);
   U9916 : NAND2_X1 port map( A1 => n23669, A2 => n29123, ZN => n3214);
   U9918 : NAND2_X1 port map( A1 => n23664, A2 => n23663, ZN => n3216);
   U9919 : OAI21_X1 port map( B1 => n13206, B2 => n12125, A => n3217, ZN => 
                           n10441);
   U9920 : NAND2_X1 port map( A1 => n11730, A2 => n11824, ZN => n3217);
   U9921 : XNOR2_X1 port map( A => n13246, B => n13243, ZN => n5166);
   U9922 : NAND2_X1 port map( A1 => n3314, A2 => n3316, ZN => n3218);
   U9923 : AND3_X1 port map( A1 => n26317, A2 => n26313, A3 => n2441, ZN => 
                           n26319);
   U9925 : OAI22_X1 port map( A1 => n26309, A2 => n27155, B1 => n401, B2 => 
                           n3220, ZN => n26312);
   U9926 : OR2_X1 port map( A1 => n17303, A2 => n3221, ZN => n17422);
   U9927 : NOR2_X1 port map( A1 => n17421, A2 => n29152, ZN => n3221);
   U9928 : NAND2_X1 port map( A1 => n5714, A2 => n17304, ZN => n17303);
   U9929 : INV_X1 port map( A => n17018, ZN => n6539);
   U9930 : NAND2_X1 port map( A1 => n15087, A2 => n14563, ZN => n14878);
   U9931 : NAND2_X1 port map( A1 => n7917, A2 => n7912, ZN => n7630);
   U9932 : NAND2_X1 port map( A1 => n5236, A2 => n23153, ZN => n24642);
   U9933 : NAND2_X1 port map( A1 => n8133, A2 => n8048, ZN => n7556);
   U9934 : MUX2_X1 port map( A => n9064, B => n8866, S => n8872, Z => n8601);
   U9936 : XNOR2_X1 port map( A => n4504, B => n16589, ZN => n15998);
   U9937 : OAI21_X1 port map( B1 => n11121, B2 => n11123, A => n6144, ZN => 
                           n10540);
   U9938 : NOR2_X1 port map( A1 => n7649, A2 => n7998, ZN => n7059);
   U9939 : NAND3_X1 port map( A1 => n7968, A2 => n7964, A3 => n3226, ZN => 
                           n5470);
   U9940 : OR2_X1 port map( A1 => n21109, A2 => n5939, ZN => n5634);
   U9941 : NAND2_X1 port map( A1 => n3595, A2 => n9565, ZN => n8947);
   U9942 : AND2_X1 port map( A1 => n23783, A2 => n23786, ZN => n23484);
   U9945 : NAND2_X1 port map( A1 => n26622, A2 => n27084, ZN => n3230);
   U9946 : INV_X1 port map( A => n26621, ZN => n3231);
   U9948 : NAND2_X1 port map( A1 => n27327, A2 => n29504, ZN => n26544);
   U9949 : NAND2_X1 port map( A1 => n3235, A2 => n3233, ZN => n17299);
   U9950 : NAND2_X1 port map( A1 => n3234, A2 => n17298, ZN => n3233);
   U9951 : INV_X1 port map( A => n17296, ZN => n3234);
   U9952 : NAND2_X1 port map( A1 => n17297, A2 => n29072, ZN => n3235);
   U9955 : OAI21_X1 port map( B1 => n25968, B2 => n27003, A => n29524, ZN => 
                           n25679);
   U9956 : OAI21_X1 port map( B1 => n5929, B2 => n21084, A => n3238, ZN => 
                           n3237);
   U9957 : INV_X1 port map( A => n14192, ZN => n3269);
   U9958 : OAI22_X1 port map( A1 => n27825, A2 => n27828, B1 => n26901, B2 => 
                           n27100, ZN => n27249);
   U9959 : AOI21_X1 port map( B1 => n6220, B2 => n28428, A => n28622, ZN => 
                           n23224);
   U9960 : INV_X1 port map( A => n23612, ZN => n4599);
   U9962 : OAI211_X1 port map( C1 => n5129, C2 => n5594, A => n9425, B => n3609
                           , ZN => n5330);
   U9963 : OR2_X1 port map( A1 => n11113, A2 => n10461, ZN => n11116);
   U9964 : NAND2_X1 port map( A1 => n3241, A2 => n3240, ZN => n22960);
   U9965 : NAND2_X1 port map( A1 => n23391, A2 => n22958, ZN => n3240);
   U9966 : NAND2_X1 port map( A1 => n22959, A2 => n6279, ZN => n3241);
   U9967 : INV_X1 port map( A => n10856, ZN => n4591);
   U9968 : INV_X1 port map( A => n19718, ZN => n5161);
   U9969 : OR2_X1 port map( A1 => n17454, A2 => n17455, ZN => n6800);
   U9970 : OR2_X1 port map( A1 => n23343, A2 => n23138, ZN => n6294);
   U9972 : INV_X1 port map( A => n18538, ZN => n18528);
   U9973 : INV_X1 port map( A => n26708, ZN => n25417);
   U9974 : INV_X1 port map( A => n12337, ZN => n11915);
   U9976 : INV_X1 port map( A => n19463, ZN => n18675);
   U9977 : OAI211_X1 port map( C1 => n25404, C2 => n28908, A => n25618, B => 
                           n280, ZN => n5831);
   U9978 : OAI22_X1 port map( A1 => n18509, A2 => n18078, B1 => n18510, B2 => 
                           n418, ZN => n17861);
   U9979 : XNOR2_X1 port map( A => n22269, B => n22268, ZN => n22284);
   U9980 : XNOR2_X1 port map( A => n12794, B => n12793, ZN => n13674);
   U9981 : OAI211_X1 port map( C1 => n10851, C2 => n11163, A => n11308, B => 
                           n9686, ZN => n3935);
   U9985 : NAND2_X1 port map( A1 => n23613, A2 => n28544, ZN => n3245);
   U9986 : NAND2_X1 port map( A1 => n20444, A2 => n6843, ZN => n3246);
   U9987 : OAI211_X1 port map( C1 => n17620, C2 => n18155, A => n18156, B => 
                           n3249, ZN => n3248);
   U9988 : NAND2_X1 port map( A1 => n17620, A2 => n18034, ZN => n3249);
   U9989 : NOR2_X1 port map( A1 => n24143, A2 => n24593, ZN => n3251);
   U9990 : INV_X1 port map( A => n24507, ZN => n3715);
   U9991 : NAND2_X1 port map( A1 => n3254, A2 => n25556, ZN => n28027);
   U9992 : NAND2_X1 port map( A1 => n25555, A2 => n27043, ZN => n3254);
   U9993 : NAND2_X1 port map( A1 => n3259, A2 => n3258, ZN => n21246);
   U9994 : NAND3_X1 port map( A1 => n21242, A2 => n21346, A3 => n21692, ZN => 
                           n3258);
   U9995 : NAND2_X1 port map( A1 => n21245, A2 => n3260, ZN => n3259);
   U9996 : OAI211_X1 port map( C1 => n28072, C2 => n28071, A => n3262, B => 
                           n3261, ZN => n28074);
   U9997 : OR2_X1 port map( A1 => n28070, A2 => n28069, ZN => n3261);
   U9998 : NAND2_X1 port map( A1 => n15100, A2 => n3315, ZN => n3314);
   U9999 : XNOR2_X1 port map( A => n3263, B => n26821, ZN => Ciphertext(33));
   U10000 : INV_X1 port map( A => n526, ZN => n3264);
   U10001 : NAND2_X1 port map( A1 => n27526, A2 => n27520, ZN => n27509);
   U10002 : NOR2_X2 port map( A1 => n19887, A2 => n19888, ZN => n21457);
   U10003 : NAND2_X1 port map( A1 => n23488, A2 => n23487, ZN => n3266);
   U10005 : NOR2_X1 port map( A1 => n495, A2 => n22013, ZN => n4380);
   U10006 : NAND2_X1 port map( A1 => n17854, A2 => n28142, ZN => n6716);
   U10010 : NAND2_X1 port map( A1 => n21645, A2 => n21642, ZN => n21399);
   U10011 : NAND3_X1 port map( A1 => n8409, A2 => n8408, A3 => n9177, ZN => 
                           n8410);
   U10013 : OAI21_X1 port map( B1 => n21304, B2 => n21150, A => n6602, ZN => 
                           n6601);
   U10014 : INV_X1 port map( A => n26990, ZN => n26323);
   U10015 : NAND2_X1 port map( A1 => n26322, A2 => n5306, ZN => n26990);
   U10016 : NAND2_X1 port map( A1 => n3269, A2 => n14193, ZN => n13868);
   U10017 : NAND3_X1 port map( A1 => n3287, A2 => n4677, A3 => n4853, ZN => 
                           n4852);
   U10019 : INV_X1 port map( A => n17822, ZN => n3875);
   U10021 : NAND2_X1 port map( A1 => n20983, A2 => n20982, ZN => n21812);
   U10022 : NOR2_X1 port map( A1 => n8014, A2 => n7742, ZN => n8019);
   U10023 : INV_X1 port map( A => n12080, ZN => n12288);
   U10025 : NAND2_X1 port map( A1 => n4278, A2 => n2023, ZN => n20289);
   U10026 : OAI21_X1 port map( B1 => n23356, B2 => n22925, A => n23461, ZN => 
                           n5269);
   U10027 : INV_X1 port map( A => n4581, ZN => n20283);
   U10028 : OAI21_X1 port map( B1 => n29183, B2 => n6203, A => n20266, ZN => 
                           n21061);
   U10029 : NAND2_X1 port map( A1 => n20451, A2 => n20647, ZN => n20266);
   U10031 : NAND2_X1 port map( A1 => n12164, A2 => n11656, ZN => n4346);
   U10035 : OR2_X1 port map( A1 => n9220, A2 => n8525, ZN => n8526);
   U10036 : INV_X1 port map( A => n5817, ZN => n20955);
   U10037 : OR2_X1 port map( A1 => n28096, A2 => n28107, ZN => n3469);
   U10038 : OAI21_X1 port map( B1 => n3270, B2 => n27984, A => n27983, ZN => 
                           n27989);
   U10039 : NAND2_X1 port map( A1 => n27981, A2 => n3271, ZN => n3270);
   U10040 : INV_X1 port map( A => n1793, ZN => n3274);
   U10041 : NAND2_X1 port map( A1 => n586, A2 => n3275, ZN => n5716);
   U10042 : AOI22_X2 port map( A1 => n18190, A2 => n16841, B1 => n16843, B2 => 
                           n16842, ZN => n19474);
   U10043 : INV_X1 port map( A => n26448, ZN => n26452);
   U10044 : XNOR2_X1 port map( A => n16646, B => n16645, ZN => n4687);
   U10045 : INV_X1 port map( A => n13914, ZN => n3798);
   U10046 : XNOR2_X1 port map( A => n10017, B => n6257, ZN => n11142);
   U10047 : INV_X1 port map( A => n15202, ZN => n15201);
   U10048 : NOR2_X1 port map( A1 => n27700, A2 => n28504, ZN => n26351);
   U10049 : XNOR2_X2 port map( A => n24931, B => n24930, ZN => n27702);
   U10050 : NAND3_X1 port map( A1 => n5494, A2 => n7890, A3 => n7774, ZN => 
                           n5493);
   U10051 : NAND2_X1 port map( A1 => n17259, A2 => n29574, ZN => n4085);
   U10052 : NAND2_X1 port map( A1 => n5133, A2 => n29209, ZN => n12024);
   U10053 : NAND2_X1 port map( A1 => n7645, A2 => n7644, ZN => n3279);
   U10054 : NOR2_X1 port map( A1 => n20587, A2 => n20585, ZN => n3974);
   U10055 : NOR2_X1 port map( A1 => n4973, A2 => n4610, ZN => n4609);
   U10056 : NAND2_X1 port map( A1 => n17797, A2 => n17639, ZN => n16841);
   U10057 : AOI21_X1 port map( B1 => n8846, B2 => n11174, A => n6289, ZN => 
                           n8847);
   U10058 : NAND3_X1 port map( A1 => n23884, A2 => n23887, A3 => n23885, ZN => 
                           n23889);
   U10060 : NAND4_X2 port map( A1 => n4911, A2 => n4909, A3 => n4910, A4 => 
                           n4912, ZN => n5953);
   U10064 : OR2_X2 port map( A1 => n7134, A2 => n7135, ZN => n8109);
   U10065 : NAND2_X1 port map( A1 => n17403, A2 => n17404, ZN => n17408);
   U10066 : XNOR2_X1 port map( A => n19606, B => n3284, ZN => n18955);
   U10067 : NAND4_X2 port map( A1 => n8068, A2 => n8067, A3 => n8066, A4 => 
                           n8065, ZN => n10144);
   U10069 : NAND2_X1 port map( A1 => n3285, A2 => n18234, ZN => n4371);
   U10071 : OR2_X1 port map( A1 => n11260, A2 => n11045, ZN => n3572);
   U10072 : INV_X1 port map( A => n5918, ZN => n13720);
   U10073 : XNOR2_X2 port map( A => Key(110), B => Plaintext(110), ZN => n8216)
                           ;
   U10074 : AOI22_X1 port map( A1 => n3286, A2 => n555, B1 => n6466, B2 => 
                           n13687, ZN => n14630);
   U10075 : NAND2_X1 port map( A1 => n13685, A2 => n13893, ZN => n3286);
   U10076 : OR2_X1 port map( A1 => n11423, A2 => n11782, ZN => n11424);
   U10078 : AND2_X1 port map( A1 => n21291, A2 => n21288, ZN => n20915);
   U10080 : NAND2_X1 port map( A1 => n3290, A2 => n3289, ZN => n17257);
   U10081 : NAND2_X1 port map( A1 => n17253, A2 => n16977, ZN => n3289);
   U10082 : NAND2_X1 port map( A1 => n17252, A2 => n16774, ZN => n3290);
   U10083 : AND2_X1 port map( A1 => n1888, A2 => n18251, ZN => n17774);
   U10084 : NAND2_X1 port map( A1 => n24975, A2 => n24258, ZN => n3291);
   U10085 : NAND2_X1 port map( A1 => n23598, A2 => n23597, ZN => n3292);
   U10086 : NAND2_X1 port map( A1 => n3294, A2 => n3293, ZN => n22176);
   U10087 : NAND2_X1 port map( A1 => n380, A2 => n23716, ZN => n3293);
   U10088 : NAND2_X1 port map( A1 => n22163, A2 => n23262, ZN => n3294);
   U10089 : INV_X1 port map( A => n18388, ZN => n5233);
   U10091 : NOR2_X2 port map( A1 => n12336, A2 => n12335, ZN => n12644);
   U10093 : OR2_X1 port map( A1 => n11113, A2 => n10490, ZN => n6241);
   U10094 : NAND2_X1 port map( A1 => n8268, A2 => n3298, ZN => n7213);
   U10095 : NAND2_X1 port map( A1 => n3299, A2 => n5888, ZN => n7226);
   U10096 : NAND2_X1 port map( A1 => n8686, A2 => n3300, ZN => n3299);
   U10097 : NAND3_X1 port map( A1 => n3302, A2 => n17458, A3 => n16810, ZN => 
                           n17461);
   U10098 : OAI21_X1 port map( B1 => n16805, B2 => n16806, A => n3303, ZN => 
                           n4914);
   U10099 : NAND2_X1 port map( A1 => n17261, A2 => n17260, ZN => n3303);
   U10100 : NAND3_X1 port map( A1 => n11111, A2 => n10492, A3 => n10461, ZN => 
                           n10462);
   U10101 : NAND2_X1 port map( A1 => n18253, A2 => n18017, ZN => n18252);
   U10102 : MUX2_X1 port map( A => n22143, B => n22142, S => n22139, Z => n3892
                           );
   U10103 : INV_X1 port map( A => n3893, ZN => n3304);
   U10104 : NAND2_X1 port map( A1 => n3894, A2 => n20580, ZN => n3305);
   U10105 : NAND3_X1 port map( A1 => n4623, A2 => n17550, A3 => n17551, ZN => 
                           n17564);
   U10106 : AND2_X1 port map( A1 => n11852, A2 => n11853, ZN => n3306);
   U10107 : AOI21_X1 port map( B1 => n10905, B2 => n11851, A => n11852, ZN => 
                           n3307);
   U10108 : OAI21_X1 port map( B1 => n12232, B2 => n1986, A => n5579, ZN => 
                           n12040);
   U10109 : OAI22_X1 port map( A1 => n5209, A2 => n18170, B1 => n18175, B2 => 
                           n28649, ZN => n18176);
   U10111 : NAND2_X1 port map( A1 => n7334, A2 => n7333, ZN => n3308);
   U10112 : NAND2_X1 port map( A1 => n27387, A2 => n27400, ZN => n27241);
   U10113 : AND2_X1 port map( A1 => n24256, A2 => n24509, ZN => n5548);
   U10114 : INV_X1 port map( A => n13979, ZN => n15113);
   U10115 : XNOR2_X1 port map( A => n1985, B => n10266, ZN => n6665);
   U10116 : NAND2_X1 port map( A1 => n5454, A2 => n3309, ZN => n24149);
   U10117 : NAND2_X1 port map( A1 => n3310, A2 => n22356, ZN => n3309);
   U10118 : OAI21_X2 port map( B1 => n412, B2 => n21006, A => n21005, ZN => 
                           n22734);
   U10119 : XNOR2_X1 port map( A => n22299, B => n22296, ZN => n6836);
   U10122 : NAND2_X1 port map( A1 => n7631, A2 => n29568, ZN => n7473);
   U10123 : OAI211_X2 port map( C1 => n19784, C2 => n21117, A => n3312, B => 
                           n3311, ZN => n22784);
   U10124 : NAND2_X1 port map( A1 => n19783, A2 => n21117, ZN => n3311);
   U10125 : NAND2_X1 port map( A1 => n19782, A2 => n21144, ZN => n3312);
   U10127 : NAND3_X1 port map( A1 => n21394, A2 => n21631, A3 => n21639, ZN => 
                           n3313);
   U10128 : NAND2_X1 port map( A1 => n3810, A2 => n7792, ZN => n7281);
   U10129 : XOR2_X1 port map( A => n19132, B => n19131, Z => n6157);
   U10130 : NAND3_X1 port map( A1 => n3320, A2 => n21716, A3 => n3319, ZN => 
                           n3318);
   U10131 : INV_X1 port map( A => n21263, ZN => n3320);
   U10133 : NAND2_X1 port map( A1 => n12363, A2 => n12359, ZN => n10611);
   U10134 : NAND2_X1 port map( A1 => n14204, A2 => n427, ZN => n13684);
   U10136 : NAND2_X1 port map( A1 => n12144, A2 => n11712, ZN => n11710);
   U10137 : NAND2_X1 port map( A1 => n11715, A2 => n12146, ZN => n12144);
   U10138 : NAND2_X1 port map( A1 => n409, A2 => n23251, ZN => n5322);
   U10140 : NAND2_X1 port map( A1 => n11262, A2 => n11266, ZN => n3325);
   U10142 : OAI21_X1 port map( B1 => n10993, B2 => n10785, A => n3328, ZN => 
                           n10996);
   U10143 : NAND2_X1 port map( A1 => n10993, A2 => n10992, ZN => n3328);
   U10144 : NAND2_X1 port map( A1 => n7630, A2 => n7633, ZN => n3330);
   U10145 : NAND2_X1 port map( A1 => n7632, A2 => n7914, ZN => n3331);
   U10146 : NAND2_X1 port map( A1 => n28660, A2 => n28545, ZN => n3332);
   U10148 : MUX2_X1 port map( A => n20743, B => n3335, S => n20857, Z => n20748
                           );
   U10149 : NOR2_X1 port map( A1 => n21155, A2 => n20744, ZN => n3335);
   U10150 : XNOR2_X1 port map( A => n3338, B => n22408, ZN => n23049);
   U10151 : NAND2_X1 port map( A1 => n3339, A2 => n20121, ZN => n18118);
   U10152 : NAND2_X1 port map( A1 => n20202, A2 => n20201, ZN => n3339);
   U10154 : OAI21_X1 port map( B1 => n8245, B2 => n7818, A => n3340, ZN => 
                           n7819);
   U10155 : NAND2_X1 port map( A1 => n8245, A2 => n7817, ZN => n3340);
   U10156 : MUX2_X1 port map( A => n29565, B => n14166, S => n29306, Z => n6143
                           );
   U10158 : INV_X1 port map( A => n12868, ZN => n12396);
   U10160 : NOR2_X1 port map( A1 => n23790, A2 => n23789, ZN => n5770);
   U10161 : INV_X1 port map( A => n5887, ZN => n5847);
   U10162 : AND2_X1 port map( A1 => n17030, A2 => n17357, ZN => n17031);
   U10163 : NAND2_X1 port map( A1 => n14693, A2 => n16995, ZN => n3342);
   U10165 : INV_X1 port map( A => n11288, ZN => n10665);
   U10166 : XNOR2_X1 port map( A => n13054, B => n13159, ZN => n13353);
   U10167 : NAND2_X1 port map( A1 => n3345, A2 => n14689, ZN => n3344);
   U10168 : NAND2_X1 port map( A1 => n13985, A2 => n551, ZN => n3345);
   U10169 : NAND2_X1 port map( A1 => n18588, A2 => n18589, ZN => n18590);
   U10170 : NAND2_X1 port map( A1 => n1835, A2 => n19955, ZN => n20112);
   U10171 : OAI211_X1 port map( C1 => n17948, C2 => n18342, A => n18344, B => 
                           n3347, ZN => n5771);
   U10172 : NAND2_X1 port map( A1 => n17663, A2 => n18342, ZN => n3347);
   U10173 : OAI211_X2 port map( C1 => n29227, C2 => n21281, A => n20994, B => 
                           n20993, ZN => n22856);
   U10174 : OAI211_X1 port map( C1 => n19032, C2 => n20476, A => n20478, B => 
                           n4556, ZN => n6451);
   U10175 : AOI21_X1 port map( B1 => n23682, B2 => n23679, A => n5882, ZN => 
                           n5881);
   U10176 : NAND2_X1 port map( A1 => n20517, A2 => n21356, ZN => n20262);
   U10177 : NAND2_X1 port map( A1 => n14132, A2 => n14342, ZN => n3348);
   U10179 : XNOR2_X1 port map( A => n19422, B => n19420, ZN => n5809);
   U10180 : XNOR2_X1 port map( A => n16229, B => n4029, ZN => n16231);
   U10181 : NAND2_X1 port map( A1 => n5535, A2 => n28649, ZN => n3350);
   U10182 : NAND2_X1 port map( A1 => n27980, A2 => n28456, ZN => n27981);
   U10183 : AND2_X2 port map( A1 => n3352, A2 => n3351, ZN => n27908);
   U10184 : NAND2_X1 port map( A1 => n27054, A2 => n27053, ZN => n3352);
   U10186 : OAI21_X1 port map( B1 => n9031, B2 => n8433, A => n3353, ZN => 
                           n8435);
   U10188 : INV_X1 port map( A => n16960, ZN => n5327);
   U10189 : NOR2_X1 port map( A1 => n14763, A2 => n15054, ZN => n6393);
   U10191 : OAI21_X1 port map( B1 => n8651, B2 => n8635, A => n3354, ZN => 
                           n8660);
   U10192 : NAND2_X1 port map( A1 => n8651, A2 => n8652, ZN => n3354);
   U10194 : AND2_X1 port map( A1 => n24772, A2 => n24697, ZN => n24699);
   U10196 : NAND2_X1 port map( A1 => n13620, A2 => n14082, ZN => n3356);
   U10197 : NAND2_X1 port map( A1 => n13621, A2 => n28625, ZN => n3357);
   U10202 : NAND2_X1 port map( A1 => n3362, A2 => n15407, ZN => n3361);
   U10203 : XNOR2_X1 port map( A => n18998, B => n19236, ZN => n19001);
   U10204 : XNOR2_X1 port map( A => n19468, B => n19555, ZN => n19236);
   U10205 : OAI22_X1 port map( A1 => n17757, A2 => n522, B1 => n17966, B2 => 
                           n18240, ZN => n17537);
   U10206 : NAND2_X1 port map( A1 => n11969, A2 => n12158, ZN => n10861);
   U10209 : INV_X1 port map( A => n27632, ZN => n3366);
   U10210 : NAND2_X1 port map( A1 => n1912, A2 => n27625, ZN => n3367);
   U10211 : OAI21_X1 port map( B1 => n11322, B2 => n11321, A => n29316, ZN => 
                           n6722);
   U10215 : INV_X1 port map( A => n7705, ZN => n3639);
   U10216 : NAND2_X1 port map( A1 => n7959, A2 => n7958, ZN => n3368);
   U10217 : NAND3_X1 port map( A1 => n3370, A2 => n6273, A3 => n6274, ZN => 
                           n22919);
   U10218 : OAI211_X1 port map( C1 => n21012, C2 => n21442, A => n3371, B => 
                           n21656, ZN => n3370);
   U10219 : NAND2_X1 port map( A1 => n21660, A2 => n20833, ZN => n3371);
   U10220 : INV_X1 port map( A => n14393, ZN => n13951);
   U10221 : OAI211_X1 port map( C1 => n28157, C2 => n581, A => n10751, B => 
                           n11197, ZN => n3373);
   U10222 : NAND2_X1 port map( A1 => n20587, A2 => n20585, ZN => n17880);
   U10223 : AND2_X1 port map( A1 => n14358, A2 => n4166, ZN => n3375);
   U10224 : NAND2_X1 port map( A1 => n6314, A2 => n29101, ZN => n21697);
   U10226 : INV_X1 port map( A => n4364, ZN => n24630);
   U10227 : INV_X1 port map( A => n17834, ZN => n18588);
   U10228 : INV_X1 port map( A => n23535, ZN => n23694);
   U10229 : MUX2_X1 port map( A => n26265, B => n26264, S => n28392, Z => n3376
                           );
   U10230 : OAI21_X1 port map( B1 => n8765, B2 => n9561, A => n3377, ZN => 
                           n8332);
   U10231 : NAND2_X1 port map( A1 => n8765, A2 => n8944, ZN => n3377);
   U10232 : NAND2_X1 port map( A1 => n4885, A2 => n4886, ZN => n4888);
   U10233 : XNOR2_X1 port map( A => n12955, B => n3382, ZN => n6831);
   U10234 : OAI21_X2 port map( B1 => n17292, B2 => n17291, A => n17295, ZN => 
                           n18033);
   U10236 : OAI21_X1 port map( B1 => n11767, B2 => n4197, A => n3383, ZN => 
                           n5019);
   U10237 : NAND2_X1 port map( A1 => n3384, A2 => n4197, ZN => n3383);
   U10238 : INV_X1 port map( A => n12305, ZN => n3384);
   U10239 : NAND2_X1 port map( A1 => n7589, A2 => n7233, ZN => n7869);
   U10240 : NAND2_X1 port map( A1 => n12976, A2 => n14091, ZN => n14092);
   U10241 : AND2_X1 port map( A1 => n20178, A2 => n20173, ZN => n19055);
   U10242 : NAND2_X1 port map( A1 => n18344, A2 => n18341, ZN => n18340);
   U10243 : NAND2_X1 port map( A1 => n3387, A2 => n20091, ZN => n20094);
   U10244 : NOR2_X1 port map( A1 => n20041, A2 => n20093, ZN => n3387);
   U10245 : XNOR2_X1 port map( A => n21756, B => n1271, ZN => n6074);
   U10248 : NAND2_X1 port map( A1 => n7978, A2 => n7979, ZN => n8073);
   U10249 : NAND3_X1 port map( A1 => n8730, A2 => n8731, A3 => n8381, ZN => 
                           n7186);
   U10251 : NAND2_X1 port map( A1 => n4916, A2 => n23447, ZN => n3391);
   U10252 : NAND2_X1 port map( A1 => n4915, A2 => n23371, ZN => n3392);
   U10253 : NAND2_X1 port map( A1 => n14064, A2 => n13652, ZN => n3393);
   U10254 : NAND2_X1 port map( A1 => n16788, A2 => n6002, ZN => n5068);
   U10256 : NAND2_X1 port map( A1 => n3396, A2 => n14264, ZN => n3395);
   U10257 : INV_X1 port map( A => n14259, ZN => n3396);
   U10258 : NAND3_X1 port map( A1 => n29132, A2 => n28536, A3 => n27177, ZN => 
                           n3397);
   U10260 : OAI21_X2 port map( B1 => n22741, B2 => n23445, A => n22740, ZN => 
                           n24552);
   U10261 : NAND2_X1 port map( A1 => n6541, A2 => n26800, ZN => n6323);
   U10262 : NAND3_X1 port map( A1 => n21158, A2 => n20744, A3 => n3401, ZN => 
                           n3400);
   U10264 : INV_X1 port map( A => n15895, ZN => n5447);
   U10265 : NAND2_X2 port map( A1 => n4239, A2 => n4238, ZN => n25836);
   U10266 : AOI21_X1 port map( B1 => n5028, B2 => n23137, A => n23694, ZN => 
                           n3405);
   U10267 : XNOR2_X1 port map( A => n3406, B => n16343, ZN => n15931);
   U10268 : XNOR2_X1 port map( A => n15926, B => n15925, ZN => n3406);
   U10269 : NAND2_X1 port map( A1 => n3409, A2 => n3408, ZN => n13743);
   U10270 : NAND2_X1 port map( A1 => n13742, A2 => n29306, ZN => n3409);
   U10272 : OAI21_X1 port map( B1 => n11852, B2 => n574, A => n3410, ZN => 
                           n10908);
   U10273 : INV_X1 port map( A => n4460, ZN => n20830);
   U10274 : NAND2_X1 port map( A1 => n20068, A2 => n20065, ZN => n3411);
   U10275 : OAI211_X1 port map( C1 => n10780, C2 => n28173, A => n3413, B => 
                           n10959, ZN => n6773);
   U10276 : AOI21_X1 port map( B1 => n24706, B2 => n29043, A => n6612, ZN => 
                           n6611);
   U10277 : XOR2_X1 port map( A => n10295, B => n9613, Z => n5032);
   U10278 : XNOR2_X1 port map( A => n25790, B => n25543, ZN => n25260);
   U10279 : INV_X1 port map( A => n4180, ZN => n4179);
   U10280 : OAI21_X1 port map( B1 => n8924, B2 => n9132, A => n9131, ZN => 
                           n9136);
   U10281 : INV_X1 port map( A => n15535, ZN => n16653);
   U10282 : INV_X1 port map( A => n17276, ZN => n16844);
   U10284 : OR2_X1 port map( A1 => n9024, A2 => n8687, ZN => n5889);
   U10286 : XNOR2_X1 port map( A => n25937, B => n25936, ZN => n27056);
   U10288 : NAND2_X1 port map( A1 => n16819, A2 => n387, ZN => n3415);
   U10289 : NAND2_X1 port map( A1 => n16820, A2 => n17463, ZN => n3416);
   U10290 : NOR2_X1 port map( A1 => n16673, A2 => n17464, ZN => n16820);
   U10292 : AND2_X1 port map( A1 => n18383, A2 => n18379, ZN => n5670);
   U10293 : XNOR2_X1 port map( A => n12830, B => n13371, ZN => n13479);
   U10295 : NAND2_X1 port map( A1 => n13411, A2 => n2075, ZN => n14881);
   U10297 : NAND2_X1 port map( A1 => n3417, A2 => n21394, ZN => n21228);
   U10298 : NAND2_X1 port map( A1 => n21226, A2 => n3418, ZN => n3417);
   U10301 : OR2_X1 port map( A1 => n20720, A2 => n21596, ZN => n20723);
   U10302 : OAI21_X1 port map( B1 => n3421, B2 => n19890, A => n3420, ZN => 
                           n19894);
   U10303 : NAND2_X1 port map( A1 => n19890, A2 => n28894, ZN => n3420);
   U10304 : INV_X1 port map( A => n14039, ZN => n13997);
   U10305 : INV_X1 port map( A => n14971, ZN => n5813);
   U10306 : NOR2_X1 port map( A1 => n20700, A2 => n21691, ZN => n6313);
   U10307 : NOR2_X1 port map( A1 => n10818, A2 => n10817, ZN => n11646);
   U10308 : INV_X1 port map( A => n14923, ZN => n15498);
   U10309 : INV_X1 port map( A => n21227, ZN => n21633);
   U10310 : XNOR2_X1 port map( A => n12421, B => n12652, ZN => n11866);
   U10312 : INV_X1 port map( A => n21632, ZN => n21637);
   U10313 : XNOR2_X1 port map( A => n22657, B => n6863, ZN => n20277);
   U10314 : XNOR2_X1 port map( A => n19408, B => n16990, ZN => n19590);
   U10315 : NAND2_X1 port map( A1 => n3427, A2 => n3424, ZN => n27437);
   U10316 : NAND3_X1 port map( A1 => n3426, A2 => n3425, A3 => n26710, ZN => 
                           n3424);
   U10317 : NAND2_X1 port map( A1 => n27442, A2 => n27433, ZN => n3425);
   U10318 : INV_X1 port map( A => n27432, ZN => n3426);
   U10319 : NAND2_X1 port map( A1 => n27435, A2 => n27434, ZN => n3427);
   U10320 : NAND2_X1 port map( A1 => n8201, A2 => n3431, ZN => n3430);
   U10321 : NAND3_X1 port map( A1 => n3433, A2 => n3748, A3 => n14917, ZN => 
                           n14503);
   U10322 : NAND2_X1 port map( A1 => n14703, A2 => n15489, ZN => n3433);
   U10323 : AOI22_X1 port map( A1 => n17108, A2 => n17472, B1 => n17107, B2 => 
                           n17470, ZN => n17112);
   U10324 : OAI21_X1 port map( B1 => n23169, B2 => n23516, A => n3434, ZN => 
                           n23521);
   U10326 : NAND2_X1 port map( A1 => n15308, A2 => n15309, ZN => n15271);
   U10328 : NAND3_X1 port map( A1 => n14086, A2 => n14088, A3 => n14087, ZN => 
                           n14089);
   U10329 : AND2_X1 port map( A1 => n12271, A2 => n12270, ZN => n11103);
   U10330 : INV_X1 port map( A => n24460, ZN => n5004);
   U10332 : OAI211_X2 port map( C1 => n6671, C2 => n3849, A => n6670, B => 
                           n18457, ZN => n19595);
   U10333 : XNOR2_X1 port map( A => n9351, B => n10188, ZN => n3437);
   U10334 : NAND2_X1 port map( A1 => n3438, A2 => n11707, ZN => n12495);
   U10336 : NAND2_X1 port map( A1 => n29559, A2 => n17283, ZN => n16066);
   U10337 : NAND2_X1 port map( A1 => n20571, A2 => n20568, ZN => n3443);
   U10338 : AND2_X2 port map( A1 => n6215, A2 => n2065, ZN => n24852);
   U10339 : NAND2_X1 port map( A1 => n8206, A2 => n3446, ZN => n8836);
   U10340 : OAI211_X1 port map( C1 => n8199, C2 => n28605, A => n3448, B => 
                           n3447, ZN => n3446);
   U10341 : NAND2_X1 port map( A1 => n8199, A2 => n8201, ZN => n3448);
   U10343 : NAND3_X1 port map( A1 => n6359, A2 => n6360, A3 => n10742, ZN => 
                           n3449);
   U10344 : NAND2_X1 port map( A1 => n28205, A2 => n10461, ZN => n10099);
   U10345 : MUX2_X2 port map( A => n14152, B => n14151, S => n14380, Z => 
                           n15359);
   U10346 : NAND3_X1 port map( A1 => n21589, A2 => n20714, A3 => n5683, ZN => 
                           n5206);
   U10348 : INV_X1 port map( A => n11751, ZN => n4712);
   U10349 : NAND2_X1 port map( A1 => n6439, A2 => n23429, ZN => n23599);
   U10350 : INV_X1 port map( A => n10971, ZN => n5267);
   U10351 : XNOR2_X1 port map( A => n3452, B => n9295, ZN => n10338);
   U10352 : XNOR2_X1 port map( A => n18727, B => n1981, ZN => n5586);
   U10353 : NAND2_X1 port map( A1 => n10994, A2 => n3454, ZN => n3453);
   U10354 : OAI22_X1 port map( A1 => n10501, A2 => n10497, B1 => n11132, B2 => 
                           n10500, ZN => n3458);
   U10355 : NAND2_X1 port map( A1 => n21193, A2 => n6936, ZN => n21197);
   U10356 : NAND2_X1 port map( A1 => n11677, A2 => n11676, ZN => n11678);
   U10357 : NAND2_X1 port map( A1 => n21551, A2 => n21519, ZN => n21552);
   U10358 : NAND2_X1 port map( A1 => n15265, A2 => n14923, ZN => n15266);
   U10361 : MUX2_X2 port map( A => n18250, B => n18249, S => n28558, Z => 
                           n19496);
   U10362 : NAND2_X1 port map( A1 => n11403, A2 => n11118, ZN => n3461);
   U10363 : NAND3_X2 port map( A1 => n9777, A2 => n9778, A3 => n11234, ZN => 
                           n12189);
   U10364 : MUX2_X2 port map( A => n19775, B => n19774, S => n20098, Z => 
                           n21119);
   U10365 : NOR2_X2 port map( A1 => n4393, A2 => n21147, ZN => n22059);
   U10366 : INV_X1 port map( A => n14366, ZN => n14094);
   U10367 : AOI22_X1 port map( A1 => n28179, A2 => n28429, B1 => n27585, B2 => 
                           n27596, ZN => n27598);
   U10368 : INV_X1 port map( A => n7641, ZN => n7457);
   U10369 : XNOR2_X1 port map( A => n16203, B => n16202, ZN => n6870);
   U10370 : NAND2_X1 port map( A1 => n7886, A2 => n7583, ZN => n7882);
   U10371 : NAND2_X1 port map( A1 => n7580, A2 => n7582, ZN => n3464);
   U10372 : OR2_X1 port map( A1 => n18688, A2 => n18687, ZN => n18703);
   U10373 : NOR2_X1 port map( A1 => n6077, A2 => n18473, ZN => n6076);
   U10375 : NAND3_X1 port map( A1 => n28489, A2 => n20511, A3 => n19785, ZN => 
                           n4912);
   U10376 : INV_X1 port map( A => n26733, ZN => n5389);
   U10377 : NAND2_X1 port map( A1 => n23318, A2 => n23648, ZN => n23192);
   U10378 : NAND2_X1 port map( A1 => n18151, A2 => n3467, ZN => n3466);
   U10379 : INV_X1 port map( A => n18149, ZN => n3467);
   U10380 : INV_X1 port map( A => n23290, ZN => n5591);
   U10381 : INV_X1 port map( A => n24380, ZN => n23906);
   U10382 : NAND2_X1 port map( A1 => n17097, A2 => n17098, ZN => n17099);
   U10383 : NAND2_X1 port map( A1 => n28094, A2 => n28107, ZN => n3470);
   U10384 : NAND2_X1 port map( A1 => n24737, A2 => n24738, ZN => n24742);
   U10386 : NAND3_X1 port map( A1 => n4391, A2 => n18135, A3 => n3471, ZN => 
                           n17636);
   U10387 : NAND2_X1 port map( A1 => n21668, A2 => n4312, ZN => n3474);
   U10388 : NAND2_X1 port map( A1 => n21667, A2 => n22404, ZN => n3475);
   U10389 : NAND2_X1 port map( A1 => n3477, A2 => n18430, ZN => n18436);
   U10390 : NAND2_X1 port map( A1 => n18429, A2 => n4762, ZN => n3477);
   U10391 : NAND2_X1 port map( A1 => n2855, A2 => n18433, ZN => n18429);
   U10392 : XNOR2_X1 port map( A => n3478, B => n27453, ZN => Ciphertext(42));
   U10393 : NAND4_X1 port map( A1 => n27450, A2 => n27451, A3 => n27448, A4 => 
                           n27449, ZN => n3478);
   U10394 : NAND2_X1 port map( A1 => n10742, A2 => n10808, ZN => n7814);
   U10395 : OAI22_X1 port map( A1 => n18887, A2 => n20150, B1 => n20099, B2 => 
                           n20098, ZN => n20156);
   U10396 : NAND2_X1 port map( A1 => n3479, A2 => n5599, ZN => n5596);
   U10397 : NAND2_X1 port map( A1 => n5597, A2 => n14551, ZN => n3479);
   U10398 : NAND2_X1 port map( A1 => n11283, A2 => n1854, ZN => n11285);
   U10399 : INV_X1 port map( A => n21425, ZN => n21085);
   U10400 : INV_X1 port map( A => n21494, ZN => n20867);
   U10401 : OAI22_X1 port map( A1 => n4025, A2 => n3480, B1 => n6406, B2 => 
                           n24324, ZN => n24326);
   U10402 : NAND2_X1 port map( A1 => n18425, A2 => n18426, ZN => n18427);
   U10403 : NOR2_X1 port map( A1 => n15389, A2 => n6517, ZN => n14631);
   U10404 : NAND2_X1 port map( A1 => n5557, A2 => n17301, ZN => n15812);
   U10405 : NOR2_X2 port map( A1 => n14666, A2 => n14660, ZN => n15444);
   U10406 : NAND2_X1 port map( A1 => n17299, A2 => n17415, ZN => n3484);
   U10410 : NAND2_X1 port map( A1 => n20946, A2 => n20945, ZN => n5879);
   U10411 : INV_X1 port map( A => n20557, ZN => n20548);
   U10412 : NAND2_X1 port map( A1 => n17172, A2 => n28501, ZN => n20557);
   U10413 : NAND3_X1 port map( A1 => n14069, A2 => n14070, A3 => n6351, ZN => 
                           n3488);
   U10414 : NAND2_X1 port map( A1 => n21258, A2 => n21714, ZN => n20977);
   U10415 : NAND2_X1 port map( A1 => n7466, A2 => n28615, ZN => n3489);
   U10416 : NAND2_X1 port map( A1 => n6782, A2 => n6783, ZN => n3490);
   U10417 : NAND2_X1 port map( A1 => n21716, A2 => n21368, ZN => n3492);
   U10419 : NAND3_X1 port map( A1 => n5072, A2 => n7519, A3 => n7518, ZN => 
                           n8592);
   U10420 : NAND2_X1 port map( A1 => n3496, A2 => n3495, ZN => n24001);
   U10421 : OR2_X1 port map( A1 => n22951, A2 => n23397, ZN => n3495);
   U10422 : OAI21_X1 port map( B1 => n23401, B2 => n22950, A => n23227, ZN => 
                           n3496);
   U10423 : OAI211_X1 port map( C1 => n29467, C2 => n3498, A => n26456, B => 
                           n3497, ZN => n6736);
   U10425 : NAND3_X1 port map( A1 => n23512, A2 => n23772, A3 => n23487, ZN => 
                           n3499);
   U10426 : NAND2_X1 port map( A1 => n3500, A2 => n12205, ZN => n11440);
   U10427 : NAND2_X1 port map( A1 => n11438, A2 => n11599, ZN => n3500);
   U10429 : OR3_X1 port map( A1 => n15290, A2 => n15217, A3 => n15036, ZN => 
                           n15219);
   U10430 : OR2_X1 port map( A1 => n4451, A2 => n14085, ZN => n14086);
   U10431 : OR2_X1 port map( A1 => n25239, A2 => n27395, ZN => n25241);
   U10432 : OR2_X1 port map( A1 => n14688, A2 => n15004, ZN => n4689);
   U10433 : NAND2_X1 port map( A1 => n20635, A2 => n20247, ZN => n3503);
   U10434 : NAND2_X1 port map( A1 => n498, A2 => n20632, ZN => n3504);
   U10435 : INV_X1 port map( A => n17772, ZN => n18018);
   U10436 : NOR2_X1 port map( A1 => n18120, A2 => n4240, ZN => n17821);
   U10437 : NAND3_X1 port map( A1 => n23263, A2 => n23713, A3 => n3505, ZN => 
                           n23264);
   U10438 : OAI21_X1 port map( B1 => n380, B2 => n23710, A => n23262, ZN => 
                           n3505);
   U10439 : NOR2_X1 port map( A1 => n26463, A2 => n2015, ZN => n26471);
   U10440 : NAND2_X1 port map( A1 => n545, A2 => n15464, ZN => n3506);
   U10441 : NAND2_X1 port map( A1 => n15159, A2 => n29153, ZN => n3507);
   U10442 : OAI21_X2 port map( B1 => n19677, B2 => n19808, A => n19676, ZN => 
                           n19732);
   U10443 : NAND2_X1 port map( A1 => n9095, A2 => n8666, ZN => n8631);
   U10444 : AOI21_X1 port map( B1 => n7231, B2 => n441, A => n7957, ZN => n7961
                           );
   U10445 : AOI21_X1 port map( B1 => n3511, B2 => n3510, A => n7692, ZN => 
                           n7694);
   U10446 : NAND2_X1 port map( A1 => n24064, A2 => n28415, ZN => n3512);
   U10447 : NAND2_X1 port map( A1 => n23269, A2 => n24138, ZN => n3514);
   U10448 : NAND2_X1 port map( A1 => n4611, A2 => n15251, ZN => n15253);
   U10449 : OAI21_X1 port map( B1 => n21192, B2 => n28611, A => n3515, ZN => 
                           n21544);
   U10450 : NAND2_X1 port map( A1 => n28611, A2 => n21539, ZN => n3515);
   U10451 : NOR2_X1 port map( A1 => n28088, A2 => n3517, ZN => Ciphertext(188))
                           ;
   U10453 : INV_X1 port map( A => n18136, ZN => n5623);
   U10454 : NOR2_X1 port map( A1 => n14752, A2 => n14153, ZN => n15358);
   U10456 : AOI21_X1 port map( B1 => n407, B2 => n28609, A => n23816, ZN => 
                           n3518);
   U10457 : OAI21_X1 port map( B1 => n17425, B2 => n2826, A => n3520, ZN => 
                           n17432);
   U10458 : NAND2_X1 port map( A1 => n17425, A2 => n5891, ZN => n3520);
   U10459 : INV_X1 port map( A => n23773, ZN => n6424);
   U10460 : OAI21_X1 port map( B1 => n11549, B2 => n574, A => n3521, ZN => 
                           n10094);
   U10461 : NAND2_X1 port map( A1 => n17598, A2 => n28558, ZN => n3523);
   U10462 : NAND2_X1 port map( A1 => n17599, A2 => n5021, ZN => n3524);
   U10463 : NAND2_X1 port map( A1 => n17600, A2 => n18709, ZN => n3525);
   U10464 : NAND2_X1 port map( A1 => n1320, A2 => n3526, ZN => n5642);
   U10465 : OR2_X1 port map( A1 => n16878, A2 => n16700, ZN => n17159);
   U10466 : INV_X1 port map( A => n14174, ZN => n15195);
   U10467 : OAI21_X1 port map( B1 => n20623, B2 => n20626, A => n20628, ZN => 
                           n5318);
   U10468 : INV_X1 port map( A => n8808, ZN => n8681);
   U10469 : XNOR2_X1 port map( A => n5984, B => n10150, ZN => n10155);
   U10470 : XNOR2_X1 port map( A => n22500, B => n26032, ZN => n5718);
   U10471 : NAND2_X1 port map( A1 => n5918, A2 => n14039, ZN => n6032);
   U10473 : AOI22_X1 port map( A1 => n17270, A2 => n17265, B1 => n17269, B2 => 
                           n17268, ZN => n17534);
   U10475 : NAND2_X1 port map( A1 => n10515, A2 => n10516, ZN => n12529);
   U10476 : NAND4_X2 port map( A1 => n11306, A2 => n11305, A3 => n11304, A4 => 
                           n11303, ZN => n13075);
   U10479 : OR2_X1 port map( A1 => n10585, A2 => n3802, ZN => n3533);
   U10480 : NAND2_X1 port map( A1 => n1941, A2 => n2026, ZN => n3534);
   U10481 : NAND2_X1 port map( A1 => n16701, A2 => n29045, ZN => n3535);
   U10482 : NAND2_X1 port map( A1 => n10823, A2 => n3536, ZN => n10822);
   U10483 : NAND2_X1 port map( A1 => n8688, A2 => n8687, ZN => n9227);
   U10484 : NAND2_X1 port map( A1 => n17730, A2 => n18455, ZN => n3538);
   U10485 : NAND2_X1 port map( A1 => n17731, A2 => n18107, ZN => n3539);
   U10486 : AND2_X1 port map( A1 => n29641, A2 => n23772, ZN => n21862);
   U10487 : NAND2_X1 port map( A1 => n3540, A2 => n17721, ZN => n17723);
   U10488 : NAND2_X1 port map( A1 => n4621, A2 => n14116, ZN => n4620);
   U10491 : OR2_X2 port map( A1 => n7356, A2 => n7355, ZN => n10193);
   U10492 : XOR2_X1 port map( A => n9388, B => n9387, Z => n4716);
   U10493 : AND2_X2 port map( A1 => n20776, A2 => n20777, ZN => n21500);
   U10494 : NAND3_X2 port map( A1 => n6660, A2 => n6659, A3 => n11539, ZN => 
                           n12830);
   U10495 : XNOR2_X2 port map( A => n5924, B => n5925, ZN => n10808);
   U10496 : AOI21_X1 port map( B1 => n3543, B2 => n11740, A => n12363, ZN => 
                           n10615);
   U10497 : NAND2_X1 port map( A1 => n11739, A2 => n12356, ZN => n3543);
   U10498 : NAND2_X1 port map( A1 => n11708, A2 => n11648, ZN => n11416);
   U10499 : NAND2_X1 port map( A1 => n3546, A2 => n3545, ZN => n14597);
   U10500 : NAND2_X1 port map( A1 => n14256, A2 => n14255, ZN => n3545);
   U10501 : NAND2_X1 port map( A1 => n14257, A2 => n14254, ZN => n3546);
   U10502 : NAND2_X1 port map( A1 => n10553, A2 => n10554, ZN => n10555);
   U10503 : NAND2_X1 port map( A1 => n10804, A2 => n10752, ZN => n10553);
   U10505 : NAND3_X1 port map( A1 => n22291, A2 => n29364, A3 => n3548, ZN => 
                           n21055);
   U10507 : NAND3_X1 port map( A1 => n29624, A2 => n24769, A3 => n24768, ZN => 
                           n24770);
   U10508 : XNOR2_X1 port map( A => n5452, B => n5453, ZN => n23353);
   U10509 : OR2_X1 port map( A1 => n20300, A2 => n6843, ZN => n3551);
   U10510 : NOR2_X1 port map( A1 => n8932, A2 => n6072, ZN => n8933);
   U10511 : OAI211_X1 port map( C1 => n20552, C2 => n6086, A => n20553, B => 
                           n6085, ZN => n6084);
   U10512 : INV_X1 port map( A => n349, ZN => n3552);
   U10513 : OR2_X1 port map( A1 => n17989, A2 => n28142, ZN => n17014);
   U10514 : AND2_X1 port map( A1 => n7864, A2 => n7092, ZN => n5191);
   U10515 : INV_X1 port map( A => n4193, ZN => n21458);
   U10516 : NOR2_X1 port map( A1 => n23303, A2 => n5530, ZN => n23105);
   U10517 : INV_X1 port map( A => n17568, ZN => n4118);
   U10520 : OAI21_X1 port map( B1 => n20844, B2 => n20843, A => n4193, ZN => 
                           n3555);
   U10522 : OR2_X1 port map( A1 => n14517, A2 => n15292, ZN => n15216);
   U10523 : NAND2_X1 port map( A1 => n12062, A2 => n3557, ZN => n3556);
   U10524 : NAND2_X1 port map( A1 => n8553, A2 => n8762, ZN => n8764);
   U10525 : NAND2_X1 port map( A1 => n20955, A2 => n20802, ZN => n3559);
   U10528 : XNOR2_X1 port map( A => n9927, B => n9926, ZN => n10097);
   U10529 : NOR2_X2 port map( A1 => n7693, A2 => n7694, ZN => n9030);
   U10530 : NAND2_X1 port map( A1 => n23319, A2 => n23493, ZN => n23323);
   U10531 : NAND2_X1 port map( A1 => n21569, A2 => n21570, ZN => n3563);
   U10532 : NAND2_X1 port map( A1 => n20314, A2 => n20585, ZN => n19828);
   U10534 : NAND2_X1 port map( A1 => n4345, A2 => n12163, ZN => n3566);
   U10535 : NAND2_X1 port map( A1 => n14846, A2 => n14845, ZN => n14847);
   U10536 : AOI21_X1 port map( B1 => n24120, B2 => n24121, A => n403, ZN => 
                           n3567);
   U10537 : AOI22_X1 port map( A1 => n11978, A2 => n11977, B1 => n6871, B2 => 
                           n28201, ZN => n4261);
   U10538 : NAND2_X1 port map( A1 => n28201, A2 => n12234, ZN => n11977);
   U10539 : OR2_X1 port map( A1 => n20047, A2 => n28187, ZN => n19987);
   U10543 : INV_X1 port map( A => n15998, ZN => n16177);
   U10544 : NAND2_X1 port map( A1 => n23979, A2 => n28519, ZN => n23980);
   U10545 : XNOR2_X1 port map( A => n21998, B => n21728, ZN => n22246);
   U10547 : NAND2_X1 port map( A1 => n18224, A2 => n17532, ZN => n18387);
   U10549 : XNOR2_X1 port map( A => n10030, B => n10027, ZN => n5400);
   U10550 : INV_X1 port map( A => n22256, ZN => n6378);
   U10551 : INV_X1 port map( A => n21457, ZN => n21125);
   U10553 : NAND2_X1 port map( A1 => n28438, A2 => n27944, ZN => n3571);
   U10554 : AOI21_X2 port map( B1 => n18310, B2 => n18309, A => n18308, ZN => 
                           n19688);
   U10555 : MUX2_X2 port map( A => n15768, B => n15767, S => n17560, Z => 
                           n18063);
   U10556 : NOR2_X1 port map( A1 => n3572, A2 => n6515, ZN => n6514);
   U10557 : NAND2_X1 port map( A1 => n3573, A2 => n4995, ZN => n23992);
   U10558 : NAND2_X1 port map( A1 => n4993, A2 => n24634, ZN => n3573);
   U10559 : XNOR2_X1 port map( A => n11805, B => n11804, ZN => n13744);
   U10561 : NAND2_X1 port map( A1 => n14792, A2 => n14881, ZN => n14584);
   U10562 : OAI21_X2 port map( B1 => n22961, B2 => n28418, A => n22960, ZN => 
                           n24020);
   U10563 : INV_X1 port map( A => n3575, ZN => n3574);
   U10564 : OAI21_X1 port map( B1 => n14765, B2 => n15262, A => n3576, ZN => 
                           n3575);
   U10565 : NAND2_X1 port map( A1 => n6393, A2 => n15053, ZN => n3576);
   U10566 : NAND2_X1 port map( A1 => n14764, A2 => n15056, ZN => n3577);
   U10569 : OAI21_X1 port map( B1 => n17067, B2 => n17066, A => n17065, ZN => 
                           n4831);
   U10570 : OR2_X1 port map( A1 => n11188, A2 => n11187, ZN => n3905);
   U10571 : NAND2_X1 port map( A1 => n12714, A2 => n4290, ZN => n3579);
   U10572 : INV_X1 port map( A => n14460, ZN => n3580);
   U10573 : NAND2_X1 port map( A1 => n12713, A2 => n14460, ZN => n3581);
   U10574 : XNOR2_X1 port map( A => n15634, B => n16131, ZN => n15635);
   U10575 : XNOR2_X1 port map( A => n16166, B => n16167, ZN => n3582);
   U10576 : OR2_X1 port map( A1 => n15420, A2 => n15101, ZN => n4547);
   U10577 : INV_X1 port map( A => n14451, ZN => n14181);
   U10578 : INV_X1 port map( A => n13118, ZN => n12637);
   U10579 : INV_X1 port map( A => n29145, ZN => n3735);
   U10581 : XNOR2_X1 port map( A => n13104, B => n13552, ZN => n6375);
   U10582 : NAND3_X1 port map( A1 => n23286, A2 => n5763, A3 => n23075, ZN => 
                           n23076);
   U10583 : AOI22_X1 port map( A1 => n5575, A2 => n6699, B1 => n15499, B2 => 
                           n14431, ZN => n3583);
   U10584 : NAND2_X1 port map( A1 => n11197, A2 => n10814, ZN => n3584);
   U10585 : NOR2_X1 port map( A1 => n17475, A2 => n3883, ZN => n4367);
   U10588 : NAND2_X1 port map( A1 => n27446, A2 => n27472, ZN => n26907);
   U10589 : NAND2_X1 port map( A1 => n7254, A2 => n3593, ZN => n7255);
   U10590 : NAND2_X1 port map( A1 => n7383, A2 => n3594, ZN => n3593);
   U10592 : XNOR2_X1 port map( A => n23961, B => n25713, ZN => n3596);
   U10594 : NAND2_X1 port map( A1 => n11273, A2 => n10522, ZN => n11039);
   U10595 : NAND2_X1 port map( A1 => n4245, A2 => n20265, ZN => n20644);
   U10596 : XNOR2_X2 port map( A => n19539, B => n19538, ZN => n4245);
   U10597 : NAND3_X1 port map( A1 => n3600, A2 => n24096, A3 => n3599, ZN => 
                           n24099);
   U10598 : NAND2_X1 port map( A1 => n24470, A2 => n24092, ZN => n3600);
   U10599 : OAI211_X1 port map( C1 => n7773, C2 => n7315, A => n3601, B => 
                           n7775, ZN => n7277);
   U10600 : NAND2_X1 port map( A1 => n7773, A2 => n7089, ZN => n3601);
   U10603 : OAI22_X1 port map( A1 => n28126, A2 => n4167, B1 => n28133, B2 => 
                           n21359, ZN => n20263);
   U10605 : NAND2_X1 port map( A1 => n13885, A2 => n14319, ZN => n3602);
   U10606 : NAND2_X1 port map( A1 => n3964, A2 => n4844, ZN => n3963);
   U10607 : OR2_X1 port map( A1 => n17719, A2 => n17859, ZN => n17721);
   U10608 : NAND2_X1 port map( A1 => n17438, A2 => n17433, ZN => n17436);
   U10609 : NAND2_X1 port map( A1 => n13694, A2 => n14323, ZN => n13695);
   U10610 : XNOR2_X1 port map( A => n13315, B => n13220, ZN => n13094);
   U10611 : INV_X1 port map( A => n23486, ZN => n3700);
   U10612 : NOR2_X2 port map( A1 => n22875, A2 => n22876, ZN => n24592);
   U10613 : INV_X2 port map( A => n16822, ZN => n17707);
   U10614 : NAND2_X1 port map( A1 => n12183, A2 => n3604, ZN => n11731);
   U10615 : MUX2_X2 port map( A => n14229, B => n14228, S => n14715, Z => 
                           n16449);
   U10617 : NAND2_X1 port map( A1 => n7176, A2 => n7900, ZN => n7803);
   U10618 : NAND2_X1 port map( A1 => n27822, A2 => n27791, ZN => n26678);
   U10619 : XNOR2_X2 port map( A => n16452, B => n16451, ZN => n17829);
   U10620 : NAND2_X1 port map( A1 => n14364, A2 => n15514, ZN => n14389);
   U10621 : XNOR2_X1 port map( A => n3611, B => n3610, ZN => Ciphertext(34));
   U10622 : NAND2_X1 port map( A1 => n485, A2 => n23419, ZN => n23096);
   U10624 : NOR2_X1 port map( A1 => n4741, A2 => n26128, ZN => n4739);
   U10625 : OAI21_X1 port map( B1 => n21019, B2 => n22023, A => n21020, ZN => 
                           n21053);
   U10626 : XNOR2_X1 port map( A => n4579, B => n19664, ZN => n4581);
   U10627 : NAND3_X1 port map( A1 => n21242, A2 => n21692, A3 => n6314, ZN => 
                           n20961);
   U10628 : NAND2_X1 port map( A1 => n13467, A2 => n14033, ZN => n3613);
   U10629 : NAND3_X2 port map( A1 => n3614, A2 => n4421, A3 => n4422, ZN => 
                           n15402);
   U10630 : NAND2_X1 port map( A1 => n4424, A2 => n4426, ZN => n3614);
   U10631 : OAI21_X1 port map( B1 => n15337, B2 => n694, A => n3615, ZN => 
                           n14528);
   U10634 : NAND2_X1 port map( A1 => n3617, A2 => n3616, ZN => n5553);
   U10635 : NAND2_X1 port map( A1 => n23387, A2 => n23220, ZN => n3617);
   U10636 : NOR2_X2 port map( A1 => n4542, A2 => n20757, ZN => n22778);
   U10638 : INV_X1 port map( A => n11198, ZN => n5917);
   U10639 : NAND2_X1 port map( A1 => n3860, A2 => n14373, ZN => n6050);
   U10640 : NAND3_X1 port map( A1 => n24422, A2 => n24420, A3 => n3618, ZN => 
                           n6547);
   U10642 : XNOR2_X1 port map( A => n4990, B => n16302, ZN => n4989);
   U10643 : OAI21_X1 port map( B1 => n14753, B2 => n15062, A => n15355, ZN => 
                           n5969);
   U10644 : INV_X1 port map( A => n18111, ZN => n17729);
   U10647 : NAND2_X1 port map( A1 => n24072, A2 => n24666, ZN => n23914);
   U10648 : NAND3_X2 port map( A1 => n3621, A2 => n3620, A3 => n21461, ZN => 
                           n22605);
   U10651 : XNOR2_X1 port map( A => n10268, B => n10267, ZN => n6666);
   U10652 : INV_X1 port map( A => n6432, ZN => n12013);
   U10654 : NAND2_X1 port map( A1 => n26496, A2 => n27366, ZN => n3623);
   U10655 : NAND2_X1 port map( A1 => n12304, A2 => n11491, ZN => n11767);
   U10656 : INV_X1 port map( A => n11003, ZN => n6779);
   U10657 : XNOR2_X1 port map( A => n13554, B => n13007, ZN => n3624);
   U10658 : NOR2_X1 port map( A1 => n27368, A2 => n27362, ZN => n27363);
   U10659 : NAND2_X1 port map( A1 => n7093, A2 => n7601, ZN => n7868);
   U10660 : NOR2_X1 port map( A1 => n27152, A2 => n27151, ZN => n27160);
   U10663 : NAND2_X1 port map( A1 => n16613, A2 => n17491, ZN => n3629);
   U10666 : NAND2_X1 port map( A1 => n23758, A2 => n23326, ZN => n23189);
   U10667 : XNOR2_X2 port map( A => n22344, B => n22345, ZN => n23758);
   U10668 : NAND2_X1 port map( A1 => n3630, A2 => n24700, ZN => n3696);
   U10669 : NAND2_X1 port map( A1 => n1856, A2 => n24765, ZN => n24700);
   U10671 : NAND2_X1 port map( A1 => n23746, A2 => n23408, ZN => n3631);
   U10672 : AOI21_X1 port map( B1 => n26501, B2 => n27069, A => n28545, ZN => 
                           n3632);
   U10673 : NAND3_X1 port map( A1 => n18015, A2 => n28633, A3 => n17674, ZN => 
                           n17675);
   U10674 : NAND2_X1 port map( A1 => n8162, A2 => n7348, ZN => n7536);
   U10675 : NAND2_X1 port map( A1 => n7303, A2 => n7582, ZN => n7883);
   U10676 : NAND2_X1 port map( A1 => n12088, A2 => n11856, ZN => n3958);
   U10678 : NAND3_X1 port map( A1 => n458, A2 => n24455, A3 => n24456, ZN => 
                           n3634);
   U10679 : NAND2_X1 port map( A1 => n5170, A2 => n11550, ZN => n6027);
   U10680 : NAND3_X1 port map( A1 => n17563, A2 => n17562, A3 => n532, ZN => 
                           n3839);
   U10681 : OR2_X1 port map( A1 => n431, A2 => n12337, ZN => n12341);
   U10682 : NAND2_X1 port map( A1 => n11351, A2 => n10847, ZN => n3636);
   U10683 : NAND3_X1 port map( A1 => n5987, A2 => n5988, A3 => n17067, ZN => 
                           n5986);
   U10684 : NAND3_X1 port map( A1 => n14806, A2 => n14769, A3 => n3638, ZN => 
                           n14772);
   U10686 : NOR2_X1 port map( A1 => n8525, A2 => n9221, ZN => n8098);
   U10687 : XOR2_X1 port map( A => n16532, B => n16533, Z => n6890);
   U10689 : AOI21_X1 port map( B1 => n17589, B2 => n18506, A => n5392, ZN => 
                           n17590);
   U10690 : XNOR2_X1 port map( A => n25757, B => n25758, ZN => n26322);
   U10691 : XNOR2_X2 port map( A => n13571, B => n13570, ZN => n14380);
   U10692 : NAND3_X1 port map( A1 => n3641, A2 => n5572, A3 => n3640, ZN => 
                           n11944);
   U10693 : NAND2_X1 port map( A1 => n10938, A2 => n10937, ZN => n3641);
   U10694 : XNOR2_X2 port map( A => n16016, B => n16015, ZN => n17249);
   U10695 : NAND2_X1 port map( A1 => n29301, A2 => n1938, ZN => n3642);
   U10696 : NAND2_X1 port map( A1 => n15107, A2 => n14937, ZN => n12370);
   U10698 : INV_X1 port map( A => n24725, ZN => n24730);
   U10699 : INV_X1 port map( A => n7675, ZN => n7963);
   U10701 : OAI211_X1 port map( C1 => n11836, C2 => n12510, A => n11835, B => 
                           n11834, ZN => n3647);
   U10706 : XNOR2_X1 port map( A => n25429, B => n25368, ZN => n3649);
   U10707 : OR2_X1 port map( A1 => n3978, A2 => n15259, ZN => n3977);
   U10709 : XNOR2_X1 port map( A => n10042, B => n10041, ZN => n3829);
   U10710 : INV_X1 port map( A => n9037, ZN => n9031);
   U10712 : INV_X1 port map( A => n10534, ZN => n11219);
   U10713 : INV_X1 port map( A => n17540, ZN => n16939);
   U10714 : INV_X1 port map( A => n14630, ZN => n15387);
   U10715 : INV_X1 port map( A => n3946, ZN => n11858);
   U10716 : OAI21_X1 port map( B1 => n1865, B2 => n10445, A => n3651, ZN => 
                           n10947);
   U10717 : NAND2_X1 port map( A1 => n10940, A2 => n28495, ZN => n3651);
   U10719 : INV_X1 port map( A => n24768, ZN => n24427);
   U10720 : INV_X1 port map( A => n17179, ZN => n4295);
   U10721 : OAI21_X1 port map( B1 => n12508, B2 => n3653, A => n3652, ZN => 
                           n10118);
   U10722 : NAND2_X1 port map( A1 => n12508, A2 => n12512, ZN => n3652);
   U10723 : OR2_X1 port map( A1 => n14301, A2 => n13646, ZN => n13817);
   U10724 : AOI21_X1 port map( B1 => n7725, B2 => n7723, A => n7721, ZN => 
                           n7339);
   U10725 : NAND2_X1 port map( A1 => n6727, A2 => n17137, ZN => n17142);
   U10726 : INV_X1 port map( A => n23377, ZN => n23202);
   U10727 : MUX2_X2 port map( A => n25197, B => n25196, S => n26775, Z => 
                           n27547);
   U10729 : NAND2_X1 port map( A1 => n3655, A2 => n7691, ZN => n5910);
   U10730 : NAND3_X1 port map( A1 => n3656, A2 => n7366, A3 => n8207, ZN => 
                           n7365);
   U10731 : NAND2_X1 port map( A1 => n8202, A2 => n7634, ZN => n3656);
   U10733 : NOR3_X1 port map( A1 => n21442, A2 => n21653, A3 => n21655, ZN => 
                           n5764);
   U10734 : INV_X1 port map( A => n18972, ZN => n19989);
   U10735 : NAND2_X1 port map( A1 => n12201, A2 => n12200, ZN => n11703);
   U10736 : OR2_X2 port map( A1 => n9257, A2 => n9256, ZN => n12201);
   U10737 : NAND3_X1 port map( A1 => n8039, A2 => n6210, A3 => n7514, ZN => 
                           n7024);
   U10738 : AOI21_X1 port map( B1 => n26969, B2 => n3657, A => n27429, ZN => 
                           n26970);
   U10739 : NAND2_X1 port map( A1 => n27420, A2 => n27428, ZN => n3657);
   U10740 : NAND2_X1 port map( A1 => n20789, A2 => n29586, ZN => n3658);
   U10741 : XNOR2_X1 port map( A => n19130, B => n18875, ZN => n3659);
   U10742 : MUX2_X1 port map( A => n28065, B => n28066, S => n28064, Z => 
                           n28059);
   U10743 : NAND2_X1 port map( A1 => n11640, A2 => n11672, ZN => n11676);
   U10744 : OR2_X1 port map( A1 => n13795, A2 => n14029, ZN => n4251);
   U10745 : AOI22_X2 port map( A1 => n23958, A2 => n23957, B1 => n23959, B2 => 
                           n24758, ZN => n25868);
   U10746 : INV_X1 port map( A => n17349, ZN => n5420);
   U10747 : XOR2_X1 port map( A => n12911, B => n12912, Z => n4961);
   U10748 : XNOR2_X1 port map( A => n21996, B => n21997, ZN => n23227);
   U10749 : NAND2_X1 port map( A1 => n29726, A2 => n24435, ZN => n23887);
   U10750 : NAND2_X1 port map( A1 => n10577, A2 => n432, ZN => n5278);
   U10752 : INV_X1 port map( A => n11094, ZN => n5279);
   U10754 : XNOR2_X1 port map( A => n16140, B => n16139, ZN => n16142);
   U10755 : NAND2_X1 port map( A1 => n13699, A2 => n14292, ZN => n14298);
   U10756 : OAI21_X2 port map( B1 => n11313, B2 => n11312, A => n11311, ZN => 
                           n4105);
   U10757 : AOI22_X1 port map( A1 => n20880, A2 => n21266, B1 => n20879, B2 => 
                           n20881, ZN => n20882);
   U10758 : INV_X1 port map( A => n10853, ZN => n5753);
   U10759 : XNOR2_X1 port map( A => n21994, B => n4861, ZN => n22918);
   U10760 : NAND2_X1 port map( A1 => n26757, A2 => n26753, ZN => n25649);
   U10762 : OAI22_X1 port map( A1 => n23196, A2 => n23799, B1 => n23319, B2 => 
                           n23795, ZN => n21929);
   U10765 : OAI21_X1 port map( B1 => n24724, B2 => n24729, A => n6377, ZN => 
                           n3725);
   U10766 : XNOR2_X1 port map( A => n9618, B => n9617, ZN => n10668);
   U10769 : INV_X1 port map( A => n3738, ZN => n3737);
   U10770 : AOI21_X1 port map( B1 => n20799, B2 => n20800, A => n28916, ZN => 
                           n6346);
   U10771 : XNOR2_X1 port map( A => n9301, B => n9596, ZN => n3663);
   U10772 : XNOR2_X1 port map( A => n25512, B => n25511, ZN => n27010);
   U10774 : INV_X1 port map( A => n23776, ZN => n23513);
   U10775 : AOI21_X1 port map( B1 => n14013, B2 => n14126, A => n13060, ZN => 
                           n14014);
   U10776 : XNOR2_X1 port map( A => n19154, B => n19153, ZN => n4747);
   U10777 : NAND2_X1 port map( A1 => n4868, A2 => n4869, ZN => n4867);
   U10778 : NAND2_X1 port map( A1 => n20532, A2 => n22013, ZN => n20934);
   U10779 : NAND2_X1 port map( A1 => n20086, A2 => n20085, ZN => n20532);
   U10780 : NAND2_X1 port map( A1 => n3665, A2 => n3664, ZN => n7095);
   U10781 : NAND2_X1 port map( A1 => n7093, A2 => n7092, ZN => n3665);
   U10782 : NAND2_X1 port map( A1 => n20935, A2 => n22012, ZN => n4378);
   U10783 : NAND2_X1 port map( A1 => n7363, A2 => n28605, ZN => n7831);
   U10784 : XNOR2_X1 port map( A => n24330, B => n26056, ZN => n24345);
   U10786 : OR3_X1 port map( A1 => n7867, A2 => n7092, A3 => n7093, ZN => n4438
                           );
   U10787 : NAND2_X1 port map( A1 => n5838, A2 => n6687, ZN => n3667);
   U10788 : NAND2_X1 port map( A1 => n5370, A2 => n11955, ZN => n3668);
   U10790 : NOR2_X1 port map( A1 => n13654, A2 => n13799, ZN => n4780);
   U10791 : XNOR2_X1 port map( A => n16119, B => n16122, ZN => n3677);
   U10792 : NAND2_X1 port map( A1 => n6657, A2 => n11537, ZN => n6660);
   U10793 : OAI21_X1 port map( B1 => n10754, B2 => n11155, A => n3669, ZN => 
                           n4971);
   U10794 : NAND2_X1 port map( A1 => n4972, A2 => n10804, ZN => n3669);
   U10795 : NOR2_X1 port map( A1 => n16820, A2 => n17463, ZN => n17090);
   U10796 : NAND2_X1 port map( A1 => n15458, A2 => n28462, ZN => n14537);
   U10798 : NAND2_X1 port map( A1 => n17067, A2 => n17450, ZN => n3672);
   U10799 : INV_X1 port map( A => n22902, ZN => n6818);
   U10801 : AOI21_X1 port map( B1 => n3674, B2 => n20496, A => n20495, ZN => 
                           n21329);
   U10802 : NAND2_X1 port map( A1 => n20494, A2 => n29616, ZN => n3674);
   U10803 : NOR3_X1 port map( A1 => n29090, A2 => n27663, A3 => n27671, ZN => 
                           n27195);
   U10804 : OAI21_X2 port map( B1 => n27160, B2 => n27159, A => n27158, ZN => 
                           n27663);
   U10805 : NAND2_X1 port map( A1 => n8765, A2 => n8763, ZN => n8943);
   U10807 : NAND2_X1 port map( A1 => n7226, A2 => n7225, ZN => n3676);
   U10809 : INV_X1 port map( A => n3679, ZN => n3678);
   U10810 : NAND2_X1 port map( A1 => n3680, A2 => n29063, ZN => n27955);
   U10811 : OAI21_X1 port map( B1 => n27970, B2 => n27997, A => n28456, ZN => 
                           n3680);
   U10813 : NAND2_X1 port map( A1 => n27854, A2 => n26641, ZN => n3681);
   U10814 : NAND2_X1 port map( A1 => n14044, A2 => n14045, ZN => n14049);
   U10815 : AOI22_X1 port map( A1 => n15357, A2 => n6674, B1 => n15358, B2 => 
                           n15359, ZN => n3682);
   U10816 : XNOR2_X1 port map( A => n2003, B => n13430, ZN => n5165);
   U10817 : NAND3_X1 port map( A1 => n26643, A2 => n6954, A3 => n26644, ZN => 
                           n26645);
   U10819 : NAND2_X1 port map( A1 => n11373, A2 => n12211, ZN => n3684);
   U10820 : NAND2_X1 port map( A1 => n11374, A2 => n6281, ZN => n3685);
   U10822 : INV_X1 port map( A => n20769, ZN => n20771);
   U10823 : AOI21_X1 port map( B1 => n17354, B2 => n2449, A => n17031, ZN => 
                           n17199);
   U10824 : OAI21_X1 port map( B1 => n21313, B2 => n21312, A => n5899, ZN => 
                           n5898);
   U10825 : XNOR2_X1 port map( A => n3689, B => n19193, ZN => n19197);
   U10826 : XNOR2_X1 port map( A => n3730, B => n5416, ZN => n3689);
   U10827 : NOR2_X1 port map( A1 => n18709, A2 => n18248, ZN => n17598);
   U10828 : NAND2_X1 port map( A1 => n3691, A2 => n28794, ZN => n3690);
   U10829 : NAND2_X1 port map( A1 => n3693, A2 => n3692, ZN => n20812);
   U10830 : NAND2_X1 port map( A1 => n3694, A2 => n21664, ZN => n3693);
   U10831 : NAND2_X1 port map( A1 => n21662, A2 => n21429, ZN => n3694);
   U10832 : INV_X1 port map( A => n19765, ZN => n3911);
   U10833 : AOI22_X1 port map( A1 => n27312, A2 => n27873, B1 => n27313, B2 => 
                           n27314, ZN => n27323);
   U10834 : NAND3_X1 port map( A1 => n20972, A2 => n20703, A3 => n21217, ZN => 
                           n19915);
   U10835 : OAI21_X1 port map( B1 => n27041, B2 => n4497, A => n4496, ZN => 
                           n4495);
   U10836 : NAND2_X1 port map( A1 => n23777, A2 => n23776, ZN => n6423);
   U10837 : NOR2_X2 port map( A1 => n3698, A2 => n23485, ZN => n24777);
   U10838 : NAND2_X1 port map( A1 => n23484, A2 => n23483, ZN => n3699);
   U10839 : OAI21_X1 port map( B1 => n18502, B2 => n18501, A => n515, ZN => 
                           n3701);
   U10841 : NAND2_X1 port map( A1 => n17137, A2 => n17138, ZN => n5471);
   U10842 : XOR2_X1 port map( A => n22055, B => n22843, Z => n6100);
   U10843 : NAND3_X2 port map( A1 => n3705, A2 => n12889, A3 => n12890, ZN => 
                           n16606);
   U10844 : INV_X1 port map( A => n4073, ZN => n4072);
   U10845 : XNOR2_X1 port map( A => n13438, B => n12410, ZN => n4198);
   U10846 : NAND2_X1 port map( A1 => n11351, A2 => n11192, ZN => n10478);
   U10847 : NAND3_X1 port map( A1 => n11914, A2 => n12030, A3 => n12340, ZN => 
                           n11917);
   U10848 : NAND2_X1 port map( A1 => n3706, A2 => n8828, ZN => n8467);
   U10849 : OAI211_X2 port map( C1 => n24108, C2 => n24107, A => n3708, B => 
                           n3707, ZN => n25385);
   U10850 : NAND2_X1 port map( A1 => n24105, A2 => n24104, ZN => n3707);
   U10851 : NAND2_X1 port map( A1 => n24106, A2 => n28416, ZN => n3708);
   U10853 : INV_X1 port map( A => n23978, ZN => n23981);
   U10854 : INV_X1 port map( A => n13816, ZN => n14300);
   U10855 : INV_X1 port map( A => n3826, ZN => n3824);
   U10856 : NAND2_X1 port map( A1 => n18495, A2 => n28745, ZN => n3709);
   U10857 : XNOR2_X1 port map( A => n16185, B => n3083, ZN => n16005);
   U10858 : NAND2_X1 port map( A1 => n15031, A2 => n14824, ZN => n15433);
   U10860 : OAI21_X1 port map( B1 => n28142, B2 => n17989, A => n3711, ZN => 
                           n17892);
   U10861 : NAND2_X1 port map( A1 => n17989, A2 => n18599, ZN => n3711);
   U10863 : XNOR2_X2 port map( A => n15710, B => n15709, ZN => n17365);
   U10865 : INV_X1 port map( A => n16526, ZN => n15706);
   U10866 : OAI21_X1 port map( B1 => n2762, B2 => n24405, A => n4081, ZN => 
                           n4176);
   U10867 : NAND2_X1 port map( A1 => n4931, A2 => n9209, ZN => n3718);
   U10868 : XNOR2_X1 port map( A => n6536, B => n6534, ZN => n20284);
   U10869 : INV_X1 port map( A => n22919, ZN => n22574);
   U10870 : NOR2_X1 port map( A1 => n23145, A2 => n23460, ZN => n23356);
   U10871 : NAND2_X1 port map( A1 => n26169, A2 => n26786, ZN => n3720);
   U10872 : XNOR2_X1 port map( A => n3721, B => n26288, ZN => Ciphertext(185));
   U10873 : NAND2_X1 port map( A1 => n5214, A2 => n5215, ZN => n3721);
   U10874 : NAND2_X1 port map( A1 => n4839, A2 => n7715, ZN => n6192);
   U10875 : NAND2_X1 port map( A1 => n4644, A2 => n26684, ZN => n26685);
   U10877 : NAND2_X1 port map( A1 => n28064, A2 => n28066, ZN => n5213);
   U10878 : NAND3_X1 port map( A1 => n23030, A2 => n23031, A3 => n23029, ZN => 
                           n23032);
   U10879 : OAI22_X1 port map( A1 => n18456, A2 => n18106, B1 => n18109, B2 => 
                           n18111, ZN => n17730);
   U10880 : XNOR2_X1 port map( A => n3724, B => n12892, ZN => n12871);
   U10881 : XNOR2_X1 port map( A => n12865, B => n12866, ZN => n3724);
   U10883 : NAND2_X1 port map( A1 => n18261, A2 => n18326, ZN => n4059);
   U10884 : INV_X1 port map( A => n21183, ZN => n21129);
   U10886 : INV_X1 port map( A => n3726, ZN => n6407);
   U10887 : OAI21_X1 port map( B1 => n23333, B2 => n6462, A => n23332, ZN => 
                           n3726);
   U10890 : NAND3_X1 port map( A1 => n17417, A2 => n17418, A3 => n17419, ZN => 
                           n18402);
   U10891 : NAND3_X1 port map( A1 => n10850, A2 => n10848, A3 => n4123, ZN => 
                           n12158);
   U10894 : NAND3_X1 port map( A1 => n17489, A2 => n17148, A3 => n17078, ZN => 
                           n4653);
   U10896 : NAND2_X1 port map( A1 => n16008, A2 => n1880, ZN => n3729);
   U10897 : NOR2_X1 port map( A1 => n294, A2 => n27213, ZN => n6809);
   U10899 : NAND2_X1 port map( A1 => n24891, A2 => n24532, ZN => n6865);
   U10900 : XNOR2_X1 port map( A => n19192, B => n3598, ZN => n3730);
   U10901 : INV_X1 port map( A => n11462, ZN => n11461);
   U10902 : OAI22_X1 port map( A1 => n10803, A2 => n28559, B1 => n10553, B2 => 
                           n11158, ZN => n10496);
   U10903 : NOR2_X1 port map( A1 => n11941, A2 => n11942, ZN => n3732);
   U10904 : NAND2_X1 port map( A1 => n29573, A2 => n26278, ZN => n26392);
   U10905 : NAND2_X1 port map( A1 => n5064, A2 => n13909, ZN => n6813);
   U10907 : INV_X1 port map( A => n3734, ZN => n3733);
   U10908 : OAI21_X1 port map( B1 => n13992, B2 => n15692, A => n13990, ZN => 
                           n3734);
   U10910 : NAND2_X1 port map( A1 => n3735, A2 => n28526, ZN => n19752);
   U10912 : NOR2_X1 port map( A1 => n27150, A2 => n6592, ZN => n6591);
   U10913 : NAND2_X1 port map( A1 => n7244, A2 => n7648, ZN => n3736);
   U10914 : OAI21_X1 port map( B1 => n1801, B2 => n16383, A => n16382, ZN => 
                           n3738);
   U10915 : NAND3_X1 port map( A1 => n4652, A2 => n4651, A3 => n29294, ZN => 
                           n3739);
   U10916 : INV_X1 port map( A => n20977, ZN => n21367);
   U10917 : INV_X1 port map( A => n8395, ZN => n8396);
   U10918 : NOR2_X1 port map( A1 => n23067, A2 => n4429, ZN => n4459);
   U10919 : XOR2_X1 port map( A => n20655, B => n20654, Z => n4430);
   U10920 : NAND3_X1 port map( A1 => n5267, A2 => n5265, A3 => n10976, ZN => 
                           n10978);
   U10921 : NAND2_X1 port map( A1 => n18354, A2 => n18312, ZN => n6030);
   U10922 : NOR2_X1 port map( A1 => n580, A2 => n12350, ZN => n5133);
   U10923 : OAI22_X1 port map( A1 => n28183, A2 => n29157, B1 => n23722, B2 => 
                           n23843, ZN => n22127);
   U10924 : OR2_X1 port map( A1 => n18340, A2 => n514, ZN => n4244);
   U10926 : NAND2_X1 port map( A1 => n3741, A2 => n14142, ZN => n14143);
   U10928 : AND2_X1 port map( A1 => n20349, A2 => n20510, ZN => n5853);
   U10929 : INV_X1 port map( A => n18520, ZN => n19262);
   U10930 : INV_X1 port map( A => n5953, ZN => n21561);
   U10931 : INV_X1 port map( A => n10502, ZN => n5672);
   U10932 : INV_X1 port map( A => n12186, ZN => n4028);
   U10934 : XNOR2_X1 port map( A => n19598, B => n18720, ZN => n5211);
   U10935 : NAND3_X1 port map( A1 => n474, A2 => n29544, A3 => n23169, ZN => 
                           n23170);
   U10936 : NAND2_X1 port map( A1 => n8511, A2 => n8914, ZN => n9105);
   U10937 : NAND2_X1 port map( A1 => n11132, A2 => n10711, ZN => n10501);
   U10939 : NAND2_X1 port map( A1 => n12264, A2 => n575, ZN => n3745);
   U10940 : NAND2_X1 port map( A1 => n8800, A2 => n8802, ZN => n8957);
   U10941 : INV_X1 port map( A => n14702, ZN => n3748);
   U10942 : NAND2_X1 port map( A1 => n14851, A2 => n15310, ZN => n5948);
   U10943 : NAND2_X1 port map( A1 => n5928, A2 => n21088, ZN => n5926);
   U10944 : MUX2_X2 port map( A => n22051, B => n22050, S => n28796, Z => 
                           n24584);
   U10945 : OR2_X1 port map( A1 => n7614, A2 => n7393, ZN => n7930);
   U10946 : OR2_X1 port map( A1 => n20784, A2 => n21177, ZN => n5087);
   U10947 : XOR2_X1 port map( A => n20797, B => n22383, Z => n5452);
   U10948 : NOR2_X1 port map( A1 => n6530, A2 => n21031, ZN => n6527);
   U10949 : XNOR2_X1 port map( A => n26103, B => n26100, ZN => n6018);
   U10950 : NAND2_X1 port map( A1 => n27186, A2 => n26397, ZN => n3754);
   U10951 : NAND2_X1 port map( A1 => n15502, A2 => n15265, ZN => n14924);
   U10952 : NAND3_X2 port map( A1 => n3757, A2 => n6402, A3 => n3756, ZN => 
                           n19726);
   U10953 : NAND2_X1 port map( A1 => n18328, A2 => n18329, ZN => n3756);
   U10955 : INV_X1 port map( A => n21563, ZN => n3759);
   U10956 : NOR2_X1 port map( A1 => n21564, A2 => n28155, ZN => n3760);
   U10957 : OAI21_X1 port map( B1 => n20500, B2 => n29601, A => n20498, ZN => 
                           n3761);
   U10958 : AOI21_X1 port map( B1 => n21156, B2 => n3762, A => n494, ZN => 
                           n4755);
   U10960 : NAND2_X1 port map( A1 => n3764, A2 => n3763, ZN => n5899);
   U10961 : INV_X1 port map( A => n21311, ZN => n3763);
   U10962 : NAND2_X1 port map( A1 => n29530, A2 => n21309, ZN => n3764);
   U10963 : NAND2_X1 port map( A1 => n6132, A2 => n12286, ZN => n3765);
   U10964 : XNOR2_X1 port map( A => n1895, B => n10184, ZN => n6136);
   U10965 : OAI21_X1 port map( B1 => n18711, B2 => n18709, A => n3766, ZN => 
                           n18714);
   U10971 : OAI21_X1 port map( B1 => n9232, B2 => n9229, A => n3773, ZN => 
                           n9046);
   U10972 : NAND2_X1 port map( A1 => n9232, A2 => n9233, ZN => n3773);
   U10973 : OAI21_X1 port map( B1 => n7695, B2 => n8227, A => n3774, ZN => 
                           n6991);
   U10974 : NAND2_X1 port map( A1 => n7695, A2 => n8222, ZN => n3774);
   U10975 : OR2_X2 port map( A1 => n10596, A2 => n10595, ZN => n12359);
   U10976 : XNOR2_X1 port map( A => n3775, B => n22504, ZN => n22991);
   U10977 : XNOR2_X1 port map( A => n6388, B => n6389, ZN => n3775);
   U10978 : AOI21_X1 port map( B1 => n11612, B2 => n11613, A => n566, ZN => 
                           n5465);
   U10980 : NOR2_X1 port map( A1 => n11140, A2 => n3829, ZN => n10721);
   U10983 : AOI21_X1 port map( B1 => n15078, B2 => n5229, A => n3778, ZN => 
                           n3777);
   U10984 : NOR2_X1 port map( A1 => n14876, A2 => n15082, ZN => n3778);
   U10985 : NAND3_X1 port map( A1 => n5546, A2 => n26768, A3 => n26771, ZN => 
                           n25158);
   U10986 : NAND2_X1 port map( A1 => n6556, A2 => n24020, ZN => n24002);
   U10987 : XOR2_X1 port map( A => n25389, B => n25388, Z => n6071);
   U10988 : XNOR2_X1 port map( A => n3779, B => n19175, ZN => n18785);
   U10989 : XNOR2_X1 port map( A => n18783, B => n19331, ZN => n3779);
   U10990 : NAND2_X1 port map( A1 => n6734, A2 => n6737, ZN => n26495);
   U10992 : NAND2_X1 port map( A1 => n26497, A2 => n27364, ZN => n25997);
   U10993 : INV_X1 port map( A => n18170, ZN => n5200);
   U10994 : NAND2_X1 port map( A1 => n23364, A2 => n23672, ZN => n23362);
   U10995 : NAND2_X2 port map( A1 => n6115, A2 => n20685, ZN => n22890);
   U10998 : XNOR2_X1 port map( A => n16059, B => n16649, ZN => n15608);
   U10999 : NAND3_X2 port map( A1 => n14022, A2 => n14023, A3 => n3782, ZN => 
                           n16059);
   U11000 : NAND2_X1 port map( A1 => n27071, A2 => n26614, ZN => n3785);
   U11001 : NAND2_X1 port map( A1 => n27070, A2 => n29520, ZN => n3786);
   U11003 : XNOR2_X1 port map( A => n16201, B => n16200, ZN => n6869);
   U11004 : XNOR2_X1 port map( A => n13355, B => n4490, ZN => n13356);
   U11005 : OAI22_X1 port map( A1 => n20397, A2 => n20396, B1 => n20395, B2 => 
                           n20394, ZN => n5871);
   U11006 : INV_X1 port map( A => n19277, ZN => n18369);
   U11007 : NAND2_X1 port map( A1 => n4429, A2 => n23067, ZN => n23348);
   U11008 : NAND2_X1 port map( A1 => n6450, A2 => n3788, ZN => n10372);
   U11009 : NAND3_X1 port map( A1 => n7659, A2 => n8305, A3 => n3790, ZN => 
                           n7402);
   U11010 : NAND2_X1 port map( A1 => n8302, A2 => n7657, ZN => n3790);
   U11011 : AND3_X2 port map( A1 => n3836, A2 => n24781, A3 => n24782, ZN => 
                           n25191);
   U11014 : NAND2_X1 port map( A1 => n17480, A2 => n17477, ZN => n3884);
   U11016 : INV_X1 port map( A => n26682, ZN => n26710);
   U11017 : INV_X1 port map( A => n28395, ZN => n14890);
   U11018 : XNOR2_X1 port map( A => n3792, B => n16024, ZN => n16555);
   U11019 : XNOR2_X1 port map( A => n28395, B => n16199, ZN => n15673);
   U11020 : AND2_X1 port map( A1 => n7792, A2 => n7793, ZN => n7795);
   U11021 : OAI21_X1 port map( B1 => n7797, B2 => n28149, A => n3793, ZN => 
                           n7798);
   U11022 : NAND3_X1 port map( A1 => n7284, A2 => n7792, A3 => n7793, ZN => 
                           n3793);
   U11023 : NAND3_X1 port map( A1 => n12990, A2 => n12090, A3 => n3796, ZN => 
                           n3794);
   U11024 : NAND2_X1 port map( A1 => n3961, A2 => n12151, ZN => n12090);
   U11025 : NAND2_X1 port map( A1 => n3797, A2 => n24405, ZN => n23503);
   U11026 : NAND2_X1 port map( A1 => n24085, A2 => n3797, ZN => n23880);
   U11028 : NAND2_X1 port map( A1 => n3799, A2 => n3798, ZN => n5834);
   U11030 : NAND2_X1 port map( A1 => n10983, A2 => n10982, ZN => n10696);
   U11032 : INV_X1 port map( A => n10980, ZN => n3804);
   U11033 : INV_X1 port map( A => n10980, ZN => n10783);
   U11034 : NAND2_X1 port map( A1 => n10988, A2 => n10985, ZN => n3805);
   U11035 : NAND2_X1 port map( A1 => n13968, A2 => n3806, ZN => n13969);
   U11036 : INV_X1 port map( A => n12711, ZN => n3806);
   U11037 : MUX2_X1 port map( A => n14459, B => n4290, S => n12711, Z => n13683
                           );
   U11039 : NAND3_X1 port map( A1 => n19947, A2 => n20200, A3 => n20305, ZN => 
                           n3808);
   U11040 : NAND3_X1 port map( A1 => n8147, A2 => n7793, A3 => n7796, ZN => 
                           n7286);
   U11041 : NAND3_X1 port map( A1 => n7541, A2 => n8148, A3 => n3810, ZN => 
                           n7354);
   U11044 : NAND2_X1 port map( A1 => n16611, A2 => n18356, ZN => n17920);
   U11045 : XNOR2_X1 port map( A => n16170, B => n16279, ZN => n3813);
   U11046 : NOR2_X2 port map( A1 => n15340, A2 => n15341, ZN => n16170);
   U11047 : INV_X1 port map( A => n11252, ZN => n3817);
   U11048 : NAND2_X1 port map( A1 => n11251, A2 => n3816, ZN => n3815);
   U11049 : NAND2_X1 port map( A1 => n11033, A2 => n11252, ZN => n3818);
   U11050 : NOR2_X1 port map( A1 => n11033, A2 => n3820, ZN => n3819);
   U11053 : NAND3_X1 port map( A1 => n6203, A2 => n5783, A3 => n4245, ZN => 
                           n21065);
   U11055 : NAND2_X1 port map( A1 => n3824, A2 => n18486, ZN => n3823);
   U11056 : NAND2_X1 port map( A1 => n18490, A2 => n18489, ZN => n3826);
   U11057 : AOI22_X1 port map( A1 => n15289, A2 => n15291, B1 => n15290, B2 => 
                           n3827, ZN => n15298);
   U11058 : NAND2_X1 port map( A1 => n3827, A2 => n14517, ZN => n15215);
   U11059 : OAI21_X1 port map( B1 => n15217, B2 => n15290, A => n3827, ZN => 
                           n15041);
   U11061 : OAI211_X1 port map( C1 => n15217, C2 => n3827, A => n15293, B => 
                           n15292, ZN => n14110);
   U11062 : OAI21_X1 port map( B1 => n15289, B2 => n3827, A => n14097, ZN => 
                           n4957);
   U11063 : NAND2_X1 port map( A1 => n11138, A2 => n3828, ZN => n10719);
   U11064 : NAND2_X1 port map( A1 => n11139, A2 => n3829, ZN => n10923);
   U11065 : NAND2_X1 port map( A1 => n10103, A2 => n3829, ZN => n10106);
   U11066 : NAND2_X1 port map( A1 => n5531, A2 => n13914, ZN => n3830);
   U11067 : NAND2_X1 port map( A1 => n17713, A2 => n18329, ZN => n3831);
   U11068 : MUX2_X1 port map( A => n27106, B => n27701, S => n27702, Z => 
                           n27107);
   U11069 : MUX2_X1 port map( A => n27162, B => n27163, S => n27702, Z => 
                           n27164);
   U11071 : INV_X1 port map( A => n25133, ZN => n3837);
   U11072 : XNOR2_X1 port map( A => n25191, B => n24897, ZN => n24898);
   U11073 : NAND2_X1 port map( A1 => n3838, A2 => n21124, ZN => n21461);
   U11074 : NOR2_X1 port map( A1 => n3838, A2 => n21459, ZN => n21460);
   U11075 : NOR2_X1 port map( A1 => n1814, A2 => n3838, ZN => n20843);
   U11076 : NAND2_X1 port map( A1 => n3784, A2 => n15008, ZN => n14867);
   U11077 : INV_X1 port map( A => n15373, ZN => n15008);
   U11078 : NOR2_X1 port map( A1 => n15373, A2 => n15374, ZN => n3841);
   U11079 : NAND2_X1 port map( A1 => n12508, A2 => n11990, ZN => n3842);
   U11080 : NAND2_X1 port map( A1 => n3842, A2 => n12507, ZN => n11521);
   U11081 : OAI21_X1 port map( B1 => n15471, B2 => n14551, A => n15472, ZN => 
                           n3845);
   U11082 : NAND2_X1 port map( A1 => n1848, A2 => n15168, ZN => n15472);
   U11085 : INV_X1 port map( A => n13866, ZN => n3846);
   U11086 : NAND2_X1 port map( A1 => n522, A2 => n17969, ZN => n3848);
   U11089 : OR2_X1 port map( A1 => n14209, A2 => n3851, ZN => n3850);
   U11090 : NAND2_X1 port map( A1 => n3853, A2 => n3852, ZN => n3855);
   U11091 : NAND2_X1 port map( A1 => n20228, A2 => n20227, ZN => n3853);
   U11092 : NAND2_X1 port map( A1 => n3854, A2 => n21439, ZN => n21441);
   U11093 : AND2_X1 port map( A1 => n3855, A2 => n21438, ZN => n3854);
   U11094 : XNOR2_X1 port map( A => n3856, B => n16585, ZN => n15631);
   U11095 : XNOR2_X1 port map( A => n3856, B => n16085, ZN => n16243);
   U11096 : OR2_X1 port map( A1 => n13725, A2 => n3860, ZN => n13724);
   U11097 : AND2_X1 port map( A1 => n3860, A2 => n13725, ZN => n13440);
   U11098 : NAND2_X1 port map( A1 => n14146, A2 => n3860, ZN => n4331);
   U11099 : NAND2_X1 port map( A1 => n5404, A2 => n3860, ZN => n5403);
   U11100 : NAND2_X1 port map( A1 => n5405, A2 => n3859, ZN => n14009);
   U11102 : OAI21_X1 port map( B1 => n3862, B2 => n11135, A => n3861, ZN => 
                           n3863);
   U11103 : NAND2_X1 port map( A1 => n11136, A2 => n11135, ZN => n3861);
   U11104 : NOR2_X2 port map( A1 => n10766, A2 => n10767, ZN => n11881);
   U11106 : OR2_X1 port map( A1 => n18109, A2 => n17902, ZN => n3866);
   U11108 : OAI21_X1 port map( B1 => n3868, B2 => n3867, A => n14157, ZN => 
                           n14550);
   U11109 : NAND2_X1 port map( A1 => n3869, A2 => n14158, ZN => n14549);
   U11110 : NAND2_X1 port map( A1 => n13847, A2 => n13936, ZN => n3869);
   U11111 : XNOR2_X1 port map( A => n13444, B => n13493, ZN => n3870);
   U11112 : XNOR2_X1 port map( A => n12699, B => n3871, ZN => n12701);
   U11113 : XNOR2_X1 port map( A => n3871, B => n3232, ZN => n13239);
   U11115 : NAND3_X1 port map( A1 => n3873, A2 => n29517, A3 => n11207, ZN => 
                           n11208);
   U11116 : NAND2_X1 port map( A1 => n11090, A2 => n3873, ZN => n10576);
   U11117 : NAND2_X1 port map( A1 => n432, A2 => n3873, ZN => n11092);
   U11118 : NAND3_X1 port map( A1 => n10431, A2 => n6164, A3 => n3873, ZN => 
                           n6163);
   U11119 : INV_X1 port map( A => n11094, ZN => n3873);
   U11120 : NAND3_X1 port map( A1 => n3875, A2 => n512, A3 => n17823, ZN => 
                           n3874);
   U11122 : NAND2_X1 port map( A1 => n1530, A2 => n29594, ZN => n3877);
   U11123 : INV_X1 port map( A => n3880, ZN => n17265);
   U11125 : NAND2_X1 port map( A1 => n3880, A2 => n29299, ZN => n17267);
   U11126 : NAND2_X1 port map( A1 => n16864, A2 => n3880, ZN => n3879);
   U11128 : NAND2_X1 port map( A1 => n6045, A2 => n14368, ZN => n3881);
   U11130 : NAND2_X1 port map( A1 => n17479, A2 => n17478, ZN => n3885);
   U11131 : INV_X1 port map( A => n3887, ZN => n23656);
   U11132 : NAND2_X1 port map( A1 => n4231, A2 => n3887, ZN => n4851);
   U11133 : OR2_X1 port map( A1 => n20840, A2 => n3887, ZN => n4770);
   U11134 : OAI22_X1 port map( A1 => n23352, A2 => n3887, B1 => n23545, B2 => 
                           n4232, ZN => n4648);
   U11135 : NAND2_X1 port map( A1 => n23142, A2 => n4772, ZN => n3886);
   U11136 : NAND2_X1 port map( A1 => n3888, A2 => n12231, ZN => n12230);
   U11137 : NAND2_X1 port map( A1 => n12227, A2 => n12226, ZN => n3888);
   U11138 : NAND2_X1 port map( A1 => n3890, A2 => n5339, ZN => n3889);
   U11139 : INV_X1 port map( A => n21030, ZN => n3890);
   U11140 : NAND2_X1 port map( A1 => n3892, A2 => n22146, ZN => n3891);
   U11141 : OAI21_X1 port map( B1 => n20418, B2 => n20192, A => n5334, ZN => 
                           n3893);
   U11142 : NAND2_X1 port map( A1 => n19748, A2 => n19749, ZN => n3894);
   U11143 : OR2_X1 port map( A1 => n308, A2 => n14366, ZN => n4812);
   U11144 : NAND2_X1 port map( A1 => n559, A2 => n6000, ZN => n3895);
   U11145 : AOI21_X1 port map( B1 => n308, B2 => n14123, A => n14366, ZN => 
                           n3896);
   U11146 : XNOR2_X2 port map( A => n12953, B => n12952, ZN => n14366);
   U11147 : XNOR2_X1 port map( A => n3898, B => n3897, ZN => Ciphertext(73));
   U11148 : INV_X1 port map( A => n27546, ZN => n3899);
   U11149 : AND2_X1 port map( A1 => n27549, A2 => n27203, ZN => n27199);
   U11150 : NAND2_X1 port map( A1 => n28604, A2 => n23673, ZN => n3902);
   U11151 : AOI22_X2 port map( A1 => n3903, A2 => n21678, B1 => n21082, B2 => 
                           n21081, ZN => n22199);
   U11152 : INV_X1 port map( A => n11322, ZN => n11187);
   U11153 : INV_X1 port map( A => n5595, ZN => n11181);
   U11154 : AOI21_X1 port map( B1 => n11162, B2 => n6411, A => n3904, ZN => 
                           n3910);
   U11155 : AOI21_X1 port map( B1 => n3909, B2 => n11053, A => n1933, ZN => 
                           n3908);
   U11156 : OAI211_X2 port map( C1 => n3907, C2 => n11322, A => n3906, B => 
                           n3905, ZN => n11195);
   U11158 : NAND2_X1 port map( A1 => n11164, A2 => n11165, ZN => n3909);
   U11159 : OR2_X1 port map( A1 => n17199, A2 => n17198, ZN => n3914);
   U11160 : NAND3_X1 port map( A1 => n18413, A2 => n3915, A3 => n28688, ZN => 
                           n6101);
   U11162 : NAND2_X1 port map( A1 => n17340, A2 => n17336, ZN => n6337);
   U11163 : NAND2_X1 port map( A1 => n3918, A2 => n3921, ZN => n3917);
   U11164 : NAND2_X1 port map( A1 => n3922, A2 => n14893, ZN => n3921);
   U11165 : INV_X1 port map( A => n14937, ZN => n15409);
   U11166 : NOR2_X1 port map( A1 => n15224, A2 => n15342, ZN => n3924);
   U11167 : MUX2_X1 port map( A => n15222, B => n15343, S => n15046, Z => n3926
                           );
   U11170 : NAND3_X1 port map( A1 => n14162, A2 => n14163, A3 => n14161, ZN => 
                           n3927);
   U11171 : NAND2_X1 port map( A1 => n14160, A2 => n14159, ZN => n3928);
   U11172 : INV_X1 port map( A => n7696, ZN => n3930);
   U11173 : NAND2_X1 port map( A1 => n7424, A2 => n7822, ZN => n7696);
   U11174 : NAND2_X1 port map( A1 => n3930, A2 => n7827, ZN => n3929);
   U11175 : NAND3_X1 port map( A1 => n18416, A2 => n18413, A3 => n3932, ZN => 
                           n3931);
   U11177 : XNOR2_X1 port map( A => n15698, B => n5798, ZN => n3938);
   U11178 : NAND2_X1 port map( A1 => n3939, A2 => n2052, ZN => n17343);
   U11179 : NAND2_X1 port map( A1 => n17155, A2 => n17204, ZN => n17156);
   U11180 : NAND2_X1 port map( A1 => n17337, A2 => n17336, ZN => n3939);
   U11181 : INV_X1 port map( A => n10945, ZN => n3941);
   U11182 : NAND2_X1 port map( A1 => n3946, A2 => n11944, ZN => n11665);
   U11183 : NAND2_X1 port map( A1 => n10947, A2 => n10946, ZN => n3942);
   U11184 : NAND3_X1 port map( A1 => n11948, A2 => n3946, A3 => n11945, ZN => 
                           n11946);
   U11185 : NAND3_X1 port map( A1 => n11947, A2 => n3946, A3 => n11948, ZN => 
                           n11949);
   U11186 : NAND2_X1 port map( A1 => n11857, A2 => n3943, ZN => n10954);
   U11187 : AND2_X1 port map( A1 => n11952, A2 => n3946, ZN => n3943);
   U11188 : NAND2_X1 port map( A1 => n11556, A2 => n3945, ZN => n3944);
   U11189 : AND2_X1 port map( A1 => n11943, A2 => n3946, ZN => n3945);
   U11190 : INV_X1 port map( A => n14346, ZN => n14136);
   U11192 : NAND2_X1 port map( A1 => n14134, A2 => n3948, ZN => n3947);
   U11193 : OR2_X1 port map( A1 => n14346, A2 => n3949, ZN => n3948);
   U11194 : NAND2_X1 port map( A1 => n13842, A2 => n14010, ZN => n3949);
   U11195 : INV_X1 port map( A => n13843, ZN => n3950);
   U11196 : NAND2_X1 port map( A1 => n20633, A2 => n28538, ZN => n3954);
   U11197 : NAND2_X1 port map( A1 => n20456, A2 => n1908, ZN => n3951);
   U11198 : INV_X1 port map( A => n20453, ZN => n20633);
   U11199 : XNOR2_X1 port map( A => n12420, B => n13175, ZN => n13287);
   U11201 : NAND2_X1 port map( A1 => n3962, A2 => n12151, ZN => n3955);
   U11202 : NAND2_X1 port map( A1 => n3957, A2 => n12991, ZN => n3956);
   U11203 : NAND2_X1 port map( A1 => n12994, A2 => n3958, ZN => n3957);
   U11205 : NAND2_X1 port map( A1 => n430, A2 => n579, ZN => n3960);
   U11206 : NOR2_X1 port map( A1 => n12150, A2 => n3961, ZN => n3962);
   U11207 : INV_X1 port map( A => n12088, ZN => n3961);
   U11208 : NAND4_X1 port map( A1 => n4843, A2 => n3966, A3 => n3965, A4 => 
                           n3963, ZN => n4842);
   U11209 : NOR2_X1 port map( A1 => n12200, A2 => n12201, ZN => n3964);
   U11210 : NAND2_X1 port map( A1 => n12202, A2 => n4844, ZN => n3965);
   U11211 : NAND2_X1 port map( A1 => n12201, A2 => n12203, ZN => n3966);
   U11212 : INV_X1 port map( A => n3968, ZN => n3967);
   U11213 : OAI21_X1 port map( B1 => n19794, B2 => n20517, A => n3969, ZN => 
                           n3968);
   U11216 : INV_X1 port map( A => n20584, ZN => n3973);
   U11217 : OAI21_X1 port map( B1 => n20590, B2 => n3975, A => n20589, ZN => 
                           n21135);
   U11218 : NAND2_X1 port map( A1 => n20590, A2 => n20589, ZN => n3971);
   U11219 : NAND2_X1 port map( A1 => n3975, A2 => n20589, ZN => n3972);
   U11220 : INV_X1 port map( A => n19828, ZN => n3975);
   U11221 : NAND2_X1 port map( A1 => n14258, A2 => n6921, ZN => n3976);
   U11222 : NAND2_X1 port map( A1 => n14761, A2 => n15260, ZN => n3978);
   U11223 : NAND3_X1 port map( A1 => n29737, A2 => n4246, A3 => n1666, ZN => 
                           n3980);
   U11225 : XNOR2_X1 port map( A => n22100, B => n3984, ZN => n3983);
   U11226 : INV_X1 port map( A => n22655, ZN => n3984);
   U11227 : NAND2_X1 port map( A1 => n23437, A2 => n23436, ZN => n3985);
   U11228 : MUX2_X1 port map( A => n24972, B => n24973, S => n24509, Z => 
                           n23600);
   U11230 : NAND3_X1 port map( A1 => n574, A2 => n11922, A3 => n11549, ZN => 
                           n3987);
   U11231 : AOI21_X1 port map( B1 => n11547, B2 => n11922, A => n11927, ZN => 
                           n3989);
   U11233 : NAND2_X1 port map( A1 => n2968, A2 => n10919, ZN => n3992);
   U11234 : OAI21_X1 port map( B1 => n18277, B2 => n3995, A => n3993, ZN => 
                           n3996);
   U11235 : NAND2_X1 port map( A1 => n3994, A2 => n18277, ZN => n3993);
   U11236 : INV_X1 port map( A => n18204, ZN => n3994);
   U11237 : AOI22_X2 port map( A1 => n18206, A2 => n3997, B1 => n3996, B2 => 
                           n18279, ZN => n19194);
   U11239 : NAND2_X1 port map( A1 => n18275, A2 => n17696, ZN => n3997);
   U11240 : NAND2_X1 port map( A1 => n578, A2 => n11869, ZN => n3998);
   U11241 : NAND2_X1 port map( A1 => n6181, A2 => n11500, ZN => n11750);
   U11242 : NAND2_X1 port map( A1 => n11868, A2 => n11867, ZN => n3999);
   U11244 : NAND2_X1 port map( A1 => n373, A2 => n4002, ZN => n5328);
   U11245 : NAND2_X1 port map( A1 => n29620, A2 => n23762, ZN => n23476);
   U11246 : NAND2_X1 port map( A1 => n23759, A2 => n29620, ZN => n5743);
   U11247 : XNOR2_X1 port map( A => n15946, B => n15945, ZN => n17276);
   U11249 : NAND3_X1 port map( A1 => n17271, A2 => n17275, A3 => n6465, ZN => 
                           n4004);
   U11250 : OAI211_X1 port map( C1 => n414, C2 => n20089, A => n4007, B => 
                           n4006, ZN => n20095);
   U11251 : NAND2_X1 port map( A1 => n4008, A2 => n29104, ZN => n4007);
   U11252 : NAND2_X1 port map( A1 => n20039, A2 => n29114, ZN => n4008);
   U11254 : XNOR2_X2 port map( A => n18717, B => n18716, ZN => n20041);
   U11255 : AOI22_X1 port map( A1 => n4012, A2 => n4010, B1 => n2549, B2 => 
                           n4009, ZN => n13708);
   U11256 : NAND2_X1 port map( A1 => n21078, A2 => n20933, ZN => n21077);
   U11257 : NAND2_X1 port map( A1 => n4015, A2 => n4014, ZN => n4013);
   U11258 : NAND3_X1 port map( A1 => n26450, A2 => n26179, A3 => n26447, ZN => 
                           n4014);
   U11259 : NAND2_X1 port map( A1 => n25625, A2 => n26456, ZN => n4015);
   U11260 : AOI22_X2 port map( A1 => n16956, A2 => n16955, B1 => n16957, B2 => 
                           n18259, ZN => n19085);
   U11261 : NAND3_X1 port map( A1 => n6706, A2 => n4341, A3 => n571, ZN => 
                           n4016);
   U11263 : NAND2_X1 port map( A1 => n11180, A2 => n11179, ZN => n11955);
   U11264 : XNOR2_X1 port map( A => n6939, B => n22667, ZN => n23305);
   U11265 : INV_X1 port map( A => n11982, ZN => n13083);
   U11266 : OAI21_X1 port map( B1 => n11811, B2 => n4021, A => n11810, ZN => 
                           n11814);
   U11269 : MUX2_X1 port map( A => n7665, B => n8264, S => n8270, Z => n4022);
   U11270 : XNOR2_X2 port map( A => Key(146), B => Plaintext(146), ZN => n8270)
                           ;
   U11271 : AOI21_X1 port map( B1 => n10507, B2 => n4023, A => n11124, ZN => 
                           n10508);
   U11272 : NAND2_X1 port map( A1 => n4024, A2 => n11120, ZN => n4023);
   U11273 : INV_X1 port map( A => n11123, ZN => n4024);
   U11274 : XNOR2_X2 port map( A => n9885, B => n9884, ZN => n11123);
   U11275 : OR2_X1 port map( A1 => n6095, A2 => n27525, ZN => n27510);
   U11277 : OAI21_X1 port map( B1 => n27510, B2 => n27531, A => n3067, ZN => 
                           n27511);
   U11278 : INV_X1 port map( A => n24677, ZN => n24322);
   U11279 : NAND2_X1 port map( A1 => n20324, A2 => n20109, ZN => n20321);
   U11280 : XNOR2_X2 port map( A => n19589, B => n19588, ZN => n20109);
   U11281 : INV_X1 port map( A => n14487, ZN => n12120);
   U11282 : OAI21_X1 port map( B1 => n14167, B2 => n14164, A => n4027, ZN => 
                           n4026);
   U11283 : NAND3_X1 port map( A1 => n12120, A2 => n14484, A3 => n29565, ZN => 
                           n4027);
   U11284 : NAND2_X1 port map( A1 => n4028, A2 => n2483, ZN => n12195);
   U11285 : NAND2_X1 port map( A1 => n4028, A2 => n12128, ZN => n11727);
   U11287 : OR2_X1 port map( A1 => n12127, A2 => n4028, ZN => n4982);
   U11288 : XNOR2_X1 port map( A => n4031, B => n2505, ZN => n12848);
   U11289 : XNOR2_X1 port map( A => n4031, B => n13414, ZN => n12908);
   U11290 : XNOR2_X1 port map( A => n4031, B => n13269, ZN => n13412);
   U11291 : XNOR2_X1 port map( A => n12826, B => n4031, ZN => n12829);
   U11292 : XNOR2_X1 port map( A => n12780, B => n4031, ZN => n12117);
   U11293 : XNOR2_X1 port map( A => n12637, B => n4031, ZN => n12385);
   U11294 : OAI211_X2 port map( C1 => n12115, C2 => n12114, A => n12113, B => 
                           n12112, ZN => n4031);
   U11297 : NOR2_X1 port map( A1 => n27380, A2 => n28394, ZN => n4035);
   U11298 : INV_X1 port map( A => n26610, ZN => n4036);
   U11299 : NOR2_X1 port map( A1 => n4038, A2 => n12211, ZN => n9655);
   U11302 : MUX2_X1 port map( A => n14808, B => n14810, S => n14775, Z => 
                           n14229);
   U11303 : NAND2_X1 port map( A1 => n11428, A2 => n11426, ZN => n4046);
   U11304 : INV_X1 port map( A => n14192, ZN => n14395);
   U11305 : OR2_X1 port map( A1 => n14393, A2 => n14192, ZN => n14195);
   U11306 : OAI211_X1 port map( C1 => n28805, C2 => n14395, A => n14393, B => 
                           n4047, ZN => n4048);
   U11308 : NOR2_X1 port map( A1 => n14192, A2 => n14194, ZN => n4049);
   U11309 : OR2_X1 port map( A1 => n7116, A2 => n7320, ZN => n4052);
   U11310 : NAND2_X1 port map( A1 => n20252, A2 => n1951, ZN => n4053);
   U11311 : NAND2_X1 port map( A1 => n21631, A2 => n21036, ZN => n21039);
   U11312 : INV_X1 port map( A => n14593, ZN => n4054);
   U11313 : NAND2_X1 port map( A1 => n13783, A2 => n4055, ZN => n4151);
   U11314 : NOR2_X1 port map( A1 => n14593, A2 => n4056, ZN => n4055);
   U11315 : INV_X1 port map( A => n14105, ZN => n4056);
   U11316 : NAND2_X1 port map( A1 => n14594, A2 => n14593, ZN => n14258);
   U11317 : NAND3_X2 port map( A1 => n4057, A2 => n10536, A3 => n10537, ZN => 
                           n13563);
   U11318 : NAND2_X1 port map( A1 => n10531, A2 => n12333, ZN => n4057);
   U11319 : INV_X1 port map( A => n13563, ZN => n13178);
   U11320 : NAND2_X1 port map( A1 => n464, A2 => n24507, ZN => n4063);
   U11321 : INV_X1 port map( A => n24269, ZN => n24789);
   U11322 : NAND2_X1 port map( A1 => n1955, A2 => n4065, ZN => n4064);
   U11323 : NAND2_X1 port map( A1 => n4576, A2 => n4066, ZN => n4065);
   U11324 : NAND2_X1 port map( A1 => n23655, A2 => n24269, ZN => n4066);
   U11325 : NAND2_X1 port map( A1 => n1854, A2 => n4067, ZN => n4068);
   U11326 : MUX2_X1 port map( A => n11282, B => n10884, S => n11281, Z => n4067
                           );
   U11327 : XNOR2_X2 port map( A => n10369, B => n10370, ZN => n10884);
   U11330 : XNOR2_X1 port map( A => n19681, B => n4069, ZN => n19432);
   U11331 : XNOR2_X1 port map( A => n18653, B => n4070, ZN => n4069);
   U11332 : NAND3_X1 port map( A1 => n4071, A2 => n21040, A3 => n21748, ZN => 
                           n5976);
   U11333 : AND2_X1 port map( A1 => n15342, A2 => n15224, ZN => n14757);
   U11335 : NAND3_X1 port map( A1 => n26131, A2 => n4079, A3 => n4078, ZN => 
                           n27724);
   U11336 : NAND3_X1 port map( A1 => n27129, A2 => n28536, A3 => n27177, ZN => 
                           n4078);
   U11337 : NAND2_X1 port map( A1 => n27173, A2 => n4080, ZN => n4079);
   U11338 : OAI21_X2 port map( B1 => n23307, B2 => n23306, A => n4081, ZN => 
                           n25884);
   U11339 : XNOR2_X1 port map( A => n25347, B => n4083, ZN => n4082);
   U11340 : XNOR2_X1 port map( A => n25346, B => n25345, ZN => n4083);
   U11341 : XNOR2_X1 port map( A => n25348, B => n25713, ZN => n4084);
   U11342 : XNOR2_X2 port map( A => n16118, B => n16117, ZN => n17259);
   U11344 : AOI21_X1 port map( B1 => n4086, B2 => n23531, A => n28164, ZN => 
                           n4124);
   U11345 : OAI21_X1 port map( B1 => n484, B2 => n23067, A => n4086, ZN => 
                           n5402);
   U11346 : NAND2_X1 port map( A1 => n28164, A2 => n4086, ZN => n6903);
   U11347 : OAI22_X1 port map( A1 => n5029, A2 => n4086, B1 => n23135, B2 => 
                           n23535, ZN => n5031);
   U11348 : NAND2_X1 port map( A1 => n10627, A2 => n11014, ZN => n4087);
   U11349 : INV_X1 port map( A => n13824, ZN => n4088);
   U11350 : XNOR2_X2 port map( A => n13053, B => n13052, ZN => n13060);
   U11351 : NAND2_X1 port map( A1 => n29373, A2 => n17491, ZN => n17063);
   U11353 : NAND2_X1 port map( A1 => n17063, A2 => n16882, ZN => n4089);
   U11354 : NAND2_X1 port map( A1 => n4092, A2 => n4091, ZN => n4090);
   U11355 : NAND3_X1 port map( A1 => n27382, A2 => n28394, A3 => n27213, ZN => 
                           n4092);
   U11356 : NAND2_X1 port map( A1 => n4093, A2 => n21304, ZN => n6733);
   U11357 : NAND2_X1 port map( A1 => n21150, A2 => n4094, ZN => n4093);
   U11358 : NAND2_X1 port map( A1 => n21311, A2 => n20938, ZN => n4094);
   U11359 : NAND2_X1 port map( A1 => n11292, A2 => n11291, ZN => n4095);
   U11360 : MUX2_X1 port map( A => n11795, B => n12081, S => n29498, Z => 
                           n11799);
   U11362 : NAND2_X1 port map( A1 => n17219, A2 => n17555, ZN => n4100);
   U11364 : NAND3_X1 port map( A1 => n4982, A2 => n12131, A3 => n4981, ZN => 
                           n4102);
   U11365 : INV_X1 port map( A => n21493, ZN => n4104);
   U11366 : OAI21_X1 port map( B1 => n21183, B2 => n21495, A => n4104, ZN => 
                           n4103);
   U11367 : NAND3_X1 port map( A1 => n21186, A2 => n6503, A3 => n4103, ZN => 
                           n6504);
   U11368 : NAND2_X1 port map( A1 => n4105, A2 => n12280, ZN => n11359);
   U11369 : OR2_X1 port map( A1 => n12408, A2 => n4106, ZN => n11627);
   U11370 : NAND2_X1 port map( A1 => n12281, A2 => n12402, ZN => n4106);
   U11371 : NAND3_X1 port map( A1 => n4105, A2 => n12400, A3 => n11801, ZN => 
                           n11626);
   U11372 : NAND3_X1 port map( A1 => n4105, A2 => n12400, A3 => n12407, ZN => 
                           n12067);
   U11373 : OAI21_X1 port map( B1 => n12286, B2 => n4105, A => n12400, ZN => 
                           n12405);
   U11374 : NOR2_X1 port map( A1 => n11333, A2 => n4107, ZN => n4461);
   U11375 : NAND2_X1 port map( A1 => n10466, A2 => n4107, ZN => n10469);
   U11378 : NAND3_X1 port map( A1 => n27193, A2 => n4243, A3 => n4109, ZN => 
                           n4108);
   U11379 : NAND2_X1 port map( A1 => n8155, A2 => n8154, ZN => n4111);
   U11380 : NAND2_X1 port map( A1 => n2056, A2 => n17393, ZN => n4113);
   U11381 : NAND2_X1 port map( A1 => n4116, A2 => n4115, ZN => n4114);
   U11382 : NAND3_X1 port map( A1 => n4117, A2 => n12201, A3 => n12202, ZN => 
                           n4115);
   U11383 : NAND2_X1 port map( A1 => n11602, A2 => n5825, ZN => n4116);
   U11384 : NAND2_X1 port map( A1 => n1966, A2 => n2063, ZN => n4117);
   U11385 : INV_X1 port map( A => n12202, ZN => n6020);
   U11386 : NAND3_X1 port map( A1 => n17986, A2 => n17985, A3 => n18268, ZN => 
                           n4120);
   U11387 : MUX2_X1 port map( A => n13842, B => n14010, S => n14131, Z => n4122
                           );
   U11389 : NAND2_X1 port map( A1 => n11348, A2 => n11192, ZN => n4123);
   U11390 : AOI21_X1 port map( B1 => n4123, B2 => n9219, A => n9218, ZN => 
                           n9257);
   U11391 : XNOR2_X2 port map( A => n19737, B => n19738, ZN => n23535);
   U11392 : INV_X1 port map( A => n10547, ZN => n4126);
   U11393 : NAND3_X1 port map( A1 => n11111, A2 => n242, A3 => n10492, ZN => 
                           n4127);
   U11394 : NAND2_X1 port map( A1 => n4056, A2 => n14107, ZN => n13608);
   U11395 : NAND2_X1 port map( A1 => n14230, A2 => n4056, ZN => n14103);
   U11396 : MUX2_X1 port map( A => n14107, B => n4056, S => n14231, Z => n11371
                           );
   U11397 : NAND3_X1 port map( A1 => n4150, A2 => n14231, A3 => n4056, ZN => 
                           n4149);
   U11398 : NAND3_X1 port map( A1 => n4129, A2 => n7728, A3 => n7727, ZN => 
                           n7731);
   U11399 : NAND2_X1 port map( A1 => n27033, A2 => n27032, ZN => n4130);
   U11400 : NAND2_X1 port map( A1 => n27030, A2 => n4133, ZN => n4132);
   U11401 : INV_X1 port map( A => n28592, ZN => n4133);
   U11402 : NAND2_X1 port map( A1 => n24713, A2 => n24716, ZN => n4135);
   U11403 : NAND2_X1 port map( A1 => n23060, A2 => n23344, ZN => n4137);
   U11404 : NAND2_X1 port map( A1 => n23059, A2 => n29108, ZN => n4138);
   U11405 : INV_X1 port map( A => n13552, ZN => n4139);
   U11406 : XNOR2_X1 port map( A => n4139, B => n12566, ZN => n11684);
   U11408 : NAND3_X2 port map( A1 => n21228, A2 => n4142, A3 => n2022, ZN => 
                           n6141);
   U11409 : INV_X1 port map( A => n21639, ZN => n4143);
   U11410 : NAND3_X1 port map( A1 => n28797, A2 => n4143, A3 => n21638, ZN => 
                           n4142);
   U11411 : INV_X1 port map( A => n12017, ZN => n12016);
   U11412 : NAND2_X1 port map( A1 => n11747, A2 => n12328, ZN => n12017);
   U11413 : OAI211_X1 port map( C1 => n10523, C2 => n11038, A => n28612, B => 
                           n11275, ZN => n4145);
   U11414 : NAND2_X1 port map( A1 => n10525, A2 => n29148, ZN => n4146);
   U11415 : INV_X1 port map( A => n4148, ZN => n21613);
   U11416 : OR2_X2 port map( A1 => n20492, A2 => n21329, ZN => n4148);
   U11417 : NAND2_X1 port map( A1 => n4148, A2 => n21327, ZN => n21618);
   U11418 : AND2_X1 port map( A1 => n28791, A2 => n21613, ZN => n20910);
   U11419 : NAND2_X1 port map( A1 => n4148, A2 => n21326, ZN => n20906);
   U11420 : NAND2_X1 port map( A1 => n4147, A2 => n21163, ZN => n20732);
   U11421 : AND2_X1 port map( A1 => n28791, A2 => n4148, ZN => n4147);
   U11422 : NAND3_X1 port map( A1 => n4151, A2 => n4149, A3 => n13784, ZN => 
                           n14928);
   U11423 : INV_X1 port map( A => n14107, ZN => n13783);
   U11424 : INV_X1 port map( A => n4152, ZN => n4153);
   U11425 : INV_X1 port map( A => n17771, ZN => n17583);
   U11427 : NAND3_X1 port map( A1 => n4157, A2 => n4158, A3 => n4156, ZN => 
                           n4154);
   U11428 : MUX2_X1 port map( A => n17575, B => n17574, S => n17707, Z => n4155
                           );
   U11429 : NAND2_X1 port map( A1 => n17707, A2 => n17570, ZN => n4158);
   U11430 : XNOR2_X1 port map( A => n4161, B => n25454, ZN => n24948);
   U11431 : XNOR2_X1 port map( A => n4161, B => n25855, ZN => n25857);
   U11432 : XNOR2_X1 port map( A => n4161, B => n4384, ZN => n25479);
   U11433 : XNOR2_X1 port map( A => n25944, B => n4161, ZN => n25094);
   U11435 : OAI21_X1 port map( B1 => n15055, B2 => n15054, A => n4162, ZN => 
                           n14764);
   U11438 : NAND2_X1 port map( A1 => n27508, A2 => n29556, ZN => n4165);
   U11439 : NAND2_X1 port map( A1 => n4166, A2 => n14278, ZN => n14274);
   U11440 : NAND2_X1 port map( A1 => n14362, A2 => n4166, ZN => n4667);
   U11442 : NAND2_X1 port map( A1 => n6188, A2 => n9037, ZN => n6190);
   U11443 : NAND3_X1 port map( A1 => n424, A2 => n16878, A3 => n29045, ZN => 
                           n4168);
   U11444 : NAND3_X1 port map( A1 => n15072, A2 => n15071, A3 => n14571, ZN => 
                           n4169);
   U11445 : NAND2_X1 port map( A1 => n4172, A2 => n20125, ZN => n18546);
   U11446 : OAI21_X1 port map( B1 => n20294, B2 => n20293, A => n4172, ZN => 
                           n20296);
   U11447 : NAND2_X1 port map( A1 => n20293, A2 => n19815, ZN => n4172);
   U11448 : AOI21_X1 port map( B1 => n26230, B2 => n26740, A => n26229, ZN => 
                           n26231);
   U11449 : NAND2_X1 port map( A1 => n25598, A2 => n26740, ZN => n25600);
   U11450 : NAND2_X1 port map( A1 => n25349, A2 => n26740, ZN => n4173);
   U11451 : NAND2_X1 port map( A1 => n4174, A2 => n18198, ZN => n16719);
   U11452 : NOR2_X1 port map( A1 => n4174, A2 => n18449, ZN => n6326);
   U11453 : INV_X1 port map( A => n23302, ZN => n4178);
   U11455 : NAND2_X1 port map( A1 => n7496, A2 => n7250, ZN => n7254);
   U11456 : NAND2_X1 port map( A1 => n7494, A2 => n7250, ZN => n7251);
   U11457 : OAI21_X1 port map( B1 => n7250, B2 => n7498, A => n7496, ZN => 
                           n4180);
   U11458 : NAND2_X1 port map( A1 => n7705, A2 => n7250, ZN => n7497);
   U11460 : NAND2_X1 port map( A1 => n4186, A2 => n14841, ZN => n4185);
   U11461 : NAND2_X1 port map( A1 => n6048, A2 => n14842, ZN => n4186);
   U11463 : NAND2_X1 port map( A1 => n4188, A2 => n16805, ZN => n16807);
   U11464 : INV_X1 port map( A => n17260, ZN => n4188);
   U11465 : NAND2_X1 port map( A1 => n6408, A2 => n414, ZN => n4189);
   U11466 : NAND2_X1 port map( A1 => n20040, A2 => n20039, ZN => n4190);
   U11467 : NAND2_X1 port map( A1 => n17958, A2 => n6914, ZN => n4192);
   U11468 : OAI211_X2 port map( C1 => n17473, C2 => n17472, A => n17471, B => 
                           n17515, ZN => n18216);
   U11469 : NAND2_X1 port map( A1 => n21567, A2 => n4193, ZN => n21462);
   U11470 : NOR2_X1 port map( A1 => n4193, A2 => n21567, ZN => n21572);
   U11471 : AND2_X1 port map( A1 => n4494, A2 => n4193, ZN => n21568);
   U11472 : NAND2_X1 port map( A1 => n5176, A2 => n4193, ZN => n5175);
   U11473 : OAI21_X1 port map( B1 => n24075, B2 => n4195, A => n4194, ZN => 
                           n24670);
   U11475 : INV_X1 port map( A => n12305, ZN => n12299);
   U11476 : OAI21_X2 port map( B1 => n6774, B2 => n10959, A => n6773, ZN => 
                           n12305);
   U11479 : NAND2_X1 port map( A1 => n21183, A2 => n21497, ZN => n4201);
   U11480 : NAND2_X1 port map( A1 => n20751, A2 => n7, ZN => n4202);
   U11481 : NAND2_X1 port map( A1 => n20752, A2 => n4104, ZN => n4206);
   U11482 : XNOR2_X2 port map( A => n13424, B => n13423, ZN => n13725);
   U11483 : NAND3_X1 port map( A1 => n14372, A2 => n5404, A3 => n14373, ZN => 
                           n6614);
   U11484 : INV_X1 port map( A => n17694, ZN => n4209);
   U11485 : NAND2_X1 port map( A1 => n17692, A2 => n18509, ZN => n4210);
   U11486 : INV_X1 port map( A => n18512, ZN => n4211);
   U11487 : NAND2_X1 port map( A1 => n17691, A2 => n18512, ZN => n4212);
   U11488 : NOR2_X1 port map( A1 => n4213, A2 => n18333, ZN => n4214);
   U11489 : XNOR2_X1 port map( A => n4216, B => n1998, ZN => n4215);
   U11490 : XNOR2_X1 port map( A => n15612, B => n1967, ZN => n4216);
   U11491 : OR2_X1 port map( A1 => n17549, A2 => n4218, ZN => n17241);
   U11492 : NOR2_X1 port map( A1 => n17239, A2 => n4218, ZN => n15685);
   U11493 : NAND3_X1 port map( A1 => n2122, A2 => n17548, A3 => n4218, ZN => 
                           n17550);
   U11494 : AOI21_X1 port map( B1 => n5398, B2 => n4218, A => n16762, ZN => 
                           n17240);
   U11495 : OR2_X2 port map( A1 => n12097, A2 => n10784, ZN => n12151);
   U11496 : NAND4_X2 port map( A1 => n6149, A2 => n4219, A3 => n26437, A4 => 
                           n6148, ZN => n27301);
   U11497 : NAND3_X1 port map( A1 => n456, A2 => n26944, A3 => n26768, ZN => 
                           n4219);
   U11501 : XNOR2_X1 port map( A => n4221, B => n19702, ZN => n19454);
   U11502 : NAND2_X1 port map( A1 => n21561, A2 => n21113, ZN => n4223);
   U11503 : NAND2_X1 port map( A1 => n6861, A2 => n1897, ZN => n4225);
   U11504 : MUX2_X1 port map( A => n4227, B => n26336, S => n27123, Z => n26337
                           );
   U11505 : INV_X1 port map( A => n27191, ZN => n4227);
   U11507 : NAND2_X1 port map( A1 => n18107, A2 => n18106, ZN => n4230);
   U11508 : NAND2_X1 port map( A1 => n18789, A2 => n29114, ZN => n6400);
   U11511 : INV_X1 port map( A => n19985, ZN => n20164);
   U11512 : NOR2_X1 port map( A1 => n24631, A2 => n24630, ZN => n24294);
   U11513 : NAND2_X1 port map( A1 => n27038, A2 => n5581, ZN => n4236);
   U11515 : NOR2_X1 port map( A1 => n5314, A2 => n27213, ZN => n27380);
   U11518 : NAND2_X1 port map( A1 => n24632, A2 => n6867, ZN => n4239);
   U11519 : INV_X1 port map( A => n21388, ZN => n4242);
   U11520 : INV_X1 port map( A => n27124, ZN => n4243);
   U11521 : NAND2_X1 port map( A1 => n20449, A2 => n4245, ZN => n19573);
   U11522 : NAND2_X1 port map( A1 => n5377, A2 => n4245, ZN => n19899);
   U11523 : NOR2_X1 port map( A1 => n19927, A2 => n4245, ZN => n19930);
   U11524 : OAI21_X1 port map( B1 => n6203, B2 => n4245, A => n20451, ZN => 
                           n5375);
   U11525 : XNOR2_X2 port map( A => n16175, B => n16174, ZN => n4246);
   U11526 : NAND2_X1 port map( A1 => n4246, A2 => n17464, ZN => n16675);
   U11527 : NOR2_X1 port map( A1 => n17467, A2 => n4246, ZN => n16819);
   U11528 : NAND2_X1 port map( A1 => n17467, A2 => n4246, ZN => n17093);
   U11529 : OAI21_X1 port map( B1 => n29022, B2 => n29118, A => n4247, ZN => 
                           n6490);
   U11530 : NAND2_X1 port map( A1 => n29022, A2 => n27772, ZN => n4247);
   U11531 : NAND2_X1 port map( A1 => n4247, A2 => n4248, ZN => n27776);
   U11533 : NAND2_X1 port map( A1 => n27784, A2 => n4250, ZN => n27770);
   U11534 : NAND2_X1 port map( A1 => n14033, A2 => n14030, ZN => n13794);
   U11535 : NAND3_X1 port map( A1 => n14033, A2 => n14030, A3 => n14029, ZN => 
                           n4252);
   U11536 : XNOR2_X1 port map( A => n4253, B => n12931, ZN => n13457);
   U11537 : XNOR2_X1 port map( A => n4253, B => n2894, ZN => n11389);
   U11538 : XNOR2_X1 port map( A => n4253, B => n6683, ZN => n12705);
   U11539 : XNOR2_X1 port map( A => n4253, B => n12960, ZN => n12962);
   U11540 : XNOR2_X1 port map( A => n13222, B => n4253, ZN => n13223);
   U11541 : NAND2_X1 port map( A1 => n21118, A2 => n29581, ZN => n20650);
   U11542 : MUX2_X1 port map( A => n21145, B => n21118, S => n21144, Z => 
                           n19784);
   U11543 : NOR2_X1 port map( A1 => n13572, A2 => n14380, ZN => n4258);
   U11544 : NAND2_X1 port map( A1 => n556, A2 => n14004, ZN => n14379);
   U11545 : XNOR2_X2 port map( A => n13560, B => n13561, ZN => n14004);
   U11546 : NAND2_X1 port map( A1 => n8642, A2 => n8984, ZN => n8456);
   U11547 : NAND3_X1 port map( A1 => n8642, A2 => n8984, A3 => n8981, ZN => 
                           n8987);
   U11548 : NAND2_X1 port map( A1 => n13729, A2 => n13914, ZN => n4260);
   U11549 : XNOR2_X1 port map( A => n4263, B => n25515, ZN => n24923);
   U11550 : XNOR2_X1 port map( A => n4263, B => n26108, ZN => n25877);
   U11551 : NAND2_X1 port map( A1 => n11677, A2 => n11515, ZN => n11517);
   U11552 : AOI21_X1 port map( B1 => n10746, B2 => n10819, A => n28208, ZN => 
                           n11633);
   U11553 : NAND3_X1 port map( A1 => n10976, A2 => n4264, A3 => n28608, ZN => 
                           n6896);
   U11554 : INV_X1 port map( A => n10972, ZN => n4264);
   U11555 : INV_X1 port map( A => n19732, ZN => n4266);
   U11556 : OAI21_X1 port map( B1 => n21379, B2 => n21810, A => n4266, ZN => 
                           n21381);
   U11557 : NAND2_X1 port map( A1 => n4270, A2 => n17484, ZN => n4269);
   U11558 : AOI21_X1 port map( B1 => n17831, B2 => n17830, A => n4272, ZN => 
                           n17832);
   U11562 : NAND3_X1 port map( A1 => n11146, A2 => n28206, A3 => n10544, ZN => 
                           n4275);
   U11563 : NAND2_X1 port map( A1 => n12071, A2 => n12070, ZN => n4276);
   U11564 : NAND2_X1 port map( A1 => n19808, A2 => n20137, ZN => n4278);
   U11565 : OAI21_X1 port map( B1 => n4283, B2 => n16953, A => n4279, ZN => 
                           n4282);
   U11567 : NAND2_X1 port map( A1 => n4282, A2 => n28793, ZN => n4280);
   U11568 : NAND2_X1 port map( A1 => n18539, A2 => n18260, ZN => n16955);
   U11569 : NAND2_X1 port map( A1 => n16952, A2 => n17354, ZN => n4281);
   U11570 : INV_X1 port map( A => n14376, ZN => n13594);
   U11571 : NAND2_X1 port map( A1 => n14533, A2 => n15190, ZN => n14531);
   U11572 : NAND2_X1 port map( A1 => n13814, A2 => n4284, ZN => n14784);
   U11573 : NAND3_X1 port map( A1 => n29737, A2 => n387, A3 => n17467, ZN => 
                           n4285);
   U11574 : XNOR2_X1 port map( A => n6080, B => n16414, ZN => n16454);
   U11575 : NAND2_X1 port map( A1 => n14577, A2 => n14936, ZN => n4287);
   U11576 : NAND2_X1 port map( A1 => n14576, A2 => n549, ZN => n4288);
   U11577 : AND2_X1 port map( A1 => n28806, A2 => n14460, ZN => n14458);
   U11578 : MUX2_X1 port map( A => n4290, B => n14204, S => n28806, Z => n13864
                           );
   U11580 : INV_X1 port map( A => n12712, ZN => n4290);
   U11581 : NAND2_X1 port map( A1 => n380, A2 => n23712, ZN => n6153);
   U11582 : NAND2_X2 port map( A1 => n4291, A2 => n4293, ZN => n18382);
   U11584 : OAI21_X1 port map( B1 => n18351, B2 => n18383, A => n18350, ZN => 
                           n5920);
   U11585 : NAND2_X1 port map( A1 => n4295, A2 => n16712, ZN => n4294);
   U11586 : INV_X1 port map( A => n11317, ZN => n4815);
   U11587 : NAND2_X1 port map( A1 => n4296, A2 => n11253, ZN => n11317);
   U11588 : XNOR2_X1 port map( A => n4298, B => n13433, ZN => n13362);
   U11589 : XNOR2_X1 port map( A => n12064, B => n4297, ZN => n12972);
   U11590 : XNOR2_X1 port map( A => n12808, B => n4298, ZN => n11563);
   U11591 : NAND2_X1 port map( A1 => n23261, A2 => n23712, ZN => n23235);
   U11592 : OAI21_X2 port map( B1 => n4299, B2 => n14994, A => n14993, ZN => 
                           n16444);
   U11594 : NAND2_X1 port map( A1 => n4303, A2 => n9202, ZN => n4302);
   U11596 : NAND2_X1 port map( A1 => n8994, A2 => n4305, ZN => n4304);
   U11597 : INV_X1 port map( A => n8995, ZN => n4305);
   U11598 : NAND2_X1 port map( A1 => n3900, A2 => n11553, ZN => n6742);
   U11599 : NAND2_X1 port map( A1 => n20458, A2 => n4306, ZN => n20459);
   U11600 : NOR2_X1 port map( A1 => n20458, A2 => n4306, ZN => n20027);
   U11603 : INV_X1 port map( A => n22401, ZN => n22398);
   U11604 : OR2_X2 port map( A1 => n20264, A2 => n20263, ZN => n22401);
   U11605 : NAND2_X1 port map( A1 => n4310, A2 => n4308, ZN => n4311);
   U11606 : NAND2_X1 port map( A1 => n5151, A2 => n22401, ZN => n4309);
   U11607 : NAND2_X1 port map( A1 => n22396, A2 => n22398, ZN => n4310);
   U11608 : NAND2_X1 port map( A1 => n17064, A2 => n538, ZN => n4315);
   U11609 : NAND2_X1 port map( A1 => n4315, A2 => n4313, ZN => n17206);
   U11610 : AOI21_X1 port map( B1 => n2549, B2 => n4509, A => n14402, ZN => 
                           n13965);
   U11611 : NAND2_X1 port map( A1 => n17566, A2 => n4316, ZN => n17227);
   U11612 : NAND2_X1 port map( A1 => n17568, A2 => n4316, ZN => n6306);
   U11613 : XNOR2_X1 port map( A => n9823, B => n9824, ZN => n10229);
   U11614 : NAND2_X1 port map( A1 => n4319, A2 => n28743, ZN => n4318);
   U11615 : NAND2_X1 port map( A1 => n4322, A2 => n8366, ZN => n4319);
   U11616 : XNOR2_X1 port map( A => n4323, B => n3378, ZN => n14868);
   U11617 : XNOR2_X1 port map( A => n16606, B => n4323, ZN => n16609);
   U11618 : XNOR2_X1 port map( A => n3661, B => n4323, ZN => n16347);
   U11619 : XNOR2_X1 port map( A => n15780, B => n4323, ZN => n15649);
   U11620 : AOI22_X1 port map( A1 => n4296, A2 => n11318, B1 => n11314, B2 => 
                           n4326, ZN => n4325);
   U11621 : NAND2_X1 port map( A1 => n4296, A2 => n11315, ZN => n4327);
   U11622 : NAND2_X1 port map( A1 => n4329, A2 => n11253, ZN => n4328);
   U11623 : NAND2_X1 port map( A1 => n29059, A2 => n14372, ZN => n14374);
   U11624 : NAND2_X1 port map( A1 => n16918, A2 => n29550, ZN => n4332);
   U11625 : NAND2_X1 port map( A1 => n4335, A2 => n24804, ZN => n4333);
   U11626 : NAND2_X1 port map( A1 => n24805, A2 => n24806, ZN => n4334);
   U11627 : NAND2_X1 port map( A1 => n23689, A2 => n1914, ZN => n23803);
   U11629 : OR2_X1 port map( A1 => n23800, A2 => n23801, ZN => n4337);
   U11630 : OAI211_X1 port map( C1 => n416, C2 => n4340, A => n5436, B => n4338
                           , ZN => n20890);
   U11631 : NAND2_X1 port map( A1 => n4340, A2 => n20302, ZN => n18117);
   U11632 : NAND2_X1 port map( A1 => n20303, A2 => n4340, ZN => n20204);
   U11633 : NAND2_X1 port map( A1 => n4341, A2 => n11194, ZN => n11956);
   U11635 : OAI21_X1 port map( B1 => n21590, B2 => n28584, A => n4342, ZN => 
                           n4343);
   U11636 : NOR2_X1 port map( A1 => n21586, A2 => n21585, ZN => n4344);
   U11638 : NAND2_X1 port map( A1 => n11843, A2 => n4346, ZN => n4345);
   U11639 : NAND2_X1 port map( A1 => n373, A2 => n17858, ZN => n6230);
   U11640 : NAND2_X1 port map( A1 => n12232, A2 => n776, ZN => n11680);
   U11641 : NAND3_X1 port map( A1 => n12232, A2 => n776, A3 => n12236, ZN => 
                           n4349);
   U11642 : INV_X1 port map( A => n10662, ZN => n4350);
   U11643 : INV_X1 port map( A => n10658, ZN => n4351);
   U11644 : AND2_X2 port map( A1 => n4353, A2 => n2078, ZN => n27855);
   U11645 : NAND2_X1 port map( A1 => n26990, A2 => n26321, ZN => n4354);
   U11646 : NAND2_X1 port map( A1 => n27079, A2 => n27074, ZN => n4355);
   U11647 : OAI211_X1 port map( C1 => n4358, C2 => n14840, A => n4357, B => 
                           n4356, ZN => n4360);
   U11648 : NAND2_X1 port map( A1 => n14840, A2 => n4359, ZN => n4356);
   U11649 : NAND2_X1 port map( A1 => n14839, A2 => n4359, ZN => n4357);
   U11650 : INV_X1 port map( A => n15887, ZN => n16436);
   U11651 : NOR2_X1 port map( A1 => n21028, A2 => n21627, ZN => n6530);
   U11652 : INV_X1 port map( A => n24629, ZN => n24293);
   U11653 : NAND2_X1 port map( A1 => n4365, A2 => n4363, ZN => n6198);
   U11654 : NAND3_X1 port map( A1 => n6867, A2 => n24891, A3 => n4364, ZN => 
                           n4363);
   U11655 : INV_X1 port map( A => n4364, ZN => n4366);
   U11657 : NAND2_X1 port map( A1 => n4369, A2 => n14075, ZN => n14830);
   U11659 : INV_X1 port map( A => n7199, ZN => n4370);
   U11660 : NAND2_X1 port map( A1 => n7406, A2 => n8280, ZN => n7199);
   U11661 : OR2_X1 port map( A1 => n17979, A2 => n18234, ZN => n4372);
   U11662 : INV_X1 port map( A => n17979, ZN => n4373);
   U11663 : NAND2_X1 port map( A1 => n18233, A2 => n18398, ZN => n17979);
   U11664 : OAI21_X1 port map( B1 => n18400, B2 => n18398, A => n18401, ZN => 
                           n4374);
   U11665 : NAND3_X1 port map( A1 => n4376, A2 => n13938, A3 => n14237, ZN => 
                           n13940);
   U11666 : OR2_X1 port map( A1 => n491, A2 => n4382, ZN => n4377);
   U11667 : INV_X1 port map( A => n22000, ZN => n22897);
   U11668 : OAI211_X2 port map( C1 => n4380, C2 => n4379, A => n4378, B => 
                           n4377, ZN => n22000);
   U11669 : NAND2_X1 port map( A1 => n4381, A2 => n21823, ZN => n4379);
   U11670 : NAND2_X1 port map( A1 => n495, A2 => n21078, ZN => n4381);
   U11671 : OR2_X1 port map( A1 => n20933, A2 => n22013, ZN => n4382);
   U11672 : AND2_X1 port map( A1 => n10114, A2 => n11124, ZN => n10505);
   U11673 : XNOR2_X1 port map( A => n4384, B => n24060, ZN => n24061);
   U11674 : XNOR2_X1 port map( A => n4384, B => n3334, ZN => n24873);
   U11675 : XNOR2_X1 port map( A => n4384, B => n25947, ZN => n25950);
   U11676 : XNOR2_X1 port map( A => n25149, B => n4384, ZN => n5432);
   U11678 : INV_X1 port map( A => n29102, ZN => n4385);
   U11679 : AND2_X1 port map( A1 => n20041, A2 => n29104, ZN => n6408);
   U11680 : XNOR2_X1 port map( A => n13180, B => n4387, ZN => n12530);
   U11681 : INV_X1 port map( A => n13284, ZN => n4387);
   U11682 : XNOR2_X1 port map( A => n4388, B => n13449, ZN => n13455);
   U11683 : INV_X1 port map( A => n13180, ZN => n4388);
   U11684 : NAND2_X1 port map( A1 => n28206, A2 => n10808, ZN => n10740);
   U11686 : INV_X1 port map( A => n17125, ZN => n4391);
   U11687 : NAND2_X1 port map( A1 => n4392, A2 => n17627, ZN => n6654);
   U11688 : NAND2_X1 port map( A1 => n17626, A2 => n17636, ZN => n4392);
   U11689 : NAND2_X1 port map( A1 => n21146, A2 => n4394, ZN => n4393);
   U11690 : NAND2_X1 port map( A1 => n21144, A2 => n21145, ZN => n4395);
   U11692 : OAI211_X1 port map( C1 => n14341, C2 => n14131, A => n14010, B => 
                           n4396, ZN => n4398);
   U11693 : NAND2_X1 port map( A1 => n14136, A2 => n14131, ZN => n4396);
   U11694 : AOI21_X1 port map( B1 => n20049, B2 => n20067, A => n6477, ZN => 
                           n4403);
   U11695 : OAI21_X1 port map( B1 => n4403, B2 => n20068, A => n6476, ZN => 
                           n20425);
   U11696 : AOI21_X1 port map( B1 => n21076, B2 => n20933, A => n21823, ZN => 
                           n20428);
   U11697 : NAND2_X1 port map( A1 => n12300, A2 => n12305, ZN => n4404);
   U11698 : NAND3_X1 port map( A1 => n11493, A2 => n12307, A3 => n11495, ZN => 
                           n11768);
   U11700 : NAND2_X1 port map( A1 => n10737, A2 => n10914, ZN => n4405);
   U11701 : NAND3_X1 port map( A1 => n18125, A2 => n18588, A3 => n18126, ZN => 
                           n4406);
   U11702 : OAI21_X1 port map( B1 => n18129, B2 => n18127, A => n4406, ZN => 
                           n18133);
   U11703 : OAI21_X1 port map( B1 => n18593, B2 => n18592, A => n4406, ZN => 
                           n18594);
   U11704 : OAI21_X2 port map( B1 => n6813, B2 => n13256, A => n6812, ZN => 
                           n15691);
   U11706 : INV_X1 port map( A => n29058, ZN => n4411);
   U11707 : AOI21_X1 port map( B1 => n28783, B2 => n4411, A => n29570, ZN => 
                           n4486);
   U11708 : NAND2_X1 port map( A1 => n2007, A2 => n28448, ZN => n6476);
   U11709 : INV_X1 port map( A => n20064, ZN => n18765);
   U11710 : INV_X1 port map( A => n17505, ZN => n17073);
   U11711 : INV_X1 port map( A => n17484, ZN => n17074);
   U11712 : NAND2_X1 port map( A1 => n17073, A2 => n17830, ZN => n4413);
   U11713 : NAND2_X1 port map( A1 => n4415, A2 => n407, ZN => n23439);
   U11714 : NAND2_X1 port map( A1 => n4418, A2 => n6207, ZN => n4417);
   U11715 : INV_X1 port map( A => n15260, ZN => n15055);
   U11717 : NAND2_X1 port map( A1 => n17891, A2 => n18600, ZN => n4420);
   U11718 : NAND2_X1 port map( A1 => n13581, A2 => n13900, ZN => n4422);
   U11719 : INV_X1 port map( A => n14144, ZN => n4423);
   U11720 : AOI21_X1 port map( B1 => n4423, B2 => n4425, A => n2974, ZN => 
                           n4424);
   U11721 : NAND2_X1 port map( A1 => n389, A2 => n13902, ZN => n4426);
   U11722 : NAND2_X1 port map( A1 => n12202, A2 => n12203, ZN => n11438);
   U11725 : XNOR2_X2 port map( A => n12838, B => n12837, ZN => n14192);
   U11727 : NAND2_X1 port map( A1 => n8326, A2 => n9425, ZN => n5132);
   U11730 : NAND2_X1 port map( A1 => n7310, A2 => n7092, ZN => n4439);
   U11732 : NAND3_X1 port map( A1 => n4442, A2 => n4441, A3 => n7419, ZN => 
                           n4440);
   U11733 : NAND2_X1 port map( A1 => n8609, A2 => n8751, ZN => n4441);
   U11734 : OAI21_X1 port map( B1 => n29395, B2 => n9532, A => n9531, ZN => 
                           n4442);
   U11735 : XNOR2_X1 port map( A => n12787, B => n12788, ZN => n12949);
   U11737 : NAND2_X1 port map( A1 => n4449, A2 => n4037, ZN => n4447);
   U11738 : NAND2_X1 port map( A1 => n12211, A2 => n12110, ZN => n4448);
   U11739 : NAND2_X1 port map( A1 => n24078, A2 => n24081, ZN => n5272);
   U11740 : OR2_X2 port map( A1 => n6277, A2 => n6278, ZN => n24078);
   U11741 : INV_X1 port map( A => n4450, ZN => n5857);
   U11742 : NOR2_X1 port map( A1 => n18504, A2 => n4450, ZN => n18505);
   U11743 : NAND3_X1 port map( A1 => n4685, A2 => n24809, A3 => n24808, ZN => 
                           n24500);
   U11744 : NOR2_X1 port map( A1 => n29500, A2 => n27069, ZN => n25720);
   U11745 : NAND2_X1 port map( A1 => n27063, A2 => n27069, ZN => n26616);
   U11746 : AOI21_X1 port map( B1 => n14288, B2 => n4451, A => n14287, ZN => 
                           n14289);
   U11747 : XNOR2_X1 port map( A => n15973, B => n15972, ZN => n4452);
   U11748 : XNOR2_X1 port map( A => n15975, B => n16198, ZN => n4453);
   U11750 : XNOR2_X1 port map( A => n16294, B => n3457, ZN => n15558);
   U11751 : NAND4_X2 port map( A1 => n14651, A2 => n4458, A3 => n4457, A4 => 
                           n4456, ZN => n16294);
   U11752 : NAND2_X1 port map( A1 => n14650, A2 => n6879, ZN => n4456);
   U11753 : NAND2_X1 port map( A1 => n15373, A2 => n14863, ZN => n4457);
   U11754 : NAND2_X1 port map( A1 => n4459, A2 => n23529, ZN => n6442);
   U11755 : NAND2_X1 port map( A1 => n21004, A2 => n4460, ZN => n20213);
   U11756 : NOR2_X1 port map( A1 => n23545, A2 => n4231, ZN => n4847);
   U11757 : NAND2_X1 port map( A1 => n5773, A2 => n23351, ZN => n23545);
   U11758 : AOI21_X1 port map( B1 => n20847, B2 => n4464, A => n5142, ZN => 
                           n4465);
   U11759 : NAND2_X1 port map( A1 => n21576, A2 => n21577, ZN => n4464);
   U11760 : NOR2_X1 port map( A1 => n21487, A2 => n21580, ZN => n4467);
   U11762 : XNOR2_X1 port map( A => n4468, B => n27850, ZN => Ciphertext(139));
   U11763 : OAI211_X1 port map( C1 => n27848, C2 => n27849, A => n4470, B => 
                           n4469, ZN => n4468);
   U11764 : NAND2_X1 port map( A1 => n27847, A2 => n2010, ZN => n4469);
   U11765 : NAND2_X1 port map( A1 => n27852, A2 => n27859, ZN => n4470);
   U11769 : NOR2_X1 port map( A1 => n28183, A2 => n23726, ZN => n23848);
   U11770 : XNOR2_X1 port map( A => n4474, B => n12608, ZN => n13510);
   U11771 : INV_X1 port map( A => n13510, ZN => n13038);
   U11772 : NAND2_X1 port map( A1 => n16759, A2 => n17232, ZN => n4476);
   U11773 : NAND2_X1 port map( A1 => n16760, A2 => n4478, ZN => n4477);
   U11774 : XNOR2_X1 port map( A => n4479, B => n3385, ZN => n9955);
   U11775 : XNOR2_X1 port map( A => n4479, B => n10356, ZN => n10015);
   U11776 : XNOR2_X1 port map( A => n4479, B => n10208, ZN => n9631);
   U11777 : NAND3_X1 port map( A1 => n28497, A2 => n17389, A3 => n16879, ZN => 
                           n4480);
   U11778 : XNOR2_X1 port map( A => n4482, B => n29548, ZN => n22581);
   U11779 : XNOR2_X1 port map( A => n22407, B => n22668, ZN => n4482);
   U11780 : NAND2_X1 port map( A1 => n24489, A2 => n24471, ZN => n24493);
   U11781 : NAND2_X1 port map( A1 => n23848, A2 => n23849, ZN => n24093);
   U11782 : OAI211_X1 port map( C1 => n28183, C2 => n23849, A => n23846, B => 
                           n23843, ZN => n4484);
   U11784 : NAND2_X1 port map( A1 => n4487, A2 => n4486, ZN => n4485);
   U11785 : OAI21_X1 port map( B1 => n1530, B2 => n18042, A => n17802, ZN => 
                           n16866);
   U11786 : XNOR2_X1 port map( A => n4489, B => n12833, ZN => n12838);
   U11787 : INV_X1 port map( A => n12834, ZN => n4489);
   U11788 : INV_X1 port map( A => n12833, ZN => n4490);
   U11789 : NAND3_X1 port map( A1 => n15024, A2 => n15023, A3 => n4491, ZN => 
                           n4493);
   U11790 : XNOR2_X1 port map( A => n15862, B => n4492, ZN => n5798);
   U11791 : XNOR2_X1 port map( A => n15862, B => n630, ZN => n16505);
   U11792 : INV_X1 port map( A => n21457, ZN => n4494);
   U11793 : NOR2_X2 port map( A1 => n4495, A2 => n4498, ZN => n27996);
   U11794 : NAND2_X1 port map( A1 => n26633, A2 => n29058, ZN => n4496);
   U11795 : MUX2_X1 port map( A => n27997, B => n27977, S => n27996, Z => 
                           n26636);
   U11796 : MUX2_X1 port map( A => n27045, B => n28130, S => n29058, Z => n4499
                           );
   U11798 : XNOR2_X1 port map( A => n13273, B => n4502, ZN => n12499);
   U11799 : XNOR2_X1 port map( A => n13273, B => n4503, ZN => n12384);
   U11800 : INV_X1 port map( A => n1248, ZN => n4503);
   U11801 : XNOR2_X1 port map( A => n10143, B => n301, ZN => n4508);
   U11802 : XNOR2_X1 port map( A => n10147, B => n10148, ZN => n4506);
   U11803 : MUX2_X1 port map( A => n28804, B => n14400, S => n13877, Z => 
                           n14213);
   U11804 : NAND2_X1 port map( A1 => n13707, A2 => n4509, ZN => n13709);
   U11805 : OAI21_X1 port map( B1 => n4801, B2 => n29148, A => n4511, ZN => 
                           n10480);
   U11806 : NAND2_X1 port map( A1 => n3820, A2 => n29149, ZN => n4511);
   U11807 : OAI211_X1 port map( C1 => n15462, C2 => n4515, A => n4513, B => 
                           n15160, ZN => n4512);
   U11808 : NAND2_X1 port map( A1 => n15462, A2 => n15463, ZN => n4514);
   U11809 : NAND2_X1 port map( A1 => n4517, A2 => n17696, ZN => n4516);
   U11810 : MUX2_X1 port map( A => n17695, B => n18275, S => n18203, Z => n4517
                           );
   U11812 : NAND3_X1 port map( A1 => n14705, A2 => n15265, A3 => n15506, ZN => 
                           n6217);
   U11813 : NAND2_X1 port map( A1 => n29558, A2 => n4520, ZN => n4519);
   U11814 : NOR2_X1 port map( A1 => n28199, A2 => n14426, ZN => n4520);
   U11815 : NAND2_X1 port map( A1 => n4523, A2 => n4522, ZN => n4521);
   U11816 : INV_X1 port map( A => n13874, ZN => n4522);
   U11817 : OAI211_X1 port map( C1 => n4526, C2 => n27224, A => n4525, B => 
                           n4524, ZN => Ciphertext(54));
   U11818 : NAND2_X1 port map( A1 => n27224, A2 => n4527, ZN => n4524);
   U11819 : OAI21_X1 port map( B1 => n27223, B2 => n4528, A => n4527, ZN => 
                           n4525);
   U11821 : INV_X1 port map( A => n27225, ZN => n4527);
   U11822 : AOI21_X1 port map( B1 => n27222, B2 => n27221, A => n27520, ZN => 
                           n4528);
   U11823 : NAND2_X1 port map( A1 => n27525, A2 => n6095, ZN => n27221);
   U11824 : XNOR2_X1 port map( A => n5621, B => n4529, ZN => n4531);
   U11825 : XNOR2_X1 port map( A => n16005, B => n4530, ZN => n4529);
   U11826 : INV_X1 port map( A => n16649, ZN => n4530);
   U11827 : NAND2_X1 port map( A1 => n24094, A2 => n24470, ZN => n24096);
   U11828 : NAND2_X1 port map( A1 => n4536, A2 => n27854, ZN => n4533);
   U11829 : XNOR2_X1 port map( A => n4535, B => n2116, ZN => Ciphertext(143));
   U11830 : NAND2_X1 port map( A1 => n10785, A2 => n10993, ZN => n10691);
   U11831 : NOR2_X1 port map( A1 => n3454, A2 => n10991, ZN => n4539);
   U11832 : XNOR2_X2 port map( A => n9798, B => n9793, ZN => n10993);
   U11833 : NAND2_X1 port map( A1 => n9179, A2 => n6828, ZN => n4540);
   U11834 : NAND2_X1 port map( A1 => n9178, A2 => n9177, ZN => n4541);
   U11835 : XNOR2_X1 port map( A => n10146, B => n9779, ZN => n10080);
   U11836 : NAND3_X1 port map( A1 => n9581, A2 => n9582, A3 => n9580, ZN => 
                           n9779);
   U11839 : OAI21_X1 port map( B1 => n18400, B2 => n18233, A => n17976, ZN => 
                           n4545);
   U11840 : INV_X1 port map( A => n18232, ZN => n4546);
   U11841 : NAND2_X1 port map( A1 => n29074, A2 => n23177, ZN => n23564);
   U11842 : NAND2_X1 port map( A1 => n4549, A2 => n15420, ZN => n4548);
   U11843 : INV_X1 port map( A => n15103, ZN => n4549);
   U11844 : NAND3_X1 port map( A1 => n7823, A2 => n8222, A3 => n1842, ZN => 
                           n4551);
   U11845 : NAND2_X1 port map( A1 => n7821, A2 => n7424, ZN => n4552);
   U11846 : NAND2_X1 port map( A1 => n10101, A2 => n11132, ZN => n4554);
   U11847 : INV_X1 port map( A => n10713, ZN => n10499);
   U11848 : INV_X1 port map( A => n10711, ZN => n4555);
   U11849 : INV_X1 port map( A => n20480, ZN => n20476);
   U11850 : INV_X1 port map( A => n20479, ZN => n4557);
   U11851 : NOR2_X2 port map( A1 => n4558, A2 => n23898, ZN => n25855);
   U11852 : AOI21_X1 port map( B1 => n24368, B2 => n24367, A => n24369, ZN => 
                           n4559);
   U11853 : NAND2_X1 port map( A1 => n379, A2 => n28581, ZN => n4561);
   U11854 : NAND2_X1 port map( A1 => n23268, A2 => n23611, ZN => n4562);
   U11855 : NAND2_X1 port map( A1 => n16541, A2 => n16812, ZN => n17117);
   U11856 : NAND2_X1 port map( A1 => n421, A2 => n4563, ZN => n17460);
   U11857 : AND2_X1 port map( A1 => n29539, A2 => n17459, ZN => n4563);
   U11858 : NOR2_X1 port map( A1 => n421, A2 => n29539, ZN => n16101);
   U11859 : OR2_X1 port map( A1 => n16813, A2 => n29539, ZN => n4564);
   U11860 : NAND2_X1 port map( A1 => n5295, A2 => n27855, ZN => n27848);
   U11861 : NAND2_X1 port map( A1 => n1916, A2 => n20601, ZN => n4567);
   U11862 : NAND2_X1 port map( A1 => n20457, A2 => n4567, ZN => n20460);
   U11863 : NAND2_X1 port map( A1 => n4570, A2 => n4569, ZN => n4568);
   U11864 : MUX2_X1 port map( A => n18305, B => n18306, S => n18476, Z => 
                           n15524);
   U11865 : NAND2_X1 port map( A1 => n24795, A2 => n24796, ZN => n4572);
   U11866 : NAND2_X1 port map( A1 => n4574, A2 => n1955, ZN => n4573);
   U11867 : NAND2_X1 port map( A1 => n4576, A2 => n28455, ZN => n4574);
   U11868 : OR2_X1 port map( A1 => n7993, A2 => n7995, ZN => n4578);
   U11869 : NAND2_X1 port map( A1 => n7650, A2 => n4578, ZN => n4577);
   U11870 : XNOR2_X1 port map( A => n4580, B => n19652, ZN => n4579);
   U11871 : INV_X1 port map( A => n19651, ZN => n4580);
   U11872 : OAI211_X1 port map( C1 => n17192, C2 => n17025, A => n17346, B => 
                           n4582, ZN => n4583);
   U11873 : NAND2_X1 port map( A1 => n17192, A2 => n17344, ZN => n4582);
   U11877 : INV_X1 port map( A => n9074, ZN => n4585);
   U11878 : XNOR2_X1 port map( A => n10005, B => n9658, ZN => n4592);
   U11879 : OAI21_X1 port map( B1 => n23611, B2 => n28582, A => n4593, ZN => 
                           n4598);
   U11880 : NAND2_X1 port map( A1 => n23611, A2 => n29115, ZN => n4593);
   U11881 : NOR2_X1 port map( A1 => n23217, A2 => n406, ZN => n4596);
   U11882 : NOR2_X1 port map( A1 => n23955, A2 => n4596, ZN => n4594);
   U11883 : NAND2_X1 port map( A1 => n4598, A2 => n4599, ZN => n4597);
   U11884 : NAND2_X1 port map( A1 => n4597, A2 => n4595, ZN => n23956);
   U11885 : MUX2_X1 port map( A => n11052, B => n10856, S => n11163, Z => 
                           n11055);
   U11886 : NAND3_X1 port map( A1 => n4604, A2 => n24667, A3 => n24666, ZN => 
                           n4603);
   U11887 : NAND2_X1 port map( A1 => n24668, A2 => n4605, ZN => n4604);
   U11888 : XNOR2_X1 port map( A => n16536, B => n4606, ZN => n15945);
   U11889 : XNOR2_X1 port map( A => n15727, B => n4607, ZN => n4606);
   U11890 : NOR2_X2 port map( A1 => n15254, A2 => n15255, ZN => n15727);
   U11891 : NAND2_X1 port map( A1 => n13692, A2 => n5584, ZN => n4608);
   U11892 : NOR2_X1 port map( A1 => n15138, A2 => n14733, ZN => n4611);
   U11893 : INV_X1 port map( A => n14733, ZN => n15249);
   U11894 : NAND3_X1 port map( A1 => n17001, A2 => n539, A3 => n16844, ZN => 
                           n4612);
   U11895 : NAND2_X1 port map( A1 => n4615, A2 => n4616, ZN => n12868);
   U11896 : INV_X1 port map( A => n12241, ZN => n12035);
   U11897 : INV_X1 port map( A => n14729, ZN => n4621);
   U11898 : NAND2_X1 port map( A1 => n17242, A2 => n16944, ZN => n4625);
   U11899 : NAND2_X1 port map( A1 => n29483, A2 => n17548, ZN => n4626);
   U11901 : NAND2_X1 port map( A1 => n28199, A2 => n13872, ZN => n4627);
   U11903 : NAND2_X1 port map( A1 => n6933, A2 => n21414, ZN => n4631);
   U11904 : OAI21_X1 port map( B1 => n490, B2 => n20663, A => n21410, ZN => 
                           n4633);
   U11905 : NAND2_X1 port map( A1 => n4635, A2 => n4828, ZN => n4634);
   U11906 : OAI21_X1 port map( B1 => n21823, B2 => n20532, A => n4636, ZN => 
                           n4635);
   U11907 : NAND2_X1 port map( A1 => n21823, A2 => n21078, ZN => n4636);
   U11909 : NAND2_X1 port map( A1 => n21819, A2 => n22013, ZN => n4638);
   U11910 : INV_X1 port map( A => n4639, ZN => n6835);
   U11911 : NAND2_X1 port map( A1 => n4642, A2 => n4641, ZN => n14547);
   U11912 : NAND3_X1 port map( A1 => n4515, A2 => n15466, A3 => n29153, ZN => 
                           n4641);
   U11913 : NAND2_X1 port map( A1 => n4515, A2 => n15466, ZN => n5016);
   U11914 : OAI21_X1 port map( B1 => n4645, B2 => n26833, A => n27442, ZN => 
                           n4644);
   U11915 : AND2_X1 port map( A1 => n27438, A2 => n26829, ZN => n4645);
   U11916 : OAI21_X2 port map( B1 => n25363, B2 => n26560, A => n25362, ZN => 
                           n27433);
   U11917 : NAND3_X1 port map( A1 => n21750, A2 => n21237, A3 => n21399, ZN => 
                           n4646);
   U11918 : NAND2_X1 port map( A1 => n11316, A2 => n594, ZN => n4650);
   U11919 : NAND2_X1 port map( A1 => n17151, A2 => n17146, ZN => n4654);
   U11920 : INV_X1 port map( A => n17489, ZN => n4655);
   U11921 : AND2_X1 port map( A1 => n20658, A2 => n4659, ZN => n20659);
   U11922 : OR2_X1 port map( A1 => n19921, A2 => n19920, ZN => n4658);
   U11923 : XNOR2_X1 port map( A => n16494, B => n16039, ZN => n16351);
   U11925 : NAND2_X1 port map( A1 => n6681, A2 => n15094, ZN => n4661);
   U11926 : NAND2_X1 port map( A1 => n4663, A2 => n24378, ZN => n4662);
   U11927 : NOR2_X1 port map( A1 => n24373, A2 => n24374, ZN => n4663);
   U11928 : NAND2_X1 port map( A1 => n24373, A2 => n24380, ZN => n4664);
   U11929 : OAI21_X1 port map( B1 => n14429, B2 => n28199, A => n4665, ZN => 
                           n12533);
   U11930 : XNOR2_X1 port map( A => n18991, B => n19347, ZN => n19353);
   U11931 : INV_X1 port map( A => n13008, ZN => n4670);
   U11932 : INV_X1 port map( A => n13244, ZN => n4669);
   U11933 : XNOR2_X1 port map( A => n4669, B => n12686, ZN => n12688);
   U11934 : XNOR2_X1 port map( A => n4670, B => n12686, ZN => n13010);
   U11935 : AOI21_X1 port map( B1 => n5120, B2 => n7875, A => n7958, ZN => 
                           n4671);
   U11937 : OR2_X1 port map( A1 => n4672, A2 => n23298, ZN => n5940);
   U11938 : INV_X1 port map( A => n8192, ZN => n4676);
   U11939 : NAND2_X1 port map( A1 => n7095, A2 => n7868, ZN => n4673);
   U11940 : NAND2_X1 port map( A1 => n7861, A2 => n7094, ZN => n4674);
   U11941 : NOR3_X1 port map( A1 => n8828, A2 => n4676, A3 => n8586, ZN => 
                           n8587);
   U11942 : NAND3_X1 port map( A1 => n8826, A2 => n8827, A3 => n4676, ZN => 
                           n8832);
   U11943 : NAND2_X1 port map( A1 => n1839, A2 => n4676, ZN => n8196);
   U11944 : OAI21_X1 port map( B1 => n26431, B2 => n26382, A => n26378, ZN => 
                           n4678);
   U11945 : INV_X1 port map( A => n26275, ZN => n4679);
   U11946 : INV_X1 port map( A => n17279, ZN => n5968);
   U11947 : NAND2_X1 port map( A1 => n539, A2 => n17272, ZN => n17279);
   U11948 : OAI21_X1 port map( B1 => n16665, B2 => n5968, A => n4681, ZN => 
                           n4680);
   U11949 : INV_X1 port map( A => n17271, ZN => n4681);
   U11950 : NAND2_X1 port map( A1 => n21253, A2 => n21811, ZN => n21808);
   U11951 : NAND2_X1 port map( A1 => n20117, A2 => n4684, ZN => n4683);
   U11952 : AND2_X1 port map( A1 => n4685, A2 => n24810, ZN => n23692);
   U11953 : INV_X1 port map( A => n24812, ZN => n4685);
   U11954 : AND2_X1 port map( A1 => n17478, A2 => n4687, ZN => n6560);
   U11955 : NAND2_X1 port map( A1 => n17481, A2 => n1816, ZN => n16690);
   U11956 : XNOR2_X1 port map( A => n4688, B => n16579, ZN => n6753);
   U11957 : XNOR2_X1 port map( A => n4688, B => n1193, ZN => n13670);
   U11958 : XNOR2_X1 port map( A => n16574, B => n4688, ZN => n15597);
   U11959 : XNOR2_X1 port map( A => n16318, B => n4688, ZN => n15703);
   U11960 : XNOR2_X1 port map( A => n16012, B => n4688, ZN => n15764);
   U11961 : XNOR2_X1 port map( A => n16255, B => n4688, ZN => n15825);
   U11962 : XNOR2_X1 port map( A => n16455, B => n4688, ZN => n16458);
   U11964 : NAND2_X1 port map( A1 => n4693, A2 => n24279, ZN => n4694);
   U11965 : INV_X1 port map( A => n7966, ZN => n4696);
   U11967 : NAND2_X1 port map( A1 => n16721, A2 => n17455, ZN => n4699);
   U11968 : NAND3_X1 port map( A1 => n4701, A2 => n4706, A3 => n28801, ZN => 
                           n4700);
   U11969 : NAND2_X1 port map( A1 => n4703, A2 => n17450, ZN => n4701);
   U11970 : INV_X1 port map( A => n17065, ZN => n4703);
   U11972 : NAND2_X1 port map( A1 => n17065, A2 => n17452, ZN => n4706);
   U11973 : NAND3_X1 port map( A1 => n390, A2 => n4712, A3 => n11458, ZN => 
                           n4711);
   U11974 : NOR2_X2 port map( A1 => n10509, A2 => n10508, ZN => n11458);
   U11976 : XNOR2_X1 port map( A => n4713, B => n10263, ZN => n9706);
   U11977 : XNOR2_X1 port map( A => n10191, B => n4713, ZN => n7329);
   U11978 : XNOR2_X1 port map( A => n4713, B => n9318, ZN => n9962);
   U11979 : XNOR2_X1 port map( A => n4714, B => n10363, ZN => n10086);
   U11980 : XNOR2_X1 port map( A => n4714, B => n2325, ZN => n9703);
   U11981 : XNOR2_X1 port map( A => n9266, B => n4714, ZN => n9268);
   U11982 : NOR2_X1 port map( A1 => n10964, A2 => n4715, ZN => n10967);
   U11984 : INV_X1 port map( A => n17569, ZN => n4717);
   U11985 : OAI22_X1 port map( A1 => n4719, A2 => n14998, B1 => n14747, B2 => 
                           n15132, ZN => n4718);
   U11986 : NAND2_X1 port map( A1 => n15132, A2 => n551, ZN => n4719);
   U11987 : NAND2_X1 port map( A1 => n14119, A2 => n4721, ZN => n13625);
   U11988 : XNOR2_X2 port map( A => n12947, B => n12946, ZN => n6000);
   U11989 : INV_X1 port map( A => n23642, ZN => n23641);
   U11990 : OAI21_X1 port map( B1 => n21002, B2 => n21220, A => n21001, ZN => 
                           n4723);
   U11991 : NOR2_X2 port map( A1 => n20702, A2 => n18753, ZN => n21220);
   U11992 : NAND2_X1 port map( A1 => n4722, A2 => n4724, ZN => n20702);
   U11993 : NAND2_X1 port map( A1 => n18574, A2 => n19844, ZN => n4722);
   U11994 : AOI21_X2 port map( B1 => n21003, B2 => n21220, A => n4723, ZN => 
                           n22912);
   U11995 : NAND2_X1 port map( A1 => n18573, A2 => n29551, ZN => n4724);
   U11996 : NAND2_X1 port map( A1 => n6379, A2 => n17286, ZN => n18236);
   U11997 : AND2_X1 port map( A1 => n1914, A2 => n23802, ZN => n5192);
   U11998 : NOR2_X1 port map( A1 => n1914, A2 => n23689, ZN => n23540);
   U11999 : AOI21_X1 port map( B1 => n23689, B2 => n23802, A => n1914, ZN => 
                           n23175);
   U12000 : NAND2_X1 port map( A1 => n29598, A2 => n16811, ZN => n17118);
   U12002 : NAND2_X1 port map( A1 => n4729, A2 => n597, ZN => n4728);
   U12003 : INV_X1 port map( A => n9825, ZN => n9603);
   U12004 : NAND2_X1 port map( A1 => n5569, A2 => n5160, ZN => n4731);
   U12006 : NAND2_X1 port map( A1 => n17846, A2 => n17847, ZN => n4732);
   U12007 : NAND2_X1 port map( A1 => n21574, A2 => n21575, ZN => n20848);
   U12009 : NAND2_X1 port map( A1 => n13891, A2 => n14444, ZN => n13685);
   U12010 : NOR2_X1 port map( A1 => n28647, A2 => n14414, ZN => n6232);
   U12011 : NAND2_X1 port map( A1 => n14419, A2 => n28648, ZN => n13687);
   U12013 : XNOR2_X1 port map( A => n8648, B => n8647, ZN => n10334);
   U12014 : NAND2_X1 port map( A1 => n4836, A2 => n13894, ZN => n15463);
   U12015 : NOR2_X2 port map( A1 => n21776, A2 => n4735, ZN => n24596);
   U12016 : NAND2_X1 port map( A1 => n4737, A2 => n4736, ZN => n4735);
   U12017 : NAND3_X1 port map( A1 => n23788, A2 => n23036, A3 => n473, ZN => 
                           n4736);
   U12018 : NAND2_X1 port map( A1 => n21769, A2 => n23482, ZN => n4737);
   U12019 : XNOR2_X1 port map( A => n21994, B => n20885, ZN => n4738);
   U12020 : XNOR2_X1 port map( A => n21761, B => n4738, ZN => n21764);
   U12021 : INV_X1 port map( A => n4738, ZN => n21760);
   U12022 : AND2_X1 port map( A1 => n455, A2 => n27701, ZN => n4741);
   U12024 : AOI21_X1 port map( B1 => n27175, B2 => n26263, A => n28480, ZN => 
                           n26265);
   U12027 : OAI21_X1 port map( B1 => n10717, B2 => n28436, A => n4744, ZN => 
                           n11791);
   U12028 : AOI22_X1 port map( A1 => n11720, A2 => n10717, B1 => n11719, B2 => 
                           n4744, ZN => n11721);
   U12030 : NAND2_X1 port map( A1 => n24596, A2 => n24597, ZN => n4748);
   U12031 : NAND2_X1 port map( A1 => n4752, A2 => n4750, ZN => n26571);
   U12032 : NAND2_X1 port map( A1 => n26566, A2 => n29610, ZN => n4752);
   U12033 : NAND2_X1 port map( A1 => n28775, A2 => n17179, ZN => n17377);
   U12035 : XNOR2_X1 port map( A => n16340, B => n1979, ZN => n4753);
   U12036 : NAND2_X1 port map( A1 => n23968, A2 => n24484, ZN => n24486);
   U12039 : NAND3_X1 port map( A1 => n4757, A2 => n17353, A3 => n28558, ZN => 
                           n4756);
   U12040 : INV_X1 port map( A => n18404, ZN => n4757);
   U12044 : XNOR2_X1 port map( A => n22008, B => n21804, ZN => n4760);
   U12045 : INV_X1 port map( A => n18431, ZN => n4762);
   U12047 : XNOR2_X1 port map( A => n4764, B => n25890, ZN => n25072);
   U12048 : XNOR2_X1 port map( A => n4764, B => n25381, ZN => n25817);
   U12049 : XNOR2_X1 port map( A => n16510, B => n16176, ZN => n4811);
   U12050 : XNOR2_X1 port map( A => n15909, B => n16000, ZN => n4767);
   U12051 : XNOR2_X1 port map( A => n16031, B => n4811, ZN => n4765);
   U12052 : NAND2_X1 port map( A1 => n23011, A2 => n4769, ZN => n4768);
   U12054 : NAND2_X1 port map( A1 => n5774, A2 => n23010, ZN => n23546);
   U12055 : NAND2_X1 port map( A1 => n6227, A2 => n23351, ZN => n4773);
   U12056 : NAND2_X1 port map( A1 => n18710, A2 => n18404, ZN => n4774);
   U12057 : OR2_X1 port map( A1 => n18248, A2 => n18708, ZN => n18710);
   U12058 : NAND2_X1 port map( A1 => n20339, A2 => n20504, ZN => n20226);
   U12059 : INV_X1 port map( A => n4776, ZN => n20909);
   U12061 : XNOR2_X1 port map( A => n16443, B => n16262, ZN => n4777);
   U12062 : XNOR2_X1 port map( A => n4777, B => n15592, ZN => n15593);
   U12063 : INV_X1 port map( A => n4777, ZN => n15720);
   U12064 : NAND2_X1 port map( A1 => n4780, A2 => n4779, ZN => n4778);
   U12065 : NAND2_X1 port map( A1 => n14325, A2 => n14323, ZN => n4779);
   U12066 : INV_X1 port map( A => n24578, ZN => n4784);
   U12067 : NAND3_X1 port map( A1 => n4784, A2 => n29025, A3 => n24581, ZN => 
                           n4783);
   U12068 : NAND2_X1 port map( A1 => n24581, A2 => n29025, ZN => n24055);
   U12069 : NOR2_X1 port map( A1 => n4786, A2 => n4953, ZN => n4785);
   U12070 : NOR2_X2 port map( A1 => n20318, A2 => n20317, ZN => n21306);
   U12071 : OAI21_X1 port map( B1 => n10804, B2 => n4788, A => n6745, ZN => 
                           n4789);
   U12072 : NAND2_X1 port map( A1 => n593, A2 => n5150, ZN => n6745);
   U12073 : NAND2_X1 port map( A1 => n11153, A2 => n11158, ZN => n4788);
   U12074 : NAND2_X1 port map( A1 => n11158, A2 => n11154, ZN => n10803);
   U12075 : XNOR2_X2 port map( A => n6184, B => n6183, ZN => n11158);
   U12077 : INV_X1 port map( A => n6745, ZN => n11159);
   U12078 : AOI21_X1 port map( B1 => n10802, B2 => n10803, A => n11153, ZN => 
                           n4790);
   U12079 : NAND2_X1 port map( A1 => n4791, A2 => n14824, ZN => n14779);
   U12080 : NAND2_X1 port map( A1 => n15433, A2 => n4791, ZN => n15894);
   U12081 : NAND2_X1 port map( A1 => n15027, A2 => n15431, ZN => n4791);
   U12082 : NAND2_X1 port map( A1 => n20242, A2 => n20241, ZN => n4793);
   U12084 : OAI21_X1 port map( B1 => n18441, B2 => n4929, A => n4796, ZN => 
                           n18185);
   U12085 : NAND2_X1 port map( A1 => n4929, A2 => n18178, ZN => n4796);
   U12086 : AND2_X1 port map( A1 => n5973, A2 => n12075, ZN => n4797);
   U12087 : OAI21_X2 port map( B1 => n4797, B2 => n5947, A => n4798, ZN => 
                           n12677);
   U12088 : NAND2_X1 port map( A1 => n12076, A2 => n12575, ZN => n4798);
   U12089 : INV_X1 port map( A => n12578, ZN => n12575);
   U12090 : AND3_X2 port map( A1 => n6438, A2 => n1996, A3 => n6437, ZN => 
                           n27520);
   U12091 : NAND2_X1 port map( A1 => n4801, A2 => n29149, ZN => n4800);
   U12092 : XNOR2_X1 port map( A => n4806, B => n9590, ZN => n9595);
   U12093 : INV_X1 port map( A => n9591, ZN => n4806);
   U12094 : XNOR2_X1 port map( A => n4807, B => n9940, ZN => n9945);
   U12095 : NOR2_X1 port map( A1 => n27502, A2 => n4808, ZN => n27223);
   U12096 : NAND2_X1 port map( A1 => n4809, A2 => n27520, ZN => n4808);
   U12097 : AOI22_X2 port map( A1 => n23931, A2 => n24591, B1 => n23930, B2 => 
                           n23929, ZN => n25249);
   U12098 : XNOR2_X1 port map( A => n4811, B => n14223, ZN => n14224);
   U12099 : INV_X1 port map( A => n16510, ZN => n16642);
   U12100 : OAI21_X1 port map( B1 => n564, B2 => n4812, A => n14367, ZN => 
                           n14371);
   U12102 : NAND2_X1 port map( A1 => n4814, A2 => n20373, ZN => n4813);
   U12103 : NAND2_X1 port map( A1 => n20070, A2 => n20071, ZN => n4814);
   U12104 : NAND2_X1 port map( A1 => n18843, A2 => n18699, ZN => n20071);
   U12106 : NOR2_X2 port map( A1 => n4817, A2 => n4816, ZN => n27447);
   U12107 : NAND2_X1 port map( A1 => n4820, A2 => n26172, ZN => n4819);
   U12108 : XNOR2_X1 port map( A => n4821, B => n26176, ZN => Ciphertext(47));
   U12109 : NAND2_X1 port map( A1 => n26175, A2 => n4822, ZN => n4821);
   U12110 : NAND2_X1 port map( A1 => n26606, A2 => n4823, ZN => n4822);
   U12112 : NAND2_X1 port map( A1 => n7643, A2 => n7981, ZN => n4826);
   U12114 : NAND2_X1 port map( A1 => n4831, A2 => n28801, ZN => n4829);
   U12115 : NAND2_X1 port map( A1 => n17069, A2 => n17068, ZN => n4830);
   U12116 : OAI21_X1 port map( B1 => n4832, B2 => n26450, A => n26179, ZN => 
                           n6124);
   U12117 : AOI21_X1 port map( B1 => n25622, B2 => n29105, A => n4832, ZN => 
                           n24039);
   U12118 : NAND3_X1 port map( A1 => n7982, A2 => n7644, A3 => n7980, ZN => 
                           n4833);
   U12119 : NAND3_X1 port map( A1 => n7642, A2 => n7644, A3 => n7641, ZN => 
                           n4834);
   U12122 : MUX2_X1 port map( A => n4515, B => n29153, S => n15463, Z => n4835)
                           ;
   U12124 : XNOR2_X1 port map( A => n19668, B => n18927, ZN => n4838);
   U12125 : XNOR2_X1 port map( A => n12726, B => n12725, ZN => n14469);
   U12126 : INV_X1 port map( A => n12743, ZN => n4840);
   U12127 : NAND2_X1 port map( A1 => n4842, A2 => n4841, ZN => n12799);
   U12128 : NAND2_X1 port map( A1 => n11702, A2 => n12201, ZN => n4841);
   U12129 : NAND2_X1 port map( A1 => n16889, A2 => n16888, ZN => n4845);
   U12130 : NAND2_X1 port map( A1 => n17088, A2 => n17137, ZN => n4846);
   U12131 : OAI21_X1 port map( B1 => n23546, B2 => n4232, A => n4851, ZN => 
                           n4850);
   U12132 : INV_X1 port map( A => n4850, ZN => n4849);
   U12133 : NAND2_X1 port map( A1 => n15162, A2 => n4515, ZN => n4853);
   U12135 : NAND3_X1 port map( A1 => n7758, A2 => n8176, A3 => n4856, ZN => 
                           n7180);
   U12136 : OR2_X1 port map( A1 => n8175, A2 => n4856, ZN => n7182);
   U12137 : INV_X1 port map( A => n7759, ZN => n4856);
   U12138 : MUX2_X1 port map( A => n24081, B => n24079, S => n24078, Z => n4857
                           );
   U12139 : NAND2_X1 port map( A1 => n4859, A2 => n29470, ZN => n4858);
   U12140 : NAND2_X1 port map( A1 => n5728, A2 => n24388, ZN => n4859);
   U12141 : INV_X1 port map( A => Key(101), ZN => n4861);
   U12142 : XNOR2_X1 port map( A => n21994, B => n4862, ZN => n21384);
   U12143 : OAI21_X1 port map( B1 => n17017, B2 => n17249, A => n17251, ZN => 
                           n4865);
   U12144 : NAND2_X1 port map( A1 => n17016, A2 => n4863, ZN => n4864);
   U12145 : AOI21_X1 port map( B1 => n12272, B2 => n12578, A => n11940, ZN => 
                           n4868);
   U12146 : NAND2_X1 port map( A1 => n4867, A2 => n4870, ZN => n12453);
   U12147 : NAND2_X1 port map( A1 => n12274, A2 => n11940, ZN => n4870);
   U12152 : NAND2_X1 port map( A1 => n20147, A2 => n4875, ZN => n4874);
   U12153 : OAI21_X1 port map( B1 => n29134, B2 => n4877, A => n4876, ZN => 
                           n4875);
   U12154 : NAND2_X1 port map( A1 => n28479, A2 => n21096, ZN => n4878);
   U12156 : XNOR2_X1 port map( A => n4880, B => n19025, ZN => n18581);
   U12157 : XNOR2_X1 port map( A => n19025, B => n4881, ZN => n17850);
   U12158 : XNOR2_X1 port map( A => n19025, B => n4882, ZN => n18640);
   U12159 : INV_X1 port map( A => n1119, ZN => n4882);
   U12160 : NOR2_X1 port map( A1 => n20054, A2 => n6114, ZN => n4885);
   U12161 : INV_X1 port map( A => n20172, ZN => n4886);
   U12162 : NAND2_X1 port map( A1 => n4888, A2 => n4889, ZN => n4887);
   U12165 : NAND2_X1 port map( A1 => n23150, A2 => n23459, ZN => n4891);
   U12166 : MUX2_X1 port map( A => n4364, B => n24629, S => n24533, Z => n23984
                           );
   U12167 : OAI21_X1 port map( B1 => n13826, B2 => n13060, A => n4893, ZN => 
                           n4895);
   U12168 : NAND2_X1 port map( A1 => n6872, A2 => n14127, ZN => n4894);
   U12170 : NAND2_X1 port map( A1 => n17382, A2 => n16878, ZN => n4900);
   U12171 : NAND2_X1 port map( A1 => n17388, A2 => n17389, ZN => n4901);
   U12172 : NAND2_X1 port map( A1 => n5532, A2 => n10847, ZN => n4904);
   U12173 : MUX2_X1 port map( A => n21698, B => n29101, S => n6314, Z => n18549
                           );
   U12174 : MUX2_X1 port map( A => n21243, B => n21244, S => n6314, Z => n21247
                           );
   U12175 : NAND2_X1 port map( A1 => n11090, A2 => n10431, ZN => n4908);
   U12176 : NAND2_X1 port map( A1 => n4908, A2 => n29517, ZN => n4907);
   U12177 : NAND2_X1 port map( A1 => n20345, A2 => n19786, ZN => n4910);
   U12178 : NAND2_X1 port map( A1 => n5853, A2 => n20014, ZN => n4911);
   U12179 : OAI21_X1 port map( B1 => n21560, B2 => n21561, A => n21113, ZN => 
                           n21114);
   U12180 : INV_X1 port map( A => n28578, ZN => n4913);
   U12181 : MUX2_X1 port map( A => n28434, B => n28385, S => n28578, Z => 
                           n25363);
   U12183 : OAI22_X1 port map( A1 => n23447, A2 => n23445, B1 => n23446, B2 => 
                           n292, ZN => n4915);
   U12184 : INV_X1 port map( A => n14797, ZN => n14980);
   U12185 : NAND2_X1 port map( A1 => n4917, A2 => n24552, ZN => n24553);
   U12186 : MUX2_X1 port map( A => n4917, B => n28519, S => n24552, Z => n22868
                           );
   U12187 : OAI22_X1 port map( A1 => n23205, A2 => n4917, B1 => n24551, B2 => 
                           n24173, ZN => n23936);
   U12188 : NAND2_X1 port map( A1 => n23937, A2 => n4917, ZN => n6121);
   U12189 : MUX2_X1 port map( A => n23976, B => n23977, S => n22869, Z => 
                           n23978);
   U12190 : XNOR2_X1 port map( A => n4918, B => n4923, ZN => Ciphertext(21));
   U12191 : NAND2_X1 port map( A1 => n4921, A2 => n4922, ZN => n4919);
   U12193 : NAND3_X1 port map( A1 => n27242, A2 => n27386, A3 => n28177, ZN => 
                           n4924);
   U12194 : AND2_X1 port map( A1 => n29138, A2 => n17229, ZN => n6292);
   U12195 : OR2_X1 port map( A1 => n18442, A2 => n18181, ZN => n4927);
   U12196 : INV_X1 port map( A => n19252, ZN => n19383);
   U12197 : NAND2_X1 port map( A1 => n2039, A2 => n16763, ZN => n4930);
   U12198 : AOI21_X1 port map( B1 => n8998, B2 => n9438, A => n9211, ZN => 
                           n4931);
   U12199 : NAND2_X1 port map( A1 => n8776, A2 => n8996, ZN => n4932);
   U12200 : INV_X1 port map( A => n9434, ZN => n8998);
   U12202 : NAND2_X1 port map( A1 => n5742, A2 => n5741, ZN => n4934);
   U12203 : NAND2_X1 port map( A1 => n23033, A2 => n4936, ZN => n4935);
   U12204 : NOR2_X1 port map( A1 => n23758, A2 => n29131, ZN => n4936);
   U12205 : INV_X1 port map( A => n4937, ZN => n21414);
   U12206 : NOR2_X1 port map( A1 => n28184, A2 => n4937, ZN => n21052);
   U12207 : NAND2_X1 port map( A1 => n21230, A2 => n4937, ZN => n21176);
   U12208 : NAND2_X1 port map( A1 => n7774, A2 => n7889, ZN => n4939);
   U12209 : INV_X1 port map( A => n8048, ZN => n4942);
   U12210 : NAND2_X1 port map( A1 => n8132, A2 => n8131, ZN => n4940);
   U12211 : NAND2_X1 port map( A1 => n4942, A2 => n7554, ZN => n4941);
   U12212 : NAND2_X1 port map( A1 => n26426, A2 => n26378, ZN => n4944);
   U12214 : NAND2_X1 port map( A1 => n17555, A2 => n16913, ZN => n16917);
   U12215 : XNOR2_X1 port map( A => n4946, B => n27550, ZN => Ciphertext(77));
   U12216 : NAND2_X1 port map( A1 => n4948, A2 => n4947, ZN => n4946);
   U12217 : OAI21_X1 port map( B1 => n5540, B2 => n27548, A => n27547, ZN => 
                           n4947);
   U12218 : NOR2_X1 port map( A1 => n27537, A2 => n27202, ZN => n5540);
   U12219 : OAI21_X1 port map( B1 => n27545, B2 => n27546, A => n394, ZN => 
                           n4948);
   U12223 : NAND2_X1 port map( A1 => n22851, A2 => n28182, ZN => n4951);
   U12224 : NOR2_X1 port map( A1 => n17792, A2 => n17793, ZN => n4953);
   U12225 : INV_X1 port map( A => n16332, ZN => n4956);
   U12226 : XNOR2_X1 port map( A => n4956, B => n15545, ZN => n16376);
   U12229 : OR2_X2 port map( A1 => n14089, A2 => n14090, ZN => n15290);
   U12230 : INV_X1 port map( A => n14285, ZN => n14282);
   U12233 : AOI21_X1 port map( B1 => n17502, B2 => n6727, A => n17501, ZN => 
                           n4963);
   U12234 : NAND2_X1 port map( A1 => n24378, A2 => n24380, ZN => n23377);
   U12235 : XNOR2_X1 port map( A => n16596, B => n15989, ZN => n4965);
   U12236 : XNOR2_X1 port map( A => n4965, B => n16193, ZN => n16194);
   U12237 : INV_X1 port map( A => n4965, ZN => n15561);
   U12238 : NAND2_X1 port map( A1 => n24592, A2 => n24591, ZN => n4966);
   U12239 : NAND3_X1 port map( A1 => n24143, A2 => n24144, A3 => n4693, ZN => 
                           n24145);
   U12240 : XNOR2_X1 port map( A => n22008, B => n22238, ZN => n4967);
   U12241 : INV_X1 port map( A => n4971, ZN => n4970);
   U12242 : NOR2_X1 port map( A1 => n11154, A2 => n11158, ZN => n4972);
   U12243 : NOR2_X1 port map( A1 => n14336, A2 => n5584, ZN => n4975);
   U12244 : NOR2_X1 port map( A1 => n1830, A2 => n4974, ZN => n4973);
   U12245 : NAND2_X1 port map( A1 => n4975, A2 => n14408, ZN => n13882);
   U12246 : XNOR2_X1 port map( A => n19305, B => n19306, ZN => n19308);
   U12247 : XNOR2_X1 port map( A => n15727, B => n4978, ZN => n4977);
   U12248 : NAND2_X1 port map( A1 => n16430, A2 => n4979, ZN => n17185);
   U12249 : NAND2_X1 port map( A1 => n2483, A2 => n12127, ZN => n4981);
   U12250 : NAND2_X1 port map( A1 => n8670, A2 => n9107, ZN => n8672);
   U12251 : NAND3_X1 port map( A1 => n8670, A2 => n8914, A3 => n9107, ZN => 
                           n8514);
   U12252 : NAND2_X1 port map( A1 => n9106, A2 => n8670, ZN => n9121);
   U12253 : OAI21_X2 port map( B1 => n28186, B2 => n4984, A => n19329, ZN => 
                           n21714);
   U12254 : OAI21_X1 port map( B1 => n20334, B2 => n20626, A => n4985, ZN => 
                           n4984);
   U12255 : NAND2_X1 port map( A1 => n20623, A2 => n20626, ZN => n4985);
   U12256 : NAND2_X1 port map( A1 => n4986, A2 => n18398, ZN => n5757);
   U12257 : NAND2_X1 port map( A1 => n18233, A2 => n18231, ZN => n4986);
   U12259 : NAND2_X1 port map( A1 => n5460, A2 => n17434, ZN => n4987);
   U12261 : NAND2_X1 port map( A1 => n6605, A2 => n20498, ZN => n4991);
   U12262 : AND2_X2 port map( A1 => n20010, A2 => n20011, ZN => n21638);
   U12263 : MUX2_X1 port map( A => n4992, B => n15243, S => n15359, Z => n14508
                           );
   U12264 : AOI22_X1 port map( A1 => n15061, A2 => n4992, B1 => n15359, B2 => 
                           n15062, ZN => n15063);
   U12265 : OAI21_X1 port map( B1 => n15358, B2 => n28197, A => n4992, ZN => 
                           n6003);
   U12266 : MUX2_X1 port map( A => n24240, B => n24559, S => n24633, Z => n4993
                           );
   U12267 : NAND2_X1 port map( A1 => n23558, A2 => n23188, ZN => n4994);
   U12268 : NAND2_X1 port map( A1 => n23989, A2 => n24557, ZN => n4995);
   U12269 : NAND2_X1 port map( A1 => n5966, A2 => n11435, ZN => n4996);
   U12270 : INV_X1 port map( A => n27938, ZN => n4998);
   U12271 : OAI211_X1 port map( C1 => n27942, C2 => n27941, A => n27940, B => 
                           n4999, ZN => n27943);
   U12272 : NAND2_X1 port map( A1 => n5000, A2 => n20899, ZN => n20141);
   U12273 : NOR2_X1 port map( A1 => n1925, A2 => n5000, ZN => n20143);
   U12274 : NOR2_X1 port map( A1 => n17254, A2 => n1880, ZN => n17256);
   U12275 : INV_X1 port map( A => n17249, ZN => n5001);
   U12276 : XNOR2_X1 port map( A => n13474, B => n12473, ZN => n5002);
   U12277 : XNOR2_X1 port map( A => n12474, B => n12471, ZN => n5003);
   U12278 : NAND3_X1 port map( A1 => n28441, A2 => n28438, A3 => n27944, ZN => 
                           n27940);
   U12279 : NAND3_X1 port map( A1 => n4998, A2 => n28439, A3 => n27941, ZN => 
                           n27928);
   U12280 : MUX2_X1 port map( A => n28438, B => n27941, S => n27925, Z => 
                           n27245);
   U12281 : MUX2_X1 port map( A => n27244, B => n27925, S => n28439, Z => 
                           n27023);
   U12282 : NAND2_X1 port map( A1 => n27932, A2 => n2060, ZN => n27933);
   U12283 : XNOR2_X1 port map( A => n19693, B => n19694, ZN => n5005);
   U12284 : AND3_X1 port map( A1 => n12234, A2 => n12236, A3 => n12233, ZN => 
                           n5007);
   U12285 : NAND2_X1 port map( A1 => n12234, A2 => n12233, ZN => n12235);
   U12286 : AOI21_X1 port map( B1 => n5009, B2 => n5008, A => n5007, ZN => 
                           n5012);
   U12287 : INV_X1 port map( A => n1986, ZN => n5009);
   U12288 : NAND2_X1 port map( A1 => n5012, A2 => n5010, ZN => n12472);
   U12289 : NAND2_X1 port map( A1 => n5011, A2 => n1986, ZN => n5010);
   U12290 : OAI21_X1 port map( B1 => n776, B2 => n12232, A => n12234, ZN => 
                           n5011);
   U12291 : NAND2_X1 port map( A1 => n20900, A2 => n21084, ZN => n5013);
   U12292 : INV_X1 port map( A => n15463, ZN => n15161);
   U12293 : INV_X1 port map( A => n15464, ZN => n14652);
   U12294 : INV_X1 port map( A => n28024, ZN => n28034);
   U12295 : NOR2_X1 port map( A1 => n28026, A2 => n5017, ZN => n28031);
   U12297 : INV_X1 port map( A => n20865, ZN => n21185);
   U12298 : INV_X1 port map( A => n22132, ZN => n22723);
   U12299 : OR2_X1 port map( A1 => n20187, A2 => n20186, ZN => n5018);
   U12300 : AOI22_X2 port map( A1 => n5020, A2 => n10701, B1 => n5019, B2 => 
                           n11768, ZN => n13014);
   U12301 : INV_X1 port map( A => n18708, ZN => n5021);
   U12302 : NAND2_X1 port map( A1 => n5025, A2 => n15404, ZN => n5024);
   U12304 : NAND2_X1 port map( A1 => n28195, A2 => n15402, ZN => n15398);
   U12306 : INV_X1 port map( A => n23067, ZN => n23693);
   U12307 : NAND2_X1 port map( A1 => n23693, A2 => n23531, ZN => n5028);
   U12308 : INV_X1 port map( A => n23531, ZN => n5030);
   U12310 : INV_X1 port map( A => n23531, ZN => n23696);
   U12311 : XNOR2_X1 port map( A => n10421, B => n2035, ZN => n9617);
   U12312 : XNOR2_X1 port map( A => n10421, B => n5032, ZN => n9386);
   U12313 : NAND2_X1 port map( A1 => n20156, A2 => n20155, ZN => n5033);
   U12314 : AOI21_X1 port map( B1 => n1121, B2 => n17347, A => n542, ZN => 
                           n16951);
   U12315 : NAND2_X1 port map( A1 => n29100, A2 => n26748, ZN => n5036);
   U12316 : NAND3_X1 port map( A1 => n12134, A2 => n12265, A3 => n12133, ZN => 
                           n5038);
   U12317 : MUX2_X1 port map( A => n12267, B => n12132, S => n11574, Z => n5040
                           );
   U12320 : NAND2_X1 port map( A1 => n5042, A2 => n23405, ZN => n5041);
   U12321 : XNOR2_X1 port map( A => n5043, B => n22584, ZN => n22032);
   U12322 : NAND3_X1 port map( A1 => n5046, A2 => n22029, A3 => n5044, ZN => 
                           n5043);
   U12323 : NAND2_X1 port map( A1 => n5045, A2 => n28108, ZN => n5044);
   U12324 : INV_X1 port map( A => n22030, ZN => n5045);
   U12325 : NAND4_X1 port map( A1 => n22294, A2 => n1927, A3 => n22030, A4 => 
                           n5047, ZN => n5046);
   U12326 : INV_X1 port map( A => n22028, ZN => n5047);
   U12328 : NAND3_X1 port map( A1 => n15512, A2 => n15514, A3 => n15515, ZN => 
                           n5051);
   U12329 : INV_X1 port map( A => n15275, ZN => n5049);
   U12330 : NAND2_X1 port map( A1 => n15274, A2 => n15275, ZN => n14920);
   U12331 : NAND2_X1 port map( A1 => n5048, A2 => n15274, ZN => n5050);
   U12332 : NOR2_X1 port map( A1 => n5049, A2 => n15514, ZN => n5048);
   U12333 : NAND2_X1 port map( A1 => n15279, A2 => n15512, ZN => n5052);
   U12334 : OAI21_X1 port map( B1 => n20152, B2 => n5053, A => n20098, ZN => 
                           n5054);
   U12335 : INV_X1 port map( A => n20150, ZN => n5053);
   U12336 : NAND2_X1 port map( A1 => n20042, A2 => n20096, ZN => n5055);
   U12337 : INV_X1 port map( A => n20098, ZN => n5056);
   U12338 : AOI21_X1 port map( B1 => n14375, B2 => n14374, A => n5057, ZN => 
                           n14378);
   U12339 : INV_X1 port map( A => n13725, ZN => n5058);
   U12340 : NAND2_X1 port map( A1 => n16852, A2 => n16853, ZN => n16854);
   U12341 : INV_X1 port map( A => n18761, ZN => n18949);
   U12342 : OAI211_X1 port map( C1 => n16868, C2 => n5059, A => n5061, B => 
                           n5060, ZN => n5062);
   U12343 : NAND3_X1 port map( A1 => n16868, A2 => n16867, A3 => n5059, ZN => 
                           n5061);
   U12344 : XNOR2_X1 port map( A => n29136, B => n5067, ZN => n5066);
   U12345 : XNOR2_X1 port map( A => n22000, B => n22896, ZN => n5067);
   U12346 : NAND2_X1 port map( A1 => n5068, A2 => n16968, ZN => n16792);
   U12347 : XNOR2_X2 port map( A => n15111, B => n15112, ZN => n17304);
   U12348 : XNOR2_X1 port map( A => n5069, B => n13055, ZN => n12833);
   U12350 : XNOR2_X1 port map( A => n12593, B => n5070, ZN => n13569);
   U12351 : INV_X1 port map( A => n13566, ZN => n5070);
   U12352 : NAND2_X1 port map( A1 => n7515, A2 => n29321, ZN => n7261);
   U12353 : OAI22_X1 port map( A1 => n29201, A2 => n1959, B1 => n3269, B2 => 
                           n14394, ZN => n5073);
   U12354 : NAND2_X1 port map( A1 => n1952, A2 => n29104, ZN => n5074);
   U12355 : NAND3_X1 port map( A1 => n28820, A2 => n20091, A3 => n20039, ZN => 
                           n5075);
   U12356 : NAND2_X1 port map( A1 => n5078, A2 => n5077, ZN => n5076);
   U12357 : NAND3_X1 port map( A1 => n11515, A2 => n11671, A3 => n29139, ZN => 
                           n5077);
   U12358 : NAND2_X1 port map( A1 => n11632, A2 => n11634, ZN => n11515);
   U12359 : NAND2_X1 port map( A1 => n11406, A2 => n5079, ZN => n5078);
   U12360 : NAND3_X1 port map( A1 => n5080, A2 => n24093, A3 => n24091, ZN => 
                           n24097);
   U12361 : NAND2_X1 port map( A1 => n17798, A2 => n18106, ZN => n18457);
   U12362 : MUX2_X1 port map( A => n23862, B => n26572, S => n25418, Z => 
                           n26573);
   U12364 : NAND2_X1 port map( A1 => n518, A2 => n18354, ZN => n5083);
   U12365 : INV_X1 port map( A => n18353, ZN => n6225);
   U12367 : NAND3_X1 port map( A1 => n21180, A2 => n21551, A3 => n20351, ZN => 
                           n5086);
   U12368 : NAND3_X1 port map( A1 => n5088, A2 => n5087, A3 => n5086, ZN => 
                           n22792);
   U12369 : NAND2_X1 port map( A1 => n2067, A2 => n21553, ZN => n5088);
   U12370 : OR2_X1 port map( A1 => n10116, A2 => n11127, ZN => n5089);
   U12371 : NAND2_X1 port map( A1 => n6833, A2 => n5090, ZN => n6832);
   U12372 : NAND2_X1 port map( A1 => n15374, A2 => n15376, ZN => n5092);
   U12373 : INV_X1 port map( A => n18034, ZN => n18158);
   U12375 : MUX2_X1 port map( A => n11970, B => n5097, S => n12159, Z => n5095)
                           ;
   U12376 : NAND2_X1 port map( A1 => n5098, A2 => n4617, ZN => n5096);
   U12377 : NAND2_X1 port map( A1 => n12244, A2 => n12158, ZN => n5097);
   U12378 : MUX2_X1 port map( A => n12156, B => n12241, S => n12244, Z => n5098
                           );
   U12379 : NAND3_X1 port map( A1 => n97, A2 => n28637, A3 => n20383, ZN => 
                           n5099);
   U12380 : NAND2_X1 port map( A1 => n5103, A2 => n5102, ZN => n5101);
   U12381 : NAND2_X1 port map( A1 => n24631, A2 => n23144, ZN => n5102);
   U12382 : INV_X1 port map( A => n24531, ZN => n5103);
   U12383 : NOR2_X1 port map( A1 => n24530, A2 => n24533, ZN => n5105);
   U12384 : XNOR2_X1 port map( A => n18321, B => n18320, ZN => n20539);
   U12385 : INV_X1 port map( A => n20539, ZN => n20389);
   U12386 : INV_X1 port map( A => n19959, ZN => n20188);
   U12387 : NAND2_X1 port map( A1 => n20223, A2 => n5106, ZN => n19861);
   U12388 : INV_X1 port map( A => n17989, ZN => n18367);
   U12391 : NAND2_X1 port map( A1 => n27077, A2 => n5113, ZN => n5112);
   U12392 : NOR2_X1 port map( A1 => n26991, A2 => n5263, ZN => n5113);
   U12393 : INV_X1 port map( A => n26994, ZN => n5114);
   U12395 : NOR2_X1 port map( A1 => n24277, A2 => n24591, ZN => n5116);
   U12396 : NAND2_X1 port map( A1 => n24593, A2 => n5116, ZN => n5115);
   U12398 : INV_X1 port map( A => n12929, ZN => n5121);
   U12399 : XNOR2_X1 port map( A => n12882, B => n5121, ZN => n5122);
   U12400 : OAI21_X1 port map( B1 => n1876, B2 => n14440, A => n14433, ZN => 
                           n14436);
   U12401 : NAND2_X1 port map( A1 => n21823, A2 => n22013, ZN => n5123);
   U12402 : NAND2_X1 port map( A1 => n4828, A2 => n5125, ZN => n5124);
   U12403 : NAND2_X1 port map( A1 => n6495, A2 => n29551, ZN => n5126);
   U12404 : MUX2_X1 port map( A => n5053, B => n20151, S => n20152, Z => n19775
                           );
   U12405 : MUX2_X1 port map( A => n20152, B => n20151, S => n20150, Z => 
                           n18888);
   U12406 : AOI21_X1 port map( B1 => n20096, B2 => n20155, A => n5053, ZN => 
                           n18833);
   U12407 : XNOR2_X1 port map( A => n17597, B => n5127, ZN => n17606);
   U12408 : INV_X1 port map( A => n18556, ZN => n5127);
   U12409 : XNOR2_X1 port map( A => n18725, B => n19139, ZN => n18556);
   U12410 : NAND3_X1 port map( A1 => n21143, A2 => n21119, A3 => n21140, ZN => 
                           n5128);
   U12411 : INV_X1 port map( A => n7569, ZN => n5129);
   U12412 : NAND2_X1 port map( A1 => n5131, A2 => n603, ZN => n5130);
   U12413 : OAI21_X1 port map( B1 => n9425, B2 => n7569, A => n5132, ZN => 
                           n5131);
   U12414 : NAND3_X1 port map( A1 => n11902, A2 => n12428, A3 => n5134, ZN => 
                           n11905);
   U12415 : XNOR2_X1 port map( A => n25876, B => n25165, ZN => n25517);
   U12416 : XNOR2_X1 port map( A => n25517, B => n25056, ZN => n24624);
   U12420 : NAND2_X1 port map( A1 => n5142, A2 => n21481, ZN => n5140);
   U12421 : NAND3_X1 port map( A1 => n21575, A2 => n20749, A3 => n21580, ZN => 
                           n5141);
   U12422 : INV_X1 port map( A => n20749, ZN => n21576);
   U12423 : INV_X1 port map( A => n21483, ZN => n21484);
   U12424 : MUX2_X1 port map( A => n10696, B => n10984, S => n10989, Z => 
                           n10584);
   U12425 : NAND2_X1 port map( A1 => n23629, A2 => n23308, ZN => n5143);
   U12428 : XNOR2_X1 port map( A => n5146, B => n28327, ZN => n24703);
   U12430 : NAND2_X1 port map( A1 => n11152, A2 => n5150, ZN => n10554);
   U12431 : AOI22_X1 port map( A1 => n593, A2 => n11153, B1 => n11154, B2 => 
                           n5150, ZN => n10093);
   U12432 : NAND2_X1 port map( A1 => n22401, A2 => n5151, ZN => n21018);
   U12433 : NOR2_X1 port map( A1 => n22401, A2 => n5151, ZN => n21067);
   U12434 : NAND3_X1 port map( A1 => n21665, A2 => n21429, A3 => n5151, ZN => 
                           n21017);
   U12438 : NAND2_X1 port map( A1 => n28802, A2 => n15334, ZN => n14781);
   U12440 : MUX2_X1 port map( A => n15047, B => n15233, S => n28802, Z => 
                           n15051);
   U12442 : NAND2_X1 port map( A1 => n18213, A2 => n18216, ZN => n5155);
   U12443 : NAND2_X1 port map( A1 => n5157, A2 => n28763, ZN => n18219);
   U12445 : INV_X1 port map( A => n9045, ZN => n9235);
   U12446 : OAI21_X1 port map( B1 => n6590, B2 => n5159, A => n5158, ZN => 
                           n9240);
   U12447 : INV_X1 port map( A => n9230, ZN => n5160);
   U12448 : XNOR2_X1 port map( A => n19315, B => n19314, ZN => n19319);
   U12450 : AND3_X2 port map( A1 => n17886, A2 => n17885, A3 => n17884, ZN => 
                           n19718);
   U12451 : INV_X1 port map( A => n19718, ZN => n18937);
   U12452 : NAND2_X1 port map( A1 => n17887, A2 => n18334, ZN => n5163);
   U12453 : INV_X1 port map( A => n13661, ZN => n14044);
   U12454 : XNOR2_X1 port map( A => n5166, B => n5165, ZN => n13661);
   U12455 : INV_X1 port map( A => n23924, ZN => n6321);
   U12456 : NAND2_X1 port map( A1 => n5167, A2 => n6746, ZN => n23924);
   U12457 : NAND2_X1 port map( A1 => n5168, A2 => n24612, ZN => n5167);
   U12458 : NAND2_X1 port map( A1 => n11159, A2 => n11158, ZN => n11783);
   U12459 : NAND2_X1 port map( A1 => n11156, A2 => n11155, ZN => n5171);
   U12460 : NAND2_X1 port map( A1 => n11157, A2 => n11154, ZN => n5172);
   U12461 : INV_X1 port map( A => n23651, ZN => n23318);
   U12462 : INV_X1 port map( A => n23261, ZN => n23584);
   U12464 : OR2_X2 port map( A1 => n5174, A2 => n5173, ZN => n9530);
   U12466 : XNOR2_X1 port map( A => n13405, B => n13461, ZN => n5177);
   U12467 : XNOR2_X1 port map( A => n13501, B => n5177, ZN => n12963);
   U12468 : INV_X1 port map( A => n5177, ZN => n13131);
   U12469 : NAND2_X1 port map( A1 => n5180, A2 => n29611, ZN => n5344);
   U12470 : NAND2_X1 port map( A1 => n5180, A2 => n14304, ZN => n5343);
   U12472 : OAI21_X1 port map( B1 => n20145, B2 => n20148, A => n5182, ZN => 
                           n5181);
   U12473 : OR2_X1 port map( A1 => n21095, A2 => n21092, ZN => n5182);
   U12475 : XNOR2_X1 port map( A => n22555, B => n22714, ZN => n5184);
   U12476 : XNOR2_X1 port map( A => n10135, B => n10055, ZN => n5185);
   U12478 : INV_X1 port map( A => n11869, ZN => n11868);
   U12480 : INV_X1 port map( A => n27771, ZN => n5188);
   U12481 : NAND2_X1 port map( A1 => n15309, A2 => n15310, ZN => n5190);
   U12486 : NOR2_X1 port map( A1 => n11501, A2 => n11874, ZN => n6305);
   U12487 : XNOR2_X2 port map( A => n8746, B => n8745, ZN => n11176);
   U12489 : OAI21_X1 port map( B1 => n23151, B2 => n5237, A => n23767, ZN => 
                           n5236);
   U12490 : XNOR2_X2 port map( A => n9776, B => n9775, ZN => n11235);
   U12491 : OR2_X1 port map( A1 => n16922, A2 => n5429, ZN => n5365);
   U12492 : XNOR2_X1 port map( A => n5996, B => n9843, ZN => n8884);
   U12493 : XNOR2_X2 port map( A => n13003, B => n13004, ZN => n14278);
   U12494 : INV_X1 port map( A => n6886, ZN => n19510);
   U12495 : OAI211_X2 port map( C1 => n28666, C2 => n15084, A => n14672, B => 
                           n14671, ZN => n16641);
   U12496 : XNOR2_X1 port map( A => n19597, B => n6193, ZN => n19344);
   U12497 : INV_X1 port map( A => n15056, ZN => n6207);
   U12498 : XNOR2_X1 port map( A => n16397, B => n13926, ZN => n6707);
   U12499 : AOI21_X2 port map( B1 => n14547, B2 => n14546, A => n14545, ZN => 
                           n16603);
   U12500 : INV_X1 port map( A => n27352, ZN => n5421);
   U12502 : OAI21_X2 port map( B1 => n11828, B2 => n11827, A => n11826, ZN => 
                           n13360);
   U12503 : OAI21_X1 port map( B1 => n27771, B2 => n6419, A => n6418, ZN => 
                           n6498);
   U12507 : NOR2_X2 port map( A1 => n14718, A2 => n14717, ZN => n16422);
   U12508 : OAI21_X1 port map( B1 => n6706, B2 => n11622, A => n6705, ZN => 
                           n11570);
   U12509 : OAI21_X1 port map( B1 => n17451, B2 => n28801, A => n17128, ZN => 
                           n17069);
   U12511 : INV_X1 port map( A => n29044, ZN => n18187);
   U12516 : OAI21_X1 port map( B1 => n23282, B2 => n1893, A => n23283, ZN => 
                           n5619);
   U12521 : XNOR2_X1 port map( A => n25557, B => n25933, ZN => n25559);
   U12522 : NAND2_X1 port map( A1 => n5191, A2 => n5149, ZN => n7602);
   U12523 : NAND3_X1 port map( A1 => n7863, A2 => n7092, A3 => n6162, ZN => 
                           n5362);
   U12526 : INV_X1 port map( A => n10079, ZN => n5195);
   U12528 : NAND2_X1 port map( A1 => n15150, A2 => n15151, ZN => n5199);
   U12529 : OAI22_X1 port map( A1 => n21333, A2 => n21332, B1 => n21613, B2 => 
                           n21612, ZN => n21336);
   U12530 : INV_X1 port map( A => n21329, ZN => n20497);
   U12531 : INV_X1 port map( A => n20492, ZN => n21331);
   U12532 : NAND3_X1 port map( A1 => n10739, A2 => n10738, A3 => n5204, ZN => 
                           n12919);
   U12533 : NAND2_X1 port map( A1 => n11489, A2 => n11431, ZN => n5204);
   U12534 : NAND2_X1 port map( A1 => n14240, A2 => n29097, ZN => n13739);
   U12535 : NOR2_X1 port map( A1 => n14240, A2 => n29097, ZN => n14173);
   U12536 : OR2_X1 port map( A1 => n14240, A2 => n15194, ZN => n5207);
   U12537 : NAND2_X1 port map( A1 => n19791, A2 => n20481, ZN => n5208);
   U12538 : NAND2_X1 port map( A1 => n18173, A2 => n18172, ZN => n5209);
   U12539 : NAND2_X1 port map( A1 => n24064, A2 => n23897, ZN => n5210);
   U12540 : AOI21_X1 port map( B1 => n28047, B2 => n28069, A => n5212, ZN => 
                           n5214);
   U12541 : AOI21_X1 port map( B1 => n5213, B2 => n28065, A => n28069, ZN => 
                           n5212);
   U12542 : INV_X1 port map( A => n28065, ZN => n28071);
   U12543 : NAND2_X1 port map( A1 => n28052, A2 => n28067, ZN => n5215);
   U12544 : NAND2_X1 port map( A1 => n5218, A2 => n5216, ZN => n5289);
   U12545 : NAND2_X1 port map( A1 => n5137, A2 => n5217, ZN => n5216);
   U12547 : NAND2_X1 port map( A1 => n22593, A2 => n23829, ZN => n5219);
   U12549 : INV_X1 port map( A => n26246, ZN => n5221);
   U12550 : AND2_X1 port map( A1 => n18172, A2 => n18174, ZN => n5222);
   U12552 : XNOR2_X1 port map( A => n19590, B => n19628, ZN => n5224);
   U12553 : NAND2_X1 port map( A1 => n20495, A2 => n5225, ZN => n20491);
   U12554 : NAND2_X1 port map( A1 => n29616, A2 => n5225, ZN => n20180);
   U12555 : NOR2_X1 port map( A1 => n29616, A2 => n5225, ZN => n19179);
   U12556 : NOR2_X1 port map( A1 => n19863, A2 => n5225, ZN => n19865);
   U12557 : NAND2_X1 port map( A1 => n6834, A2 => n5225, ZN => n20183);
   U12559 : NAND2_X1 port map( A1 => n5229, A2 => n14874, ZN => n13128);
   U12560 : OAI21_X1 port map( B1 => n12053, B2 => n12320, A => n5230, ZN => 
                           n6679);
   U12561 : NAND2_X1 port map( A1 => n12320, A2 => n12051, ZN => n5230);
   U12563 : INV_X1 port map( A => n18393, ZN => n17767);
   U12564 : NAND2_X1 port map( A1 => n5234, A2 => n17766, ZN => n5231);
   U12565 : OR2_X1 port map( A1 => n17769, A2 => n18388, ZN => n5235);
   U12566 : NAND2_X1 port map( A1 => n15046, A2 => n15225, ZN => n15353);
   U12567 : INV_X1 port map( A => n7116, ZN => n7340);
   U12569 : NAND2_X1 port map( A1 => n7118, A2 => n5240, ZN => n5239);
   U12570 : NAND2_X1 port map( A1 => n5241, A2 => n7767, ZN => n5240);
   U12571 : NAND2_X1 port map( A1 => n7116, A2 => n5242, ZN => n5241);
   U12572 : NAND2_X1 port map( A1 => n5244, A2 => n7164, ZN => n5243);
   U12573 : XNOR2_X1 port map( A => n5245, B => n18799, ZN => n19290);
   U12575 : NAND2_X1 port map( A1 => n28506, A2 => n23800, ZN => n23538);
   U12576 : OAI21_X1 port map( B1 => n23172, B2 => n23540, A => n28506, ZN => 
                           n23173);
   U12577 : NAND2_X1 port map( A1 => n20417, A2 => n20578, ZN => n6508);
   U12578 : AND2_X1 port map( A1 => n5248, A2 => n24768, ZN => n23548);
   U12579 : INV_X1 port map( A => n24697, ZN => n5248);
   U12581 : NAND2_X1 port map( A1 => n6830, A2 => n5251, ZN => n5250);
   U12582 : NAND2_X1 port map( A1 => n11812, A2 => n12231, ZN => n5488);
   U12583 : OAI22_X1 port map( A1 => n21590, A2 => n21591, B1 => n5684, B2 => 
                           n21589, ZN => n21592);
   U12586 : NAND3_X1 port map( A1 => n386, A2 => n20275, A3 => n20597, ZN => 
                           n5253);
   U12587 : XNOR2_X2 port map( A => n7047, B => Key(161), ZN => n7967);
   U12588 : NAND2_X1 port map( A1 => n7967, A2 => n29300, ZN => n7962);
   U12589 : OAI21_X2 port map( B1 => n10578, B2 => n5258, A => n5257, ZN => 
                           n12428);
   U12590 : NAND3_X1 port map( A1 => n11092, A2 => n10577, A3 => n5258, ZN => 
                           n5257);
   U12591 : OAI21_X1 port map( B1 => n17192, B2 => n17347, A => n5259, ZN => 
                           n5260);
   U12592 : NAND2_X1 port map( A1 => n17192, A2 => n17346, ZN => n5259);
   U12593 : NAND2_X1 port map( A1 => n14146, A2 => n13725, ZN => n5261);
   U12594 : OAI21_X1 port map( B1 => n29059, B2 => n13725, A => n5261, ZN => 
                           n13593);
   U12595 : NOR2_X1 port map( A1 => n28521, A2 => n5263, ZN => n27075);
   U12596 : NAND2_X1 port map( A1 => n28521, A2 => n5263, ZN => n26862);
   U12597 : INV_X1 port map( A => n10973, ZN => n5265);
   U12598 : INV_X1 port map( A => n10972, ZN => n10681);
   U12600 : NOR2_X1 port map( A1 => n5267, A2 => n10970, ZN => n5266);
   U12601 : XNOR2_X2 port map( A => n5268, B => n9297, ZN => n10970);
   U12602 : INV_X1 port map( A => n337, ZN => n17309);
   U12603 : NAND2_X1 port map( A1 => n15307, A2 => n15311, ZN => n15272);
   U12606 : NAND2_X1 port map( A1 => n1921, A2 => n29569, ZN => n20888);
   U12607 : OAI21_X1 port map( B1 => n5728, B2 => n24079, A => n5272, ZN => 
                           n5307);
   U12608 : OAI22_X1 port map( A1 => n20230, A2 => n4557, B1 => n20353, B2 => 
                           n20475, ZN => n21437);
   U12609 : XNOR2_X1 port map( A => n5275, B => n25869, ZN => n25215);
   U12610 : XNOR2_X1 port map( A => n25868, B => n5275, ZN => n25145);
   U12611 : XNOR2_X1 port map( A => n5275, B => n25922, ZN => n25923);
   U12612 : XNOR2_X1 port map( A => n5275, B => n2523, ZN => n24137);
   U12613 : XNOR2_X1 port map( A => n26095, B => n5275, ZN => n25475);
   U12614 : NAND3_X1 port map( A1 => n7340, A2 => n7770, A3 => n7320, ZN => 
                           n5282);
   U12615 : NAND2_X1 port map( A1 => n2017, A2 => n5956, ZN => n5284);
   U12616 : MUX2_X1 port map( A => n14300, B => n28478, S => n14299, Z => n5285
                           );
   U12617 : INV_X1 port map( A => n15069, ZN => n5287);
   U12619 : NAND3_X1 port map( A1 => n16962, A2 => n17309, A3 => n17440, ZN => 
                           n5288);
   U12621 : NAND2_X1 port map( A1 => n23078, A2 => n28460, ZN => n23283);
   U12622 : NAND2_X1 port map( A1 => n23839, A2 => n23390, ZN => n5291);
   U12623 : OR2_X1 port map( A1 => n29536, A2 => n29497, ZN => n5297);
   U12624 : NAND2_X1 port map( A1 => n5295, A2 => n5294, ZN => n27856);
   U12626 : NAND2_X1 port map( A1 => n27902, A2 => n29575, ZN => n5301);
   U12627 : NAND2_X1 port map( A1 => n5304, A2 => n5303, ZN => n5302);
   U12628 : MUX2_X1 port map( A => n20182, B => n20493, S => n20495, Z => n5304
                           );
   U12629 : INV_X1 port map( A => n17313, ZN => n17317);
   U12630 : NAND2_X1 port map( A1 => n13060, A2 => n14354, ZN => n14356);
   U12631 : NAND2_X1 port map( A1 => n13060, A2 => n13824, ZN => n14349);
   U12632 : NAND3_X1 port map( A1 => n4088, A2 => n13060, A3 => n14351, ZN => 
                           n14128);
   U12633 : NAND2_X1 port map( A1 => n13825, A2 => n13060, ZN => n13627);
   U12635 : INV_X2 port map( A => n5306, ZN => n27076);
   U12636 : NAND2_X1 port map( A1 => n26178, A2 => n26177, ZN => n6125);
   U12637 : OAI22_X1 port map( A1 => n6947, A2 => n26447, B1 => n26452, B2 => 
                           n26179, ZN => n26178);
   U12638 : AOI21_X1 port map( B1 => n6828, B2 => n8643, A => n9396, ZN => 
                           n5308);
   U12639 : NAND2_X1 port map( A1 => n436, A2 => n8981, ZN => n6828);
   U12640 : NAND2_X1 port map( A1 => n409, A2 => n23405, ZN => n5310);
   U12643 : NAND2_X1 port map( A1 => n27209, A2 => n446, ZN => n5312);
   U12644 : NAND2_X1 port map( A1 => n5313, A2 => n295, ZN => n27212);
   U12645 : INV_X1 port map( A => n27208, ZN => n5313);
   U12646 : OAI21_X1 port map( B1 => n12049, B2 => n12050, A => n5315, ZN => 
                           n11770);
   U12647 : NAND2_X1 port map( A1 => n12049, A2 => n12320, ZN => n5315);
   U12648 : NAND2_X1 port map( A1 => n10490, A2 => n29627, ZN => n10098);
   U12649 : NAND2_X1 port map( A1 => n10549, A2 => n29627, ZN => n10548);
   U12650 : AOI21_X1 port map( B1 => n11114, B2 => n11115, A => n29627, ZN => 
                           n6250);
   U12651 : OAI211_X2 port map( C1 => n1881, C2 => n20631, A => n20629, B => 
                           n5317, ZN => n21601);
   U12652 : NAND2_X1 port map( A1 => n5318, A2 => n28186, ZN => n5317);
   U12653 : NAND2_X1 port map( A1 => n5322, A2 => n5321, ZN => n5320);
   U12654 : NAND2_X1 port map( A1 => n23254, A2 => n28796, ZN => n5321);
   U12655 : AND2_X1 port map( A1 => n11685, A2 => n11996, ZN => n5323);
   U12657 : OAI21_X2 port map( B1 => n5323, B2 => n11757, A => n11687, ZN => 
                           n12686);
   U12658 : OAI21_X2 port map( B1 => n5328, B2 => n18521, A => n5324, ZN => 
                           n19577);
   U12659 : NAND3_X1 port map( A1 => n27287, A2 => n27282, A3 => n27286, ZN => 
                           n5331);
   U12660 : MUX2_X1 port map( A => n5332, B => n24558, S => n25794, Z => n24563
                           );
   U12661 : NAND2_X1 port map( A1 => n20577, A2 => n20413, ZN => n5334);
   U12662 : OAI211_X1 port map( C1 => n5336, C2 => n5335, A => n27103, B => 
                           n27104, ZN => n5337);
   U12663 : XNOR2_X1 port map( A => n5337, B => n27105, ZN => Ciphertext(134));
   U12664 : OAI21_X2 port map( B1 => n21628, B2 => n22141, A => n5338, ZN => 
                           n22606);
   U12666 : NAND3_X1 port map( A1 => n5344, A2 => n5343, A3 => n14302, ZN => 
                           n5342);
   U12667 : OAI21_X1 port map( B1 => n23603, B2 => n23247, A => n5347, ZN => 
                           n5346);
   U12668 : NAND2_X1 port map( A1 => n21512, A2 => n21530, ZN => n21515);
   U12669 : NOR2_X1 port map( A1 => n14278, A2 => n14362, ZN => n5352);
   U12670 : NAND2_X1 port map( A1 => n5355, A2 => n23329, ZN => n5353);
   U12671 : NAND2_X1 port map( A1 => n5358, A2 => n5356, ZN => n21432);
   U12672 : NAND2_X1 port map( A1 => n5357, A2 => n4569, ZN => n5356);
   U12674 : NOR2_X1 port map( A1 => n6507, A2 => n29541, ZN => n26496);
   U12676 : INV_X1 port map( A => n7871, ZN => n5360);
   U12677 : NAND3_X1 port map( A1 => n5362, A2 => n7866, A3 => n5361, ZN => 
                           n8499);
   U12679 : OAI21_X1 port map( B1 => n8656, B2 => n8116, A => n8500, ZN => 
                           n8117);
   U12680 : NAND2_X1 port map( A1 => n7880, A2 => n5364, ZN => n5363);
   U12681 : OAI21_X1 port map( B1 => n7879, B2 => n7999, A => n7878, ZN => 
                           n5364);
   U12682 : XNOR2_X1 port map( A => n19568, B => n1246, ZN => n19569);
   U12683 : OR2_X1 port map( A1 => n10467, A2 => n5366, ZN => n6885);
   U12684 : AND2_X1 port map( A1 => n5377, A2 => n20644, ZN => n20646);
   U12685 : NAND3_X1 port map( A1 => n5368, A2 => n27497, A3 => n29523, ZN => 
                           n5367);
   U12686 : INV_X1 port map( A => n27492, ZN => n5368);
   U12687 : INV_X1 port map( A => n27497, ZN => n27480);
   U12688 : NAND2_X1 port map( A1 => n29522, A2 => n27496, ZN => n5369);
   U12689 : OAI22_X1 port map( A1 => n6706, A2 => n11194, B1 => n6687, B2 => 
                           n11622, ZN => n5370);
   U12690 : NAND2_X1 port map( A1 => n5603, A2 => n11953, ZN => n5371);
   U12691 : NAND2_X1 port map( A1 => n8320, A2 => n9531, ZN => n8576);
   U12692 : OAI21_X1 port map( B1 => n8320, B2 => n8610, A => n9529, ZN => 
                           n8611);
   U12693 : OAI21_X1 port map( B1 => n29662, B2 => n8320, A => n8747, ZN => 
                           n8748);
   U12694 : NAND2_X1 port map( A1 => n27038, A2 => n27213, ZN => n5372);
   U12695 : NAND2_X1 port map( A1 => n20452, A2 => n5377, ZN => n5376);
   U12696 : AOI21_X1 port map( B1 => n14394, B2 => n5378, A => n14193, ZN => 
                           n12846);
   U12698 : MUX2_X1 port map( A => n15423, B => n15101, S => n15102, Z => n5382
                           );
   U12699 : AND2_X2 port map( A1 => n12805, A2 => n12804, ZN => n15102);
   U12700 : INV_X1 port map( A => n18379, ZN => n17647);
   U12701 : OAI21_X2 port map( B1 => n17154, B2 => n17153, A => n17152, ZN => 
                           n18379);
   U12702 : NOR2_X1 port map( A1 => n28791, A2 => n21326, ZN => n20907);
   U12703 : NAND3_X1 port map( A1 => n13907, A2 => n13906, A3 => n14051, ZN => 
                           n5386);
   U12704 : NAND3_X1 port map( A1 => n23487, A2 => n6424, A3 => n23776, ZN => 
                           n5387);
   U12706 : XNOR2_X1 port map( A => n19124, B => n5393, ZN => n19128);
   U12707 : XNOR2_X1 port map( A => n19123, B => n19122, ZN => n5393);
   U12709 : INV_X1 port map( A => n8608, ZN => n5396);
   U12710 : NAND2_X1 port map( A1 => n17548, A2 => n5398, ZN => n5397);
   U12711 : XNOR2_X1 port map( A => n10393, B => n10081, ZN => n5401);
   U12712 : NAND2_X1 port map( A1 => n23694, A2 => n5402, ZN => n6441);
   U12713 : NAND2_X1 port map( A1 => n29059, A2 => n14146, ZN => n5405);
   U12715 : NAND2_X1 port map( A1 => n13958, A2 => n5409, ZN => n13961);
   U12716 : NAND2_X1 port map( A1 => n562, A2 => n14433, ZN => n5409);
   U12717 : XNOR2_X1 port map( A => n5416, B => n1046, ZN => n19543);
   U12718 : XNOR2_X1 port map( A => n5416, B => n891, ZN => n19003);
   U12719 : XNOR2_X1 port map( A => n5416, B => n2916, ZN => n18256);
   U12720 : XNOR2_X1 port map( A => n19403, B => n5416, ZN => n19607);
   U12721 : OR2_X1 port map( A1 => n18706, A2 => n18404, ZN => n18405);
   U12722 : NAND2_X1 port map( A1 => n6693, A2 => n8819, ZN => n6692);
   U12723 : NAND3_X1 port map( A1 => n17352, A2 => n17351, A3 => n5418, ZN => 
                           n17353);
   U12724 : NAND3_X1 port map( A1 => n17348, A2 => n17347, A3 => n5419, ZN => 
                           n5418);
   U12725 : NAND2_X1 port map( A1 => n5420, A2 => n17344, ZN => n5419);
   U12727 : AND3_X1 port map( A1 => n5421, A2 => n27358, A3 => n27355, ZN => 
                           n6287);
   U12728 : INV_X1 port map( A => n14362, ZN => n14359);
   U12729 : NAND2_X1 port map( A1 => n27259, A2 => n5425, ZN => n26881);
   U12730 : INV_X1 port map( A => n27255, ZN => n5425);
   U12731 : AOI22_X1 port map( A1 => n26887, A2 => n5426, B1 => n26885, B2 => 
                           n26886, ZN => n26888);
   U12732 : NAND2_X1 port map( A1 => n24028, A2 => n6664, ZN => n5427);
   U12733 : NOR2_X1 port map( A1 => n17297, A2 => n17414, ZN => n16922);
   U12734 : NAND2_X1 port map( A1 => n5430, A2 => n3234, ZN => n5429);
   U12735 : XNOR2_X1 port map( A => n25336, B => n5431, ZN => n5433);
   U12736 : XNOR2_X1 port map( A => n25150, B => n5432, ZN => n5434);
   U12738 : NAND2_X1 port map( A1 => n19807, A2 => n5436, ZN => n5435);
   U12739 : NAND2_X1 port map( A1 => n19806, A2 => n20302, ZN => n5437);
   U12741 : NAND2_X1 port map( A1 => n5234, A2 => n18227, ZN => n18389);
   U12742 : NOR2_X1 port map( A1 => n5234, A2 => n17592, ZN => n18220);
   U12743 : XNOR2_X1 port map( A => n22334, B => n22896, ZN => n22362);
   U12744 : AOI21_X1 port map( B1 => n21311, B2 => n21309, A => n21308, ZN => 
                           n5443);
   U12745 : XNOR2_X1 port map( A => n15828, B => n16071, ZN => n6637);
   U12746 : OAI21_X2 port map( B1 => n5447, B2 => n15434, A => n5446, ZN => 
                           n16071);
   U12747 : NAND2_X1 port map( A1 => n15894, A2 => n15434, ZN => n5446);
   U12748 : MUX2_X1 port map( A => n15431, B => n15432, S => n14826, Z => 
                           n15895);
   U12749 : NOR2_X1 port map( A1 => n23474, A2 => n23762, ZN => n5448);
   U12750 : NAND2_X1 port map( A1 => n2042, A2 => n8354, ZN => n5449);
   U12751 : NAND3_X1 port map( A1 => n5450, A2 => n279, A3 => n11272, ZN => 
                           n10842);
   U12752 : MUX2_X1 port map( A => n279, B => n10523, S => n5450, Z => n9555);
   U12753 : INV_X1 port map( A => n11275, ZN => n5450);
   U12754 : MUX2_X1 port map( A => n29131, B => n23762, S => n23761, Z => 
                           n23328);
   U12755 : NAND3_X1 port map( A1 => n4617, A2 => n11969, A3 => n12156, ZN => 
                           n11973);
   U12756 : NAND2_X1 port map( A1 => n12241, A2 => n4617, ZN => n11514);
   U12757 : NOR2_X1 port map( A1 => n5839, A2 => n4617, ZN => n10862);
   U12758 : NAND2_X1 port map( A1 => n5693, A2 => n14452, ZN => n5451);
   U12760 : XNOR2_X1 port map( A => n22461, B => n21856, ZN => n5453);
   U12761 : INV_X1 port map( A => n24602, ZN => n24738);
   U12763 : NAND2_X1 port map( A1 => n22355, A2 => n22354, ZN => n5456);
   U12764 : NAND2_X1 port map( A1 => n22310, A2 => n23636, ZN => n5457);
   U12765 : AND2_X1 port map( A1 => n29566, A2 => n17435, ZN => n5460);
   U12766 : NAND2_X1 port map( A1 => n5461, A2 => n17440, ZN => n5459);
   U12767 : AND2_X1 port map( A1 => n336, A2 => n17439, ZN => n5461);
   U12768 : INV_X1 port map( A => n21306, ZN => n21307);
   U12769 : NAND2_X1 port map( A1 => n20768, A2 => n29530, ZN => n20774);
   U12770 : XNOR2_X1 port map( A => n13054, B => n5463, ZN => n12551);
   U12771 : NAND2_X1 port map( A1 => n12239, A2 => n5839, ZN => n5462);
   U12772 : NAND2_X1 port map( A1 => n11612, A2 => n11613, ZN => n5464);
   U12773 : NAND2_X1 port map( A1 => n12316, A2 => n12049, ZN => n11612);
   U12774 : INV_X1 port map( A => n13054, ZN => n12790);
   U12775 : OAI21_X1 port map( B1 => n12028, B2 => n5466, A => n12026, ZN => 
                           n5467);
   U12776 : NAND2_X1 port map( A1 => n10489, A2 => n431, ZN => n5468);
   U12777 : NAND2_X1 port map( A1 => n5473, A2 => n5472, ZN => n5474);
   U12778 : NAND2_X1 port map( A1 => n18130, A2 => n18591, ZN => n5472);
   U12779 : NAND3_X1 port map( A1 => n5475, A2 => n17835, A3 => n18129, ZN => 
                           n5473);
   U12780 : OAI21_X2 port map( B1 => n5476, B2 => n17632, A => n5474, ZN => 
                           n19256);
   U12781 : NAND2_X1 port map( A1 => n17835, A2 => n18589, ZN => n17632);
   U12783 : NAND2_X1 port map( A1 => n24814, A2 => n24809, ZN => n5478);
   U12784 : OAI21_X2 port map( B1 => n14052, B2 => n14051, A => n14050, ZN => 
                           n14695);
   U12785 : NAND2_X1 port map( A1 => n7869, A2 => n5483, ZN => n7959);
   U12787 : NAND3_X1 port map( A1 => n5486, A2 => n5484, A3 => n29585, ZN => 
                           n5485);
   U12788 : NAND2_X1 port map( A1 => n27193, A2 => n27124, ZN => n5484);
   U12789 : OAI211_X1 port map( C1 => n17394, C2 => n17393, A => n5487, B => 
                           n17400, ZN => n17399);
   U12790 : NAND3_X2 port map( A1 => n11530, A2 => n11531, A3 => n5488, ZN => 
                           n13533);
   U12791 : NAND3_X1 port map( A1 => n12230, A2 => n12229, A3 => n5489, ZN => 
                           n13448);
   U12792 : NAND2_X1 port map( A1 => n11812, A2 => n13087, ZN => n5489);
   U12794 : NAND2_X1 port map( A1 => n18043, A2 => n18042, ZN => n5496);
   U12796 : OAI21_X1 port map( B1 => n27025, B2 => n28592, A => n5497, ZN => 
                           n5498);
   U12797 : NAND2_X1 port map( A1 => n393, A2 => n27029, ZN => n5497);
   U12798 : NAND2_X1 port map( A1 => n5501, A2 => n5499, ZN => n26593);
   U12799 : NAND2_X1 port map( A1 => n5500, A2 => n306, ZN => n5499);
   U12800 : MUX2_X1 port map( A => n29588, B => n27032, S => n27025, Z => n5500
                           );
   U12801 : NAND2_X1 port map( A1 => n24576, A2 => n28482, ZN => n5502);
   U12802 : NAND2_X1 port map( A1 => n26933, A2 => n5505, ZN => n26166);
   U12803 : INV_X1 port map( A => n26579, ZN => n5505);
   U12805 : INV_X1 port map( A => n26581, ZN => n26930);
   U12806 : INV_X1 port map( A => n24916, ZN => n5873);
   U12807 : NAND2_X1 port map( A1 => n5511, A2 => n5512, ZN => n5507);
   U12808 : XNOR2_X1 port map( A => n5873, B => n26083, ZN => n24753);
   U12809 : NAND3_X1 port map( A1 => n24550, A2 => n5509, A3 => n22869, ZN => 
                           n5508);
   U12810 : NAND2_X1 port map( A1 => n24554, A2 => n24555, ZN => n5510);
   U12811 : NAND2_X1 port map( A1 => n24052, A2 => n24468, ZN => n5511);
   U12812 : NAND2_X1 port map( A1 => n24467, A2 => n24053, ZN => n5512);
   U12813 : INV_X1 port map( A => n12891, ZN => n5514);
   U12814 : OAI21_X1 port map( B1 => n15209, B2 => n14960, A => n5515, ZN => 
                           n14927);
   U12815 : NAND2_X1 port map( A1 => n11608, A2 => n4197, ZN => n11492);
   U12816 : NAND2_X1 port map( A1 => n18397, A2 => n18396, ZN => n18403);
   U12817 : NAND2_X1 port map( A1 => n18232, A2 => n17977, ZN => n18396);
   U12818 : NAND2_X1 port map( A1 => n17407, A2 => n423, ZN => n5517);
   U12819 : NAND2_X1 port map( A1 => n17408, A2 => n17570, ZN => n5518);
   U12820 : AND2_X2 port map( A1 => n6765, A2 => n6900, ZN => n18232);
   U12821 : INV_X1 port map( A => n14494, ZN => n14154);
   U12823 : NAND3_X1 port map( A1 => n14154, A2 => n14498, A3 => n14493, ZN => 
                           n5519);
   U12824 : XNOR2_X1 port map( A => n18802, B => n1248, ZN => n5521);
   U12825 : XNOR2_X1 port map( A => n18761, B => n5759, ZN => n5522);
   U12826 : XNOR2_X1 port map( A => n18409, B => n18987, ZN => n5523);
   U12827 : NAND2_X1 port map( A1 => n11599, A2 => n12202, ZN => n5526);
   U12828 : NOR2_X1 port map( A1 => n10988, A2 => n10983, ZN => n10697);
   U12829 : NAND2_X1 port map( A1 => n10630, A2 => n10983, ZN => n10634);
   U12830 : OAI21_X1 port map( B1 => n16888, B2 => n17143, A => n5527, ZN => 
                           n16228);
   U12831 : NAND2_X1 port map( A1 => n17143, A2 => n17137, ZN => n5527);
   U12833 : NAND2_X1 port map( A1 => n5408, A2 => n383, ZN => n5529);
   U12834 : XNOR2_X2 port map( A => n13321, B => n13320, ZN => n5531);
   U12835 : NAND3_X1 port map( A1 => n13910, A2 => n13729, A3 => n5531, ZN => 
                           n5886);
   U12836 : NOR2_X1 port map( A1 => n28171, A2 => n5531, ZN => n13915);
   U12837 : NAND3_X1 port map( A1 => n3798, A2 => n13730, A3 => n5531, ZN => 
                           n6352);
   U12838 : AOI21_X1 port map( B1 => n13643, B2 => n13912, A => n5531, ZN => 
                           n13644);
   U12839 : NAND2_X1 port map( A1 => n5534, A2 => n11190, ZN => n5532);
   U12840 : NAND3_X1 port map( A1 => n11191, A2 => n11355, A3 => n11352, ZN => 
                           n5533);
   U12841 : NAND2_X1 port map( A1 => n11355, A2 => n11351, ZN => n5534);
   U12842 : NOR2_X1 port map( A1 => n18172, A2 => n18168, ZN => n5535);
   U12844 : XNOR2_X1 port map( A => n19590, B => n19269, ZN => n5539);
   U12845 : XNOR2_X1 port map( A => n19591, B => n19593, ZN => n5538);
   U12846 : INV_X1 port map( A => n17255, ZN => n17251);
   U12850 : NAND2_X1 port map( A1 => n12399, A2 => n14411, ZN => n5542);
   U12851 : XNOR2_X1 port map( A => n13447, B => n13227, ZN => n12834);
   U12852 : OAI22_X1 port map( A1 => n5544, A2 => n28155, B1 => n21563, B2 => 
                           n21560, ZN => n20757);
   U12853 : NAND2_X1 port map( A1 => n20418, A2 => n5545, ZN => n20419);
   U12854 : OAI22_X1 port map( A1 => n25152, A2 => n5546, B1 => n26936, B2 => 
                           n26944, ZN => n25159);
   U12855 : NAND2_X1 port map( A1 => n23420, A2 => n483, ZN => n5547);
   U12856 : NAND2_X1 port map( A1 => n29507, A2 => n17802, ZN => n18426);
   U12857 : INV_X1 port map( A => n5551, ZN => n5550);
   U12859 : NAND2_X1 port map( A1 => n23625, A2 => n23624, ZN => n5554);
   U12860 : NAND2_X1 port map( A1 => n23623, A2 => n23622, ZN => n5556);
   U12861 : OR2_X1 port map( A1 => n17298, A2 => n3234, ZN => n5557);
   U12862 : NAND2_X1 port map( A1 => n7885, A2 => n7886, ZN => n5559);
   U12863 : NAND2_X1 port map( A1 => n28479, A2 => n21091, ZN => n5560);
   U12865 : NAND2_X1 port map( A1 => n17933, A2 => n18480, ZN => n5561);
   U12867 : XNOR2_X1 port map( A => n22705, B => n27534, ZN => n22769);
   U12868 : NAND2_X1 port map( A1 => n20985, A2 => n19013, ZN => n5564);
   U12869 : NAND2_X1 port map( A1 => n20913, A2 => n19014, ZN => n5565);
   U12870 : XNOR2_X1 port map( A => n15893, B => n14523, ZN => n5566);
   U12871 : INV_X1 port map( A => n9045, ZN => n5568);
   U12872 : INV_X1 port map( A => n9233, ZN => n5567);
   U12873 : NOR2_X1 port map( A1 => n9235, A2 => n9233, ZN => n5569);
   U12874 : OAI21_X1 port map( B1 => n9233, B2 => n5945, A => n5570, ZN => 
                           n7001);
   U12875 : NAND2_X1 port map( A1 => n5160, A2 => n5945, ZN => n5570);
   U12876 : INV_X1 port map( A => n24704, ZN => n24708);
   U12877 : OAI211_X1 port map( C1 => n592, C2 => n28405, A => n5574, B => 
                           n5573, ZN => n5572);
   U12878 : NAND2_X1 port map( A1 => n592, A2 => n10936, ZN => n5574);
   U12879 : OAI21_X1 port map( B1 => n14622, B2 => n15500, A => n5577, ZN => 
                           n5576);
   U12880 : AND2_X1 port map( A1 => n14705, A2 => n15498, ZN => n14622);
   U12881 : NAND2_X1 port map( A1 => n12236, A2 => n375, ZN => n5578);
   U12882 : NAND2_X1 port map( A1 => n1986, A2 => n12236, ZN => n5579);
   U12883 : INV_X1 port map( A => n294, ZN => n5581);
   U12884 : NAND2_X1 port map( A1 => n11077, A2 => n11076, ZN => n10663);
   U12885 : INV_X1 port map( A => n11294, ZN => n11077);
   U12886 : NAND2_X1 port map( A1 => n1830, A2 => n5584, ZN => n13815);
   U12887 : NAND2_X1 port map( A1 => n13880, A2 => n5584, ZN => n13883);
   U12888 : NAND2_X1 port map( A1 => n16722, A2 => n16803, ZN => n5585);
   U12889 : NAND2_X1 port map( A1 => n16725, A2 => n3883, ZN => n16802);
   U12891 : NAND2_X1 port map( A1 => n11335, A2 => n11176, ZN => n11175);
   U12894 : NAND2_X1 port map( A1 => n6849, A2 => n5590, ZN => n6848);
   U12895 : NAND3_X1 port map( A1 => n571, A2 => n6687, A3 => n5838, ZN => 
                           n5590);
   U12896 : INV_X1 port map( A => n14972, ZN => n14583);
   U12897 : NOR2_X1 port map( A1 => n8575, A2 => n5594, ZN => n9420);
   U12898 : MUX2_X1 port map( A => n606, B => n5594, S => n7569, Z => n8582);
   U12899 : NAND3_X1 port map( A1 => n5129, A2 => n5594, A3 => n603, ZN => 
                           n8768);
   U12900 : OAI21_X1 port map( B1 => n5129, B2 => n5594, A => n5592, ZN => 
                           n9422);
   U12901 : OAI21_X1 port map( B1 => n8327, B2 => n606, A => n9425, ZN => n5593
                           );
   U12903 : NAND2_X1 port map( A1 => n11184, A2 => n29316, ZN => n11185);
   U12904 : OAI211_X1 port map( C1 => n11321, C2 => n29316, A => n10473, B => 
                           n11183, ZN => n10475);
   U12906 : MUX2_X1 port map( A => n15167, B => n15166, S => n15165, Z => n5597
                           );
   U12907 : NAND2_X1 port map( A1 => n15169, A2 => n15168, ZN => n5599);
   U12908 : NOR2_X1 port map( A1 => n27409, A2 => n1175, ZN => n5601);
   U12909 : INV_X1 port map( A => n27403, ZN => n5600);
   U12910 : NAND2_X1 port map( A1 => n5601, A2 => n5600, ZN => n25638);
   U12911 : NOR2_X1 port map( A1 => n27403, A2 => n27409, ZN => n5602);
   U12912 : NOR2_X1 port map( A1 => n25634, A2 => n5602, ZN => n25640);
   U12913 : XNOR2_X1 port map( A => n13226, B => n13451, ZN => n11629);
   U12914 : INV_X1 port map( A => n27496, ZN => n5607);
   U12915 : INV_X1 port map( A => n5605, ZN => n27476);
   U12916 : INV_X1 port map( A => n27494, ZN => n5604);
   U12917 : NAND2_X1 port map( A1 => n5608, A2 => n5607, ZN => n5606);
   U12918 : NOR2_X1 port map( A1 => n29523, A2 => n27497, ZN => n5608);
   U12919 : NAND2_X1 port map( A1 => n16953, A2 => n17359, ZN => n16714);
   U12920 : OAI21_X1 port map( B1 => n23759, B2 => n23760, A => n23758, ZN => 
                           n5611);
   U12922 : XNOR2_X2 port map( A => n5613, B => n5612, ZN => n6114);
   U12923 : XNOR2_X1 port map( A => n18989, B => n18990, ZN => n5612);
   U12924 : XNOR2_X1 port map( A => n18987, B => n18988, ZN => n5613);
   U12925 : NAND2_X1 port map( A1 => n14127, A2 => n5615, ZN => n14129);
   U12926 : NOR2_X1 port map( A1 => n14353, A2 => n14126, ZN => n5615);
   U12927 : NAND2_X1 port map( A1 => n5617, A2 => n14126, ZN => n5616);
   U12928 : INV_X1 port map( A => n14354, ZN => n5617);
   U12930 : NAND2_X1 port map( A1 => n16601, A2 => n17109, ZN => n5620);
   U12931 : XNOR2_X1 port map( A => n14983, B => n5621, ZN => n14984);
   U12932 : XNOR2_X1 port map( A => n16650, B => n5621, ZN => n16651);
   U12933 : OAI211_X2 port map( C1 => n24524, C2 => n24525, A => n24528, B => 
                           n6223, ZN => n25948);
   U12934 : OAI21_X2 port map( B1 => n5622, B2 => n20143, A => n20142, ZN => 
                           n22270);
   U12936 : NAND2_X1 port map( A1 => n6656, A2 => n5623, ZN => n6655);
   U12937 : INV_X1 port map( A => n27433, ZN => n27441);
   U12939 : NAND2_X1 port map( A1 => n437, A2 => n7993, ZN => n7241);
   U12940 : XNOR2_X2 port map( A => n7056, B => Key(165), ZN => n7993);
   U12941 : OAI21_X1 port map( B1 => n23171, B2 => n23516, A => n23170, ZN => 
                           n5626);
   U12942 : AOI21_X1 port map( B1 => n23681, B2 => n5883, A => n29544, ZN => 
                           n5627);
   U12943 : OAI211_X1 port map( C1 => n5632, C2 => n6420, A => n5631, B => 
                           n5628, ZN => n5629);
   U12944 : NAND2_X1 port map( A1 => n6420, A2 => n5633, ZN => n5628);
   U12945 : XNOR2_X1 port map( A => n25820, B => n5629, ZN => n5630);
   U12946 : XNOR2_X1 port map( A => n25071, B => n5630, ZN => n25073);
   U12948 : NAND2_X1 port map( A1 => n6422, A2 => n5633, ZN => n5631);
   U12950 : XNOR2_X2 port map( A => n13356, B => n13357, ZN => n13914);
   U12951 : NAND2_X1 port map( A1 => n5637, A2 => n12512, ZN => n11837);
   U12953 : NAND3_X1 port map( A1 => n15892, A2 => n18299, A3 => n18298, ZN => 
                           n18300);
   U12954 : AOI21_X1 port map( B1 => n5645, B2 => n5644, A => n15494, ZN => 
                           n5640);
   U12956 : NAND2_X1 port map( A1 => n22955, A2 => n28484, ZN => n5646);
   U12957 : NAND2_X1 port map( A1 => n22956, A2 => n28183, ZN => n5647);
   U12958 : XNOR2_X1 port map( A => n5650, B => n5649, ZN => Ciphertext(16));
   U12961 : NAND2_X1 port map( A1 => n26612, A2 => n26613, ZN => n5652);
   U12963 : NAND2_X1 port map( A1 => n24729, A2 => n24598, ZN => n5653);
   U12965 : NAND2_X1 port map( A1 => n5656, A2 => n460, ZN => n5655);
   U12966 : NOR2_X1 port map( A1 => n24730, A2 => n24726, ZN => n5656);
   U12967 : NAND2_X1 port map( A1 => n19832, A2 => n5657, ZN => n21758);
   U12968 : MUX2_X1 port map( A => n20864, B => n21497, S => n21493, Z => n5658
                           );
   U12969 : INV_X1 port map( A => n18344, ZN => n5659);
   U12970 : OAI21_X1 port map( B1 => n11954, B2 => n11580, A => n5661, ZN => 
                           n5660);
   U12971 : AOI22_X1 port map( A1 => n1924, A2 => n21420, B1 => n5664, B2 => 
                           n21087, ZN => n5663);
   U12972 : NOR2_X1 port map( A1 => n21425, A2 => n21424, ZN => n5664);
   U12973 : NAND2_X1 port map( A1 => n21427, A2 => n28602, ZN => n5665);
   U12974 : NOR2_X1 port map( A1 => n7114, A2 => n8828, ZN => n7447);
   U12975 : INV_X1 port map( A => n8828, ZN => n8193);
   U12976 : NAND2_X1 port map( A1 => n5667, A2 => n14177, ZN => n5666);
   U12977 : OAI21_X1 port map( B1 => n14451, B2 => n13753, A => n14450, ZN => 
                           n5667);
   U12978 : OR2_X1 port map( A1 => n20181, A2 => n20182, ZN => n5668);
   U12979 : NAND2_X1 port map( A1 => n20163, A2 => n20162, ZN => n5669);
   U12980 : AND2_X1 port map( A1 => n17883, A2 => n18379, ZN => n5671);
   U12981 : NAND2_X1 port map( A1 => n3283, A2 => n5671, ZN => n17884);
   U12984 : NAND2_X1 port map( A1 => n8661, A2 => n8910, ZN => n5677);
   U12985 : NAND2_X1 port map( A1 => n9015, A2 => n8908, ZN => n8661);
   U12986 : INV_X1 port map( A => n14916, ZN => n5679);
   U12987 : NAND2_X1 port map( A1 => n14500, A2 => n14501, ZN => n5678);
   U12988 : NAND3_X1 port map( A1 => n15488, A2 => n15487, A3 => n5679, ZN => 
                           n15493);
   U12989 : NAND2_X1 port map( A1 => n21495, A2 => n21493, ZN => n21126);
   U12990 : NAND2_X1 port map( A1 => n19850, A2 => n19851, ZN => n5680);
   U12991 : NAND3_X1 port map( A1 => n5680, A2 => n20394, A3 => n20560, ZN => 
                           n19853);
   U12992 : NAND2_X1 port map( A1 => n14657, A2 => n548, ZN => n5681);
   U12994 : NAND2_X1 port map( A1 => n12977, A2 => n5682, ZN => n14874);
   U12995 : NOR2_X1 port map( A1 => n21322, A2 => n5684, ZN => n20575);
   U12996 : NAND2_X1 port map( A1 => n28584, A2 => n5684, ZN => n6043);
   U13000 : NAND2_X1 port map( A1 => n26625, A2 => n27013, ZN => n5687);
   U13001 : NAND2_X1 port map( A1 => n5691, A2 => n5689, ZN => n5688);
   U13002 : NAND3_X1 port map( A1 => n5690, A2 => n18216, A3 => n18500, ZN => 
                           n5689);
   U13003 : INV_X1 port map( A => n13753, ZN => n5693);
   U13004 : INV_X1 port map( A => n17543, ZN => n5695);
   U13005 : INV_X1 port map( A => n17543, ZN => n17217);
   U13006 : XNOR2_X2 port map( A => n15800, B => n15799, ZN => n17540);
   U13007 : NAND2_X1 port map( A1 => n22676, A2 => n5699, ZN => n5698);
   U13008 : NAND3_X1 port map( A1 => n18346, A2 => n17948, A3 => n514, ZN => 
                           n5700);
   U13009 : XNOR2_X1 port map( A => n21876, B => n22809, ZN => n5702);
   U13010 : XNOR2_X1 port map( A => n21877, B => n21878, ZN => n5703);
   U13012 : OR2_X1 port map( A1 => n11237, A2 => n11235, ZN => n5707);
   U13014 : XNOR2_X2 port map( A => n9738, B => n9739, ZN => n11237);
   U13015 : NAND2_X1 port map( A1 => n23296, A2 => n22864, ZN => n23298);
   U13019 : OAI211_X1 port map( C1 => n12288, C2 => n12289, A => n3558, B => 
                           n5715, ZN => n12295);
   U13020 : XNOR2_X1 port map( A => n5718, B => n22501, ZN => n22503);
   U13022 : NAND2_X1 port map( A1 => n5725, A2 => n5726, ZN => n5723);
   U13023 : INV_X1 port map( A => n15502, ZN => n5726);
   U13024 : NOR2_X1 port map( A1 => n15506, A2 => n15265, ZN => n5724);
   U13025 : NOR2_X1 port map( A1 => n15500, A2 => n15265, ZN => n5725);
   U13026 : INV_X1 port map( A => n24077, ZN => n5728);
   U13027 : NAND2_X1 port map( A1 => n5729, A2 => n28401, ZN => n23508);
   U13028 : AND2_X1 port map( A1 => n24081, A2 => n24133, ZN => n5729);
   U13029 : NAND3_X1 port map( A1 => n23911, A2 => n24079, A3 => n28401, ZN => 
                           n23912);
   U13030 : OAI211_X1 port map( C1 => n14774, C2 => n14775, A => n14773, B => 
                           n14812, ZN => n14776);
   U13031 : NAND2_X1 port map( A1 => n14772, A2 => n14807, ZN => n14812);
   U13032 : INV_X1 port map( A => n14051, ZN => n5731);
   U13035 : NAND2_X1 port map( A1 => n16538, A2 => n4703, ZN => n5734);
   U13036 : NOR2_X1 port map( A1 => n393, A2 => n306, ZN => n24826);
   U13037 : AOI21_X1 port map( B1 => n393, B2 => n306, A => n27032, ZN => 
                           n26692);
   U13038 : AOI21_X1 port map( B1 => n26691, B2 => n26819, A => n393, ZN => 
                           n26694);
   U13040 : NOR2_X1 port map( A1 => n24823, A2 => n1978, ZN => n5735);
   U13041 : OAI211_X1 port map( C1 => n17078, C2 => n5738, A => n4655, B => 
                           n5736, ZN => n5739);
   U13042 : INV_X1 port map( A => n17148, ZN => n5737);
   U13043 : INV_X1 port map( A => n17485, ZN => n5738);
   U13044 : NAND2_X1 port map( A1 => n17490, A2 => n17489, ZN => n5740);
   U13045 : NAND2_X1 port map( A1 => n23759, A2 => n23760, ZN => n5741);
   U13047 : NAND2_X1 port map( A1 => n13953, A2 => n14194, ZN => n5745);
   U13048 : XNOR2_X1 port map( A => n19520, B => n5746, ZN => n18929);
   U13049 : AND3_X2 port map( A1 => n5747, A2 => n17594, A3 => n17595, ZN => 
                           n19139);
   U13050 : XNOR2_X1 port map( A => n25440, B => n25819, ZN => n25113);
   U13052 : NAND2_X1 port map( A1 => n5751, A2 => n5752, ZN => n5748);
   U13053 : NAND2_X1 port map( A1 => n5753, A2 => n11308, ZN => n5835);
   U13054 : MUX2_X1 port map( A => n11309, B => n11310, S => n1933, Z => n11311
                           );
   U13055 : MUX2_X1 port map( A => n23445, B => n23442, S => n23448, Z => 
                           n23111);
   U13056 : XNOR2_X1 port map( A => n24924, B => n24926, ZN => n5755);
   U13058 : XNOR2_X1 port map( A => n19289, B => n19290, ZN => n19295);
   U13060 : NAND2_X1 port map( A1 => n5757, A2 => n18401, ZN => n5756);
   U13061 : NAND2_X1 port map( A1 => n18403, A2 => n18402, ZN => n5758);
   U13062 : OR2_X1 port map( A1 => n5760, A2 => n26748, ZN => n25644);
   U13063 : AND2_X1 port map( A1 => n26748, A2 => n5760, ZN => n25979);
   U13064 : NAND2_X1 port map( A1 => n29099, A2 => n28563, ZN => n5761);
   U13065 : NOR2_X1 port map( A1 => n28583, A2 => n5760, ZN => n25978);
   U13066 : MUX2_X1 port map( A => n28583, B => n26224, S => n28563, Z => 
                           n26225);
   U13071 : NAND2_X1 port map( A1 => n7116, A2 => n7320, ZN => n7768);
   U13072 : NAND2_X1 port map( A1 => n7321, A2 => n7116, ZN => n7322);
   U13073 : AOI21_X1 port map( B1 => n7769, B2 => n7116, A => n614, ZN => n7325
                           );
   U13074 : NAND2_X1 port map( A1 => n24729, A2 => n5767, ZN => n24290);
   U13075 : NAND2_X1 port map( A1 => n460, A2 => n5768, ZN => n24147);
   U13076 : INV_X1 port map( A => n5769, ZN => n6310);
   U13077 : OAI21_X1 port map( B1 => n5770, B2 => n23492, A => n23799, ZN => 
                           n5769);
   U13078 : OAI22_X1 port map( A1 => n23011, A2 => n23351, B1 => n5773, B2 => 
                           n23657, ZN => n23659);
   U13079 : INV_X1 port map( A => n23351, ZN => n5774);
   U13080 : NAND2_X1 port map( A1 => n11377, A2 => n12166, ZN => n11843);
   U13081 : INV_X1 port map( A => n22284, ZN => n23628);
   U13082 : NAND2_X1 port map( A1 => n23040, A2 => n23309, ZN => n23041);
   U13083 : INV_X1 port map( A => n23633, ZN => n5775);
   U13084 : OR2_X1 port map( A1 => n27771, A2 => n5776, ZN => n27775);
   U13085 : NAND2_X1 port map( A1 => n15047, A2 => n15238, ZN => n5777);
   U13087 : INV_X1 port map( A => n20041, ZN => n5778);
   U13088 : NAND2_X1 port map( A1 => n5781, A2 => n20646, ZN => n5779);
   U13090 : XNOR2_X1 port map( A => n16481, B => n16479, ZN => n5784);
   U13091 : XNOR2_X1 port map( A => n16399, B => n16398, ZN => n16488);
   U13092 : OAI211_X2 port map( C1 => n3362, C2 => n5788, A => n5786, B => 
                           n5785, ZN => n16398);
   U13093 : NAND3_X1 port map( A1 => n3362, A2 => n15407, A3 => n15406, ZN => 
                           n5786);
   U13095 : NAND2_X1 port map( A1 => n29312, A2 => n14250, ZN => n5936);
   U13096 : NAND2_X1 port map( A1 => n5789, A2 => n29312, ZN => n5790);
   U13097 : NAND2_X1 port map( A1 => n16491, A2 => n17829, ZN => n5792);
   U13098 : NAND2_X1 port map( A1 => n17073, A2 => n17506, ZN => n16550);
   U13099 : NAND2_X1 port map( A1 => n19768, A2 => n5793, ZN => n21145);
   U13100 : NAND3_X1 port map( A1 => n18919, A2 => n5794, A3 => n20106, ZN => 
                           n5793);
   U13101 : NOR2_X1 port map( A1 => n20704, A2 => n20967, ZN => n20705);
   U13102 : NAND2_X1 port map( A1 => n381, A2 => n20972, ZN => n20704);
   U13103 : AND2_X1 port map( A1 => n14697, A2 => n15513, ZN => n15276);
   U13104 : NAND2_X1 port map( A1 => n5168, A2 => n24017, ZN => n5799);
   U13105 : XNOR2_X1 port map( A => n5801, B => n21903, ZN => n22620);
   U13106 : INV_X1 port map( A => n21987, ZN => n5801);
   U13107 : XNOR2_X1 port map( A => n21903, B => n5802, ZN => n22101);
   U13108 : INV_X1 port map( A => n21903, ZN => n5803);
   U13109 : NAND2_X1 port map( A1 => n558, A2 => n14158, ZN => n14159);
   U13111 : NOR2_X1 port map( A1 => n29320, A2 => n14479, ZN => n5804);
   U13113 : NAND2_X1 port map( A1 => n17070, A2 => n17830, ZN => n17513);
   U13114 : NAND2_X1 port map( A1 => n5808, A2 => n17070, ZN => n5807);
   U13115 : NAND2_X1 port map( A1 => n5812, A2 => n5810, ZN => n13791);
   U13117 : INV_X1 port map( A => n14882, ZN => n5811);
   U13118 : NAND2_X1 port map( A1 => n13790, A2 => n5813, ZN => n5812);
   U13119 : NAND2_X1 port map( A1 => n1896, A2 => n14044, ZN => n6010);
   U13120 : NOR2_X1 port map( A1 => n28626, A2 => n23416, ZN => n22928);
   U13121 : MUX2_X1 port map( A => n23417, B => n28626, S => n23416, Z => n6091
                           );
   U13122 : MUX2_X1 port map( A => n23419, B => n28626, S => n5856, Z => n22808
                           );
   U13123 : XNOR2_X1 port map( A => n22459, B => n22123, ZN => n20923);
   U13126 : OAI21_X1 port map( B1 => n20802, B2 => n5817, A => n20801, ZN => 
                           n20803);
   U13127 : OAI21_X1 port map( B1 => n20955, B2 => n29586, A => n5816, ZN => 
                           n21101);
   U13128 : NAND2_X1 port map( A1 => n21930, A2 => n21099, ZN => n5816);
   U13129 : OR2_X1 port map( A1 => n21934, A2 => n5817, ZN => n6345);
   U13131 : XOR2_X1 port map( A => n10087, B => n10426, Z => n5818);
   U13132 : AND2_X1 port map( A1 => n8117, A2 => n8502, ZN => n5819);
   U13134 : NAND2_X1 port map( A1 => n13757, A2 => n14158, ZN => n5822);
   U13135 : NAND2_X1 port map( A1 => n14162, A2 => n13756, ZN => n5823);
   U13136 : NAND2_X1 port map( A1 => n14474, A2 => n13754, ZN => n14162);
   U13137 : XNOR2_X1 port map( A => n9924, B => n5824, ZN => n8520);
   U13138 : INV_X1 port map( A => n5824, ZN => n10320);
   U13139 : XNOR2_X1 port map( A => n10250, B => n10386, ZN => n5824);
   U13140 : NAND2_X1 port map( A1 => n5825, A2 => n12203, ZN => n6073);
   U13141 : NAND2_X1 port map( A1 => n20587, A2 => n20584, ZN => n6914);
   U13144 : NAND2_X1 port map( A1 => n5827, A2 => n21424, ZN => n21422);
   U13145 : NAND2_X1 port map( A1 => n5827, A2 => n20899, ZN => n20804);
   U13146 : NOR2_X1 port map( A1 => n21425, A2 => n5827, ZN => n20140);
   U13147 : INV_X1 port map( A => n16588, ZN => n5828);
   U13149 : NAND3_X1 port map( A1 => n5832, A2 => n25405, A3 => n5831, ZN => 
                           n26708);
   U13150 : NAND2_X1 port map( A1 => n26463, A2 => n26469, ZN => n5832);
   U13151 : NAND2_X1 port map( A1 => n25008, A2 => n25005, ZN => n24305);
   U13152 : NOR2_X1 port map( A1 => n388, A2 => n14882, ZN => n6061);
   U13154 : NAND2_X1 port map( A1 => n24338, A2 => n24341, ZN => n24128);
   U13155 : NAND3_X1 port map( A1 => n24708, A2 => n24338, A3 => n24707, ZN => 
                           n24342);
   U13156 : OAI21_X1 port map( B1 => n6611, B2 => n24338, A => n5836, ZN => 
                           n25543);
   U13157 : XNOR2_X1 port map( A => n5841, B => n5840, ZN => n22283);
   U13158 : NAND2_X1 port map( A1 => n16615, A2 => n5844, ZN => n5843);
   U13159 : NAND2_X1 port map( A1 => n518, A2 => n18356, ZN => n5844);
   U13160 : NAND2_X1 port map( A1 => n5847, A2 => n5846, ZN => n5845);
   U13161 : NOR2_X1 port map( A1 => n13912, A2 => n13914, ZN => n5846);
   U13162 : NAND2_X1 port map( A1 => n13914, A2 => n13915, ZN => n5848);
   U13163 : XNOR2_X1 port map( A => n5849, B => n26409, ZN => Ciphertext(178));
   U13164 : OAI211_X1 port map( C1 => n26408, C2 => n29031, A => n5851, B => 
                           n5850, ZN => n5849);
   U13165 : OAI21_X1 port map( B1 => n5852, B2 => n28040, A => n6859, ZN => 
                           n5851);
   U13166 : AND2_X1 port map( A1 => n28024, A2 => n28027, ZN => n28040);
   U13167 : AND2_X1 port map( A1 => n28025, A2 => n29031, ZN => n5852);
   U13168 : NOR2_X1 port map( A1 => n21213, A2 => n21211, ZN => n5855);
   U13169 : MUX2_X1 port map( A => n25750, B => n27074, S => n27076, Z => 
                           n25770);
   U13170 : MUX2_X1 port map( A => n27074, B => n27075, S => n27076, Z => 
                           n27900);
   U13171 : MUX2_X1 port map( A => n25767, B => n25768, S => n27076, Z => 
                           n25769);
   U13172 : INV_X1 port map( A => n23073, ZN => n5856);
   U13173 : XNOR2_X1 port map( A => n14997, B => n5858, ZN => n5859);
   U13176 : NAND2_X1 port map( A1 => n20340, A2 => n20504, ZN => n5865);
   U13177 : NAND2_X1 port map( A1 => n15006, A2 => n5866, ZN => n15772);
   U13178 : INV_X1 port map( A => n8521, ZN => n8812);
   U13181 : NOR2_X1 port map( A1 => n5869, A2 => n8810, ZN => n5868);
   U13182 : OR2_X1 port map( A1 => n8808, A2 => n8521, ZN => n5870);
   U13183 : XNOR2_X1 port map( A => n5872, B => n24916, ZN => n25722);
   U13184 : INV_X1 port map( A => n24949, ZN => n5872);
   U13185 : XNOR2_X1 port map( A => n25244, B => n5873, ZN => n25245);
   U13186 : NAND3_X1 port map( A1 => n5877, A2 => n27653, A3 => n5874, ZN => 
                           n27654);
   U13190 : MUX2_X1 port map( A => n29090, B => n27663, S => n27672, Z => 
                           n27196);
   U13191 : XNOR2_X1 port map( A => n22481, B => n22502, ZN => n22022);
   U13192 : NAND4_X2 port map( A1 => n5880, A2 => n5878, A3 => n20949, A4 => 
                           n5879, ZN => n22692);
   U13193 : NAND2_X1 port map( A1 => n20947, A2 => n28185, ZN => n5880);
   U13194 : INV_X1 port map( A => n28457, ZN => n5882);
   U13195 : NAND2_X1 port map( A1 => n23517, A2 => n474, ZN => n23518);
   U13197 : INV_X1 port map( A => n23682, ZN => n5883);
   U13198 : INV_X1 port map( A => n13912, ZN => n14068);
   U13199 : INV_X1 port map( A => n13913, ZN => n5887);
   U13200 : NAND2_X1 port map( A1 => n8526, A2 => n5888, ZN => n5961);
   U13201 : INV_X1 port map( A => n8687, ZN => n5888);
   U13204 : NAND2_X1 port map( A1 => n17005, A2 => n5891, ZN => n16974);
   U13205 : OAI21_X1 port map( B1 => n17720, B2 => n17425, A => n5891, ZN => 
                           n14227);
   U13206 : NAND2_X1 port map( A1 => n14712, A2 => n13922, ZN => n5894);
   U13207 : XNOR2_X1 port map( A => n21982, B => n22152, ZN => n22596);
   U13208 : NAND2_X1 port map( A1 => n21304, A2 => n21305, ZN => n5897);
   U13209 : NAND3_X1 port map( A1 => n11947, A2 => n11952, A3 => n11951, ZN => 
                           n5901);
   U13210 : NAND2_X1 port map( A1 => n10917, A2 => n10605, ZN => n5902);
   U13211 : NAND2_X1 port map( A1 => n10914, A2 => n10913, ZN => n5903);
   U13212 : XNOR2_X1 port map( A => n19472, B => n19473, ZN => n19479);
   U13214 : NAND2_X1 port map( A1 => n17860, A2 => n17859, ZN => n5906);
   U13215 : NAND2_X1 port map( A1 => n18526, A2 => n18081, ZN => n5907);
   U13216 : NAND2_X1 port map( A1 => n18525, A2 => n5909, ZN => n5908);
   U13217 : NAND3_X1 port map( A1 => n5913, A2 => n5915, A3 => n5912, ZN => 
                           n12257);
   U13218 : NAND2_X1 port map( A1 => n5914, A2 => n5916, ZN => n5912);
   U13219 : NAND3_X1 port map( A1 => n5917, A2 => n28157, A3 => n5914, ZN => 
                           n5913);
   U13220 : OAI21_X1 port map( B1 => n10749, B2 => n3585, A => n28638, ZN => 
                           n5915);
   U13221 : NOR2_X1 port map( A1 => n28569, A2 => n5918, ZN => n13718);
   U13222 : NAND2_X1 port map( A1 => n13587, A2 => n5918, ZN => n14037);
   U13223 : NAND2_X1 port map( A1 => n13997, A2 => n5918, ZN => n13998);
   U13224 : NAND2_X1 port map( A1 => n17182, A2 => n17183, ZN => n5921);
   U13225 : XNOR2_X1 port map( A => n25436, B => n26007, ZN => n25395);
   U13226 : NAND2_X1 port map( A1 => n24149, A2 => n5923, ZN => n5922);
   U13227 : INV_X1 port map( A => n24740, ZN => n5923);
   U13228 : XNOR2_X1 port map( A => n7415, B => n7329, ZN => n5925);
   U13229 : INV_X1 port map( A => n21084, ZN => n5927);
   U13230 : INV_X1 port map( A => n20141, ZN => n5929);
   U13231 : INV_X1 port map( A => n16575, ZN => n15701);
   U13235 : NAND2_X1 port map( A1 => n14237, A2 => n5936, ZN => n13939);
   U13236 : NAND2_X1 port map( A1 => n18838, A2 => n20077, ZN => n5937);
   U13238 : NAND3_X1 port map( A1 => n21028, A2 => n21029, A3 => n22142, ZN => 
                           n5938);
   U13239 : INV_X1 port map( A => n22140, ZN => n5939);
   U13240 : XNOR2_X1 port map( A => n16526, B => n16605, ZN => n16138);
   U13241 : INV_X1 port map( A => n16138, ZN => n16139);
   U13242 : XNOR2_X1 port map( A => n14850, B => n16138, ZN => n14870);
   U13243 : INV_X1 port map( A => n17847, ZN => n18138);
   U13244 : OAI211_X2 port map( C1 => n21579, C2 => n5142, A => n5942, B => 
                           n5941, ZN => n22033);
   U13245 : NAND2_X1 port map( A1 => n20849, A2 => n5142, ZN => n5941);
   U13246 : INV_X1 port map( A => n23126, ZN => n6556);
   U13247 : NAND2_X1 port map( A1 => n9045, A2 => n9230, ZN => n5944);
   U13248 : NAND2_X1 port map( A1 => n14315, A2 => n14320, ZN => n5949);
   U13249 : XNOR2_X1 port map( A => n5950, B => n17779, ZN => n19949);
   U13250 : XNOR2_X1 port map( A => n5951, B => n18670, ZN => n5950);
   U13251 : XNOR2_X1 port map( A => n17770, B => n5952, ZN => n5951);
   U13253 : OAI21_X1 port map( B1 => n21463, B2 => n5953, A => n6636, ZN => 
                           n20863);
   U13254 : NAND2_X1 port map( A1 => n5955, A2 => n5954, ZN => n21469);
   U13255 : OR2_X1 port map( A1 => n21465, A2 => n21561, ZN => n5954);
   U13256 : NAND2_X1 port map( A1 => n29236, A2 => n21465, ZN => n5955);
   U13257 : NAND2_X1 port map( A1 => n6072, A2 => n9146, ZN => n9373);
   U13258 : NAND3_X1 port map( A1 => n6072, A2 => n9146, A3 => n5958, ZN => 
                           n5957);
   U13260 : NAND2_X1 port map( A1 => n8592, A2 => n8817, ZN => n5962);
   U13261 : OAI21_X1 port map( B1 => n12133, B2 => n11574, A => n5963, ZN => 
                           n5966);
   U13263 : OR2_X1 port map( A1 => n16768, A2 => n5968, ZN => n5967);
   U13264 : AND2_X2 port map( A1 => n6252, A2 => n6254, ZN => n15361);
   U13265 : NAND2_X1 port map( A1 => n14508, A2 => n15360, ZN => n5970);
   U13266 : NAND2_X1 port map( A1 => n23407, A2 => n5971, ZN => n24387);
   U13267 : INV_X1 port map( A => n12516, ZN => n5974);
   U13268 : NAND2_X1 port map( A1 => n5974, A2 => n12578, ZN => n5973);
   U13269 : NAND3_X1 port map( A1 => n5978, A2 => n14393, A3 => n14192, ZN => 
                           n5977);
   U13270 : NAND2_X1 port map( A1 => n13952, A2 => n13953, ZN => n5979);
   U13271 : NAND2_X1 port map( A1 => n14192, A2 => n14194, ZN => n5980);
   U13272 : INV_X1 port map( A => n14194, ZN => n5981);
   U13273 : NAND2_X1 port map( A1 => n17266, A2 => n17267, ZN => n17268);
   U13274 : INV_X1 port map( A => n5984, ZN => n6644);
   U13275 : XNOR2_X1 port map( A => n5984, B => n9242, ZN => n10063);
   U13276 : XNOR2_X1 port map( A => n29136, B => n1984, ZN => n22637);
   U13277 : NAND2_X1 port map( A1 => n17065, A2 => n16797, ZN => n5988);
   U13278 : NAND2_X1 port map( A1 => n7700, A2 => n5990, ZN => n5989);
   U13279 : NAND2_X1 port map( A1 => n7368, A2 => n7367, ZN => n5990);
   U13280 : NAND2_X1 port map( A1 => n5991, A2 => n28509, ZN => n23958);
   U13281 : NAND2_X1 port map( A1 => n17987, A2 => n29603, ZN => n5992);
   U13282 : XNOR2_X1 port map( A => n19568, B => n27298, ZN => n19017);
   U13283 : NAND2_X1 port map( A1 => n27673, A2 => n27671, ZN => n27664);
   U13284 : NAND2_X1 port map( A1 => n2011, A2 => n5994, ZN => n5993);
   U13285 : XNOR2_X1 port map( A => n5995, B => n1853, ZN => n9843);
   U13286 : INV_X1 port map( A => n8883, ZN => n5996);
   U13287 : INV_X1 port map( A => n12151, ZN => n12149);
   U13291 : NAND2_X1 port map( A1 => n6000, A2 => n14091, ZN => n14120);
   U13292 : NOR2_X1 port map( A1 => n14366, A2 => n6000, ZN => n6045);
   U13293 : NAND3_X1 port map( A1 => n14366, A2 => n6000, A3 => n14365, ZN => 
                           n14367);
   U13294 : NAND2_X1 port map( A1 => n13834, A2 => n6000, ZN => n6046);
   U13295 : NAND2_X1 port map( A1 => n17304, A2 => n6002, ZN => n17013);
   U13297 : NAND3_X1 port map( A1 => n15361, A2 => n14752, A3 => n6674, ZN => 
                           n6004);
   U13298 : NAND2_X1 port map( A1 => n6007, A2 => n6005, ZN => n27691);
   U13299 : NAND2_X1 port map( A1 => n6009, A2 => n6006, ZN => n6005);
   U13300 : NAND2_X1 port map( A1 => n6008, A2 => n455, ZN => n6006);
   U13301 : NAND2_X1 port map( A1 => n26127, A2 => n27702, ZN => n6007);
   U13302 : AOI21_X1 port map( B1 => n27700, B2 => n27701, A => n27702, ZN => 
                           n6009);
   U13303 : MUX2_X1 port map( A => n14044, B => n14046, S => n14047, Z => 
                           n13908);
   U13304 : NAND2_X1 port map( A1 => n13468, A2 => n6010, ZN => n13470);
   U13305 : MUX2_X1 port map( A => n14046, B => n13576, S => n1896, Z => n13580
                           );
   U13306 : OAI21_X1 port map( B1 => n17008, B2 => n17431, A => n6012, ZN => 
                           n17010);
   U13307 : NAND2_X1 port map( A1 => n16846, A2 => n17426, ZN => n6012);
   U13308 : INV_X1 port map( A => n17716, ZN => n6013);
   U13309 : XNOR2_X1 port map( A => n6018, B => n26101, ZN => n26105);
   U13310 : NOR2_X1 port map( A1 => n2656, A2 => n6526, ZN => n6019);
   U13311 : NAND2_X1 port map( A1 => n11053, A2 => n11165, ZN => n6411);
   U13312 : OR2_X1 port map( A1 => n12202, A2 => n2063, ZN => n8650);
   U13313 : NAND2_X1 port map( A1 => n11599, A2 => n6020, ZN => n11601);
   U13314 : OAI21_X1 port map( B1 => n11127, B2 => n11119, A => n11118, ZN => 
                           n6021);
   U13315 : NAND2_X1 port map( A1 => n15102, A2 => n14575, ZN => n6023);
   U13316 : OAI21_X1 port map( B1 => n26296, B2 => n26351, A => n26295, ZN => 
                           n6025);
   U13318 : AOI22_X1 port map( A1 => n26326, A2 => n27142, B1 => n26519, B2 => 
                           n29633, ZN => n6026);
   U13319 : AND2_X1 port map( A1 => n29070, A2 => n27772, ZN => n26298);
   U13320 : NAND2_X1 port map( A1 => n19999, A2 => n20353, ZN => n6028);
   U13321 : NAND2_X1 port map( A1 => n19997, A2 => n20480, ZN => n20353);
   U13323 : NAND2_X1 port map( A1 => n6029, A2 => n18357, ZN => n18358);
   U13324 : OAI21_X1 port map( B1 => n518, B2 => n18356, A => n6030, ZN => 
                           n6029);
   U13325 : NAND3_X1 port map( A1 => n6033, A2 => n29544, A3 => n23679, ZN => 
                           n23017);
   U13326 : NAND2_X1 port map( A1 => n23167, A2 => n23680, ZN => n6033);
   U13327 : INV_X1 port map( A => n23016, ZN => n6034);
   U13328 : INV_X1 port map( A => n23167, ZN => n6035);
   U13329 : AOI22_X1 port map( A1 => n29120, A2 => n24800, B1 => n24804, B2 => 
                           n24806, ZN => n24506);
   U13330 : NAND3_X1 port map( A1 => n6038, A2 => n6037, A3 => n18457, ZN => 
                           n6036);
   U13331 : OAI21_X1 port map( B1 => n17902, B2 => n18111, A => n18456, ZN => 
                           n6037);
   U13332 : NAND2_X1 port map( A1 => n20887, A2 => n21591, ZN => n6040);
   U13333 : MUX2_X1 port map( A => n6043, B => n6042, S => n21591, Z => n6041);
   U13334 : OAI21_X1 port map( B1 => n20580, B2 => n28779, A => n20941, ZN => 
                           n20582);
   U13335 : OAI21_X1 port map( B1 => n14146, B2 => n14008, A => n6050, ZN => 
                           n14148);
   U13336 : XNOR2_X1 port map( A => n13426, B => n13427, ZN => n6051);
   U13337 : NAND2_X1 port map( A1 => n20755, A2 => n21463, ZN => n6053);
   U13338 : INV_X1 port map( A => n23735, ZN => n22949);
   U13339 : NAND2_X1 port map( A1 => n23733, A2 => n23736, ZN => n6054);
   U13341 : NAND2_X1 port map( A1 => n24467, A2 => n29025, ZN => n24579);
   U13342 : INV_X1 port map( A => n20334, ZN => n6057);
   U13343 : NAND2_X1 port map( A1 => n6057, A2 => n1881, ZN => n20012);
   U13344 : INV_X1 port map( A => n9073, ZN => n9071);
   U13347 : OAI21_X1 port map( B1 => n6066, B2 => n14031, A => n6062, ZN => 
                           n6065);
   U13348 : NAND2_X1 port map( A1 => n6063, A2 => n29107, ZN => n6062);
   U13349 : INV_X1 port map( A => n13917, ZN => n6063);
   U13350 : NAND2_X1 port map( A1 => n6064, A2 => n13667, ZN => n13979);
   U13351 : MUX2_X1 port map( A => n6065, B => n13794, S => n13921, Z => n6064)
                           ;
   U13352 : INV_X1 port map( A => n13917, ZN => n6066);
   U13353 : OAI21_X1 port map( B1 => n26567, B2 => n29610, A => n6068, ZN => 
                           n26915);
   U13354 : INV_X1 port map( A => n26565, ZN => n6069);
   U13355 : NOR2_X1 port map( A1 => n1872, A2 => n26568, ZN => n6070);
   U13356 : INV_X1 port map( A => n9148, ZN => n6072);
   U13357 : NAND2_X1 port map( A1 => n578, A2 => n11867, ZN => n6075);
   U13358 : NAND2_X1 port map( A1 => n18470, A2 => n6079, ZN => n6078);
   U13359 : NAND3_X1 port map( A1 => n20206, A2 => n6083, A3 => n28501, ZN => 
                           n6082);
   U13360 : NAND2_X1 port map( A1 => n20552, A2 => n20404, ZN => n6083);
   U13362 : NAND2_X1 port map( A1 => n505, A2 => n20549, ZN => n20206);
   U13363 : OAI21_X1 port map( B1 => n28642, B2 => n26387, A => n28572, ZN => 
                           n6087);
   U13364 : XNOR2_X1 port map( A => n16505, B => n16506, ZN => n16507);
   U13365 : XNOR2_X1 port map( A => n15618, B => n15992, ZN => n16506);
   U13366 : NAND2_X1 port map( A1 => n14742, A2 => n544, ZN => n6088);
   U13367 : NAND3_X1 port map( A1 => n14745, A2 => n15117, A3 => n14744, ZN => 
                           n6089);
   U13368 : NAND2_X1 port map( A1 => n14741, A2 => n15115, ZN => n6090);
   U13369 : NAND2_X1 port map( A1 => n6973, A2 => n7358, ZN => n7357);
   U13370 : MUX2_X1 port map( A => n6973, B => n29110, S => n8231, Z => n8233);
   U13371 : MUX2_X1 port map( A => n7620, B => n29110, S => n6973, Z => n7623);
   U13372 : MUX2_X1 port map( A => n7431, B => n6974, S => n6973, Z => n6975);
   U13373 : INV_X1 port map( A => n11350, ZN => n11348);
   U13374 : XNOR2_X2 port map( A => n9130, B => n9129, ZN => n11350);
   U13375 : INV_X1 port map( A => n14484, ZN => n14170);
   U13377 : INV_X1 port map( A => n14483, ZN => n12122);
   U13380 : NAND2_X1 port map( A1 => n8795, A2 => n8794, ZN => n6092);
   U13381 : NAND2_X1 port map( A1 => n7689, A2 => n7688, ZN => n6093);
   U13382 : NAND2_X1 port map( A1 => n7686, A2 => n7687, ZN => n6094);
   U13383 : NAND2_X1 port map( A1 => n6095, A2 => n27528, ZN => n27096);
   U13384 : NOR2_X1 port map( A1 => n6095, A2 => n27531, ZN => n27508);
   U13387 : NAND2_X1 port map( A1 => n24489, A2 => n29051, ZN => n6098);
   U13388 : INV_X1 port map( A => n24100, ZN => n6097);
   U13389 : NOR2_X1 port map( A1 => n6099, A2 => n23706, ZN => n23707);
   U13390 : NOR2_X1 port map( A1 => n23220, A2 => n6099, ZN => n6582);
   U13391 : OAI21_X1 port map( B1 => n22451, B2 => n22452, A => n6099, ZN => 
                           n22454);
   U13393 : NAND2_X1 port map( A1 => n17625, A2 => n18411, ZN => n6103);
   U13394 : NAND2_X1 port map( A1 => n6104, A2 => n21702, ZN => n20994);
   U13399 : INV_X1 port map( A => n10919, ZN => n11138);
   U13401 : INV_X1 port map( A => n10415, ZN => n6107);
   U13402 : NAND2_X1 port map( A1 => n6111, A2 => n24078, ZN => n6109);
   U13403 : XNOR2_X1 port map( A => n6110, B => n12503, ZN => n25180);
   U13404 : NAND2_X1 port map( A1 => n29584, A2 => n6114, ZN => n19977);
   U13405 : OAI21_X1 port map( B1 => n20178, B2 => n20173, A => n6112, ZN => 
                           n19868);
   U13406 : NAND2_X1 port map( A1 => n6114, A2 => n20173, ZN => n6112);
   U13407 : INV_X1 port map( A => n504, ZN => n6113);
   U13408 : MUX2_X1 port map( A => n20177, B => n20171, S => n6114, Z => n6341)
                           ;
   U13410 : NAND2_X1 port map( A1 => n6117, A2 => n6116, ZN => n6115);
   U13411 : NAND2_X1 port map( A1 => n21289, A2 => n21288, ZN => n6118);
   U13412 : XNOR2_X1 port map( A => n22845, B => n21872, ZN => n22599);
   U13413 : XNOR2_X1 port map( A => n22845, B => n6119, ZN => n21786);
   U13414 : XNOR2_X1 port map( A => n25807, B => n24890, ZN => n6122);
   U13415 : NAND2_X1 port map( A1 => n23936, A2 => n24556, ZN => n6120);
   U13416 : NAND2_X1 port map( A1 => n6123, A2 => n6097, ZN => n23944);
   U13420 : OR2_X1 port map( A1 => n17304, A2 => n28768, ZN => n6128);
   U13422 : OAI211_X2 port map( C1 => n6132, C2 => n11507, A => n12283, B => 
                           n11506, ZN => n13150);
   U13423 : XNOR2_X1 port map( A => n9601, B => n10231, ZN => n9985);
   U13424 : XNOR2_X1 port map( A => n6134, B => n6136, ZN => n6133);
   U13425 : INV_X1 port map( A => n9985, ZN => n6134);
   U13426 : NAND2_X1 port map( A1 => n6140, A2 => n6139, ZN => n17856);
   U13427 : OR2_X1 port map( A1 => n6927, A2 => n17989, ZN => n6139);
   U13428 : NAND2_X1 port map( A1 => n17990, A2 => n6927, ZN => n6140);
   U13429 : XNOR2_X1 port map( A => n22919, B => n6141, ZN => n22838);
   U13430 : XNOR2_X1 port map( A => n6141, B => n22441, ZN => n22443);
   U13432 : NAND2_X1 port map( A1 => n13948, A2 => n14170, ZN => n6142);
   U13433 : NAND2_X1 port map( A1 => n10114, A2 => n11120, ZN => n6144);
   U13434 : NAND2_X1 port map( A1 => n11477, A2 => n11998, ZN => n6145);
   U13435 : NAND2_X1 port map( A1 => n12000, A2 => n11755, ZN => n11540);
   U13436 : INV_X1 port map( A => n8908, ZN => n6147);
   U13437 : INV_X1 port map( A => n27300, ZN => n6150);
   U13438 : NAND2_X1 port map( A1 => n6948, A2 => n26935, ZN => n6148);
   U13439 : NAND2_X1 port map( A1 => n26558, A2 => n26940, ZN => n6149);
   U13440 : MUX2_X1 port map( A => n24760, B => n24215, S => n24756, Z => 
                           n24216);
   U13443 : NAND2_X1 port map( A1 => n20500, A2 => n29601, ZN => n6156);
   U13444 : INV_X1 port map( A => n22139, ZN => n21624);
   U13445 : XNOR2_X1 port map( A => n16198, B => n16197, ZN => n6160);
   U13446 : MUX2_X1 port map( A => n16706, B => n16884, S => n17526, Z => 
                           n16885);
   U13447 : INV_X1 port map( A => n6162, ZN => n7861);
   U13448 : NAND2_X1 port map( A1 => n7308, A2 => n7172, ZN => n6162);
   U13449 : NAND2_X1 port map( A1 => n587, A2 => n29517, ZN => n6164);
   U13450 : INV_X1 port map( A => n18856, ZN => n18922);
   U13451 : OAI21_X1 port map( B1 => n14334, B2 => n14410, A => n14333, ZN => 
                           n14335);
   U13452 : NAND2_X1 port map( A1 => n6166, A2 => n29607, ZN => n14333);
   U13454 : INV_X1 port map( A => n14408, ZN => n6166);
   U13455 : OR2_X1 port map( A1 => n24430, A2 => n19041, ZN => n6171);
   U13456 : XNOR2_X1 port map( A => n25145, B => n6167, ZN => n25148);
   U13457 : XNOR2_X1 port map( A => n6168, B => n365, ZN => n6167);
   U13458 : OAI211_X1 port map( C1 => n6171, C2 => n24429, A => n6169, B => 
                           n6170, ZN => n6168);
   U13459 : NAND2_X1 port map( A1 => n24429, A2 => n19041, ZN => n6169);
   U13460 : NAND2_X1 port map( A1 => n24430, A2 => n19041, ZN => n6170);
   U13461 : NOR2_X2 port map( A1 => n24429, A2 => n24430, ZN => n25867);
   U13462 : XNOR2_X1 port map( A => n15575, B => n26656, ZN => n15763);
   U13463 : INV_X1 port map( A => n16579, ZN => n6173);
   U13464 : XNOR2_X1 port map( A => n15575, B => n6173, ZN => n15658);
   U13465 : XNOR2_X1 port map( A => n15575, B => n6174, ZN => n15904);
   U13467 : NAND2_X1 port map( A1 => n17547, A2 => n16947, ZN => n6175);
   U13468 : NAND2_X1 port map( A1 => n18529, A2 => n17864, ZN => n6177);
   U13469 : AND2_X2 port map( A1 => n6179, A2 => n6178, ZN => n17864);
   U13470 : NAND2_X1 port map( A1 => n16933, A2 => n17046, ZN => n6178);
   U13471 : NAND2_X1 port map( A1 => n16934, A2 => n6180, ZN => n6179);
   U13472 : INV_X1 port map( A => n11458, ZN => n6181);
   U13473 : INV_X1 port map( A => n11457, ZN => n11460);
   U13474 : INV_X1 port map( A => n11152, ZN => n6182);
   U13475 : NAND2_X1 port map( A1 => n6182, A2 => n11158, ZN => n10494);
   U13476 : OAI21_X2 port map( B1 => n27171, B2 => n6185, A => n27170, ZN => 
                           n27672);
   U13477 : NAND2_X1 port map( A1 => n6567, A2 => n20618, ZN => n19921);
   U13478 : INV_X1 port map( A => n9030, ZN => n8433);
   U13479 : NOR2_X1 port map( A1 => n28210, A2 => n9030, ZN => n6188);
   U13480 : NAND3_X1 port map( A1 => n9027, A2 => n9030, A3 => n7714, ZN => 
                           n6191);
   U13481 : INV_X1 port map( A => n6193, ZN => n19338);
   U13482 : XNOR2_X1 port map( A => n19220, B => n19111, ZN => n6193);
   U13483 : NOR2_X1 port map( A1 => n6294, A2 => n28122, ZN => n6196);
   U13484 : INV_X1 port map( A => n23139, ZN => n6194);
   U13485 : NAND2_X1 port map( A1 => n23427, A2 => n23138, ZN => n23139);
   U13487 : INV_X1 port map( A => n6200, ZN => n6199);
   U13488 : OAI22_X1 port map( A1 => n7241, A2 => n7995, B1 => n7993, B2 => 
                           n6201, ZN => n6200);
   U13489 : OR2_X1 port map( A1 => n7992, A2 => n7876, ZN => n6201);
   U13490 : MUX2_X1 port map( A => n27300, B => n5425, S => n27301, Z => n26689
                           );
   U13492 : NAND2_X1 port map( A1 => n6203, A2 => n28417, ZN => n6202);
   U13493 : INV_X1 port map( A => n19928, ZN => n6203);
   U13494 : NAND2_X1 port map( A1 => n20451, A2 => n20449, ZN => n6204);
   U13495 : AND2_X1 port map( A1 => n28417, A2 => n20265, ZN => n6205);
   U13496 : MUX2_X1 port map( A => n20449, B => n28552, S => n28417, Z => 
                           n20452);
   U13497 : INV_X1 port map( A => n21749, ZN => n21643);
   U13498 : NAND2_X1 port map( A1 => n20659, A2 => n21748, ZN => n6206);
   U13499 : XOR2_X1 port map( A => n16090, B => n16233, Z => n15366);
   U13500 : NAND2_X1 port map( A1 => n7231, A2 => n7591, ZN => n7318);
   U13501 : NAND2_X1 port map( A1 => n6210, A2 => n29629, ZN => n7727);
   U13502 : NAND2_X1 port map( A1 => n6211, A2 => n22944, ZN => n22593);
   U13503 : NAND2_X1 port map( A1 => n28181, A2 => n23738, ZN => n6211);
   U13504 : INV_X1 port map( A => n21738, ZN => n6212);
   U13505 : NAND3_X1 port map( A1 => n1814, A2 => n20841, A3 => n21458, ZN => 
                           n6213);
   U13506 : XNOR2_X1 port map( A => n24852, B => n2306, ZN => n24453);
   U13508 : NAND2_X1 port map( A1 => n28552, A2 => n21063, ZN => n6219);
   U13509 : AOI21_X1 port map( B1 => n9686, B2 => n1933, A => n29637, ZN => 
                           n10485);
   U13510 : AOI22_X1 port map( A1 => n10486, A2 => n29637, B1 => n10487, B2 => 
                           n1933, ZN => n10488);
   U13511 : OAI21_X1 port map( B1 => n9248, B2 => n9245, A => n28211, ZN => 
                           n7161);
   U13512 : XNOR2_X1 port map( A => n16588, B => n1980, ZN => n15280);
   U13514 : AOI211_X1 port map( C1 => n28482, C2 => n377, A => n6222, B => 
                           n26461, ZN => n6221);
   U13515 : AND2_X1 port map( A1 => n28476, A2 => n26559, ZN => n6222);
   U13517 : NAND2_X1 port map( A1 => n6225, A2 => n18354, ZN => n17919);
   U13518 : NAND2_X1 port map( A1 => n17666, A2 => n6225, ZN => n17668);
   U13519 : INV_X1 port map( A => n13458, ZN => n13460);
   U13520 : NAND3_X1 port map( A1 => n2012, A2 => n11592, A3 => n12581, ZN => 
                           n13458);
   U13521 : NAND4_X1 port map( A1 => n1864, A2 => n6226, A3 => n27302, A4 => 
                           n27301, ZN => n27307);
   U13522 : XNOR2_X1 port map( A => n20735, B => n20734, ZN => n6227);
   U13523 : XNOR2_X1 port map( A => n19717, B => n19668, ZN => n19399);
   U13525 : NAND2_X1 port map( A1 => n13728, A2 => n14135, ZN => n6233);
   U13526 : NAND2_X1 port map( A1 => n20381, A2 => n28637, ZN => n6236);
   U13527 : NAND2_X1 port map( A1 => n20779, A2 => n20778, ZN => n6240);
   U13528 : OAI211_X1 port map( C1 => n10549, C2 => n10492, A => n11115, B => 
                           n6241, ZN => n6242);
   U13529 : NOR2_X1 port map( A1 => n17854, A2 => n6526, ZN => n17988);
   U13530 : NAND2_X1 port map( A1 => n17988, A2 => n18367, ZN => n6243);
   U13531 : XNOR2_X1 port map( A => n16291, B => n14709, ZN => n16270);
   U13532 : NAND2_X1 port map( A1 => n14704, A2 => n6244, ZN => n16291);
   U13533 : NAND3_X1 port map( A1 => n6245, A2 => n6246, A3 => n15268, ZN => 
                           n6244);
   U13534 : NAND2_X1 port map( A1 => n6250, A2 => n6249, ZN => n6248);
   U13535 : NAND2_X1 port map( A1 => n242, A2 => n10549, ZN => n6249);
   U13536 : NAND2_X1 port map( A1 => n6253, A2 => n13724, ZN => n6252);
   U13537 : NAND2_X1 port map( A1 => n14148, A2 => n14374, ZN => n6253);
   U13540 : XNOR2_X1 port map( A => n10018, B => n10016, ZN => n6257);
   U13541 : NAND2_X1 port map( A1 => n11136, A2 => n11142, ZN => n11139);
   U13542 : INV_X1 port map( A => n11139, ZN => n10463);
   U13544 : NAND2_X1 port map( A1 => n20190, A2 => n20547, ZN => n6259);
   U13549 : INV_X1 port map( A => n24408, ZN => n6265);
   U13550 : INV_X1 port map( A => n24404, ZN => n6266);
   U13551 : OAI21_X1 port map( B1 => n27539, B2 => n27548, A => n27538, ZN => 
                           n6268);
   U13552 : XNOR2_X1 port map( A => n6647, B => n13208, ZN => n13542);
   U13553 : NAND2_X1 port map( A1 => n10749, A2 => n11198, ZN => n6271);
   U13554 : NAND2_X1 port map( A1 => n21658, A2 => n21657, ZN => n6273);
   U13555 : NAND2_X1 port map( A1 => n21659, A2 => n6275, ZN => n6274);
   U13556 : INV_X1 port map( A => n6276, ZN => n19144);
   U13557 : XNOR2_X1 port map( A => n19145, B => n6276, ZN => n6606);
   U13558 : INV_X1 port map( A => n18948, ZN => n19199);
   U13559 : NOR2_X1 port map( A1 => n23393, A2 => n23392, ZN => n6277);
   U13560 : AOI21_X1 port map( B1 => n23838, B2 => n6610, A => n6279, ZN => 
                           n6278);
   U13561 : INV_X1 port map( A => n23391, ZN => n6279);
   U13562 : NAND2_X1 port map( A1 => n7662, A2 => n8265, ZN => n9084);
   U13563 : OR2_X2 port map( A1 => n12846, A2 => n6283, ZN => n14575);
   U13564 : NAND2_X1 port map( A1 => n18540, A2 => n18539, ZN => n6284);
   U13565 : NAND2_X1 port map( A1 => n18541, A2 => n18529, ZN => n6285);
   U13566 : NAND2_X1 port map( A1 => n7233, A2 => n7231, ZN => n7594);
   U13568 : INV_X1 port map( A => n28549, ZN => n27353);
   U13569 : INV_X1 port map( A => n11176, ZN => n11334);
   U13570 : NOR2_X1 port map( A1 => n6292, A2 => n6290, ZN => n16755);
   U13571 : NOR2_X1 port map( A1 => n17229, A2 => n6291, ZN => n6290);
   U13572 : NAND2_X1 port map( A1 => n17567, A2 => n17568, ZN => n6291);
   U13573 : NAND2_X1 port map( A1 => n15279, A2 => n6293, ZN => n6493);
   U13574 : XNOR2_X1 port map( A => n15545, B => n6296, ZN => n15836);
   U13575 : INV_X1 port map( A => n13456, ZN => n6297);
   U13576 : AOI21_X1 port map( B1 => n6299, B2 => n8024, A => n29130, ZN => 
                           n8025);
   U13578 : NAND2_X1 port map( A1 => n26860, A2 => n29633, ZN => n6300);
   U13579 : NAND3_X1 port map( A1 => n26855, A2 => n27142, A3 => n28487, ZN => 
                           n6301);
   U13580 : NAND2_X1 port map( A1 => n26325, A2 => n27139, ZN => n6302);
   U13581 : INV_X1 port map( A => n27141, ZN => n27139);
   U13585 : OAI21_X1 port map( B1 => n24288, B2 => n24597, A => n24148, ZN => 
                           n23933);
   U13586 : XNOR2_X1 port map( A => n22248, B => n2350, ZN => n21902);
   U13587 : OAI21_X2 port map( B1 => n6321, B2 => n6835, A => n23954, ZN => 
                           n25773);
   U13588 : NAND3_X1 port map( A1 => n6325, A2 => n16711, A3 => n6324, ZN => 
                           n16718);
   U13589 : NAND2_X1 port map( A1 => n16709, A2 => n17335, ZN => n6324);
   U13590 : NAND2_X1 port map( A1 => n16710, A2 => n17342, ZN => n6325);
   U13591 : INV_X1 port map( A => n19534, ZN => n6327);
   U13592 : XNOR2_X1 port map( A => n6327, B => n19220, ZN => n18984);
   U13593 : NAND2_X1 port map( A1 => n12240, A2 => n11969, ZN => n12242);
   U13594 : NAND2_X1 port map( A1 => n12156, A2 => n12158, ZN => n12240);
   U13595 : NAND2_X1 port map( A1 => n10453, A2 => n11876, ZN => n10869);
   U13596 : NAND2_X1 port map( A1 => n11879, A2 => n567, ZN => n6329);
   U13597 : NAND3_X1 port map( A1 => n1926, A2 => n15013, A3 => n15014, ZN => 
                           n6332);
   U13600 : NAND2_X1 port map( A1 => n6338, A2 => n23830, ZN => n6579);
   U13602 : INV_X1 port map( A => n20053, ZN => n20172);
   U13603 : XNOR2_X1 port map( A => n13350, B => n12822, ZN => n6343);
   U13604 : NAND2_X1 port map( A1 => n6348, A2 => n23842, ZN => n24492);
   U13605 : NAND2_X1 port map( A1 => n6348, A2 => n24471, ZN => n23850);
   U13606 : NOR2_X1 port map( A1 => n29033, A2 => n6348, ZN => n24473);
   U13607 : NAND3_X1 port map( A1 => n24100, A2 => n29033, A3 => n6348, ZN => 
                           n24101);
   U13608 : AOI21_X1 port map( B1 => n24490, B2 => n24489, A => n6348, ZN => 
                           n24495);
   U13609 : OAI211_X1 port map( C1 => n21442, C2 => n6275, A => n21441, B => 
                           n21440, ZN => n6350);
   U13610 : NAND2_X1 port map( A1 => n13729, A2 => n13912, ZN => n14070);
   U13611 : NAND3_X1 port map( A1 => n6462, A2 => n6354, A3 => n6353, ZN => 
                           n6356);
   U13612 : NAND2_X1 port map( A1 => n28554, A2 => n23765, ZN => n6353);
   U13613 : NAND2_X1 port map( A1 => n23764, A2 => n23763, ZN => n6354);
   U13614 : NAND3_X1 port map( A1 => n6356, A2 => n6357, A3 => n6355, ZN => 
                           n24502);
   U13615 : NAND2_X1 port map( A1 => n23766, A2 => n6358, ZN => n6357);
   U13616 : NAND2_X1 port map( A1 => n7813, A2 => n10806, ZN => n6359);
   U13617 : NAND2_X1 port map( A1 => n10512, A2 => n10544, ZN => n6361);
   U13618 : INV_X1 port map( A => n21304, ZN => n6362);
   U13619 : INV_X1 port map( A => n22301, ZN => n22757);
   U13620 : NAND2_X1 port map( A1 => n6363, A2 => n20327, ZN => n22301);
   U13621 : NAND2_X1 port map( A1 => n8825, A2 => n29147, ZN => n8584);
   U13622 : NAND3_X1 port map( A1 => n8825, A2 => n8586, A3 => n8824, ZN => 
                           n8834);
   U13623 : NAND2_X1 port map( A1 => n6365, A2 => n6086, ZN => n19856);
   U13624 : NAND2_X1 port map( A1 => n20206, A2 => n20404, ZN => n6365);
   U13625 : NAND2_X1 port map( A1 => n10972, A2 => n10976, ZN => n6367);
   U13626 : NAND3_X1 port map( A1 => n21484, A2 => n21581, A3 => n21481, ZN => 
                           n6369);
   U13627 : NAND2_X1 port map( A1 => n6371, A2 => n16814, ZN => n16817);
   U13628 : OR2_X1 port map( A1 => n17097, A2 => n16815, ZN => n17104);
   U13629 : NAND3_X1 port map( A1 => n6371, A2 => n1466, A3 => n16860, ZN => 
                           n16680);
   U13630 : INV_X1 port map( A => n17097, ZN => n6371);
   U13631 : NAND2_X1 port map( A1 => n12510, A2 => n6372, ZN => n11993);
   U13633 : INV_X1 port map( A => n6375, ZN => n12685);
   U13634 : XNOR2_X1 port map( A => n6375, B => n12389, ZN => n12393);
   U13635 : NAND2_X1 port map( A1 => n18341, A2 => n18342, ZN => n6376);
   U13636 : NAND2_X1 port map( A1 => n24727, A2 => n29695, ZN => n6377);
   U13637 : NAND2_X1 port map( A1 => n24596, A2 => n24288, ZN => n24724);
   U13638 : XNOR2_X1 port map( A => n22691, B => n22437, ZN => n21739);
   U13639 : NAND2_X1 port map( A1 => n7234, A2 => n7591, ZN => n6381);
   U13640 : NOR2_X1 port map( A1 => n11048, A2 => n11266, ZN => n6385);
   U13641 : INV_X1 port map( A => n29122, ZN => n11044);
   U13642 : NAND3_X1 port map( A1 => n17906, A2 => n17947, A3 => n18341, ZN => 
                           n6387);
   U13643 : XNOR2_X1 port map( A => n22246, B => n22265, ZN => n6388);
   U13644 : NAND2_X1 port map( A1 => n6392, A2 => n6390, ZN => n16388);
   U13645 : NAND2_X1 port map( A1 => n15263, A2 => n6391, ZN => n6390);
   U13646 : OAI21_X1 port map( B1 => n6393, B2 => n14761, A => n15264, ZN => 
                           n6392);
   U13648 : NAND2_X1 port map( A1 => n21270, A2 => n21271, ZN => n6394);
   U13650 : NAND2_X1 port map( A1 => n20815, A2 => n21269, ZN => n21272);
   U13651 : NAND2_X1 port map( A1 => n6398, A2 => n29488, ZN => n6397);
   U13652 : NAND2_X1 port map( A1 => n21267, A2 => n21268, ZN => n6398);
   U13653 : NAND2_X1 port map( A1 => n16930, A2 => n6403, ZN => n6402);
   U13654 : NAND3_X1 port map( A1 => n8610, A2 => n8749, A3 => n9533, ZN => 
                           n6404);
   U13655 : NAND2_X1 port map( A1 => n6413, A2 => n694, ZN => n6412);
   U13656 : NAND2_X1 port map( A1 => n14781, A2 => n15338, ZN => n6413);
   U13657 : XNOR2_X1 port map( A => n21791, B => n21792, ZN => n6414);
   U13658 : XNOR2_X2 port map( A => n6414, B => n21795, ZN => n23764);
   U13659 : XNOR2_X1 port map( A => n16518, B => n15941, ZN => n6415);
   U13660 : XNOR2_X1 port map( A => n15942, B => n5858, ZN => n6416);
   U13661 : AOI21_X1 port map( B1 => n17037, B2 => n6417, A => n17569, ZN => 
                           n17042);
   U13662 : OAI21_X1 port map( B1 => n4784, B2 => n24466, A => n6421, ZN => 
                           n6420);
   U13665 : NAND2_X1 port map( A1 => n12481, A2 => n14215, ZN => n14214);
   U13666 : NAND2_X1 port map( A1 => n555, A2 => n12481, ZN => n12470);
   U13670 : NAND3_X1 port map( A1 => n6432, A2 => n12332, A3 => n12327, ZN => 
                           n10537);
   U13671 : NAND2_X1 port map( A1 => n12018, A2 => n6432, ZN => n12334);
   U13672 : NAND2_X1 port map( A1 => n12016, A2 => n6432, ZN => n10536);
   U13673 : NAND2_X1 port map( A1 => n12015, A2 => n6432, ZN => n11890);
   U13674 : NAND3_X1 port map( A1 => n11449, A2 => n12332, A3 => n6432, ZN => 
                           n6431);
   U13675 : NAND3_X1 port map( A1 => n4118, A2 => n17569, A3 => n17227, ZN => 
                           n16756);
   U13677 : NAND2_X1 port map( A1 => n14313, A2 => n14314, ZN => n6434);
   U13679 : XNOR2_X1 port map( A => n25061, B => n25060, ZN => n6436);
   U13680 : NAND2_X1 port map( A1 => n26918, A2 => n457, ZN => n6438);
   U13681 : XNOR2_X1 port map( A => n10146, B => n9934, ZN => n6440);
   U13683 : XNOR2_X1 port map( A => n16076, B => n6448, ZN => n6447);
   U13684 : XNOR2_X1 port map( A => n6449, B => n29319, ZN => n6448);
   U13685 : NAND2_X1 port map( A1 => n8871, A2 => n7568, ZN => n6450);
   U13686 : NAND2_X1 port map( A1 => n9059, A2 => n9064, ZN => n8868);
   U13687 : INV_X1 port map( A => n16323, ZN => n6454);
   U13688 : INV_X1 port map( A => n16323, ZN => n16455);
   U13689 : OR2_X1 port map( A1 => n15318, A2 => n15319, ZN => n6457);
   U13690 : XNOR2_X1 port map( A => n6458, B => n1928, ZN => n20837);
   U13691 : XNOR2_X1 port map( A => n6458, B => n3369, ZN => n22368);
   U13692 : XNOR2_X1 port map( A => n21805, B => n6458, ZN => n21816);
   U13693 : XNOR2_X1 port map( A => n22180, B => n6458, ZN => n22902);
   U13694 : XNOR2_X1 port map( A => n22609, B => n6458, ZN => n22612);
   U13697 : NAND2_X1 port map( A1 => n21829, A2 => n6462, ZN => n6461);
   U13698 : XNOR2_X2 port map( A => n8991, B => n8990, ZN => n11322);
   U13701 : OAI21_X1 port map( B1 => n27592, B2 => n26285, A => n27597, ZN => 
                           n6464);
   U13702 : INV_X1 port map( A => n17272, ZN => n6465);
   U13703 : INV_X1 port map( A => n14416, ZN => n6466);
   U13705 : NAND2_X1 port map( A1 => n14420, A2 => n14421, ZN => n14448);
   U13706 : OR2_X1 port map( A1 => n14416, A2 => n14414, ZN => n14421);
   U13707 : XNOR2_X1 port map( A => n19290, B => n6468, ZN => n6467);
   U13711 : NAND2_X1 port map( A1 => n885, A2 => n29564, ZN => n6474);
   U13714 : NAND2_X1 port map( A1 => n6480, A2 => n6479, ZN => n6478);
   U13715 : NOR2_X1 port map( A1 => n16539, A2 => n28801, ZN => n6485);
   U13716 : NAND2_X1 port map( A1 => n17899, A2 => n6484, ZN => n6483);
   U13717 : INV_X1 port map( A => n18356, ZN => n6484);
   U13720 : XNOR2_X1 port map( A => n6487, B => n19276, ZN => n20597);
   U13721 : INV_X2 port map( A => n6488, ZN => n19487);
   U13722 : XNOR2_X1 port map( A => n19313, B => n19487, ZN => n18210);
   U13723 : NAND3_X1 port map( A1 => n27772, A2 => n29537, A3 => n29022, ZN => 
                           n27774);
   U13724 : OAI22_X1 port map( A1 => n27233, A2 => n6490, B1 => n27762, B2 => 
                           n29022, ZN => n27234);
   U13725 : OR2_X1 port map( A1 => n26289, A2 => n29633, ZN => n6492);
   U13727 : INV_X1 port map( A => n20081, ZN => n6495);
   U13728 : NAND2_X1 port map( A1 => n19846, A2 => n29145, ZN => n6494);
   U13730 : XNOR2_X1 port map( A => n6496, B => n15576, ZN => Ciphertext(123));
   U13731 : NAND3_X1 port map( A1 => n6498, A2 => n27770, A3 => n6497, ZN => 
                           n6496);
   U13732 : NAND2_X1 port map( A1 => n29117, A2 => n27769, ZN => n6497);
   U13733 : XNOR2_X1 port map( A => n16379, B => n16378, ZN => n6502);
   U13734 : NAND3_X1 port map( A1 => n21493, A2 => n21185, A3 => n21496, ZN => 
                           n6503);
   U13735 : NAND2_X1 port map( A1 => n9042, A2 => n9247, ZN => n6505);
   U13736 : NAND2_X1 port map( A1 => n24417, A2 => n24341, ZN => n6506);
   U13737 : INV_X1 port map( A => n25998, ZN => n6507);
   U13738 : NAND2_X1 port map( A1 => n19858, A2 => n20412, ZN => n6509);
   U13739 : OAI21_X1 port map( B1 => n11188, B2 => n11322, A => n6510, ZN => 
                           n10813);
   U13741 : INV_X1 port map( A => n15274, ZN => n14698);
   U13742 : NAND2_X1 port map( A1 => n20481, A2 => n20485, ZN => n6512);
   U13743 : NAND2_X1 port map( A1 => n10669, A2 => n10670, ZN => n6516);
   U13744 : XNOR2_X1 port map( A => n13482, B => n13273, ZN => n12944);
   U13745 : NAND3_X1 port map( A1 => n11680, A2 => n5009, A3 => n11541, ZN => 
                           n6518);
   U13746 : XNOR2_X1 port map( A => n6520, B => n29549, ZN => n21884);
   U13747 : XNOR2_X1 port map( A => n6520, B => n22110, ZN => n22111);
   U13749 : NAND2_X1 port map( A1 => n6522, A2 => n6521, ZN => n15449);
   U13750 : OAI21_X1 port map( B1 => n15327, B2 => n15322, A => n6522, ZN => 
                           n13978);
   U13751 : NAND2_X1 port map( A1 => n15327, A2 => n15323, ZN => n6522);
   U13752 : AND2_X1 port map( A1 => n23290, A2 => n23816, ZN => n23821);
   U13754 : INV_X1 port map( A => n12775, ZN => n12476);
   U13755 : NAND2_X1 port map( A1 => n17000, A2 => n17402, ZN => n6524);
   U13757 : XNOR2_X1 port map( A => n22271, B => n22248, ZN => n22728);
   U13758 : XNOR2_X1 port map( A => n22728, B => n22727, ZN => n22729);
   U13759 : XNOR2_X1 port map( A => n19631, B => n19632, ZN => n6535);
   U13760 : XNOR2_X1 port map( A => n19634, B => n19635, ZN => n6536);
   U13761 : NAND3_X1 port map( A1 => n24712, A2 => n28524, A3 => n24713, ZN => 
                           n24352);
   U13762 : NAND2_X1 port map( A1 => n23055, A2 => n23054, ZN => n6537);
   U13763 : MUX2_X1 port map( A => n29573, B => n26799, S => n26278, Z => n6541
                           );
   U13765 : OAI22_X1 port map( A1 => n6542, A2 => n10593, B1 => n10705, B2 => 
                           n10944, ZN => n10596);
   U13767 : NAND2_X1 port map( A1 => n9581, A2 => n9580, ZN => n9579);
   U13768 : OAI211_X2 port map( C1 => n7314, C2 => n7900, A => n6546, B => 
                           n6545, ZN => n7569);
   U13769 : NAND3_X1 port map( A1 => n7804, A2 => n7800, A3 => n7898, ZN => 
                           n6546);
   U13770 : NAND2_X1 port map( A1 => n24423, A2 => n24422, ZN => n6548);
   U13771 : INV_X1 port map( A => n12359, ZN => n12361);
   U13772 : NAND2_X1 port map( A1 => n11739, A2 => n11740, ZN => n12360);
   U13773 : NAND3_X1 port map( A1 => n11742, A2 => n11740, A3 => n12359, ZN => 
                           n6549);
   U13774 : NAND3_X1 port map( A1 => n12363, A2 => n12362, A3 => n12361, ZN => 
                           n6550);
   U13775 : NAND2_X1 port map( A1 => n12357, A2 => n12356, ZN => n6552);
   U13776 : NAND2_X1 port map( A1 => n17544, A2 => n17543, ZN => n6553);
   U13777 : NAND2_X1 port map( A1 => n6555, A2 => n17217, ZN => n6554);
   U13778 : MUX2_X1 port map( A => n17540, B => n17539, S => n17545, Z => n6555
                           );
   U13779 : NAND2_X1 port map( A1 => n16939, A2 => n28454, ZN => n17546);
   U13782 : NAND2_X1 port map( A1 => n24547, A2 => n6556, ZN => n6868);
   U13783 : NOR2_X1 port map( A1 => n24547, A2 => n6556, ZN => n23129);
   U13784 : AOI21_X1 port map( B1 => n24543, B2 => n24544, A => n6556, ZN => 
                           n24545);
   U13785 : NAND2_X1 port map( A1 => n22965, A2 => n29020, ZN => n6558);
   U13786 : NOR2_X1 port map( A1 => n6559, A2 => n16723, ZN => n16726);
   U13787 : NAND2_X1 port map( A1 => n17476, A2 => n6560, ZN => n16801);
   U13788 : OR2_X1 port map( A1 => n14107, A2 => n6563, ZN => n6562);
   U13790 : INV_X1 port map( A => n20617, ZN => n20432);
   U13791 : NOR2_X2 port map( A1 => n20434, A2 => n6564, ZN => n21514);
   U13792 : OAI21_X1 port map( B1 => n20617, B2 => n6567, A => n6566, ZN => 
                           n6565);
   U13793 : NAND2_X1 port map( A1 => n6567, A2 => n20619, ZN => n6566);
   U13794 : INV_X1 port map( A => n20431, ZN => n6567);
   U13795 : NOR2_X1 port map( A1 => n20635, A2 => n20248, ZN => n20032);
   U13797 : NAND2_X1 port map( A1 => n13943, A2 => n15194, ZN => n14175);
   U13798 : NAND2_X1 port map( A1 => n6571, A2 => n13943, ZN => n6572);
   U13799 : INV_X1 port map( A => n15415, ZN => n15410);
   U13800 : XNOR2_X1 port map( A => n18802, B => n19643, ZN => n19039);
   U13801 : NAND2_X1 port map( A1 => n18479, A2 => n18011, ZN => n6574);
   U13802 : NAND2_X1 port map( A1 => n6576, A2 => n18475, ZN => n6575);
   U13803 : INV_X1 port map( A => n20219, ZN => n19992);
   U13804 : INV_X1 port map( A => n18972, ZN => n6578);
   U13806 : NOR2_X1 port map( A1 => n28551, A2 => n23281, ZN => n6580);
   U13807 : NAND3_X1 port map( A1 => n27433, A2 => n25417, A3 => n26830, ZN => 
                           n25424);
   U13808 : NAND2_X1 port map( A1 => n28622, A2 => n6582, ZN => n6584);
   U13809 : NAND2_X1 port map( A1 => n22084, A2 => n23700, ZN => n6587);
   U13811 : NAND2_X1 port map( A1 => n22085, A2 => n6587, ZN => n6586);
   U13812 : NAND2_X1 port map( A1 => n17717, A2 => n17720, ZN => n6588);
   U13813 : NAND3_X1 port map( A1 => n9235, A2 => n9047, A3 => n6590, ZN => 
                           n9048);
   U13814 : XNOR2_X1 port map( A => n6591, B => n3654, ZN => Ciphertext(81));
   U13815 : NAND2_X1 port map( A1 => n6594, A2 => n6593, ZN => n6592);
   U13816 : NAND2_X1 port map( A1 => n27554, A2 => n29085, ZN => n6593);
   U13817 : NAND2_X1 port map( A1 => n27149, A2 => n29578, ZN => n6594);
   U13818 : NAND2_X1 port map( A1 => n24503, A2 => n6596, ZN => n6595);
   U13820 : OAI21_X1 port map( B1 => n10572, B2 => n10883, A => n6603, ZN => 
                           n10655);
   U13821 : NAND2_X1 port map( A1 => n11212, A2 => n10883, ZN => n6603);
   U13822 : AND2_X1 port map( A1 => n6605, A2 => n20504, ZN => n19799);
   U13823 : XNOR2_X2 port map( A => n19148, B => n6606, ZN => n20504);
   U13824 : INV_X1 port map( A => n20339, ZN => n6605);
   U13825 : NAND2_X1 port map( A1 => n23791, A2 => n23789, ZN => n6607);
   U13826 : INV_X1 port map( A => n23280, ZN => n6610);
   U13827 : INV_X1 port map( A => n24707, ZN => n24124);
   U13828 : NOR2_X1 port map( A1 => n24704, A2 => n24707, ZN => n6612);
   U13829 : INV_X1 port map( A => n7997, ZN => n7998);
   U13830 : OAI211_X1 port map( C1 => n6623, C2 => n6622, A => n6616, B => 
                           n6618, ZN => Ciphertext(9));
   U13831 : INV_X1 port map( A => n27367, ZN => n6617);
   U13832 : INV_X1 port map( A => n6619, ZN => n6618);
   U13833 : OAI21_X1 port map( B1 => n3751, B2 => n27375, A => n6620, ZN => 
                           n6619);
   U13834 : NAND3_X1 port map( A1 => n27375, A2 => n27374, A3 => n3751, ZN => 
                           n6622);
   U13835 : AOI21_X1 port map( B1 => n27369, B2 => n6624, A => n27364, ZN => 
                           n6623);
   U13836 : OR2_X1 port map( A1 => n27370, A2 => n29541, ZN => n6624);
   U13837 : NAND2_X1 port map( A1 => n26237, A2 => n26757, ZN => n26760);
   U13838 : NAND2_X1 port map( A1 => n6625, A2 => n26237, ZN => n6626);
   U13839 : NAND2_X1 port map( A1 => n26756, A2 => n26241, ZN => n6627);
   U13841 : OAI21_X1 port map( B1 => n23458, B2 => n23461, A => n23357, ZN => 
                           n6628);
   U13842 : INV_X1 port map( A => n23148, ZN => n23455);
   U13843 : NAND2_X1 port map( A1 => n11266, A2 => n29122, ZN => n6631);
   U13845 : NAND2_X1 port map( A1 => n25079, A2 => n26422, ZN => n6634);
   U13846 : INV_X1 port map( A => n21565, ZN => n6636);
   U13847 : XNOR2_X1 port map( A => n15635, B => n6637, ZN => n15638);
   U13848 : INV_X1 port map( A => n6637, ZN => n16266);
   U13849 : NAND2_X1 port map( A1 => n17273, A2 => n539, ZN => n6638);
   U13850 : NAND2_X1 port map( A1 => n13916, A2 => n6066, ZN => n6639);
   U13851 : XNOR2_X1 port map( A => n6644, B => n9787, ZN => n9792);
   U13852 : NAND2_X1 port map( A1 => n11361, A2 => n15576, ZN => n6646);
   U13853 : XNOR2_X1 port map( A => n13061, B => n6647, ZN => n12349);
   U13854 : XNOR2_X1 port map( A => n12746, B => n6647, ZN => n11368);
   U13855 : XNOR2_X1 port map( A => n15779, B => n16617, ZN => n6650);
   U13856 : NAND2_X1 port map( A1 => n15402, A2 => n13639, ZN => n13602);
   U13857 : NAND2_X1 port map( A1 => n13579, A2 => n13580, ZN => n13639);
   U13858 : XNOR2_X1 port map( A => n13481, B => n6652, ZN => n6651);
   U13859 : NAND2_X1 port map( A1 => n17848, A2 => n17847, ZN => n6656);
   U13860 : INV_X1 port map( A => n17269, ZN => n16863);
   U13861 : NAND2_X1 port map( A1 => n2985, A2 => n29299, ZN => n16773);
   U13862 : INV_X1 port map( A => n12000, ZN => n6658);
   U13863 : OAI21_X1 port map( B1 => n12004, B2 => n11996, A => n6658, ZN => 
                           n6657);
   U13864 : INV_X1 port map( A => n12004, ZN => n11538);
   U13865 : INV_X1 port map( A => n11755, ZN => n6661);
   U13866 : NAND2_X1 port map( A1 => n8957, A2 => n6662, ZN => n8959);
   U13867 : OR2_X1 port map( A1 => n18195, A2 => n6663, ZN => n18103);
   U13868 : NAND2_X1 port map( A1 => n10876, A2 => n29593, ZN => n11217);
   U13869 : INV_X1 port map( A => n18774, ZN => n19154);
   U13870 : XNOR2_X1 port map( A => n18774, B => n1982, ZN => n6667);
   U13872 : AND2_X1 port map( A1 => n29537, A2 => n27777, ZN => n27784);
   U13873 : INV_X1 port map( A => n15361, ZN => n6675);
   U13877 : NOR2_X1 port map( A1 => n10815, A2 => n6677, ZN => n10565);
   U13878 : NAND2_X1 port map( A1 => n11246, A2 => n12316, ZN => n6680);
   U13880 : INV_X1 port map( A => n16797, ZN => n17451);
   U13883 : XNOR2_X1 port map( A => n6683, B => n13543, ZN => n13456);
   U13884 : XNOR2_X1 port map( A => n6683, B => n5490, ZN => n11604);
   U13885 : XNOR2_X1 port map( A => n6683, B => n13459, ZN => n13296);
   U13886 : XNOR2_X1 port map( A => n6683, B => n13133, ZN => n12417);
   U13887 : OAI211_X1 port map( C1 => n28648, C2 => n14215, A => n14413, B => 
                           n6466, ZN => n13955);
   U13889 : NAND2_X1 port map( A1 => n24020, A2 => n23126, ZN => n24019);
   U13890 : AND2_X1 port map( A1 => n24020, A2 => n2054, ZN => n24543);
   U13891 : INV_X1 port map( A => n24020, ZN => n6686);
   U13892 : NAND2_X1 port map( A1 => n6693, A2 => n8977, ZN => n6691);
   U13893 : NAND2_X1 port map( A1 => n8978, A2 => n8976, ZN => n6693);
   U13894 : XNOR2_X1 port map( A => n22437, B => n22501, ZN => n22172);
   U13895 : NAND3_X1 port map( A1 => n6698, A2 => n5142, A3 => n6697, ZN => 
                           n6695);
   U13896 : NAND2_X1 port map( A1 => n20849, A2 => n21576, ZN => n6696);
   U13897 : NAND2_X1 port map( A1 => n21577, A2 => n21485, ZN => n6697);
   U13899 : NAND2_X1 port map( A1 => n17278, A2 => n539, ZN => n16766);
   U13901 : XNOR2_X1 port map( A => n18929, B => n19181, ZN => n6702);
   U13902 : XNOR2_X2 port map( A => n6702, B => n6701, ZN => n20148);
   U13903 : NAND2_X1 port map( A1 => n8427, A2 => n8351, ZN => n7809);
   U13904 : NAND2_X1 port map( A1 => n11195, A2 => n6687, ZN => n11568);
   U13905 : XNOR2_X1 port map( A => n6708, B => n26910, ZN => Ciphertext(46));
   U13906 : OR2_X1 port map( A1 => n26908, A2 => n27458, ZN => n6709);
   U13907 : OAI21_X1 port map( B1 => n6712, B2 => n6711, A => n27458, ZN => 
                           n6710);
   U13908 : NOR2_X1 port map( A1 => n28435, A2 => n29468, ZN => n6711);
   U13909 : NAND2_X1 port map( A1 => n23862, A2 => n25418, ZN => n26151);
   U13910 : NOR2_X1 port map( A1 => n17988, A2 => n17890, ZN => n6715);
   U13911 : NAND2_X1 port map( A1 => n6716, A2 => n6715, ZN => n6714);
   U13912 : XNOR2_X1 port map( A => n20761, B => n20760, ZN => n23010);
   U13913 : INV_X1 port map( A => n23010, ZN => n23657);
   U13914 : INV_X1 port map( A => n23140, ZN => n23141);
   U13915 : XNOR2_X1 port map( A => n19015, B => n19016, ZN => n6717);
   U13916 : INV_X1 port map( A => n28142, ZN => n18366);
   U13918 : XNOR2_X1 port map( A => n22363, B => n22434, ZN => n21620);
   U13919 : OAI21_X1 port map( B1 => n11328, B2 => n10858, A => n6721, ZN => 
                           n6720);
   U13920 : INV_X1 port map( A => n6722, ZN => n6721);
   U13921 : NAND2_X1 port map( A1 => n26940, A2 => n26943, ZN => n6724);
   U13922 : NAND2_X1 port map( A1 => n15407, A2 => n15108, ZN => n12371);
   U13924 : NAND2_X1 port map( A1 => n17500, A2 => n6727, ZN => n17503);
   U13926 : NOR2_X1 port map( A1 => n1835, A2 => n19956, ZN => n6729);
   U13927 : INV_X1 port map( A => n20321, ZN => n6730);
   U13928 : NOR2_X1 port map( A1 => n21248, A2 => n6730, ZN => n21249);
   U13929 : NOR2_X1 port map( A1 => n20695, A2 => n6730, ZN => n21254);
   U13930 : OR3_X1 port map( A1 => n21304, A2 => n21311, A3 => n29328, ZN => 
                           n6731);
   U13932 : NAND2_X1 port map( A1 => n6735, A2 => n27425, ZN => n6734);
   U13933 : MUX2_X1 port map( A => n27428, B => n27427, S => n29542, Z => n6735
                           );
   U13934 : NAND2_X1 port map( A1 => n26494, A2 => n29515, ZN => n6737);
   U13937 : NAND2_X1 port map( A1 => n6741, A2 => n24582, ZN => n6740);
   U13938 : NAND2_X1 port map( A1 => n11554, A2 => n6742, ZN => n6743);
   U13939 : OAI21_X1 port map( B1 => n11152, B2 => n593, A => n6745, ZN => 
                           n11157);
   U13940 : INV_X1 port map( A => n9146, ZN => n6747);
   U13941 : INV_X1 port map( A => n9146, ZN => n9150);
   U13942 : OAI211_X2 port map( C1 => n4104, C2 => n6751, A => n6750, B => 
                           n6749, ZN => n22619);
   U13943 : NAND2_X1 port map( A1 => n21494, A2 => n6752, ZN => n6751);
   U13944 : INV_X1 port map( A => n21496, ZN => n6752);
   U13945 : XNOR2_X1 port map( A => n6753, B => n16041, ZN => n6754);
   U13946 : XNOR2_X1 port map( A => n6754, B => n16042, ZN => n16679);
   U13947 : NAND2_X1 port map( A1 => n8227, A2 => n7424, ZN => n8224);
   U13948 : NAND2_X1 port map( A1 => n6756, A2 => n26995, ZN => n6755);
   U13949 : NAND2_X1 port map( A1 => n6757, A2 => n26632, ZN => n6756);
   U13950 : INV_X1 port map( A => n26632, ZN => n26996);
   U13951 : NAND2_X1 port map( A1 => n26997, A2 => n26998, ZN => n6757);
   U13953 : NAND2_X1 port map( A1 => n6759, A2 => n14796, ZN => n6758);
   U13954 : NAND2_X1 port map( A1 => n15204, A2 => n14961, ZN => n6759);
   U13955 : NAND2_X1 port map( A1 => n14927, A2 => n14968, ZN => n6760);
   U13956 : INV_X1 port map( A => n14961, ZN => n14967);
   U13957 : NAND2_X1 port map( A1 => n6762, A2 => n29531, ZN => n6761);
   U13958 : INV_X1 port map( A => n21308, ZN => n6762);
   U13959 : NAND2_X1 port map( A1 => n17399, A2 => n17398, ZN => n6765);
   U13960 : NAND2_X1 port map( A1 => n14238, A2 => n14171, ZN => n14174);
   U13961 : NAND2_X1 port map( A1 => n26435, A2 => n6768, ZN => n6767);
   U13962 : XNOR2_X1 port map( A => n22270, B => n22418, ZN => n22100);
   U13963 : INV_X1 port map( A => n16797, ZN => n6772);
   U13964 : NAND2_X1 port map( A1 => n6772, A2 => n17129, ZN => n17454);
   U13966 : NAND2_X1 port map( A1 => n10683, A2 => n5573, ZN => n6777);
   U13967 : NAND2_X1 port map( A1 => n10684, A2 => n6779, ZN => n6778);
   U13968 : NOR2_X1 port map( A1 => n8258, A2 => n28615, ZN => n6783);
   U13972 : AOI22_X1 port map( A1 => n8257, A2 => n6782, B1 => n28614, B2 => 
                           n28618, ZN => n6785);
   U13974 : NAND2_X1 port map( A1 => n24976, A2 => n23467, ZN => n6786);
   U13975 : NAND2_X1 port map( A1 => n24256, A2 => n24972, ZN => n24012);
   U13978 : OAI21_X1 port map( B1 => n26723, B2 => n26716, A => n6790, ZN => 
                           n25316);
   U13979 : NAND2_X1 port map( A1 => n26716, A2 => n283, ZN => n6790);
   U13983 : OAI21_X1 port map( B1 => n26216, B2 => n26217, A => n6793, ZN => 
                           n26218);
   U13984 : INV_X1 port map( A => n26723, ZN => n6793);
   U13985 : XNOR2_X2 port map( A => n6795, B => n9623, ZN => n11045);
   U13986 : XNOR2_X1 port map( A => n29509, B => n6796, ZN => n6795);
   U13987 : NAND2_X1 port map( A1 => n17453, A2 => n28193, ZN => n6799);
   U13988 : OAI21_X1 port map( B1 => n1814, B2 => n21459, A => n6803, ZN => 
                           n21570);
   U13989 : XNOR2_X1 port map( A => n19724, B => n19723, ZN => n6804);
   U13991 : MUX2_X1 port map( A => n20440, B => n20609, S => n20437, Z => 
                           n19886);
   U13993 : AOI22_X1 port map( A1 => n27372, A2 => n27366, B1 => n25360, B2 => 
                           n25359, ZN => n6806);
   U13994 : NOR2_X1 port map( A1 => n295, A2 => n28394, ZN => n27376);
   U13995 : OAI21_X1 port map( B1 => n27212, B2 => n27382, A => n6808, ZN => 
                           n6810);
   U13996 : NAND2_X1 port map( A1 => n6809, A2 => n5313, ZN => n6808);
   U13997 : NOR2_X1 port map( A1 => n27214, A2 => n6810, ZN => n27215);
   U13998 : OAI211_X1 port map( C1 => n524, C2 => n17771, A => n18254, B => 
                           n18252, ZN => n6811);
   U13999 : NAND2_X1 port map( A1 => n11867, A2 => n11869, ZN => n11462);
   U14002 : NOR2_X1 port map( A1 => n6814, A2 => n333, ZN => n10568);
   U14003 : INV_X1 port map( A => n10797, ZN => n6814);
   U14004 : NAND2_X1 port map( A1 => n11227, A2 => n11225, ZN => n6815);
   U14005 : NAND2_X1 port map( A1 => n11232, A2 => n6816, ZN => n11894);
   U14006 : XNOR2_X1 port map( A => n6817, B => n22238, ZN => n22244);
   U14007 : INV_X1 port map( A => n22748, ZN => n6817);
   U14008 : XNOR2_X1 port map( A => n22238, B => n6818, ZN => n22907);
   U14009 : XNOR2_X1 port map( A => n13221, B => n13220, ZN => n6820);
   U14010 : XNOR2_X2 port map( A => n6820, B => n6819, ZN => n14045);
   U14011 : NAND2_X1 port map( A1 => n23644, A2 => n23180, ZN => n6822);
   U14012 : NAND2_X1 port map( A1 => n6827, A2 => n26793, ZN => n6823);
   U14013 : NAND2_X1 port map( A1 => n25419, A2 => n6826, ZN => n6825);
   U14014 : INV_X1 port map( A => n26793, ZN => n6826);
   U14015 : NAND2_X1 port map( A1 => n26792, A2 => n26789, ZN => n6827);
   U14016 : INV_X1 port map( A => n16973, ZN => n6829);
   U14017 : INV_X1 port map( A => n12955, ZN => n12514);
   U14018 : INV_X1 port map( A => n13014, ZN => n13524);
   U14019 : XNOR2_X1 port map( A => n6831, B => n13014, ZN => n13442);
   U14020 : INV_X1 port map( A => n20495, ZN => n6834);
   U14021 : INV_X1 port map( A => n20494, ZN => n20218);
   U14022 : NAND2_X1 port map( A1 => n6841, A2 => n6838, ZN => n21251);
   U14023 : NAND2_X1 port map( A1 => n19506, A2 => n6843, ZN => n6841);
   U14024 : OAI22_X2 port map( A1 => n6841, A2 => n21248, B1 => n6839, B2 => 
                           n6842, ZN => n21809);
   U14025 : NAND2_X1 port map( A1 => n21251, A2 => n6840, ZN => n21807);
   U14026 : NAND4_X1 port map( A1 => n27500, A2 => n27499, A3 => n6845, A4 => 
                           n6844, ZN => n27501);
   U14027 : NAND3_X1 port map( A1 => n27487, A2 => n29093, A3 => n27496, ZN => 
                           n6844);
   U14028 : NAND2_X1 port map( A1 => n27495, A2 => n29093, ZN => n6845);
   U14029 : NAND3_X1 port map( A1 => n5811, A2 => n14969, A3 => n13789, ZN => 
                           n13788);
   U14030 : XNOR2_X1 port map( A => n22495, B => n22497, ZN => n6846);
   U14031 : XNOR2_X1 port map( A => n22498, B => n22496, ZN => n6847);
   U14032 : NAND2_X1 port map( A1 => n6850, A2 => n12257, ZN => n6849);
   U14033 : NAND2_X1 port map( A1 => n6855, A2 => n6853, ZN => n6852);
   U14034 : NAND2_X1 port map( A1 => n14943, A2 => n14944, ZN => n6855);
   U14035 : NAND2_X1 port map( A1 => n25506, A2 => n25505, ZN => n27054);
   U14036 : XNOR2_X1 port map( A => n6858, B => n26604, ZN => Ciphertext(177));
   U14037 : NAND2_X1 port map( A1 => n9028, A2 => n9030, ZN => n7715);
   U14038 : NOR2_X1 port map( A1 => n6636, A2 => n21465, ZN => n20755);
   U14039 : NOR2_X1 port map( A1 => n28155, A2 => n29236, ZN => n6861);
   U14041 : INV_X1 port map( A => n20277, ZN => n22041);
   U14042 : INV_X1 port map( A => n24631, ZN => n6867);
   U14043 : NOR2_X1 port map( A1 => n6866, A2 => n6867, ZN => n6864);
   U14044 : NOR2_X1 port map( A1 => n4366, A2 => n24532, ZN => n6866);
   U14045 : XNOR2_X1 port map( A => n13133, B => n12768, ZN => n13325);
   U14046 : INV_X1 port map( A => n14351, ZN => n13825);
   U14047 : NOR2_X1 port map( A1 => n13826, A2 => n14351, ZN => n6872);
   U14048 : NAND2_X1 port map( A1 => n596, A2 => n8642, ZN => n6875);
   U14049 : MUX2_X1 port map( A => n23849, B => n23721, S => n23726, Z => 
                           n22956);
   U14050 : NAND2_X1 port map( A1 => n23723, A2 => n29157, ZN => n23731);
   U14051 : NAND3_X1 port map( A1 => n6880, A2 => n6878, A3 => n6877, ZN => 
                           n15940);
   U14052 : NAND3_X1 port map( A1 => n6879, A2 => n3784, A3 => n426, ZN => 
                           n6878);
   U14053 : INV_X1 port map( A => n15371, ZN => n6879);
   U14054 : NAND3_X1 port map( A1 => n20628, A2 => n20334, A3 => n20258, ZN => 
                           n6882);
   U14055 : NAND2_X1 port map( A1 => n6884, A2 => n28186, ZN => n6881);
   U14056 : AND2_X1 port map( A1 => n20625, A2 => n20626, ZN => n6884);
   U14057 : XNOR2_X1 port map( A => n19322, B => n6886, ZN => n19326);
   U14058 : XNOR2_X1 port map( A => n19320, B => n19321, ZN => n6886);
   U14059 : NAND2_X1 port map( A1 => n26168, A2 => n29610, ZN => n6887);
   U14060 : NAND3_X1 port map( A1 => n4751, A2 => n26914, A3 => n1872, ZN => 
                           n6888);
   U14061 : NAND2_X1 port map( A1 => n17518, A2 => n17106, ZN => n6889);
   U14062 : XNOR2_X1 port map( A => n10303, B => n1983, ZN => n6891);
   U14064 : XNOR2_X1 port map( A => n13322, B => n2025, ZN => n6895);
   U14065 : NOR2_X1 port map( A1 => n14310, A2 => n14309, ZN => n14311);
   U14066 : NAND3_X2 port map( A1 => n10979, A2 => n10978, A3 => n6896, ZN => 
                           n12252);
   U14067 : INV_X1 port map( A => n12252, ZN => n11933);
   U14068 : XNOR2_X1 port map( A => n12522, B => n13434, ZN => n12526);
   U14069 : XNOR2_X1 port map( A => n25178, B => n25177, ZN => n26374);
   U14070 : OR2_X1 port map( A1 => n1030, A2 => n26380, ZN => n26430);
   U14071 : AOI21_X1 port map( B1 => n26991, B2 => n25770, A => n25769, ZN => 
                           n26537);
   U14072 : OR2_X1 port map( A1 => n26254, A2 => n28053, ZN => n26255);
   U14075 : BUF_X1 port map( A => n12762, Z => n12735);
   U14076 : OAI211_X1 port map( C1 => n28012, C2 => n443, A => n28011, B => 
                           n28010, ZN => n28014);
   U14078 : OR2_X1 port map( A1 => n29036, A2 => n28601, ZN => n12796);
   U14079 : INV_X1 port map( A => n15738, ZN => n16483);
   U14080 : XNOR2_X2 port map( A => n25085, B => n25084, ZN => n26917);
   U14081 : MUX2_X2 port map( A => n26916, B => n26915, S => n26914, Z => 
                           n27531);
   U14082 : OR2_X1 port map( A1 => n25957, A2 => n27357, ZN => n25671);
   U14083 : OR2_X1 port map( A1 => n25997, A2 => n28562, ZN => n26002);
   U14084 : AOI22_X1 port map( A1 => n27091, A2 => n27090, B1 => n27089, B2 => 
                           n27088, ZN => n27271);
   U14085 : NAND2_X1 port map( A1 => n23949, A2 => n23948, ZN => n25922);
   U14086 : OAI22_X1 port map( A1 => n28003, A2 => n28019, B1 => n28001, B2 => 
                           n28015, ZN => n28022);
   U14087 : NOR2_X1 port map( A1 => n17729, A2 => n18456, ZN => n17731);
   U14088 : OR2_X1 port map( A1 => n24556, A2 => n24551, ZN => n24175);
   U14089 : AND3_X1 port map( A1 => n27521, A2 => n27527, A3 => n27520, ZN => 
                           n27522);
   U14091 : AND2_X1 port map( A1 => n27843, A2 => n27101, ZN => n27099);
   U14092 : NOR2_X1 port map( A1 => n23906, A2 => n24373, ZN => n24377);
   U14093 : AND2_X1 port map( A1 => n13844, A2 => n15456, ZN => n13845);
   U14094 : OR2_X1 port map( A1 => n22451, A2 => n23387, ZN => n23222);
   U14095 : OR2_X1 port map( A1 => n21591, A2 => n21322, ZN => n21323);
   U14096 : AND2_X1 port map( A1 => n24427, A2 => n28531, ZN => n24428);
   U14097 : AND2_X1 port map( A1 => n25660, A2 => n26721, ZN => n26217);
   U14101 : NOR2_X2 port map( A1 => n23910, A2 => n23909, ZN => n25375);
   U14102 : XNOR2_X1 port map( A => n25248, B => n25830, ZN => n26754);
   U14103 : OR2_X1 port map( A1 => n14215, A2 => n13686, ZN => n14419);
   U14104 : AND2_X1 port map( A1 => n27562, A2 => n27551, ZN => n27149);
   U14105 : OR2_X1 port map( A1 => n27101, A2 => n27100, ZN => n27248);
   U14106 : AOI21_X1 port map( B1 => n27637, B2 => n26980, A => n26672, ZN => 
                           n26675);
   U14108 : OR2_X1 port map( A1 => n339, A2 => n23776, ZN => n23780);
   U14109 : XNOR2_X2 port map( A => n25326, B => n25327, ZN => n26204);
   U14110 : XNOR2_X2 port map( A => n7137, B => Key(53), ZN => n8014);
   U14112 : INV_X1 port map( A => n27638, ZN => n27637);
   U14114 : INV_X1 port map( A => n26933, ZN => n24788);
   U14115 : AND2_X1 port map( A1 => n24390, A2 => n24391, ZN => n23900);
   U14116 : OAI21_X1 port map( B1 => n24364, B2 => n28592, A => n24363, ZN => 
                           n26705);
   U14117 : NOR2_X1 port map( A1 => n449, A2 => n29468, ZN => n26605);
   U14118 : XNOR2_X1 port map( A => n22511, B => n22510, ZN => n22512);
   U14119 : OR2_X1 port map( A1 => n20444, A2 => n415, ZN => n19505);
   U14121 : XNOR2_X1 port map( A => n25507, B => n25210, ZN => n25212);
   U14122 : INV_X1 port map( A => n24858, ZN => n25848);
   U14126 : XNOR2_X1 port map( A => n25351, B => n25352, ZN => n26077);
   U14127 : XNOR2_X2 port map( A => n16188, B => n16187, ZN => n17467);
   U14128 : OAI21_X1 port map( B1 => n26159, B2 => n26457, A => n25616, ZN => 
                           n25633);
   U14132 : NOR2_X2 port map( A1 => n17538, A2 => n17537, ZN => n19555);
   U14133 : OAI211_X2 port map( C1 => n18445, C2 => n18185, A => n18184, B => 
                           n18183, ZN => n19397);
   U14134 : OR2_X1 port map( A1 => n28524, A2 => n24716, ZN => n24353);
   U14136 : AND2_X1 port map( A1 => n9194, A2 => n329, ZN => n6897);
   U14137 : XOR2_X1 port map( A => n10248, B => n10247, Z => n6898);
   U14138 : OR2_X1 port map( A1 => n17561, A2 => n17560, ZN => n6899);
   U14139 : OR3_X1 port map( A1 => n17402, A2 => n29572, A3 => n17400, ZN => 
                           n6900);
   U14140 : AND2_X1 port map( A1 => n8381, A2 => n8384, ZN => n6901);
   U14141 : OR2_X1 port map( A1 => n29314, A2 => n1930, ZN => n6904);
   U14142 : OR2_X1 port map( A1 => n7626, A2 => n8217, ZN => n6905);
   U14143 : AND2_X1 port map( A1 => n2209, A2 => n29643, ZN => n6906);
   U14144 : AND2_X1 port map( A1 => n27859, A2 => n27847, ZN => n6907);
   U14145 : OR2_X1 port map( A1 => n8487, A2 => n8486, ZN => n6908);
   U14146 : AOI21_X1 port map( B1 => n25975, B2 => n26236, A => n25974, ZN => 
                           n28009);
   U14148 : AND2_X1 port map( A1 => n8384, A2 => n8729, ZN => n6909);
   U14149 : AND2_X1 port map( A1 => n5425, A2 => n26880, ZN => n6910);
   U14150 : AND2_X1 port map( A1 => n21292, A2 => n20726, ZN => n6911);
   U14152 : NAND2_X1 port map( A1 => n26274, A2 => n26273, ZN => n27582);
   U14153 : INV_X1 port map( A => n27582, ZN => n26346);
   U14154 : INV_X1 port map( A => n2274, ZN => n22755);
   U14155 : AND2_X1 port map( A1 => n9033, A2 => n9032, ZN => n6915);
   U14156 : AND2_X1 port map( A1 => n11723, A2 => n11722, ZN => n6917);
   U14157 : AND2_X1 port map( A1 => n10761, A2 => n11119, ZN => n6918);
   U14158 : OR2_X1 port map( A1 => n12339, A2 => n12338, ZN => n6919);
   U14159 : AND2_X1 port map( A1 => n12049, A2 => n12050, ZN => n6920);
   U14160 : OR2_X1 port map( A1 => n14233, A2 => n14593, ZN => n6921);
   U14161 : XOR2_X1 port map( A => n13099, B => n13098, Z => n6922);
   U14162 : XOR2_X1 port map( A => n12570, B => n12569, Z => n6923);
   U14163 : INV_X1 port map( A => n15420, ZN => n15422);
   U14164 : OR2_X1 port map( A1 => n17264, A2 => n16996, ZN => n6926);
   U14165 : AND3_X2 port map( A1 => n16998, A2 => n16997, A3 => n6926, ZN => 
                           n6927);
   U14166 : AND2_X1 port map( A1 => n16884, A2 => n16883, ZN => n6928);
   U14167 : XOR2_X1 port map( A => n15563, B => n15562, Z => n6929);
   U14168 : AND2_X1 port map( A1 => n17637, A2 => n17636, ZN => n6930);
   U14170 : XNOR2_X1 port map( A => n18617, B => n18616, ZN => n20568);
   U14171 : OR2_X1 port map( A1 => n20567, A2 => n20573, ZN => n6932);
   U14172 : AND2_X1 port map( A1 => n21412, A2 => n20663, ZN => n6933);
   U14173 : AND2_X1 port map( A1 => n20201, A2 => n20200, ZN => n6935);
   U14174 : OR2_X1 port map( A1 => n21500, A2 => n21192, ZN => n6936);
   U14175 : AND2_X1 port map( A1 => n20118, A2 => n21424, ZN => n6937);
   U14176 : XOR2_X1 port map( A => n22591, B => n22590, Z => n6938);
   U14177 : XOR2_X1 port map( A => n22666, B => n22665, Z => n6939);
   U14178 : OR2_X1 port map( A1 => n22402, A2 => n22401, ZN => n6940);
   U14179 : AND2_X1 port map( A1 => n23145, A2 => n23461, ZN => n6941);
   U14180 : XNOR2_X1 port map( A => n17752, B => n17751, ZN => n20412);
   U14182 : OR2_X1 port map( A1 => n1955, A2 => n28512, ZN => n6943);
   U14183 : OR2_X1 port map( A1 => n24672, A2 => n28635, ZN => n6944);
   U14184 : OR3_X1 port map( A1 => n24347, A2 => n24437, A3 => n24433, ZN => 
                           n6945);
   U14185 : OR2_X1 port map( A1 => n24806, A2 => n24261, ZN => n6946);
   U14186 : XOR2_X1 port map( A => n25414, B => n25413, Z => n6947);
   U14187 : AND2_X1 port map( A1 => n6768, A2 => n26940, ZN => n6948);
   U14188 : AND2_X1 port map( A1 => n27852, A2 => n27854, ZN => n6949);
   U14189 : OR2_X1 port map( A1 => n5505, A2 => n26933, ZN => n6950);
   U14190 : OR2_X1 port map( A1 => n27118, A2 => n26835, ZN => n6951);
   U14191 : OR2_X1 port map( A1 => n26146, A2 => n325, ZN => n6952);
   U14192 : AND2_X1 port map( A1 => n326, A2 => n26126, ZN => n6953);
   U14193 : OR3_X1 port map( A1 => n27855, A2 => n26641, A3 => n27847, ZN => 
                           n6954);
   U14194 : AND2_X1 port map( A1 => n28021, A2 => n28003, ZN => n6955);
   U14195 : AND2_X1 port map( A1 => n14230, A2 => n14101, ZN => n6956);
   U14196 : OR2_X1 port map( A1 => n7759, A2 => n8176, ZN => n7345);
   U14197 : OR2_X1 port map( A1 => n7958, A2 => n7589, ZN => n7590);
   U14198 : INV_X1 port map( A => n8161, ZN => n8166);
   U14199 : INV_X1 port map( A => Plaintext(159), ZN => n7049);
   U14200 : OR2_X1 port map( A1 => n8270, A2 => n8267, ZN => n7211);
   U14201 : OR2_X1 port map( A1 => n8280, A2 => n8275, ZN => n7407);
   U14202 : BUF_X1 port map( A => n7069, Z => n7582);
   U14203 : XNOR2_X1 port map( A => Key(125), B => Plaintext(125), ZN => n8290)
                           ;
   U14204 : OR2_X1 port map( A1 => n8336, A2 => n8886, ZN => n8007);
   U14205 : INV_X1 port map( A => n8462, ZN => n7445);
   U14206 : OR2_X1 port map( A1 => n7618, A2 => n8256, ZN => n7389);
   U14207 : INV_X1 port map( A => Plaintext(167), ZN => n7058);
   U14208 : OR2_X1 port map( A1 => n7763, A2 => n613, ZN => n7764);
   U14209 : OR2_X1 port map( A1 => n8300, A2 => n7400, ZN => n7940);
   U14210 : INV_X1 port map( A => n29081, ZN => n8002);
   U14211 : INV_X1 port map( A => n8397, ZN => n8864);
   U14212 : INV_X1 port map( A => n8873, ZN => n8876);
   U14213 : OR2_X1 port map( A1 => n8917, A2 => n9108, ZN => n8915);
   U14214 : OR2_X1 port map( A1 => n8955, A2 => n8801, ZN => n9162);
   U14215 : AOI22_X1 port map( A1 => n7720, A2 => n8049, B1 => n7719, B2 => 
                           n7718, ZN => n7726);
   U14216 : INV_X1 port map( A => n9060, ZN => n8866);
   U14217 : INV_X1 port map( A => n9562, ZN => n8765);
   U14218 : OR2_X1 port map( A1 => n8549, A2 => n7410, ZN => n7412);
   U14219 : OR2_X1 port map( A1 => n9060, A2 => n8872, ZN => n8395);
   U14220 : OR2_X1 port map( A1 => n9582, A2 => n1196, ZN => n9583);
   U14221 : OR2_X1 port map( A1 => n8965, A2 => n8963, ZN => n8640);
   U14222 : INV_X1 port map( A => n8763, ZN => n8945);
   U14223 : INV_X1 port map( A => n8608, ZN => n9529);
   U14224 : INV_X1 port map( A => n10956, ZN => n9858);
   U14225 : XNOR2_X1 port map( A => n10271, B => n10350, ZN => n9849);
   U14226 : OAI211_X1 port map( C1 => n9160, C2 => n8625, A => n8624, B => 
                           n8804, ZN => n9306);
   U14227 : XNOR2_X1 port map( A => n9838, B => n9495, ZN => n9496);
   U14228 : INV_X1 port map( A => n9701, ZN => n9666);
   U14229 : XNOR2_X1 port map( A => n10249, B => n6898, ZN => n10534);
   U14230 : XNOR2_X1 port map( A => n10175, B => n10174, ZN => n11067);
   U14231 : XNOR2_X1 port map( A => n7571, B => n7570, ZN => n7572);
   U14232 : OR2_X1 port map( A1 => n11223, A2 => n29593, ZN => n10660);
   U14233 : XNOR2_X1 port map( A => n9336, B => n9780, ZN => n9337);
   U14234 : NOR2_X1 port map( A1 => n9860, A2 => n9859, ZN => n9861);
   U14237 : AND2_X1 port map( A1 => n11147, A2 => n10742, ZN => n11148);
   U14238 : BUF_X1 port map( A => n10518, Z => n11027);
   U14239 : XNOR2_X1 port map( A => n10299, B => n10417, ZN => n10301);
   U14240 : XNOR2_X1 port map( A => n10279, B => n10278, ZN => n11223);
   U14241 : XNOR2_X1 port map( A => n9337, B => n9338, ZN => n10912);
   U14242 : XNOR2_X1 port map( A => n8090, B => n8089, ZN => n10820);
   U14243 : AOI21_X1 port map( B1 => n10807, B2 => n11149, A => n11148, ZN => 
                           n11419);
   U14244 : OR2_X1 port map( A1 => n11039, A2 => n28612, ZN => n11040);
   U14245 : OAI21_X1 port map( B1 => n10894, B2 => n10893, A => n10892, ZN => 
                           n11660);
   U14246 : INV_X1 port map( A => n11739, ZN => n11908);
   U14247 : NOR2_X1 port map( A1 => n11940, A2 => n12517, ZN => n12579);
   U14248 : INV_X1 port map( A => n12188, ZN => n12192);
   U14249 : OR2_X1 port map( A1 => n10908, A2 => n11927, ZN => n10909);
   U14250 : AND2_X1 port map( A1 => n12022, A2 => n12354, ZN => n12429);
   U14251 : OR2_X1 port map( A1 => n11395, A2 => n11951, ZN => n11396);
   U14252 : AOI22_X1 port map( A1 => n10782, A2 => n9858, B1 => n10781, B2 => 
                           n10780, ZN => n10793);
   U14253 : OAI21_X1 port map( B1 => n12100, B2 => n12099, A => n12098, ZN => 
                           n12101);
   U14254 : OAI21_X1 port map( B1 => n12579, B2 => n12575, A => n11591, ZN => 
                           n11592);
   U14255 : AOI21_X1 port map( B1 => n10645, B2 => n12219, A => n10644, ZN => 
                           n12608);
   U14256 : INV_X1 port map( A => n13012, ZN => n13013);
   U14258 : OR2_X1 port map( A1 => n11655, A2 => n11378, ZN => n11379);
   U14259 : INV_X1 port map( A => n14830, ZN => n14831);
   U14260 : AND2_X1 port map( A1 => n14400, A2 => n14399, ZN => n14403);
   U14261 : XNOR2_X1 port map( A => n12904, B => n12298, ZN => n11734);
   U14263 : OR2_X1 port map( A1 => n14264, A2 => n14259, ZN => n13762);
   U14264 : INV_X1 port map( A => n14287, ZN => n14085);
   U14265 : XNOR2_X1 port map( A => n13520, B => n12634, ZN => n12635);
   U14266 : XNOR2_X1 port map( A => n13241, B => n13242, ZN => n14046);
   U14267 : XNOR2_X1 port map( A => n10444, B => n10443, ZN => n13606);
   U14268 : INV_X1 port map( A => n14314, ZN => n13884);
   U14269 : XNOR2_X1 port map( A => n12386, B => n12387, ZN => n14407);
   U14270 : AND2_X1 port map( A1 => n13629, A2 => n13628, ZN => n13630);
   U14271 : OR2_X1 port map( A1 => n14298, A2 => n13803, ZN => n13658);
   U14272 : OR2_X1 port map( A1 => n15127, A2 => n15001, ZN => n14999);
   U14273 : INV_X1 port map( A => n15000, ZN => n13632);
   U14275 : AND2_X1 port map( A1 => n14563, A2 => n15083, ZN => n14670);
   U14277 : INV_X1 port map( A => n14706, ZN => n14431);
   U14279 : AND2_X1 port map( A1 => n13632, A2 => n15123, ZN => n14686);
   U14280 : OR2_X1 port map( A1 => n14874, A2 => n15071, ZN => n14876);
   U14281 : INV_X1 port map( A => n15015, ZN => n15327);
   U14282 : AND2_X1 port map( A1 => n17474, A2 => n17124, ZN => n17480);
   U14283 : XNOR2_X1 port map( A => n16638, B => n16637, ZN => n16724);
   U14284 : BUF_X1 port map( A => n16477, Z => n15777);
   U14286 : XNOR2_X1 port map( A => n15771, B => n15770, ZN => n15776);
   U14287 : XNOR2_X1 port map( A => n16218, B => n16145, ZN => n15820);
   U14288 : INV_X1 port map( A => n17350, ZN => n17351);
   U14289 : INV_X1 port map( A => n18124, ZN => n18125);
   U14290 : OR2_X1 port map( A1 => n18513, A2 => n18516, ZN => n18514);
   U14291 : INV_X1 port map( A => n18707, ZN => n17980);
   U14292 : OR2_X1 port map( A1 => n16726, A2 => n16725, ZN => n16727);
   U14293 : XNOR2_X1 port map( A => n16350, B => n16349, ZN => n16712);
   U14295 : OAI211_X1 port map( C1 => n17217, C2 => n16940, A => n15809, B => 
                           n15808, ZN => n15810);
   U14296 : AND2_X1 port map( A1 => n18042, A2 => n18422, ZN => n17822);
   U14297 : INV_X1 port map( A => n18433, ZN => n18149);
   U14298 : INV_X1 port map( A => n18314, ZN => n16442);
   U14299 : INV_X1 port map( A => n18528, ZN => n17699);
   U14300 : AND2_X1 port map( A1 => n18261, A2 => n18262, ZN => n17896);
   U14301 : INV_X1 port map( A => n17353, ZN => n18706);
   U14302 : AND2_X1 port map( A1 => n18190, A2 => n19562, ZN => n17796);
   U14304 : NOR2_X1 port map( A1 => n17775, A2 => n17774, ZN => n17776);
   U14305 : NOR2_X1 port map( A1 => n17703, A2 => n17702, ZN => n17704);
   U14307 : XNOR2_X1 port map( A => n19718, B => n3423, ZN => n19180);
   U14308 : XNOR2_X1 port map( A => n19413, B => n19412, ZN => n19624);
   U14309 : OR2_X1 port map( A1 => n20480, A2 => n20475, ZN => n20355);
   U14310 : XNOR2_X1 port map( A => n17630, B => n17631, ZN => n17687);
   U14311 : XNOR2_X1 port map( A => n19074, B => n19073, ZN => n19093);
   U14312 : AND2_X1 port map( A1 => n28140, A2 => n20413, ZN => n20583);
   U14313 : XNOR2_X1 port map( A => n19444, B => n19443, ZN => n19795);
   U14314 : AND2_X1 port map( A1 => n20157, A2 => n20159, ZN => n19983);
   U14315 : INV_X1 port map( A => n21653, ZN => n21012);
   U14317 : XNOR2_X1 port map( A => n18905, B => n18904, ZN => n19766);
   U14318 : XNOR2_X1 port map( A => n19239, B => n19238, ZN => n20013);
   U14319 : XNOR2_X1 port map( A => n18686, B => n18685, ZN => n18699);
   U14320 : NAND2_X1 port map( A1 => n19950, A2 => n20314, ZN => n19951);
   U14321 : INV_X1 port map( A => n21429, ZN => n22397);
   U14323 : OR2_X1 port map( A1 => n21435, A2 => n20339, ZN => n20011);
   U14324 : OAI21_X1 port map( B1 => n20392, B2 => n20545, A => n20391, ZN => 
                           n20393);
   U14325 : OR2_X1 port map( A1 => n21401, A2 => n20658, ZN => n21043);
   U14326 : AND2_X1 port map( A1 => n20857, A2 => n21156, ZN => n20527);
   U14327 : OAI22_X1 port map( A1 => n20622, A2 => n20621, B1 => n20620, B2 => 
                           n20619, ZN => n20722);
   U14328 : AND2_X1 port map( A1 => n20241, A2 => n29527, ZN => n19792);
   U14329 : INV_X1 port map( A => n21014, ZN => n21664);
   U14330 : OAI211_X1 port map( C1 => n20205, C2 => n20307, A => n20204, B => 
                           n20203, ZN => n20207);
   U14331 : OR2_X1 port map( A1 => n21347, A2 => n28440, ZN => n21344);
   U14332 : XNOR2_X1 port map( A => n22677, B => n5513, ZN => n22680);
   U14333 : AND2_X1 port map( A1 => n20951, A2 => n20184, ZN => n20185);
   U14334 : INV_X1 port map( A => n21286, ZN => n21297);
   U14335 : AOI21_X1 port map( B1 => n3763, B2 => n21307, A => n20772, ZN => 
                           n20773);
   U14336 : AND2_X1 port map( A1 => n21194, A2 => n21500, ZN => n21195);
   U14337 : OR2_X1 port map( A1 => n22404, A2 => n22398, ZN => n20276);
   U14338 : INV_X1 port map( A => n28327, ZN => n22534);
   U14339 : INV_X1 port map( A => n22677, ZN => n22556);
   U14341 : OR2_X1 port map( A1 => n23245, A2 => n23246, ZN => n22984);
   U14342 : XNOR2_X1 port map( A => n22697, B => n22879, ZN => n22468);
   U14343 : XNOR2_X1 port map( A => n22615, B => n22656, ZN => n22350);
   U14344 : OR2_X1 port map( A1 => n23456, A2 => n23148, ZN => n23149);
   U14345 : AND2_X1 port map( A1 => n23416, A2 => n23419, ZN => n23098);
   U14346 : XNOR2_X1 port map( A => n22157, B => n20470, ZN => n20471);
   U14347 : XNOR2_X1 port map( A => n21937, B => n22500, ZN => n22205);
   U14348 : XNOR2_X1 port map( A => n22468, B => n22467, ZN => n22471);
   U14349 : XNOR2_X1 port map( A => n22478, B => n22477, ZN => n22494);
   U14350 : XNOR2_X1 port map( A => n22654, B => n22653, ZN => n23102);
   U14351 : XNOR2_X1 port map( A => n21546, B => n21545, ZN => n21559);
   U14352 : OR2_X1 port map( A1 => n23427, A2 => n1873, ZN => n23341);
   U14353 : XNOR2_X1 port map( A => n21852, B => n21851, ZN => n23156);
   U14354 : INV_X1 port map( A => n24502, ZN => n24503);
   U14355 : XNOR2_X1 port map( A => n21341, B => n21340, ZN => n23422);
   U14357 : BUF_X1 port map( A => n22284, Z => n23558);
   U14358 : AND2_X1 port map( A1 => n23727, A2 => n23726, ZN => n23728);
   U14359 : XNOR2_X1 port map( A => n22512, B => n22513, ZN => n23077);
   U14360 : OR2_X1 port map( A1 => n24682, A2 => n24688, ZN => n24311);
   U14363 : OR2_X1 port map( A1 => n24891, A2 => n24631, ZN => n24297);
   U14364 : NOR2_X1 port map( A1 => n23036, A2 => n23482, ZN => n23486);
   U14365 : OR2_X1 port map( A1 => n21898, A2 => n23662, ZN => n21724);
   U14366 : INV_X1 port map( A => n24600, ZN => n24607);
   U14367 : NOR2_X1 port map( A1 => n23729, A2 => n23728, ZN => n23730);
   U14368 : AND2_X1 port map( A1 => n404, A2 => n24678, ZN => n24067);
   U14369 : AND2_X1 port map( A1 => n29050, A2 => n24603, ZN => n24285);
   U14371 : OR2_X1 port map( A1 => n1883, A2 => n23378, ZN => n23379);
   U14372 : AND2_X1 port map( A1 => n24772, A2 => n24766, ZN => n24774);
   U14373 : AND2_X1 port map( A1 => n26240, A2 => n26761, ZN => n25602);
   U14374 : AND2_X1 port map( A1 => n26450, A2 => n26449, ZN => n26451);
   U14375 : AOI21_X1 port map( B1 => n26427, B2 => n26426, A => n26425, ZN => 
                           n26428);
   U14376 : XNOR2_X1 port map( A => n25138, B => n25137, ZN => n26436);
   U14377 : XNOR2_X1 port map( A => n26008, B => n24955, ZN => n24958);
   U14378 : INV_X1 port map( A => n25270, ZN => n25056);
   U14379 : XNOR2_X1 port map( A => n25886, B => n1225, ZN => n25557);
   U14380 : OR2_X1 port map( A1 => n28660, A2 => n27069, ZN => n25963);
   U14382 : INV_X1 port map( A => n26240, ZN => n25603);
   U14383 : OR2_X1 port map( A1 => n26194, A2 => n26191, ZN => n25240);
   U14384 : AND2_X1 port map( A1 => n26949, A2 => n26266, ZN => n26267);
   U14385 : XNOR2_X1 port map( A => n24882, B => n24881, ZN => n26263);
   U14386 : XNOR2_X1 port map( A => n26007, B => n26008, ZN => n26009);
   U14387 : XNOR2_X1 port map( A => n26077, B => n26076, ZN => n26078);
   U14389 : NOR2_X1 port map( A1 => n26748, A2 => n25453, ZN => n25461);
   U14390 : XNOR2_X1 port map( A => n25229, B => n25228, ZN => n26729);
   U14392 : OR2_X1 port map( A1 => n28561, A2 => n28525, ZN => n24200);
   U14393 : XNOR2_X1 port map( A => n25917, B => n25918, ZN => n26850);
   U14394 : AOI21_X1 port map( B1 => n29482, B2 => n26998, A => n26995, ZN => 
                           n25972);
   U14395 : OR2_X1 port map( A1 => n27388, A2 => n27402, ZN => n25627);
   U14396 : AND3_X1 port map( A1 => n24202, A2 => n24201, A3 => n24200, ZN => 
                           n24203);
   U14397 : INV_X1 port map( A => n27282, ZN => n27278);
   U14398 : NAND2_X1 port map( A1 => n26434, A2 => n26433, ZN => n26880);
   U14399 : AND2_X1 port map( A1 => n26846, A2 => n27827, ZN => n26902);
   U14400 : INV_X1 port map( A => n27852, ZN => n27847);
   U14401 : AND2_X1 port map( A1 => n27872, A2 => n27865, ZN => n25897);
   U14402 : OR2_X1 port map( A1 => n26984, A2 => n28001, ZN => n28002);
   U14403 : BUF_X1 port map( A => n28009, Z => n28003);
   U14404 : OR2_X1 port map( A1 => n25957, A2 => n27328, ZN => n25958);
   U14405 : OR2_X1 port map( A1 => n26816, A2 => n24826, ZN => n24827);
   U14407 : AOI22_X1 port map( A1 => n26809, A2 => n25997, B1 => n25995, B2 => 
                           n27363, ZN => n25996);
   U14408 : AND3_X1 port map( A1 => n27615, A2 => n26973, A3 => n3154, ZN => 
                           n27624);
   U14409 : INV_X1 port map( A => n25991, ZN => n25992);
   U14410 : INV_X1 port map( A => Plaintext(113), ZN => n6957);
   U14411 : XNOR2_X1 port map( A => n6957, B => Key(113), ZN => n6958);
   U14413 : XNOR2_X1 port map( A => Key(109), B => Plaintext(109), ZN => n7924)
                           ;
   U14414 : NAND2_X1 port map( A1 => n8214, A2 => n626, ZN => n6963);
   U14415 : INV_X1 port map( A => n8216, ZN => n7437);
   U14416 : OAI21_X1 port map( B1 => n7437, B2 => n7626, A => n7924, ZN => 
                           n6962);
   U14419 : OAI21_X1 port map( B1 => n8216, B2 => n8213, A => n7625, ZN => 
                           n6960);
   U14420 : INV_X1 port map( A => Plaintext(114), ZN => n6964);
   U14421 : XNOR2_X1 port map( A => n6964, B => Key(114), ZN => n7613);
   U14422 : INV_X1 port map( A => n7614, ZN => n7932);
   U14424 : INV_X1 port map( A => n7933, ZN => n8308);
   U14425 : NAND2_X1 port map( A1 => n8308, A2 => n7935, ZN => n6965);
   U14426 : MUX2_X1 port map( A => n8310, B => n6965, S => n29135, Z => n6967);
   U14427 : XNOR2_X1 port map( A => Key(115), B => Plaintext(115), ZN => n7393)
                           ;
   U14428 : OAI211_X1 port map( C1 => n7613, C2 => n7393, A => n8310, B => 
                           n7934, ZN => n6966);
   U14429 : AND2_X1 port map( A1 => n6967, A2 => n6966, ZN => n9230);
   U14430 : INV_X1 port map( A => n9230, ZN => n9047);
   U14431 : INV_X1 port map( A => Plaintext(103), ZN => n6968);
   U14432 : INV_X1 port map( A => n7619, ZN => n8235);
   U14433 : INV_X1 port map( A => Plaintext(104), ZN => n6969);
   U14434 : INV_X1 port map( A => Plaintext(107), ZN => n6970);
   U14435 : INV_X1 port map( A => Plaintext(106), ZN => n6971);
   U14437 : NAND2_X1 port map( A1 => n7358, A2 => n8237, ZN => n7431);
   U14438 : INV_X1 port map( A => Plaintext(102), ZN => n6972);
   U14439 : NAND2_X1 port map( A1 => n8232, A2 => n8231, ZN => n6974);
   U14440 : XNOR2_X1 port map( A => Key(100), B => Plaintext(100), ZN => n7362)
                           ;
   U14441 : INV_X1 port map( A => Plaintext(101), ZN => n6977);
   U14442 : AND2_X1 port map( A1 => n8205, A2 => n7362, ZN => n6983);
   U14443 : INV_X1 port map( A => Plaintext(97), ZN => n6978);
   U14445 : INV_X1 port map( A => n7634, ZN => n8199);
   U14446 : INV_X1 port map( A => Plaintext(99), ZN => n6979);
   U14447 : INV_X1 port map( A => n7635, ZN => n8201);
   U14448 : NAND2_X1 port map( A1 => n8199, A2 => n8201, ZN => n6982);
   U14449 : INV_X1 port map( A => Plaintext(96), ZN => n6980);
   U14451 : INV_X1 port map( A => n7363, ZN => n8207);
   U14452 : MUX2_X1 port map( A => n7832, B => n8207, S => n28605, Z => n6981);
   U14454 : INV_X1 port map( A => Plaintext(93), ZN => n6984);
   U14455 : XNOR2_X1 port map( A => n6984, B => Key(93), ZN => n6988);
   U14456 : INV_X1 port map( A => Plaintext(94), ZN => n6985);
   U14457 : XNOR2_X1 port map( A => n6985, B => Key(94), ZN => n7825);
   U14458 : INV_X1 port map( A => n7825, ZN => n7695);
   U14459 : INV_X1 port map( A => Plaintext(90), ZN => n6986);
   U14460 : OAI21_X1 port map( B1 => n7821, B2 => n7695, A => n6987, ZN => 
                           n6994);
   U14461 : INV_X1 port map( A => Plaintext(91), ZN => n6989);
   U14463 : INV_X1 port map( A => Plaintext(92), ZN => n6990);
   U14464 : XNOR2_X1 port map( A => n6990, B => Key(92), ZN => n7371);
   U14465 : XNOR2_X1 port map( A => Key(95), B => Plaintext(95), ZN => n8221);
   U14466 : INV_X1 port map( A => n8221, ZN => n8223);
   U14467 : NAND2_X1 port map( A1 => n6991, A2 => n8223, ZN => n6992);
   U14468 : INV_X1 port map( A => Plaintext(120), ZN => n6995);
   U14470 : INV_X1 port map( A => Plaintext(121), ZN => n6996);
   U14471 : INV_X1 port map( A => n8290, ZN => n7910);
   U14472 : INV_X1 port map( A => Plaintext(122), ZN => n6997);
   U14474 : INV_X1 port map( A => n7909, ZN => n7914);
   U14475 : XNOR2_X1 port map( A => Key(124), B => Plaintext(124), ZN => n8287)
                           ;
   U14476 : INV_X1 port map( A => Plaintext(123), ZN => n6998);
   U14477 : XNOR2_X1 port map( A => n6998, B => Key(123), ZN => n7911);
   U14478 : XNOR2_X1 port map( A => Key(73), B => Plaintext(73), ZN => n7498);
   U14479 : INV_X1 port map( A => n7498, ZN => n7708);
   U14480 : XNOR2_X1 port map( A => Key(75), B => Plaintext(75), ZN => n7382);
   U14481 : AND2_X1 port map( A1 => n7498, A2 => n7382, ZN => n7855);
   U14482 : INV_X1 port map( A => n7855, ZN => n7002);
   U14483 : XNOR2_X1 port map( A => Key(74), B => Plaintext(74), ZN => n7852);
   U14484 : NAND3_X1 port map( A1 => n7856, A2 => n7002, A3 => n3594, ZN => 
                           n7006);
   U14485 : XNOR2_X1 port map( A => Key(76), B => Plaintext(76), ZN => n7384);
   U14486 : INV_X1 port map( A => n7384, ZN => n7494);
   U14487 : INV_X1 port map( A => n7852, ZN => n7496);
   U14488 : INV_X1 port map( A => Plaintext(72), ZN => n7003);
   U14489 : NAND2_X1 port map( A1 => n617, A2 => n7382, ZN => n7707);
   U14490 : NAND2_X1 port map( A1 => n7707, A2 => n371, ZN => n7004);
   U14491 : XNOR2_X1 port map( A => Key(67), B => Plaintext(67), ZN => n7850);
   U14492 : INV_X1 port map( A => Plaintext(69), ZN => n7007);
   U14493 : INV_X1 port map( A => Plaintext(71), ZN => n7008);
   U14494 : INV_X1 port map( A => Plaintext(66), ZN => n7009);
   U14495 : INV_X1 port map( A => n7846, ZN => n7843);
   U14497 : NAND2_X1 port map( A1 => n7846, A2 => n8023, ZN => n7520);
   U14498 : INV_X1 port map( A => n7011, ZN => n7685);
   U14500 : INV_X1 port map( A => n7844, ZN => n7517);
   U14501 : INV_X1 port map( A => n8023, ZN => n7684);
   U14505 : INV_X1 port map( A => Plaintext(86), ZN => n7015);
   U14506 : XNOR2_X1 port map( A => n7015, B => Key(86), ZN => n7838);
   U14507 : INV_X1 port map( A => n7838, ZN => n7835);
   U14508 : XNOR2_X1 port map( A => Key(85), B => Plaintext(85), ZN => n7836);
   U14509 : INV_X1 port map( A => Plaintext(88), ZN => n7016);
   U14512 : INV_X1 port map( A => n7690, ZN => n8244);
   U14513 : XNOR2_X1 port map( A => Key(79), B => Plaintext(79), ZN => n7377);
   U14514 : INV_X1 port map( A => n7377, ZN => n8246);
   U14515 : XNOR2_X1 port map( A => Key(81), B => Plaintext(81), ZN => n7017);
   U14516 : NAND2_X1 port map( A1 => n7017, A2 => n7690, ZN => n7816);
   U14517 : INV_X1 port map( A => n7017, ZN => n7691);
   U14518 : NAND2_X1 port map( A1 => n7691, A2 => n7692, ZN => n7018);
   U14519 : NAND3_X1 port map( A1 => n7816, A2 => n7817, A3 => n7018, ZN => 
                           n7021);
   U14520 : XNOR2_X1 port map( A => Key(82), B => Plaintext(82), ZN => n7376);
   U14521 : INV_X1 port map( A => n7376, ZN => n8247);
   U14523 : NAND3_X1 port map( A1 => n8247, A2 => n7690, A3 => n7692, ZN => 
                           n7020);
   U14524 : OAI211_X1 port map( C1 => n7501, C2 => n8246, A => n7021, B => 
                           n7020, ZN => n8877);
   U14525 : INV_X1 port map( A => n8881, ZN => n8709);
   U14526 : INV_X1 port map( A => Plaintext(56), ZN => n7022);
   U14527 : XNOR2_X1 port map( A => Key(58), B => Plaintext(58), ZN => n7508);
   U14528 : NAND2_X1 port map( A1 => n7257, A2 => n7508, ZN => n7258);
   U14530 : INV_X1 port map( A => n7508, ZN => n7729);
   U14532 : OAI21_X1 port map( B1 => n7729, B2 => n7507, A => n7506, ZN => 
                           n7023);
   U14533 : NAND2_X1 port map( A1 => n7024, A2 => n7023, ZN => n7025);
   U14534 : OAI21_X1 port map( B1 => n7258, B2 => n29629, A => n7025, ZN => 
                           n8404);
   U14535 : INV_X1 port map( A => n8404, ZN => n8875);
   U14536 : INV_X1 port map( A => Plaintext(62), ZN => n7026);
   U14538 : INV_X1 port map( A => n7265, ZN => n8030);
   U14539 : INV_X1 port map( A => Plaintext(65), ZN => n7027);
   U14540 : NAND2_X1 port map( A1 => n8030, A2 => n7268, ZN => n7735);
   U14541 : INV_X1 port map( A => Plaintext(64), ZN => n7028);
   U14543 : INV_X1 port map( A => Plaintext(61), ZN => n7029);
   U14545 : INV_X1 port map( A => n8032, ZN => n7267);
   U14546 : INV_X1 port map( A => Plaintext(63), ZN => n7030);
   U14547 : NAND3_X1 port map( A1 => n7521, A2 => n7267, A3 => n7709, ZN => 
                           n7031);
   U14548 : XNOR2_X1 port map( A => Key(60), B => Plaintext(60), ZN => n7737);
   U14549 : INV_X1 port map( A => n7737, ZN => n8028);
   U14550 : NAND3_X1 port map( A1 => n7268, A2 => n7267, A3 => n7709, ZN => 
                           n7032);
   U14551 : OAI21_X1 port map( B1 => n8875, B2 => n8699, A => n8710, ZN => 
                           n7033);
   U14552 : NOR2_X1 port map( A1 => n7033, A2 => n8876, ZN => n7034);
   U14553 : XNOR2_X1 port map( A => n9732, B => n10297, ZN => n10343);
   U14554 : INV_X1 port map( A => Plaintext(153), ZN => n7036);
   U14555 : XNOR2_X1 port map( A => n7036, B => Key(153), ZN => n7040);
   U14556 : INV_X1 port map( A => Plaintext(150), ZN => n7037);
   U14557 : NAND2_X1 port map( A1 => n7982, A2 => n7456, ZN => n7194);
   U14558 : INV_X1 port map( A => Plaintext(154), ZN => n7038);
   U14559 : INV_X1 port map( A => Plaintext(155), ZN => n7039);
   U14560 : XNOR2_X1 port map( A => n7039, B => Key(155), ZN => n7192);
   U14561 : NAND2_X1 port map( A1 => n7641, A2 => n7985, ZN => n7041);
   U14562 : INV_X1 port map( A => n7040, ZN => n7643);
   U14563 : AOI21_X1 port map( B1 => n7194, B2 => n7041, A => n7643, ZN => 
                           n7044);
   U14564 : INV_X1 port map( A => Plaintext(152), ZN => n7042);
   U14565 : XNOR2_X1 port map( A => n7042, B => Key(152), ZN => n7191);
   U14566 : INV_X1 port map( A => Plaintext(151), ZN => n7043);
   U14567 : INV_X1 port map( A => Plaintext(157), ZN => n7045);
   U14569 : NAND2_X1 port map( A1 => n7965, A2 => n7675, ZN => n7188);
   U14570 : INV_X1 port map( A => Plaintext(161), ZN => n7047);
   U14571 : INV_X1 port map( A => Plaintext(160), ZN => n7048);
   U14572 : XNOR2_X1 port map( A => n7048, B => Key(160), ZN => n7966);
   U14573 : INV_X1 port map( A => n7965, ZN => n7968);
   U14574 : INV_X1 port map( A => n8809, ZN => n8523);
   U14575 : XNOR2_X1 port map( A => Key(170), B => Plaintext(170), ZN => n7589)
                           ;
   U14576 : INV_X1 port map( A => Plaintext(173), ZN => n7050);
   U14577 : XNOR2_X1 port map( A => n7050, B => Key(173), ZN => n7233);
   U14578 : INV_X1 port map( A => Plaintext(172), ZN => n7051);
   U14579 : XNOR2_X1 port map( A => n7051, B => Key(172), ZN => n7958);
   U14580 : INV_X1 port map( A => n7958, ZN => n7872);
   U14582 : NAND2_X1 port map( A1 => n7869, A2 => n441, ZN => n7053);
   U14583 : INV_X1 port map( A => Plaintext(171), ZN => n7052);
   U14584 : INV_X1 port map( A => n7592, ZN => n7873);
   U14585 : OAI211_X2 port map( C1 => n7875, C2 => n7872, A => n7055, B => 
                           n7054, ZN => n8810);
   U14586 : MUX2_X1 port map( A => n8808, B => n8523, S => n8810, Z => n7081);
   U14587 : INV_X1 port map( A => Plaintext(165), ZN => n7056);
   U14588 : INV_X1 port map( A => n7241, ZN => n7060);
   U14589 : INV_X1 port map( A => Plaintext(166), ZN => n7057);
   U14591 : INV_X1 port map( A => n7999, ZN => n7649);
   U14592 : OAI21_X1 port map( B1 => n7060, B2 => n7059, A => n8002, ZN => 
                           n7066);
   U14593 : INV_X1 port map( A => Plaintext(163), ZN => n7061);
   U14595 : NAND2_X1 port map( A1 => n7995, A2 => n7993, ZN => n7652);
   U14596 : INV_X1 port map( A => n7652, ZN => n7064);
   U14597 : INV_X1 port map( A => Plaintext(162), ZN => n7062);
   U14599 : INV_X1 port map( A => n7992, ZN => n7994);
   U14600 : NOR2_X1 port map( A1 => n7993, A2 => n7994, ZN => n7063);
   U14601 : OAI21_X1 port map( B1 => n7064, B2 => n7063, A => n29081, ZN => 
                           n7065);
   U14602 : INV_X1 port map( A => Plaintext(176), ZN => n7067);
   U14603 : XNOR2_X1 port map( A => n7067, B => Key(176), ZN => n7069);
   U14604 : NAND2_X1 port map( A1 => n7582, A2 => n7071, ZN => n7237);
   U14605 : INV_X1 port map( A => Plaintext(175), ZN => n7068);
   U14606 : INV_X1 port map( A => n7069, ZN => n7583);
   U14607 : INV_X1 port map( A => Plaintext(177), ZN => n7070);
   U14608 : XNOR2_X1 port map( A => n7070, B => Key(177), ZN => n7072);
   U14610 : INV_X1 port map( A => n7071, ZN => n7884);
   U14611 : INV_X1 port map( A => Plaintext(179), ZN => n7073);
   U14612 : XNOR2_X1 port map( A => Key(178), B => Plaintext(178), ZN => n7082)
                           ;
   U14613 : INV_X1 port map( A => n7082, ZN => n7581);
   U14614 : NAND3_X1 port map( A1 => n7581, A2 => n7585, A3 => n7583, ZN => 
                           n7075);
   U14615 : OAI211_X1 port map( C1 => n7237, C2 => n7584, A => n7076, B => 
                           n7075, ZN => n8811);
   U14616 : INV_X1 port map( A => n8811, ZN => n8680);
   U14617 : OAI21_X1 port map( B1 => n29241, B2 => n8810, A => n8679, ZN => 
                           n7080);
   U14618 : INV_X1 port map( A => n7172, ZN => n7310);
   U14619 : XNOR2_X1 port map( A => Key(181), B => Plaintext(181), ZN => n7308)
                           ;
   U14620 : INV_X1 port map( A => n7308, ZN => n7862);
   U14621 : XNOR2_X1 port map( A => Key(180), B => Plaintext(180), ZN => n7865)
                           ;
   U14622 : AOI21_X1 port map( B1 => n7310, B2 => n7862, A => n7865, ZN => 
                           n7079);
   U14623 : INV_X1 port map( A => Plaintext(185), ZN => n7077);
   U14626 : XNOR2_X1 port map( A => Key(184), B => Plaintext(184), ZN => n7867)
                           ;
   U14627 : NAND2_X1 port map( A1 => n7095, A2 => n5149, ZN => n7078);
   U14628 : OAI21_X1 port map( B1 => n7883, B2 => n7585, A => n7083, ZN => 
                           n7084);
   U14629 : INV_X1 port map( A => Plaintext(4), ZN => n7085);
   U14630 : INV_X1 port map( A => Plaintext(3), ZN => n7086);
   U14631 : INV_X1 port map( A => n7315, ZN => n7774);
   U14632 : INV_X1 port map( A => Plaintext(5), ZN => n7087);
   U14634 : NAND2_X1 port map( A1 => n7090, A2 => n1350, ZN => n7091);
   U14635 : INV_X1 port map( A => n7092, ZN => n7601);
   U14636 : INV_X1 port map( A => n7093, ZN => n7864);
   U14637 : NAND2_X1 port map( A1 => n7864, A2 => n7867, ZN => n7094);
   U14638 : NAND2_X1 port map( A1 => n8586, A2 => n8192, ZN => n7102);
   U14639 : XNOR2_X1 port map( A => Key(12), B => Plaintext(12), ZN => n7100);
   U14640 : INV_X1 port map( A => n7100, ZN => n7289);
   U14641 : INV_X1 port map( A => Plaintext(13), ZN => n7096);
   U14642 : XNOR2_X1 port map( A => n7096, B => Key(13), ZN => n8173);
   U14643 : INV_X1 port map( A => Plaintext(14), ZN => n7097);
   U14644 : XNOR2_X1 port map( A => n7097, B => Key(14), ZN => n7101);
   U14645 : INV_X1 port map( A => n7101, ZN => n7758);
   U14646 : INV_X1 port map( A => Plaintext(17), ZN => n7098);
   U14647 : NAND2_X1 port map( A1 => n7758, A2 => n7759, ZN => n7763);
   U14648 : INV_X1 port map( A => Plaintext(16), ZN => n7099);
   U14649 : XNOR2_X1 port map( A => n7099, B => Key(16), ZN => n8176);
   U14650 : NAND2_X1 port map( A1 => n7102, A2 => n8824, ZN => n7120);
   U14651 : INV_X1 port map( A => Plaintext(187), ZN => n7103);
   U14653 : INV_X1 port map( A => Plaintext(189), ZN => n7104);
   U14654 : XNOR2_X1 port map( A => n7104, B => Key(189), ZN => n7106);
   U14655 : NAND2_X1 port map( A1 => n7801, A2 => n7895, ZN => n7597);
   U14656 : INV_X1 port map( A => Plaintext(186), ZN => n7105);
   U14657 : INV_X1 port map( A => n7106, ZN => n7800);
   U14658 : NAND2_X1 port map( A1 => n7312, A2 => n7800, ZN => n7107);
   U14659 : XNOR2_X1 port map( A => Key(191), B => Plaintext(191), ZN => n7110)
                           ;
   U14660 : AOI21_X1 port map( B1 => n7597, B2 => n7107, A => n7898, ZN => 
                           n7113);
   U14661 : INV_X1 port map( A => Plaintext(188), ZN => n7108);
   U14662 : INV_X1 port map( A => Plaintext(190), ZN => n7109);
   U14663 : NAND2_X1 port map( A1 => n7900, A2 => n7897, ZN => n7313);
   U14664 : INV_X1 port map( A => n7900, ZN => n7896);
   U14665 : INV_X1 port map( A => n7110, ZN => n7176);
   U14668 : INV_X1 port map( A => n8826, ZN => n8830);
   U14669 : INV_X1 port map( A => Plaintext(6), ZN => n7115);
   U14671 : XNOR2_X1 port map( A => Key(7), B => Plaintext(7), ZN => n7162);
   U14672 : INV_X1 port map( A => Plaintext(8), ZN => n7117);
   U14674 : OAI21_X1 port map( B1 => n7164, B2 => n7342, A => n7770, ZN => 
                           n7118);
   U14675 : NAND2_X1 port map( A1 => n7447, A2 => n8826, ZN => n7119);
   U14676 : INV_X1 port map( A => n9799, ZN => n7121);
   U14677 : XNOR2_X1 port map( A => n7121, B => n10037, ZN => n8953);
   U14678 : XNOR2_X1 port map( A => n8953, B => n10343, ZN => n7230);
   U14679 : XNOR2_X1 port map( A => Key(37), B => Plaintext(37), ZN => n7722);
   U14680 : INV_X1 port map( A => n7722, ZN => n8139);
   U14681 : XNOR2_X1 port map( A => Key(36), B => Plaintext(36), ZN => n8138);
   U14682 : INV_X1 port map( A => n8138, ZN => n8041);
   U14683 : XNOR2_X1 port map( A => Key(39), B => Plaintext(39), ZN => n7560);
   U14685 : INV_X1 port map( A => Plaintext(38), ZN => n7122);
   U14686 : INV_X1 port map( A => Plaintext(40), ZN => n7123);
   U14688 : NAND2_X1 port map( A1 => n8141, A2 => n8143, ZN => n7562);
   U14690 : INV_X1 port map( A => n8141, ZN => n8142);
   U14691 : MUX2_X2 port map( A => n7125, B => n7124, S => n7336, Z => n9245);
   U14693 : INV_X1 port map( A => n8048, ZN => n8134);
   U14694 : XNOR2_X1 port map( A => Key(45), B => Plaintext(45), ZN => n8047);
   U14695 : INV_X1 port map( A => n8047, ZN => n8135);
   U14696 : INV_X1 port map( A => Plaintext(42), ZN => n7126);
   U14697 : XNOR2_X1 port map( A => n7126, B => Key(42), ZN => n7554);
   U14698 : INV_X1 port map( A => Plaintext(46), ZN => n7128);
   U14700 : NAND2_X1 port map( A1 => n7127, A2 => n8131, ZN => n7717);
   U14701 : NAND2_X1 port map( A1 => n8134, A2 => n29119, ZN => n7130);
   U14702 : AOI21_X1 port map( B1 => n7717, B2 => n7130, A => n8049, ZN => 
                           n7131);
   U14703 : INV_X1 port map( A => n9041, ZN => n9248);
   U14704 : NAND2_X1 port map( A1 => n7257, A2 => n7514, ZN => n7733);
   U14705 : OAI21_X1 port map( B1 => n8039, B2 => n7257, A => n7733, ZN => 
                           n7135);
   U14706 : INV_X1 port map( A => n7514, ZN => n7728);
   U14707 : AOI21_X1 port map( B1 => n7133, B2 => n7132, A => n7507, ZN => 
                           n7134);
   U14708 : INV_X1 port map( A => Plaintext(51), ZN => n7136);
   U14709 : AND2_X1 port map( A1 => n7744, A2 => n28161, ZN => n7146);
   U14710 : INV_X1 port map( A => Plaintext(53), ZN => n7137);
   U14711 : INV_X1 port map( A => Plaintext(48), ZN => n7138);
   U14712 : OAI21_X1 port map( B1 => n8014, B2 => n7744, A => n8013, ZN => 
                           n7145);
   U14713 : INV_X1 port map( A => Plaintext(52), ZN => n7139);
   U14715 : INV_X1 port map( A => n8014, ZN => n7746);
   U14716 : INV_X1 port map( A => Plaintext(49), ZN => n7140);
   U14717 : INV_X1 port map( A => n7743, ZN => n7745);
   U14718 : INV_X1 port map( A => n8013, ZN => n7747);
   U14719 : NAND2_X1 port map( A1 => n7745, A2 => n7747, ZN => n7142);
   U14720 : INV_X1 port map( A => n7141, ZN => n7523);
   U14722 : INV_X1 port map( A => n8693, ZN => n9039);
   U14723 : NOR2_X1 port map( A1 => n9410, A2 => n9039, ZN => n7160);
   U14724 : XNOR2_X1 port map( A => Key(27), B => Plaintext(27), ZN => n7150);
   U14725 : INV_X1 port map( A => Plaintext(26), ZN => n7147);
   U14726 : XNOR2_X1 port map( A => n7147, B => Key(26), ZN => n7283);
   U14727 : MUX2_X1 port map( A => n7541, B => n8150, S => n8151, Z => n7152);
   U14728 : INV_X1 port map( A => Plaintext(29), ZN => n7148);
   U14729 : XNOR2_X1 port map( A => n7148, B => Key(29), ZN => n7285);
   U14730 : INV_X1 port map( A => n7285, ZN => n8148);
   U14731 : INV_X1 port map( A => Plaintext(24), ZN => n7149);
   U14732 : INV_X1 port map( A => n7150, ZN => n8147);
   U14733 : INV_X1 port map( A => Plaintext(31), ZN => n7153);
   U14735 : INV_X1 port map( A => Plaintext(30), ZN => n7154);
   U14736 : NAND2_X1 port map( A1 => n8165, A2 => n7348, ZN => n7297);
   U14737 : INV_X1 port map( A => n8161, ZN => n8159);
   U14738 : INV_X1 port map( A => Plaintext(34), ZN => n7155);
   U14739 : XNOR2_X1 port map( A => n7155, B => Key(34), ZN => n8158);
   U14740 : INV_X1 port map( A => n8158, ZN => n7750);
   U14742 : INV_X1 port map( A => Plaintext(33), ZN => n7156);
   U14743 : XNOR2_X1 port map( A => n7156, B => Key(33), ZN => n7298);
   U14744 : INV_X1 port map( A => n8165, ZN => n8167);
   U14745 : NAND3_X1 port map( A1 => n7157, A2 => n8162, A3 => n8167, ZN => 
                           n7158);
   U14746 : NAND2_X1 port map( A1 => n8166, A2 => n7349, ZN => n7296);
   U14748 : NAND2_X1 port map( A1 => n9041, A2 => n9243, ZN => n8110);
   U14749 : INV_X1 port map( A => n7890, ZN => n7778);
   U14750 : INV_X1 port map( A => n7889, ZN => n7777);
   U14751 : INV_X1 port map( A => n7162, ZN => n7321);
   U14752 : INV_X1 port map( A => n7342, ZN => n7163);
   U14753 : INV_X1 port map( A => Plaintext(20), ZN => n7166);
   U14754 : INV_X1 port map( A => n7291, ZN => n7781);
   U14755 : NAND2_X1 port map( A1 => n7781, A2 => n7330, ZN => n7168);
   U14756 : XNOR2_X1 port map( A => Key(19), B => Plaintext(19), ZN => n7787);
   U14757 : XNOR2_X1 port map( A => Key(18), B => Plaintext(18), ZN => n7786);
   U14758 : XNOR2_X1 port map( A => Key(22), B => Plaintext(22), ZN => n7550);
   U14759 : INV_X1 port map( A => n7550, ZN => n7785);
   U14760 : XNOR2_X1 port map( A => Key(21), B => Plaintext(21), ZN => n7292);
   U14761 : INV_X1 port map( A => n7292, ZN => n7782);
   U14762 : INV_X1 port map( A => n7787, ZN => n7331);
   U14763 : AOI21_X1 port map( B1 => n7782, B2 => n7331, A => n7786, ZN => 
                           n7169);
   U14764 : OR2_X1 port map( A1 => n7169, A2 => n7781, ZN => n7170);
   U14765 : NAND2_X2 port map( A1 => n7171, A2 => n7170, ZN => n8381);
   U14766 : INV_X1 port map( A => n8381, ZN => n8536);
   U14767 : NAND2_X1 port map( A1 => n7862, A2 => n7172, ZN => n7173);
   U14768 : INV_X1 port map( A => n7865, ZN => n7174);
   U14769 : NAND2_X1 port map( A1 => n7310, A2 => n7174, ZN => n7604);
   U14770 : NAND2_X1 port map( A1 => n7801, A2 => n7312, ZN => n7595);
   U14771 : INV_X1 port map( A => n7595, ZN => n7177);
   U14772 : OAI21_X1 port map( B1 => n7177, B2 => n7176, A => n7803, ZN => 
                           n7179);
   U14773 : INV_X1 port map( A => n7801, ZN => n7902);
   U14774 : OAI211_X1 port map( C1 => n7897, C2 => n7176, A => n7800, B => 
                           n7902, ZN => n7178);
   U14775 : AND2_X1 port map( A1 => n7179, A2 => n7178, ZN => n8729);
   U14776 : NAND3_X1 port map( A1 => n8537, A2 => n8729, A3 => n8381, ZN => 
                           n7185);
   U14777 : NAND2_X1 port map( A1 => n7289, A2 => n8177, ZN => n8175);
   U14778 : NAND3_X1 port map( A1 => n8175, A2 => n8179, A3 => n7289, ZN => 
                           n7183);
   U14779 : NAND3_X1 port map( A1 => n8175, A2 => n8179, A3 => n613, ZN => 
                           n7181);
   U14780 : NOR2_X1 port map( A1 => n8381, A2 => n8733, ZN => n8538);
   U14781 : NAND2_X1 port map( A1 => n8538, A2 => n8739, ZN => n7184);
   U14782 : XNOR2_X1 port map( A => n10346, B => n9542, ZN => n10169);
   U14783 : AOI21_X1 port map( B1 => n7188, B2 => n7962, A => n4696, ZN => 
                           n7190);
   U14784 : NAND2_X1 port map( A1 => n7965, A2 => n1938, ZN => n7236);
   U14785 : AOI21_X1 port map( B1 => n7236, B2 => n7675, A => n29302, ZN => 
                           n7189);
   U14787 : INV_X1 port map( A => n7191, ZN => n7980);
   U14789 : INV_X1 port map( A => n7981, ZN => n7243);
   U14790 : OAI211_X1 port map( C1 => n7456, C2 => n7243, A => n7194, B => 
                           n7642, ZN => n7195);
   U14791 : INV_X1 port map( A => n8685, ZN => n8688);
   U14792 : XNOR2_X1 port map( A => Key(139), B => Plaintext(139), ZN => n7480)
                           ;
   U14793 : INV_X1 port map( A => n7480, ZN => n8284);
   U14794 : INV_X1 port map( A => Plaintext(141), ZN => n7196);
   U14795 : XNOR2_X1 port map( A => n7196, B => Key(141), ZN => n7405);
   U14796 : INV_X1 port map( A => n7405, ZN => n7975);
   U14799 : OAI21_X1 port map( B1 => n8284, B2 => n7975, A => n7477, ZN => 
                           n7217);
   U14800 : INV_X1 port map( A => Plaintext(140), ZN => n7197);
   U14801 : XNOR2_X1 port map( A => n7197, B => Key(140), ZN => n7198);
   U14803 : NAND2_X1 port map( A1 => n8281, A2 => n7975, ZN => n8279);
   U14804 : NAND2_X1 port map( A1 => n7199, A2 => n8279, ZN => n7214);
   U14805 : INV_X1 port map( A => Plaintext(143), ZN => n7200);
   U14806 : XNOR2_X1 port map( A => n7200, B => Key(143), ZN => n7404);
   U14807 : INV_X1 port map( A => Plaintext(132), ZN => n7201);
   U14808 : XNOR2_X1 port map( A => n7201, B => Key(132), ZN => n7942);
   U14809 : INV_X1 port map( A => Plaintext(133), ZN => n7202);
   U14811 : NAND2_X1 port map( A1 => n7942, A2 => n7657, ZN => n7941);
   U14812 : NAND2_X1 port map( A1 => n7941, A2 => n29317, ZN => n7209);
   U14813 : INV_X1 port map( A => Plaintext(134), ZN => n7203);
   U14815 : NAND2_X1 port map( A1 => n8305, A2 => n8297, ZN => n7208);
   U14816 : INV_X1 port map( A => Plaintext(135), ZN => n7204);
   U14817 : XNOR2_X1 port map( A => n7204, B => Key(135), ZN => n7399);
   U14818 : INV_X1 port map( A => n7399, ZN => n8301);
   U14819 : INV_X1 port map( A => n7657, ZN => n8303);
   U14820 : INV_X1 port map( A => Plaintext(136), ZN => n7205);
   U14821 : INV_X1 port map( A => n7655, ZN => n7939);
   U14822 : NAND2_X1 port map( A1 => n7939, A2 => n29317, ZN => n7206);
   U14823 : INV_X1 port map( A => n8525, ZN => n9222);
   U14824 : XNOR2_X1 port map( A => Key(148), B => Plaintext(148), ZN => n8267)
                           ;
   U14825 : XNOR2_X1 port map( A => Key(145), B => Plaintext(145), ZN => n7485)
                           ;
   U14826 : INV_X1 port map( A => n7485, ZN => n8271);
   U14827 : XNOR2_X1 port map( A => Key(149), B => Plaintext(149), ZN => n7488)
                           ;
   U14828 : INV_X1 port map( A => Plaintext(144), ZN => n7212);
   U14829 : XNOR2_X1 port map( A => n7212, B => Key(144), ZN => n7665);
   U14830 : INV_X1 port map( A => n7665, ZN => n8268);
   U14831 : INV_X1 port map( A => n9221, ZN => n8686);
   U14832 : NAND2_X1 port map( A1 => n8098, A2 => n8687, ZN => n7227);
   U14833 : INV_X1 port map( A => n7214, ZN => n7215);
   U14834 : INV_X1 port map( A => Plaintext(130), ZN => n7218);
   U14836 : INV_X1 port map( A => Plaintext(128), ZN => n7219);
   U14837 : NAND2_X1 port map( A1 => n29590, A2 => n8256, ZN => n8259);
   U14838 : INV_X1 port map( A => Plaintext(129), ZN => n7220);
   U14839 : NAND2_X1 port map( A1 => n6782, A2 => n28617, ZN => n7221);
   U14840 : NAND2_X1 port map( A1 => n8259, A2 => n7221, ZN => n7224);
   U14841 : XNOR2_X2 port map( A => Key(131), B => Plaintext(131), ZN => n8258)
                           ;
   U14842 : INV_X1 port map( A => n8258, ZN => n7465);
   U14844 : INV_X1 port map( A => n8263, ZN => n7463);
   U14845 : OAI21_X1 port map( B1 => n6782, B2 => n7618, A => n7463, ZN => 
                           n7223);
   U14846 : XNOR2_X1 port map( A => Key(126), B => Plaintext(126), ZN => n7466)
                           ;
   U14847 : NAND2_X1 port map( A1 => n28618, A2 => n7946, ZN => n7222);
   U14849 : OAI21_X1 port map( B1 => n9220, B2 => n8686, A => n8687, ZN => 
                           n7225);
   U14850 : XNOR2_X1 port map( A => n9971, B => n26214, ZN => n7228);
   U14851 : XNOR2_X1 port map( A => n10169, B => n7228, ZN => n7229);
   U14852 : NOR2_X1 port map( A1 => n7591, A2 => n7870, ZN => n7232);
   U14853 : OAI21_X1 port map( B1 => n7592, B2 => n7872, A => n7960, ZN => 
                           n7235);
   U14854 : INV_X1 port map( A => n7594, ZN => n7234);
   U14855 : NAND2_X1 port map( A1 => n7887, A2 => n7583, ZN => n7305);
   U14856 : NAND2_X1 port map( A1 => n7581, A2 => n7884, ZN => n7238);
   U14857 : NAND2_X1 port map( A1 => n7999, A2 => n7876, ZN => n7877);
   U14858 : INV_X1 port map( A => n7877, ZN => n7240);
   U14859 : INV_X1 port map( A => n7995, ZN => n7879);
   U14860 : AOI21_X1 port map( B1 => n7998, B2 => n7879, A => n6615, ZN => 
                           n7239);
   U14861 : OAI21_X1 port map( B1 => n7240, B2 => n7998, A => n7239, ZN => 
                           n7242);
   U14863 : NAND2_X1 port map( A1 => n7644, A2 => n7457, ZN => n7244);
   U14865 : NAND2_X1 port map( A1 => n7485, A2 => n8269, ZN => n7990);
   U14866 : INV_X1 port map( A => n7488, ZN => n7986);
   U14867 : NOR2_X1 port map( A1 => n29639, A2 => n8264, ZN => n7245);
   U14868 : NAND2_X1 port map( A1 => n8270, A2 => n8267, ZN => n8266);
   U14869 : OAI21_X1 port map( B1 => n7662, B2 => n7245, A => n8266, ZN => 
                           n7246);
   U14871 : NAND2_X1 port map( A1 => n8134, A2 => n8047, ZN => n7248);
   U14872 : OAI21_X1 port map( B1 => n8049, B2 => n615, A => n8133, ZN => n7249
                           );
   U14873 : NAND2_X1 port map( A1 => n7251, A2 => n3594, ZN => n7253);
   U14874 : NAND2_X1 port map( A1 => n7251, A2 => n3639, ZN => n7252);
   U14875 : NAND3_X1 port map( A1 => n7253, A2 => n7252, A3 => n7708, ZN => 
                           n7256);
   U14876 : INV_X1 port map( A => n7851, ZN => n7853);
   U14877 : NAND2_X1 port map( A1 => n7256, A2 => n7255, ZN => n8763);
   U14878 : INV_X1 port map( A => n7257, ZN => n8038);
   U14879 : INV_X1 port map( A => n29629, ZN => n7511);
   U14880 : NAND2_X1 port map( A1 => n8763, A2 => n9562, ZN => n9565);
   U14883 : NAND2_X1 port map( A1 => n7260, A2 => n29106, ZN => n7264);
   U14884 : INV_X1 port map( A => n8024, ZN => n7515);
   U14885 : NAND3_X1 port map( A1 => n7847, A2 => n7684, A3 => n7261, ZN => 
                           n7263);
   U14886 : NAND3_X1 port map( A1 => n7517, A2 => n7685, A3 => n29130, ZN => 
                           n7262);
   U14888 : INV_X1 port map( A => n8944, ZN => n10401);
   U14889 : NAND3_X1 port map( A1 => n7268, A2 => n8032, A3 => n8030, ZN => 
                           n7272);
   U14890 : NAND3_X1 port map( A1 => n7268, A2 => n7265, A3 => n7521, ZN => 
                           n7271);
   U14891 : NAND3_X1 port map( A1 => n7266, A2 => n7267, A3 => n8030, ZN => 
                           n7270);
   U14892 : NAND3_X1 port map( A1 => n618, A2 => n7709, A3 => n7737, ZN => 
                           n7269);
   U14893 : AOI21_X2 port map( B1 => n8947, B2 => n10401, A => n7274, ZN => 
                           n10191);
   U14894 : INV_X1 port map( A => n7891, ZN => n7773);
   U14895 : MUX2_X1 port map( A => n7275, B => n7889, S => n7315, Z => n7276);
   U14896 : NAND2_X1 port map( A1 => n7770, A2 => n7342, ZN => n7278);
   U14897 : NAND2_X1 port map( A1 => n7279, A2 => n7278, ZN => n7280);
   U14898 : NAND2_X1 port map( A1 => n8334, A2 => n8889, ZN => n8079);
   U14899 : NAND2_X1 port map( A1 => n8147, A2 => n7793, ZN => n7282);
   U14900 : INV_X1 port map( A => n8151, ZN => n7284);
   U14901 : AOI21_X1 port map( B1 => n7284, B2 => n8148, A => n7542, ZN => 
                           n7287);
   U14903 : NAND2_X1 port map( A1 => n8177, A2 => n7758, ZN => n7288);
   U14904 : INV_X1 port map( A => n8177, ZN => n7760);
   U14905 : NAND2_X1 port map( A1 => n7330, A2 => n7291, ZN => n8154);
   U14906 : NAND2_X1 port map( A1 => n1899, A2 => n7787, ZN => n8156);
   U14908 : INV_X1 port map( A => n7330, ZN => n8153);
   U14909 : NAND3_X1 port map( A1 => n1899, A2 => n8153, A3 => n7786, ZN => 
                           n7294);
   U14910 : AOI21_X1 port map( B1 => n7297, B2 => n7296, A => n7750, ZN => 
                           n7300);
   U14911 : NAND2_X1 port map( A1 => n8165, A2 => n7298, ZN => n7535);
   U14912 : AOI21_X1 port map( B1 => n7535, B2 => n7348, A => n7349, ZN => 
                           n7299);
   U14913 : OR2_X2 port map( A1 => n7300, A2 => n7299, ZN => n8009);
   U14914 : NAND3_X1 port map( A1 => n8891, A2 => n8009, A3 => n8335, ZN => 
                           n7301);
   U14915 : OAI211_X1 port map( C1 => n8079, C2 => n8887, A => n7302, B => 
                           n7301, ZN => n9795);
   U14916 : INV_X1 port map( A => n9795, ZN => n9266);
   U14917 : NAND2_X1 port map( A1 => n7172, A2 => n7865, ZN => n7306);
   U14918 : NAND3_X1 port map( A1 => n7310, A2 => n7309, A3 => n7308, ZN => 
                           n7311);
   U14920 : NAND2_X1 port map( A1 => n7315, A2 => n7777, ZN => n7317);
   U14921 : NAND2_X1 port map( A1 => n29112, A2 => n7089, ZN => n7316);
   U14922 : OAI21_X1 port map( B1 => n7594, B2 => n7872, A => n7318, ZN => 
                           n7319);
   U14923 : AOI22_X1 port map( A1 => n9425, A2 => n7569, B1 => n8574, B2 => 
                           n8327, ZN => n7328);
   U14924 : AOI21_X1 port map( B1 => n7323, B2 => n7322, A => n7342, ZN => 
                           n7324);
   U14925 : NAND2_X1 port map( A1 => n8327, A2 => n9425, ZN => n7326);
   U14926 : NAND2_X1 port map( A1 => n8580, A2 => n7326, ZN => n7327);
   U14927 : XNOR2_X1 port map( A => n9266, B => n10007, ZN => n9003);
   U14928 : OAI211_X1 port map( C1 => n7781, C2 => n7550, A => n7332, B => 
                           n8153, ZN => n7334);
   U14929 : OAI21_X1 port map( B1 => n7782, B2 => n7786, A => n7330, ZN => 
                           n7333);
   U14930 : NAND2_X1 port map( A1 => n8041, A2 => n8139, ZN => n7725);
   U14931 : INV_X1 port map( A => n7336, ZN => n8043);
   U14932 : INV_X1 port map( A => n8143, ZN => n7721);
   U14933 : NAND2_X1 port map( A1 => n29751, A2 => n8139, ZN => n7337);
   U14934 : AOI21_X1 port map( B1 => n7337, B2 => n8041, A => n8142, ZN => 
                           n7338);
   U14936 : NAND2_X1 port map( A1 => n614, A2 => n7342, ZN => n7341);
   U14937 : NAND2_X1 port map( A1 => n7341, A2 => n7767, ZN => n7344);
   U14938 : NOR2_X1 port map( A1 => n5242, A2 => n7342, ZN => n7343);
   U14939 : NAND3_X1 port map( A1 => n7345, A2 => n613, A3 => n7760, ZN => 
                           n7346);
   U14940 : NAND2_X1 port map( A1 => n8563, A2 => n8185, ZN => n8939);
   U14941 : INV_X1 port map( A => n7348, ZN => n8160);
   U14942 : OAI21_X1 port map( B1 => n8162, B2 => n8160, A => n8159, ZN => 
                           n7351);
   U14943 : OAI21_X1 port map( B1 => n8168, B2 => n7750, A => n8161, ZN => 
                           n7350);
   U14944 : NAND2_X1 port map( A1 => n8167, A2 => n8160, ZN => n7352);
   U14945 : AOI21_X1 port map( B1 => n8937, B2 => n8939, A => n9140, ZN => 
                           n7356);
   U14946 : OAI21_X1 port map( B1 => n8148, B2 => n28149, A => n7542, ZN => 
                           n7353);
   U14947 : NAND2_X1 port map( A1 => n9139, A2 => n8185, ZN => n8330);
   U14948 : AOI21_X1 port map( B1 => n8330, B2 => n8563, A => n8562, ZN => 
                           n7355);
   U14949 : MUX2_X1 port map( A => n7357, B => n8232, S => n29110, Z => n7361);
   U14950 : INV_X1 port map( A => n8237, ZN => n7919);
   U14951 : INV_X1 port map( A => n8232, ZN => n8236);
   U14952 : INV_X1 port map( A => n7358, ZN => n7920);
   U14955 : NAND2_X1 port map( A1 => n7635, A2 => n7828, ZN => n7366);
   U14956 : INV_X1 port map( A => n7828, ZN => n8202);
   U14957 : NAND3_X1 port map( A1 => n3431, A2 => n8205, A3 => n7363, ZN => 
                           n7364);
   U14958 : OAI211_X1 port map( C1 => n7366, C2 => n8205, A => n7365, B => 
                           n7364, ZN => n9149);
   U14959 : INV_X1 port map( A => n7837, ZN => n8208);
   U14960 : NAND2_X1 port map( A1 => n7371, A2 => n7825, ZN => n8225);
   U14961 : INV_X1 port map( A => n7371, ZN => n7824);
   U14962 : NAND2_X1 port map( A1 => n7822, A2 => n7824, ZN => n7372);
   U14963 : AOI21_X1 port map( B1 => n8225, B2 => n7372, A => n8221, ZN => 
                           n7375);
   U14964 : NAND3_X1 port map( A1 => n7821, A2 => n7824, A3 => n3821, ZN => 
                           n7373);
   U14965 : NAND2_X1 port map( A1 => n7376, A2 => n7692, ZN => n7378);
   U14966 : NAND3_X1 port map( A1 => n7378, A2 => n8245, A3 => n7818, ZN => 
                           n7381);
   U14967 : NAND2_X1 port map( A1 => n8243, A2 => n7690, ZN => n7380);
   U14968 : NAND3_X1 port map( A1 => n8246, A2 => n7817, A3 => n7692, ZN => 
                           n7379);
   U14969 : INV_X1 port map( A => n7382, ZN => n7705);
   U14970 : NAND3_X1 port map( A1 => n9374, A2 => n9149, A3 => n5958, ZN => 
                           n7386);
   U14971 : XNOR2_X1 port map( A => n10364, B => n10193, ZN => n9094);
   U14972 : NAND2_X1 port map( A1 => n8263, A2 => n7618, ZN => n8260);
   U14973 : NAND3_X1 port map( A1 => n7463, A2 => n8258, A3 => n7946, ZN => 
                           n7388);
   U14974 : NAND2_X1 port map( A1 => n6782, A2 => n28615, ZN => n7390);
   U14975 : AOI21_X1 port map( B1 => n7390, B2 => n7389, A => n8258, ZN => 
                           n7391);
   U14977 : INV_X1 port map( A => n7393, ZN => n8311);
   U14978 : NAND2_X1 port map( A1 => n7613, A2 => n8311, ZN => n7427);
   U14979 : AND2_X1 port map( A1 => n7393, A2 => n7614, ZN => n7610);
   U14980 : NAND2_X1 port map( A1 => n7933, A2 => n29135, ZN => n7394);
   U14981 : NAND2_X1 port map( A1 => n7610, A2 => n7394, ZN => n7395);
   U14982 : OAI211_X2 port map( C1 => n28810, C2 => n7427, A => n7395, B => 
                           n7609, ZN => n9340);
   U14983 : NAND2_X1 port map( A1 => n9132, A2 => n9340, ZN => n8340);
   U14984 : INV_X1 port map( A => n8340, ZN => n7397);
   U14985 : INV_X1 port map( A => n7911, ZN => n7916);
   U14986 : AOI21_X1 port map( B1 => n7628, B2 => n7916, A => n8290, ZN => 
                           n7396);
   U14987 : NAND2_X1 port map( A1 => n7924, A2 => n7626, ZN => n7926);
   U14988 : NAND2_X1 port map( A1 => n8216, A2 => n8213, ZN => n7398);
   U14989 : INV_X1 port map( A => n8213, ZN => n7438);
   U14990 : INV_X1 port map( A => n7942, ZN => n8302);
   U14991 : INV_X1 port map( A => n7400, ZN => n8296);
   U14992 : NAND3_X1 port map( A1 => n7655, A2 => n8296, A3 => n29317, ZN => 
                           n7401);
   U14993 : NAND2_X1 port map( A1 => n7403, A2 => n9134, ZN => n7413);
   U14994 : NAND2_X1 port map( A1 => n8342, A2 => n9134, ZN => n8549);
   U14995 : NAND2_X1 port map( A1 => n7976, A2 => n8281, ZN => n7671);
   U14996 : NAND2_X1 port map( A1 => n7406, A2 => n8275, ZN => n8285);
   U14997 : OAI21_X1 port map( B1 => n7671, B2 => n8280, A => n8285, ZN => 
                           n7409);
   U14998 : NAND2_X1 port map( A1 => n7406, A2 => n8276, ZN => n7408);
   U14999 : INV_X1 port map( A => n9133, ZN => n7410);
   U15000 : INV_X1 port map( A => n29247, ZN => n27952);
   U15001 : NOR2_X1 port map( A1 => n8608, A2 => n9533, ZN => n7416);
   U15002 : NAND3_X1 port map( A1 => n29662, A2 => n8749, A3 => n9533, ZN => 
                           n7417);
   U15003 : OAI21_X1 port map( B1 => n370, B2 => n8208, A => n7839, ZN => n7421
                           );
   U15004 : NAND3_X1 port map( A1 => n619, A2 => n7840, A3 => n8208, ZN => 
                           n7422);
   U15005 : INV_X1 port map( A => n8741, ZN => n9074);
   U15006 : AND2_X1 port map( A1 => n7827, A2 => n7695, ZN => n7425);
   U15007 : INV_X1 port map( A => n8740, ZN => n8378);
   U15008 : AOI21_X1 port map( B1 => n7427, B2 => n7609, A => n7933, ZN => 
                           n7429);
   U15009 : AOI21_X1 port map( B1 => n7930, B2 => n7613, A => n7935, ZN => 
                           n7428);
   U15012 : NOR2_X1 port map( A1 => n9073, A2 => n8740, ZN => n8855);
   U15013 : NAND2_X1 port map( A1 => n7634, A2 => n7635, ZN => n7829);
   U15014 : NAND2_X1 port map( A1 => n7635, A2 => n7363, ZN => n7433);
   U15015 : AOI21_X1 port map( B1 => n8200, B2 => n7433, A => n7830, ZN => 
                           n7434);
   U15016 : INV_X1 port map( A => n9070, ZN => n8856);
   U15017 : OAI21_X1 port map( B1 => n8855, B2 => n8856, A => n9075, ZN => 
                           n7443);
   U15018 : NAND2_X1 port map( A1 => n8217, A2 => n627, ZN => n7441);
   U15019 : NAND3_X1 port map( A1 => n7441, A2 => n7437, A3 => n7436, ZN => 
                           n7440);
   U15020 : NAND3_X1 port map( A1 => n7438, A2 => n8216, A3 => n7925, ZN => 
                           n7439);
   U15021 : OAI211_X1 port map( C1 => n7441, C2 => n7925, A => n7440, B => 
                           n7439, ZN => n8857);
   U15022 : NAND2_X1 port map( A1 => n8855, A2 => n8857, ZN => n7442);
   U15023 : XNOR2_X1 port map( A => n9996, B => n9754, ZN => n7449);
   U15024 : NAND2_X1 port map( A1 => n8824, A2 => n8826, ZN => n7444);
   U15025 : OAI21_X1 port map( B1 => n7445, B2 => n8824, A => n7444, ZN => 
                           n7446);
   U15026 : OAI21_X1 port map( B1 => n7447, B2 => n8196, A => n7446, ZN => 
                           n9447);
   U15027 : XNOR2_X1 port map( A => n9447, B => n3212, ZN => n7448);
   U15028 : XNOR2_X1 port map( A => n7449, B => n7448, ZN => n7573);
   U15029 : NAND2_X1 port map( A1 => n7399, A2 => n7657, ZN => n7943);
   U15030 : NAND2_X1 port map( A1 => n8305, A2 => n7655, ZN => n7452);
   U15031 : NAND2_X1 port map( A1 => n8296, A2 => n8304, ZN => n7451);
   U15034 : NAND2_X1 port map( A1 => n7456, A2 => n7981, ZN => n7458);
   U15035 : AOI21_X1 port map( B1 => n7459, B2 => n7458, A => n7457, ZN => 
                           n7460);
   U15036 : NAND2_X1 port map( A1 => n29590, A2 => n8258, ZN => n7464);
   U15038 : INV_X1 port map( A => n28614, ZN => n7948);
   U15039 : INV_X1 port map( A => n7466, ZN => n8257);
   U15040 : INV_X1 port map( A => n7618, ZN => n7947);
   U15042 : INV_X1 port map( A => n8287, ZN => n7631);
   U15043 : INV_X1 port map( A => n7912, ZN => n7470);
   U15044 : OAI21_X1 port map( B1 => n7631, B2 => n7470, A => n7916, ZN => 
                           n7472);
   U15045 : INV_X1 port map( A => n7628, ZN => n7917);
   U15046 : NAND2_X1 port map( A1 => n29568, A2 => n7917, ZN => n7471);
   U15047 : AND2_X1 port map( A1 => n7472, A2 => n7471, ZN => n7476);
   U15048 : AOI21_X1 port map( B1 => n7474, B2 => n7473, A => n7915, ZN => 
                           n7475);
   U15050 : OAI21_X1 port map( B1 => n8280, B2 => n8281, A => n7976, ZN => 
                           n7478);
   U15052 : AND2_X1 port map( A1 => n7480, A2 => n7975, ZN => n7670);
   U15053 : INV_X1 port map( A => n7670, ZN => n7481);
   U15054 : INV_X1 port map( A => n9080, ZN => n7484);
   U15055 : NAND3_X1 port map( A1 => n7484, A2 => n8605, A3 => n8603, ZN => 
                           n7492);
   U15056 : OR2_X1 port map( A1 => n9080, A2 => n8726, ZN => n8851);
   U15057 : OAI21_X1 port map( B1 => n341, B2 => n8268, A => n7486, ZN => n7487
                           );
   U15058 : INV_X1 port map( A => n8270, ZN => n7663);
   U15059 : NAND2_X1 port map( A1 => n7487, A2 => n7663, ZN => n9082);
   U15061 : INV_X1 port map( A => n9313, ZN => n7530);
   U15062 : NAND2_X1 port map( A1 => n7494, A2 => n7852, ZN => n7495);
   U15063 : MUX2_X1 port map( A => n7497, B => n7495, S => n7851, Z => n7500);
   U15064 : OAI21_X1 port map( B1 => n8242, B2 => n8244, A => n7501, ZN => 
                           n7505);
   U15065 : NAND2_X1 port map( A1 => n8247, A2 => n7817, ZN => n7503);
   U15067 : AOI21_X1 port map( B1 => n7503, B2 => n7502, A => n7818, ZN => 
                           n7504);
   U15068 : INV_X1 port map( A => n7507, ZN => n7732);
   U15069 : NAND2_X1 port map( A1 => n7732, A2 => n8034, ZN => n8036);
   U15070 : NAND2_X1 port map( A1 => n7507, A2 => n7506, ZN => n8035);
   U15071 : NAND2_X1 port map( A1 => n8034, A2 => n7508, ZN => n7509);
   U15072 : NAND2_X1 port map( A1 => n7510, A2 => n7509, ZN => n7513);
   U15075 : NAND2_X1 port map( A1 => n7850, A2 => n29130, ZN => n7516);
   U15076 : OAI211_X1 port map( C1 => n7517, C2 => n29130, A => n7516, B => 
                           n29106, ZN => n7518);
   U15077 : NOR2_X1 port map( A1 => n8817, A2 => n8592, ZN => n8129);
   U15078 : INV_X1 port map( A => n8129, ZN => n7529);
   U15079 : INV_X1 port map( A => n7521, ZN => n7734);
   U15081 : NAND2_X1 port map( A1 => n7266, A2 => n8032, ZN => n7738);
   U15082 : OAI21_X1 port map( B1 => n7266, B2 => n7737, A => n7738, ZN => 
                           n7522);
   U15083 : NAND2_X1 port map( A1 => n7523, A2 => n8014, ZN => n7748);
   U15086 : AOI21_X1 port map( B1 => n7525, B2 => n7747, A => n7744, ZN => 
                           n7526);
   U15087 : NAND2_X1 port map( A1 => n2024, A2 => n607, ZN => n7528);
   U15088 : XNOR2_X1 port map( A => n7530, B => n10395, ZN => n10288);
   U15089 : INV_X1 port map( A => n10288, ZN => n7571);
   U15090 : NAND2_X1 port map( A1 => n7743, A2 => n7742, ZN => n8015);
   U15091 : NAND2_X1 port map( A1 => n8015, A2 => n8013, ZN => n7532);
   U15092 : INV_X1 port map( A => n7533, ZN => n7749);
   U15093 : INV_X1 port map( A => n9062, ZN => n8393);
   U15094 : NAND3_X1 port map( A1 => n7536, A2 => n8159, A3 => n7535, ZN => 
                           n7539);
   U15095 : NAND2_X1 port map( A1 => n7537, A2 => n8161, ZN => n7538);
   U15096 : NAND2_X1 port map( A1 => n8393, A2 => n9060, ZN => n8871);
   U15097 : AND2_X1 port map( A1 => n28149, A2 => n8148, ZN => n7546);
   U15098 : INV_X1 port map( A => n7792, ZN => n7540);
   U15099 : NAND2_X1 port map( A1 => n7541, A2 => n7540, ZN => n7545);
   U15102 : OAI21_X1 port map( B1 => n7546, B2 => n7545, A => n7544, ZN => 
                           n8865);
   U15103 : OAI21_X1 port map( B1 => n7785, B2 => n7787, A => n1899, ZN => 
                           n7548);
   U15104 : NAND2_X1 port map( A1 => n7782, A2 => n7786, ZN => n7547);
   U15105 : NAND2_X1 port map( A1 => n7548, A2 => n7547, ZN => n7553);
   U15106 : NAND2_X1 port map( A1 => n7291, A2 => n7550, ZN => n7549);
   U15107 : OAI21_X1 port map( B1 => n7550, B2 => n1899, A => n7549, ZN => 
                           n7551);
   U15108 : NAND2_X1 port map( A1 => n7551, A2 => n7330, ZN => n7552);
   U15109 : NAND2_X1 port map( A1 => n7553, A2 => n7552, ZN => n8397);
   U15110 : NAND2_X1 port map( A1 => n8865, A2 => n8397, ZN => n8104);
   U15111 : NAND2_X1 port map( A1 => n9062, A2 => n8104, ZN => n7568);
   U15112 : MUX2_X1 port map( A => n29646, B => n7127, S => n8047, Z => n7555);
   U15113 : NAND2_X1 port map( A1 => n7555, A2 => n7554, ZN => n7559);
   U15115 : NAND2_X1 port map( A1 => n8044, A2 => n8138, ZN => n7561);
   U15116 : NAND2_X1 port map( A1 => n7561, A2 => n7336, ZN => n7564);
   U15117 : NAND2_X1 port map( A1 => n8043, A2 => n7562, ZN => n7563);
   U15118 : NAND2_X1 port map( A1 => n7564, A2 => n7563, ZN => n7567);
   U15119 : MUX2_X1 port map( A => n7723, B => n7565, S => n7722, Z => n7566);
   U15120 : INV_X1 port map( A => n8865, ZN => n9059);
   U15121 : NAND2_X1 port map( A1 => n8581, A2 => n606, ZN => n9581);
   U15122 : NOR2_X1 port map( A1 => n7569, A2 => n9421, ZN => n8770);
   U15123 : XNOR2_X1 port map( A => n9779, B => n10201, ZN => n7570);
   U15124 : INV_X1 port map( A => n11146, ZN => n7813);
   U15125 : INV_X1 port map( A => n8729, ZN => n8734);
   U15126 : AND2_X1 port map( A1 => n8381, A2 => n8733, ZN => n8369);
   U15127 : NAND2_X1 port map( A1 => n6909, A2 => n8537, ZN => n7574);
   U15129 : AOI21_X1 port map( B1 => n4696, B2 => n29301, A => n1568, ZN => 
                           n7577);
   U15130 : NAND2_X1 port map( A1 => n7966, A2 => n7964, ZN => n7576);
   U15133 : NAND2_X1 port map( A1 => n7995, A2 => n7992, ZN => n7651);
   U15134 : NAND2_X1 port map( A1 => n8002, A2 => n7649, ZN => n7579);
   U15135 : NAND2_X1 port map( A1 => n7582, A2 => n7581, ZN => n7587);
   U15136 : NAND2_X1 port map( A1 => n7584, A2 => n7583, ZN => n7586);
   U15137 : AOI21_X1 port map( B1 => n7587, B2 => n7586, A => n7585, ZN => 
                           n7588);
   U15139 : INV_X1 port map( A => n8718, ZN => n8785);
   U15140 : INV_X1 port map( A => n7897, ZN => n7805);
   U15141 : AOI21_X1 port map( B1 => n7596, B2 => n7595, A => n7805, ZN => 
                           n7599);
   U15142 : AOI21_X1 port map( B1 => n7597, B2 => n7312, A => n7896, ZN => 
                           n7598);
   U15143 : NAND2_X1 port map( A1 => n7862, A2 => n7865, ZN => n7600);
   U15144 : NAND3_X1 port map( A1 => n7604, A2 => n7601, A3 => n7600, ZN => 
                           n7603);
   U15145 : NOR2_X1 port map( A1 => n8788, A2 => n8718, ZN => n7605);
   U15146 : AOI22_X1 port map( A1 => n7606, A2 => n8787, B1 => n7605, B2 => 
                           n8717, ZN => n7608);
   U15147 : OAI211_X2 port map( C1 => n8438, C2 => n8442, A => n7608, B => 
                           n7607, ZN => n10019);
   U15148 : OAI21_X1 port map( B1 => n8311, B2 => n7934, A => n7609, ZN => 
                           n7612);
   U15149 : INV_X1 port map( A => n7610, ZN => n7611);
   U15151 : INV_X1 port map( A => n7613, ZN => n7931);
   U15152 : NAND2_X1 port map( A1 => n7931, A2 => n7614, ZN => n7615);
   U15153 : INV_X1 port map( A => n9196, ZN => n8779);
   U15154 : INV_X1 port map( A => n329, ZN => n9201);
   U15155 : NAND2_X1 port map( A1 => n2089, A2 => n7920, ZN => n7621);
   U15156 : NAND3_X1 port map( A1 => n7621, A2 => n8231, A3 => n8235, ZN => 
                           n7622);
   U15158 : NAND2_X1 port map( A1 => n7925, A2 => n8213, ZN => n7927);
   U15159 : NAND2_X1 port map( A1 => n8217, A2 => n7626, ZN => n7624);
   U15160 : NAND3_X1 port map( A1 => n7626, A2 => n8216, A3 => n7925, ZN => 
                           n7627);
   U15161 : INV_X1 port map( A => n9200, ZN => n9194);
   U15162 : NAND2_X1 port map( A1 => n29568, A2 => n7628, ZN => n7633);
   U15163 : NAND2_X1 port map( A1 => n7631, A2 => n7915, ZN => n7632);
   U15164 : MUX2_X1 port map( A => n7636, B => n8202, S => n7635, Z => n7637);
   U15165 : INV_X1 port map( A => n9197, ZN => n9195);
   U15166 : NAND3_X1 port map( A1 => n9195, A2 => n8779, A3 => n9201, ZN => 
                           n7638);
   U15168 : INV_X1 port map( A => n9211, ZN => n9435);
   U15170 : AOI21_X1 port map( B1 => n7652, B2 => n7992, A => n7998, ZN => 
                           n7653);
   U15172 : NAND2_X1 port map( A1 => n8304, A2 => n7655, ZN => n7656);
   U15173 : AOI21_X1 port map( B1 => n8298, B2 => n7656, A => n29317, ZN => 
                           n7661);
   U15177 : NAND2_X1 port map( A1 => n7664, A2 => n7663, ZN => n7668);
   U15178 : NAND3_X1 port map( A1 => n631, A2 => n8270, A3 => n8264, ZN => 
                           n7667);
   U15179 : NAND3_X1 port map( A1 => n8265, A2 => n7986, A3 => n341, ZN => 
                           n7666);
   U15180 : INV_X1 port map( A => n8777, ZN => n9436);
   U15181 : INV_X1 port map( A => n8996, ZN => n9209);
   U15182 : INV_X1 port map( A => n29301, ZN => n7674);
   U15183 : OAI21_X1 port map( B1 => n7675, B2 => n7968, A => n7674, ZN => 
                           n7677);
   U15184 : NAND2_X1 port map( A1 => n7966, A2 => n29302, ZN => n7676);
   U15185 : NAND3_X1 port map( A1 => n9434, A2 => n8777, A3 => n9210, ZN => 
                           n7681);
   U15186 : XNOR2_X1 port map( A => n9772, B => n10322, ZN => n9675);
   U15187 : XNOR2_X1 port map( A => n8883, B => n9675, ZN => n7812);
   U15188 : NAND2_X1 port map( A1 => n8022, A2 => n7685, ZN => n7689);
   U15189 : NAND2_X1 port map( A1 => n7684, A2 => n29106, ZN => n7688);
   U15190 : AND2_X1 port map( A1 => n7850, A2 => n7843, ZN => n7687);
   U15192 : NAND2_X1 port map( A1 => n7821, A2 => n7822, ZN => n7697);
   U15193 : NAND2_X1 port map( A1 => n439, A2 => n7367, ZN => n7704);
   U15194 : NAND2_X1 port map( A1 => n619, A2 => n7839, ZN => n7701);
   U15195 : OAI211_X1 port map( C1 => n7840, C2 => n7839, A => n7701, B => 
                           n7700, ZN => n7703);
   U15196 : NAND3_X1 port map( A1 => n7837, A2 => n7835, A3 => n370, ZN => 
                           n7702);
   U15197 : NAND2_X1 port map( A1 => n9034, A2 => n8792, ZN => n8360);
   U15198 : AOI21_X1 port map( B1 => n7711, B2 => n7710, A => n618, ZN => n7712
                           );
   U15199 : XNOR2_X1 port map( A => n10384, B => n2511, ZN => n7810);
   U15200 : AOI21_X1 port map( B1 => n8135, B2 => n8048, A => n8049, ZN => 
                           n7719);
   U15201 : NAND2_X1 port map( A1 => n9188, A2 => n9007, ZN => n7741);
   U15202 : INV_X1 port map( A => n7726, ZN => n8445);
   U15203 : NAND3_X1 port map( A1 => n7729, A2 => n8038, A3 => n29629, ZN => 
                           n7730);
   U15205 : NAND2_X1 port map( A1 => n8445, A2 => n9186, ZN => n7740);
   U15206 : NAND2_X1 port map( A1 => n7265, A2 => n7737, ZN => n8033);
   U15207 : OAI21_X1 port map( B1 => n7738, B2 => n8030, A => n8033, ZN => 
                           n7739);
   U15208 : INV_X1 port map( A => n8782, ZN => n9187);
   U15209 : AOI21_X1 port map( B1 => n7741, B2 => n7740, A => n9187, ZN => 
                           n7757);
   U15210 : MUX2_X1 port map( A => n8160, B => n8167, S => n8162, Z => n7754);
   U15211 : NAND2_X1 port map( A1 => n7751, A2 => n8159, ZN => n7753);
   U15212 : AND2_X1 port map( A1 => n8162, A2 => n8158, ZN => n7752);
   U15213 : AOI21_X2 port map( B1 => n7754, B2 => n7753, A => n7752, ZN => 
                           n9009);
   U15214 : INV_X1 port map( A => n9007, ZN => n9185);
   U15215 : NAND2_X1 port map( A1 => n613, A2 => n7758, ZN => n7762);
   U15217 : AND2_X1 port map( A1 => n7775, A2 => n7089, ZN => n7893);
   U15218 : INV_X1 port map( A => n7893, ZN => n7780);
   U15219 : NAND3_X1 port map( A1 => n7778, A2 => n7777, A3 => n438, ZN => 
                           n7779);
   U15221 : INV_X1 port map( A => n7786, ZN => n7783);
   U15222 : NAND2_X1 port map( A1 => n7787, A2 => n7786, ZN => n7788);
   U15223 : MUX2_X1 port map( A => n7789, B => n7788, S => n7291, Z => n7790);
   U15224 : AOI21_X1 port map( B1 => n7794, B2 => n7793, A => n8150, ZN => 
                           n7799);
   U15225 : NAND2_X1 port map( A1 => n7796, A2 => n8150, ZN => n7797);
   U15226 : OAI211_X1 port map( C1 => n8353, C2 => n8351, A => n7809, B => 
                           n8077, ZN => n7808);
   U15229 : XNOR2_X1 port map( A => n7810, B => n10179, ZN => n7811);
   U15230 : NAND2_X1 port map( A1 => n8244, A2 => n7376, ZN => n7815);
   U15231 : AND2_X1 port map( A1 => n7815, A2 => n7816, ZN => n7820);
   U15232 : NAND2_X1 port map( A1 => n608, A2 => n9012, ZN => n9019);
   U15233 : AOI21_X1 port map( B1 => n7829, B2 => n7828, A => n7363, ZN => 
                           n7834);
   U15234 : AOI21_X1 port map( B1 => n7832, B2 => n7831, A => n7362, ZN => 
                           n7833);
   U15235 : INV_X1 port map( A => n8910, ZN => n9018);
   U15236 : NAND2_X1 port map( A1 => n9019, A2 => n5674, ZN => n7860);
   U15237 : AND2_X1 port map( A1 => n7836, A2 => n7840, ZN => n8209);
   U15239 : NAND2_X1 port map( A1 => n7844, A2 => n8023, ZN => n7845);
   U15240 : OAI211_X1 port map( C1 => n7846, C2 => n7844, A => n7845, B => 
                           n29106, ZN => n7848);
   U15241 : NAND2_X1 port map( A1 => n8908, A2 => n9014, ZN => n8906);
   U15242 : NAND2_X1 port map( A1 => n8906, A2 => n8910, ZN => n7859);
   U15243 : NAND2_X1 port map( A1 => n7851, A2 => n7384, ZN => n7854);
   U15244 : AOI22_X1 port map( A1 => n7855, A2 => n7854, B1 => n7853, B2 => 
                           n7852, ZN => n7858);
   U15245 : INV_X1 port map( A => n9015, ZN => n9013);
   U15246 : NAND3_X1 port map( A1 => n7865, A2 => n7172, A3 => n7864, ZN => 
                           n7866);
   U15247 : NAND2_X1 port map( A1 => n7873, A2 => n7872, ZN => n7874);
   U15248 : INV_X1 port map( A => n8116, ZN => n8655);
   U15249 : NAND2_X1 port map( A1 => n29082, A2 => n7997, ZN => n7881);
   U15250 : NAND3_X1 port map( A1 => n7877, A2 => n7993, A3 => n7994, ZN => 
                           n7880);
   U15251 : INV_X1 port map( A => n7993, ZN => n7878);
   U15252 : INV_X1 port map( A => n8502, ZN => n8651);
   U15253 : NOR2_X1 port map( A1 => n7890, A2 => n7889, ZN => n7892);
   U15254 : OAI21_X1 port map( B1 => n7893, B2 => n7892, A => n29112, ZN => 
                           n7894);
   U15255 : NOR2_X1 port map( A1 => n8658, A2 => n8502, ZN => n7905);
   U15256 : NAND2_X1 port map( A1 => n7895, A2 => n7312, ZN => n7901);
   U15257 : MUX2_X1 port map( A => n7901, B => n7899, S => n7898, Z => n7904);
   U15258 : OAI211_X1 port map( C1 => n7312, C2 => n7902, A => n7901, B => 
                           n7900, ZN => n7903);
   U15259 : AOI22_X1 port map( A1 => n7906, A2 => n8658, B1 => n7905, B2 => 
                           n8653, ZN => n7907);
   U15260 : NAND2_X1 port map( A1 => n7910, A2 => n7909, ZN => n8292);
   U15261 : INV_X1 port map( A => n9116, ZN => n8917);
   U15262 : MUX2_X1 port map( A => n8231, B => n7919, S => n7920, Z => n7923);
   U15263 : MUX2_X1 port map( A => n7921, B => n8236, S => n5946, Z => n7922);
   U15264 : NAND2_X1 port map( A1 => n8917, A2 => n9108, ZN => n8671);
   U15265 : INV_X1 port map( A => n9108, ZN => n9106);
   U15266 : NAND2_X1 port map( A1 => n8212, A2 => n7925, ZN => n7929);
   U15267 : INV_X1 port map( A => n7926, ZN => n7928);
   U15268 : NAND2_X1 port map( A1 => n9106, A2 => n8669, ZN => n7938);
   U15269 : OAI21_X1 port map( B1 => n7932, B2 => n7931, A => n7930, ZN => 
                           n9109);
   U15270 : INV_X1 port map( A => n7935, ZN => n7934);
   U15271 : NAND2_X1 port map( A1 => n7934, A2 => n7933, ZN => n7937);
   U15272 : NAND2_X1 port map( A1 => n7935, A2 => n7614, ZN => n7936);
   U15273 : AND2_X1 port map( A1 => n7937, A2 => n7936, ZN => n9112);
   U15274 : MUX2_X2 port map( A => n9109, B => n9112, S => n29135, Z => n8670);
   U15275 : AOI21_X1 port map( B1 => n8671, B2 => n7938, A => n8511, ZN => 
                           n7956);
   U15276 : AOI21_X1 port map( B1 => n7941, B2 => n7940, A => n7939, ZN => 
                           n7945);
   U15277 : AOI21_X1 port map( B1 => n7943, B2 => n7942, A => n8296, ZN => 
                           n7944);
   U15278 : INV_X1 port map( A => n8914, ZN => n8513);
   U15279 : NAND2_X1 port map( A1 => n28618, A2 => n8257, ZN => n7952);
   U15280 : NAND3_X1 port map( A1 => n6782, A2 => n7948, A3 => n8258, ZN => 
                           n7950);
   U15281 : NAND2_X1 port map( A1 => n8513, A2 => n9107, ZN => n7954);
   U15282 : NAND3_X1 port map( A1 => n9108, A2 => n9116, A3 => n8914, ZN => 
                           n7953);
   U15284 : INV_X1 port map( A => n8666, ZN => n8492);
   U15285 : NAND2_X1 port map( A1 => n7967, A2 => n7966, ZN => n7971);
   U15287 : MUX2_X1 port map( A => n7971, B => n7970, S => n29302, Z => n7972);
   U15288 : NAND2_X1 port map( A1 => n8284, A2 => n8280, ZN => n7974);
   U15289 : MUX2_X1 port map( A => n7974, B => n8275, S => n8276, Z => n7979);
   U15290 : NOR2_X1 port map( A1 => n7975, A2 => n8280, ZN => n7977);
   U15291 : NAND2_X1 port map( A1 => n8665, A2 => n8073, ZN => n8006);
   U15292 : NAND2_X1 port map( A1 => n7982, A2 => n7981, ZN => n7983);
   U15293 : AND2_X1 port map( A1 => n8267, A2 => n8264, ZN => n7989);
   U15294 : NAND2_X1 port map( A1 => n7986, A2 => n8270, ZN => n7988);
   U15295 : NAND3_X1 port map( A1 => n8271, A2 => n8265, A3 => n8264, ZN => 
                           n7987);
   U15296 : NAND2_X1 port map( A1 => n7993, A2 => n7992, ZN => n8003);
   U15297 : NAND2_X1 port map( A1 => n7995, A2 => n7994, ZN => n7996);
   U15298 : NAND3_X1 port map( A1 => n8003, A2 => n7997, A3 => n7996, ZN => 
                           n8001);
   U15299 : NAND3_X1 port map( A1 => n7999, A2 => n8002, A3 => n7998, ZN => 
                           n8000);
   U15300 : OAI211_X1 port map( C1 => n8003, C2 => n8002, A => n8001, B => 
                           n8000, ZN => n9095);
   U15301 : OAI211_X1 port map( C1 => n8492, C2 => n8006, A => n8005, B => 
                           n8004, ZN => n10310);
   U15302 : XNOR2_X1 port map( A => n10310, B => n10357, ZN => n9672);
   U15303 : XNOR2_X1 port map( A => n10433, B => n9672, ZN => n8063);
   U15304 : OAI21_X1 port map( B1 => n8334, B2 => n8889, A => n8007, ZN => 
                           n8008);
   U15306 : INV_X1 port map( A => n8009, ZN => n8507);
   U15307 : NAND3_X1 port map( A1 => n8507, A2 => n8891, A3 => n8335, ZN => 
                           n8011);
   U15308 : NAND2_X1 port map( A1 => n8009, A2 => n8336, ZN => n8888);
   U15310 : NAND3_X1 port map( A1 => n8016, A2 => n8015, A3 => n8014, ZN => 
                           n8017);
   U15311 : NAND2_X1 port map( A1 => n8019, A2 => n28161, ZN => n8020);
   U15312 : NAND2_X1 port map( A1 => n29106, A2 => n29130, ZN => n8021);
   U15313 : AOI21_X1 port map( B1 => n8022, B2 => n8021, A => n7844, ZN => 
                           n8026);
   U15314 : INV_X1 port map( A => n8899, ZN => n8898);
   U15316 : NAND2_X1 port map( A1 => n8898, A2 => n9124, ZN => n9364);
   U15317 : NAND3_X1 port map( A1 => n8036, A2 => n8035, A3 => n8038, ZN => 
                           n8037);
   U15318 : AND2_X1 port map( A1 => n29304, A2 => n8899, ZN => n8663);
   U15319 : NAND2_X1 port map( A1 => n8041, A2 => n29751, ZN => n8146);
   U15320 : NAND2_X1 port map( A1 => n8043, A2 => n8143, ZN => n8042);
   U15321 : AOI21_X1 port map( B1 => n8146, B2 => n8042, A => n8044, ZN => 
                           n8487);
   U15322 : NAND2_X1 port map( A1 => n8043, A2 => n8141, ZN => n8046);
   U15324 : AOI21_X1 port map( B1 => n8046, B2 => n8045, A => n8143, ZN => 
                           n8486);
   U15325 : NAND2_X1 port map( A1 => n8663, A2 => n9125, ZN => n9365);
   U15326 : AND2_X1 port map( A1 => n8048, A2 => n8047, ZN => n8051);
   U15327 : NAND2_X1 port map( A1 => n9125, A2 => n29304, ZN => n8053);
   U15328 : OAI211_X1 port map( C1 => n284, C2 => n9125, A => n8053, B => n3274
                           , ZN => n8054);
   U15329 : OAI211_X1 port map( C1 => n3274, C2 => n9364, A => n9365, B => 
                           n8054, ZN => n8055);
   U15330 : XNOR2_X1 port map( A => n9504, B => n8055, ZN => n10209);
   U15331 : NAND3_X1 port map( A1 => n8431, A2 => n8351, A3 => n8353, ZN => 
                           n8057);
   U15332 : INV_X1 port map( A => n8351, ZN => n8428);
   U15333 : NAND3_X1 port map( A1 => n8426, A2 => n8427, A3 => n8428, ZN => 
                           n8056);
   U15334 : AND2_X1 port map( A1 => n8056, A2 => n8057, ZN => n8060);
   U15335 : NAND3_X1 port map( A1 => n8430, A2 => n8428, A3 => n8058, ZN => 
                           n8059);
   U15336 : XNOR2_X1 port map( A => n10071, B => n1172, ZN => n8061);
   U15337 : XNOR2_X1 port map( A => n10209, B => n8061, ZN => n8062);
   U15338 : INV_X1 port map( A => n284, ZN => n8488);
   U15339 : NAND3_X1 port map( A1 => n8898, A2 => n9125, A3 => n8488, ZN => 
                           n8068);
   U15340 : NAND3_X1 port map( A1 => n610, A2 => n284, A3 => n8899, ZN => n8067
                           );
   U15341 : NAND3_X1 port map( A1 => n610, A2 => n284, A3 => n9124, ZN => n8066
                           );
   U15342 : NAND2_X1 port map( A1 => n8899, A2 => n1793, ZN => n8065);
   U15343 : NAND2_X1 port map( A1 => n8656, A2 => n8116, ZN => n8498);
   U15344 : NAND2_X1 port map( A1 => n8498, A2 => n8502, ZN => n8070);
   U15345 : OAI21_X1 port map( B1 => n8498, B2 => n8635, A => n8115, ZN => 
                           n8069);
   U15346 : XNOR2_X1 port map( A => n10144, B => n10219, ZN => n9892);
   U15347 : INV_X1 port map( A => n9892, ZN => n9336);
   U15348 : INV_X1 port map( A => n8669, ZN => n9118);
   U15349 : AND2_X1 port map( A1 => n8073, A2 => n8664, ZN => n9096);
   U15350 : NAND2_X1 port map( A1 => n9096, A2 => n8492, ZN => n8076);
   U15351 : INV_X1 port map( A => n8665, ZN => n8630);
   U15352 : INV_X1 port map( A => n8664, ZN => n8491);
   U15353 : NAND3_X1 port map( A1 => n8630, A2 => n8491, A3 => n9095, ZN => 
                           n8075);
   U15354 : NAND3_X1 port map( A1 => n8630, A2 => n8491, A3 => n8666, ZN => 
                           n8074);
   U15355 : XNOR2_X1 port map( A => n28634, B => n10028, ZN => n9782);
   U15356 : XNOR2_X1 port map( A => n9336, B => n9782, ZN => n8090);
   U15357 : NAND2_X1 port map( A1 => n8079, A2 => n8507, ZN => n8080);
   U15358 : NAND2_X1 port map( A1 => n8080, A2 => n8892, ZN => n8083);
   U15359 : INV_X1 port map( A => n8889, ZN => n8081);
   U15360 : INV_X1 port map( A => n8336, ZN => n8890);
   U15361 : OAI211_X1 port map( C1 => n8891, C2 => n8009, A => n8081, B => 
                           n8890, ZN => n8082);
   U15362 : INV_X1 port map( A => n10289, ZN => n9757);
   U15363 : XNOR2_X1 port map( A => n9992, B => n9757, ZN => n8088);
   U15364 : INV_X1 port map( A => n8481, ZN => n8086);
   U15365 : NAND3_X1 port map( A1 => n5674, A2 => n9013, A3 => n9014, ZN => 
                           n8084);
   U15366 : AND3_X1 port map( A1 => n8086, A2 => n8085, A3 => n8084, ZN => 
                           n10143);
   U15367 : XNOR2_X1 port map( A => n10143, B => n3087, ZN => n8087);
   U15368 : XNOR2_X1 port map( A => n8088, B => n8087, ZN => n8089);
   U15369 : INV_X1 port map( A => n10820, ZN => n11169);
   U15370 : NAND2_X1 port map( A1 => n9238, A2 => n8544, ZN => n8092);
   U15371 : INV_X1 port map( A => n9229, ZN => n9237);
   U15372 : OAI21_X1 port map( B1 => n9237, B2 => n9233, A => n9232, ZN => 
                           n8091);
   U15374 : AOI21_X1 port map( B1 => n8433, B2 => n28210, A => n9027, ZN => 
                           n8094);
   U15375 : INV_X1 port map( A => n8526, ZN => n8097);
   U15376 : NAND2_X1 port map( A1 => n8097, A2 => n8688, ZN => n8101);
   U15377 : NAND2_X1 port map( A1 => n597, A2 => n9220, ZN => n8100);
   U15378 : NAND2_X1 port map( A1 => n8098, A2 => n597, ZN => n8099);
   U15379 : NAND4_X2 port map( A1 => n8102, A2 => n8101, A3 => n8099, A4 => 
                           n8100, ZN => n9929);
   U15382 : INV_X1 port map( A => n8104, ZN => n8105);
   U15383 : NAND2_X1 port map( A1 => n8105, A2 => n9061, ZN => n8106);
   U15384 : OAI211_X1 port map( C1 => n8395, C2 => n9062, A => n8107, B => 
                           n8106, ZN => n9963);
   U15385 : XNOR2_X1 port map( A => n9963, B => n9929, ZN => n8108);
   U15386 : XNOR2_X1 port map( A => n10123, B => n8108, ZN => n8126);
   U15387 : AND2_X1 port map( A1 => n8109, A2 => n8693, ZN => n9246);
   U15388 : INV_X1 port map( A => n9246, ZN => n8114);
   U15389 : NAND2_X1 port map( A1 => n8110, A2 => n9247, ZN => n8111);
   U15390 : NAND2_X1 port map( A1 => n8111, A2 => n9245, ZN => n8113);
   U15391 : AND2_X1 port map( A1 => n9247, A2 => n9243, ZN => n9412);
   U15392 : NAND2_X1 port map( A1 => n9412, A2 => n8693, ZN => n8112);
   U15393 : OAI211_X2 port map( C1 => n8114, C2 => n9245, A => n8113, B => 
                           n8112, ZN => n10304);
   U15394 : XNOR2_X1 port map( A => n10009, B => n10304, ZN => n8124);
   U15395 : INV_X1 port map( A => n8427, ZN => n8119);
   U15396 : AOI21_X1 port map( B1 => n8119, B2 => n1910, A => n8426, ZN => 
                           n8122);
   U15397 : NAND2_X1 port map( A1 => n8120, A2 => n8353, ZN => n8121);
   U15398 : XNOR2_X1 port map( A => n10088, B => n2602, ZN => n8123);
   U15399 : XNOR2_X1 port map( A => n8124, B => n8123, ZN => n8125);
   U15400 : INV_X1 port map( A => n11330, ZN => n11331);
   U15402 : INV_X1 port map( A => n8817, ZN => n8976);
   U15403 : INV_X1 port map( A => n8593, ZN => n8974);
   U15404 : INV_X1 port map( A => n8592, ZN => n8591);
   U15405 : NAND3_X1 port map( A1 => n8974, A2 => n607, A3 => n8591, ZN => 
                           n8128);
   U15406 : NAND3_X1 port map( A1 => n8977, A2 => n8819, A3 => n8594, ZN => 
                           n8127);
   U15407 : AOI21_X1 port map( B1 => n8135, B2 => n8134, A => n8133, ZN => 
                           n8137);
   U15408 : NAND2_X1 port map( A1 => n8139, A2 => n8138, ZN => n8140);
   U15409 : NAND3_X1 port map( A1 => n8146, A2 => n8141, A3 => n8140, ZN => 
                           n8145);
   U15410 : NAND3_X1 port map( A1 => n8143, A2 => n7336, A3 => n8142, ZN => 
                           n8144);
   U15411 : OAI211_X1 port map( C1 => n8146, C2 => n7336, A => n8145, B => 
                           n8144, ZN => n9396);
   U15412 : NAND2_X1 port map( A1 => n8981, A2 => n9396, ZN => n9398);
   U15413 : NAND2_X1 port map( A1 => n8147, A2 => n8150, ZN => n8149);
   U15414 : OAI211_X1 port map( C1 => n28149, C2 => n1607, A => n8149, B => 
                           n8148, ZN => n8152);
   U15415 : AND2_X1 port map( A1 => n8153, A2 => n7550, ZN => n8157);
   U15416 : NAND3_X1 port map( A1 => n8162, A2 => n8161, A3 => n8160, ZN => 
                           n8163);
   U15418 : NAND2_X1 port map( A1 => n8166, A2 => n8165, ZN => n8170);
   U15420 : AOI21_X1 port map( B1 => n8170, B2 => n8169, A => n8168, ZN => 
                           n8171);
   U15421 : INV_X1 port map( A => n8176, ZN => n8178);
   U15422 : NAND3_X1 port map( A1 => n8173, A2 => n7760, A3 => n8178, ZN => 
                           n8174);
   U15423 : NAND2_X1 port map( A1 => n8175, A2 => n8174, ZN => n8183);
   U15424 : NAND2_X1 port map( A1 => n8177, A2 => n8176, ZN => n8181);
   U15425 : INV_X1 port map( A => n8980, ZN => n8644);
   U15426 : NAND3_X1 port map( A1 => n8644, A2 => n596, A3 => n8982, ZN => 
                           n8184);
   U15427 : INV_X1 port map( A => n9144, ZN => n8561);
   U15428 : NAND2_X1 port map( A1 => n8561, A2 => n8185, ZN => n8186);
   U15429 : INV_X1 port map( A => n8563, ZN => n9142);
   U15430 : NAND3_X1 port map( A1 => n8561, A2 => n598, A3 => n9142, ZN => 
                           n8188);
   U15431 : XNOR2_X1 port map( A => n9295, B => n3770, ZN => n8191);
   U15432 : XNOR2_X1 port map( A => n9770, B => n8191, ZN => n8319);
   U15433 : NAND2_X1 port map( A1 => n8829, A2 => n8827, ZN => n8198);
   U15434 : NAND2_X1 port map( A1 => n8829, A2 => n8192, ZN => n8195);
   U15435 : OAI21_X1 port map( B1 => n8829, B2 => n8193, A => n8826, ZN => 
                           n8194);
   U15436 : OAI211_X1 port map( C1 => n8196, C2 => n8826, A => n8195, B => 
                           n8194, ZN => n8197);
   U15437 : NAND2_X1 port map( A1 => n8203, A2 => n8205, ZN => n8204);
   U15438 : NOR2_X1 port map( A1 => n8836, A2 => n8838, ZN => n9169);
   U15439 : INV_X1 port map( A => n8838, ZN => n8229);
   U15441 : AOI21_X1 port map( B1 => n8218, B2 => n8217, A => n8216, ZN => 
                           n8219);
   U15442 : OR2_X2 port map( A1 => n8220, A2 => n8219, ZN => n9171);
   U15443 : MUX2_X1 port map( A => n3821, B => n8222, S => n8221, Z => n8228);
   U15444 : INV_X1 port map( A => n8230, ZN => n8964);
   U15445 : OAI21_X1 port map( B1 => n8229, B2 => n9171, A => n8964, ZN => 
                           n8250);
   U15446 : NAND2_X1 port map( A1 => n8233, A2 => n8232, ZN => n8241);
   U15448 : NAND2_X1 port map( A1 => n8236, A2 => n8235, ZN => n8238);
   U15449 : MUX2_X1 port map( A => n8239, B => n8238, S => n29110, Z => n8240);
   U15450 : NAND3_X1 port map( A1 => n8961, A2 => n9171, A3 => n9170, ZN => 
                           n8249);
   U15451 : INV_X1 port map( A => n8836, ZN => n8962);
   U15452 : NAND3_X1 port map( A1 => n8962, A2 => n605, A3 => n8837, ZN => 
                           n8248);
   U15453 : XNOR2_X1 port map( A => n10060, B => n10178, ZN => n9845);
   U15454 : NAND2_X1 port map( A1 => n8521, A2 => n8811, ZN => n8251);
   U15455 : AND2_X1 port map( A1 => n8253, A2 => n8252, ZN => n8254);
   U15456 : MUX2_X1 port map( A => n8257, B => n28615, S => n8258, Z => n8262);
   U15457 : MUX2_X1 port map( A => n8260, B => n8259, S => n8258, Z => n8261);
   U15459 : INV_X1 port map( A => n8954, ZN => n8471);
   U15460 : INV_X1 port map( A => n8266, ZN => n8274);
   U15461 : NAND2_X1 port map( A1 => n8272, A2 => n8271, ZN => n8273);
   U15462 : NAND2_X1 port map( A1 => n8471, A2 => n8958, ZN => n9167);
   U15463 : INV_X1 port map( A => n8275, ZN => n8278);
   U15464 : INV_X1 port map( A => n8280, ZN => n8282);
   U15465 : INV_X1 port map( A => n8956, ZN => n9163);
   U15466 : INV_X1 port map( A => n8286, ZN => n8289);
   U15467 : NAND2_X1 port map( A1 => n7915, A2 => n8287, ZN => n8288);
   U15469 : NAND2_X1 port map( A1 => n8291, A2 => n7915, ZN => n8293);
   U15472 : NAND3_X1 port map( A1 => n8302, A2 => n8301, A3 => n29317, ZN => 
                           n8307);
   U15473 : OAI211_X1 port map( C1 => n9160, C2 => n8958, A => n9162, B => 
                           n29096, ZN => n8317);
   U15474 : INV_X1 port map( A => n8958, ZN => n9164);
   U15475 : NAND2_X1 port map( A1 => n8308, A2 => n28810, ZN => n8309);
   U15476 : AOI21_X1 port map( B1 => n8310, B2 => n8309, A => n7614, ZN => 
                           n8315);
   U15477 : NAND3_X1 port map( A1 => n7934, A2 => n28810, A3 => n7933, ZN => 
                           n8313);
   U15478 : NAND3_X1 port map( A1 => n8311, A2 => n7614, A3 => n7933, ZN => 
                           n8312);
   U15479 : NAND2_X1 port map( A1 => n8313, A2 => n8312, ZN => n8314);
   U15480 : INV_X1 port map( A => n8802, ZN => n9161);
   U15481 : INV_X1 port map( A => n8955, ZN => n8800);
   U15482 : XNOR2_X1 port map( A => n28488, B => n10059, ZN => n9549);
   U15483 : XNOR2_X1 port map( A => n9845, B => n9549, ZN => n8318);
   U15485 : NOR2_X1 port map( A1 => n9531, A2 => n9532, ZN => n8322);
   U15486 : OAI21_X1 port map( B1 => n9532, B2 => n8749, A => n8747, ZN => 
                           n8321);
   U15488 : NOR2_X1 port map( A1 => n8610, A2 => n9530, ZN => n8323);
   U15489 : NAND2_X1 port map( A1 => n8323, A2 => n9531, ZN => n9537);
   U15491 : NAND2_X1 port map( A1 => n7569, A2 => n8579, ZN => n8575);
   U15494 : INV_X1 port map( A => n9323, ZN => n9870);
   U15495 : XNOR2_X1 port map( A => n10033, B => n9870, ZN => n10055);
   U15496 : NAND2_X1 port map( A1 => n598, A2 => n8563, ZN => n8560);
   U15497 : OAI21_X1 port map( B1 => n8762, B2 => n8941, A => n8764, ZN => 
                           n8331);
   U15498 : XNOR2_X1 port map( A => n10055, B => n9736, ZN => n8348);
   U15499 : NAND3_X1 port map( A1 => n8760, A2 => n9148, A3 => n9146, ZN => 
                           n8333);
   U15500 : OAI21_X1 port map( B1 => n8334, B2 => n8336, A => n8009, ZN => 
                           n8339);
   U15501 : NAND3_X1 port map( A1 => n8507, A2 => n8336, A3 => n8335, ZN => 
                           n8338);
   U15502 : NAND3_X1 port map( A1 => n8507, A2 => n8504, A3 => n8891, ZN => 
                           n8337);
   U15503 : XNOR2_X1 port map( A => n10171, B => n9698, ZN => n8346);
   U15504 : AOI21_X1 port map( B1 => n8341, B2 => n8340, A => n7410, ZN => 
                           n8344);
   U15505 : XNOR2_X1 port map( A => n10138, B => n5059, ZN => n8345);
   U15506 : XNOR2_X1 port map( A => n8346, B => n8345, ZN => n8347);
   U15507 : XNOR2_X1 port map( A => n8348, B => n8347, ZN => n10467);
   U15509 : INV_X1 port map( A => n9186, ZN => n9004);
   U15510 : OAI21_X1 port map( B1 => n8445, B2 => n9186, A => n8782, ZN => 
                           n8350);
   U15512 : NOR2_X1 port map( A1 => n8353, A2 => n1909, ZN => n8355);
   U15513 : INV_X1 port map( A => n9202, ZN => n8448);
   U15514 : NOR2_X1 port map( A1 => n9196, A2 => n28862, ZN => n8357);
   U15515 : OAI21_X1 port map( B1 => n6897, B2 => n8357, A => n8448, ZN => 
                           n8359);
   U15517 : OAI21_X1 port map( B1 => n9028, B2 => n8792, A => n9030, ZN => 
                           n8361);
   U15518 : XNOR2_X1 port map( A => n10183, B => n9948, ZN => n10157);
   U15519 : XNOR2_X1 port map( A => n9748, B => n10157, ZN => n8377);
   U15521 : NAND2_X1 port map( A1 => n9435, A2 => n9434, ZN => n8364);
   U15522 : OAI211_X1 port map( C1 => n9434, C2 => n9208, A => n8364, B => 
                           n9210, ZN => n8365);
   U15523 : NAND2_X1 port map( A1 => n9437, A2 => n8365, ZN => n8368);
   U15524 : NAND2_X1 port map( A1 => n8718, A2 => n8787, ZN => n8366);
   U15525 : INV_X1 port map( A => n8787, ZN => n8439);
   U15526 : XNOR2_X1 port map( A => n9823, B => n8368, ZN => n10068);
   U15527 : INV_X1 port map( A => n8369, ZN => n8738);
   U15529 : INV_X1 port map( A => n8733, ZN => n8370);
   U15530 : NAND3_X1 port map( A1 => n8730, A2 => n8370, A3 => n8734, ZN => 
                           n8372);
   U15531 : NAND3_X1 port map( A1 => n8739, A2 => n8370, A3 => n8381, ZN => 
                           n8371);
   U15532 : XNOR2_X1 port map( A => n1895, B => n3607, ZN => n8375);
   U15533 : XNOR2_X1 port map( A => n8375, B => n10068, ZN => n8376);
   U15534 : NAND3_X1 port map( A1 => n11331, A2 => n11166, A3 => n11168, ZN => 
                           n8424);
   U15536 : OAI21_X1 port map( B1 => n8378, B2 => n8741, A => n9070, ZN => 
                           n8379);
   U15537 : NAND2_X1 port map( A1 => n8537, A2 => n8381, ZN => n8382);
   U15538 : OAI21_X1 port map( B1 => n8384, B2 => n8537, A => n8382, ZN => 
                           n8383);
   U15539 : NAND2_X1 port map( A1 => n8383, A2 => n8735, ZN => n8387);
   U15540 : NAND3_X1 port map( A1 => n8384, A2 => n8536, A3 => n8733, ZN => 
                           n8386);
   U15541 : NAND3_X1 port map( A1 => n8731, A2 => n8739, A3 => n8729, ZN => 
                           n8385);
   U15542 : XNOR2_X1 port map( A => n10074, B => n10207, ZN => n9850);
   U15543 : NAND2_X1 port map( A1 => n29311, A2 => n2320, ZN => n8391);
   U15544 : NAND2_X1 port map( A1 => n9080, A2 => n8605, ZN => n10240);
   U15545 : OAI211_X1 port map( C1 => n29311, C2 => n28500, A => n10240, B => 
                           n8848, ZN => n8389);
   U15546 : INV_X1 port map( A => n8848, ZN => n9079);
   U15547 : OAI21_X1 port map( B1 => n29311, B2 => n8726, A => n9079, ZN => 
                           n8388);
   U15548 : NAND2_X1 port map( A1 => n8389, A2 => n8388, ZN => n8390);
   U15549 : OAI21_X1 port map( B1 => n8724, B2 => n8391, A => n8390, ZN => 
                           n9509);
   U15550 : INV_X1 port map( A => n9509, ZN => n9368);
   U15551 : INV_X1 port map( A => n9064, ZN => n8392);
   U15552 : NAND2_X1 port map( A1 => n8392, A2 => n8397, ZN => n8598);
   U15555 : NAND2_X1 port map( A1 => n8396, A2 => n9062, ZN => n8401);
   U15556 : NAND3_X1 port map( A1 => n9060, A2 => n8864, A3 => n9059, ZN => 
                           n8400);
   U15557 : NAND2_X1 port map( A1 => n9064, A2 => n8397, ZN => n9063);
   U15558 : INV_X1 port map( A => n9063, ZN => n8398);
   U15559 : NAND2_X1 port map( A1 => n8398, A2 => n9060, ZN => n8399);
   U15560 : NAND4_X1 port map( A1 => n8402, A2 => n8401, A3 => n8400, A4 => 
                           n8399, ZN => n9592);
   U15561 : XNOR2_X1 port map( A => n9592, B => n9368, ZN => n9943);
   U15562 : XNOR2_X1 port map( A => n9850, B => n9943, ZN => n8421);
   U15563 : NAND2_X1 port map( A1 => n8709, A2 => n8877, ZN => n8708);
   U15564 : OR2_X1 port map( A1 => n8708, A2 => n8873, ZN => n8406);
   U15565 : NAND2_X1 port map( A1 => n8875, A2 => n8881, ZN => n8712);
   U15566 : OR2_X1 port map( A1 => n8712, A2 => n8874, ZN => n8405);
   U15567 : XNOR2_X1 port map( A => n10128, B => n3493, ZN => n8419);
   U15568 : MUX2_X1 port map( A => n8642, B => n8984, S => n8980, Z => n8411);
   U15569 : OR2_X1 port map( A1 => n9396, A2 => n8981, ZN => n9177);
   U15570 : OAI21_X1 port map( B1 => n8644, B2 => n8982, A => n8981, ZN => 
                           n8409);
   U15573 : NAND2_X1 port map( A1 => n8413, A2 => n4321, ZN => n8417);
   U15574 : INV_X1 port map( A => n8788, ZN => n8440);
   U15575 : NAND3_X1 port map( A1 => n8440, A2 => n8720, A3 => n8787, ZN => 
                           n8416);
   U15576 : INV_X1 port map( A => n8719, ZN => n8786);
   U15577 : NAND3_X1 port map( A1 => n8717, A2 => n8786, A3 => n8414, ZN => 
                           n8415);
   U15578 : XNOR2_X1 port map( A => n8419, B => n8418, ZN => n8420);
   U15579 : XNOR2_X1 port map( A => n8421, B => n8420, ZN => n10821);
   U15580 : INV_X1 port map( A => n9392, ZN => n9614);
   U15581 : MUX2_X1 port map( A => n9027, B => n9028, S => n8433, Z => n8434);
   U15582 : INV_X1 port map( A => n10295, ZN => n10034);
   U15583 : XNOR2_X1 port map( A => n10034, B => n9614, ZN => n8444);
   U15584 : MUX2_X1 port map( A => n9211, B => n9434, S => n8777, Z => n8437);
   U15586 : XNOR2_X1 port map( A => n9735, B => n1920, ZN => n8443);
   U15587 : XNOR2_X1 port map( A => n8444, B => n8443, ZN => n8455);
   U15588 : MUX2_X1 port map( A => n9009, B => n9007, S => n9184, Z => n8447);
   U15589 : MUX2_X1 port map( A => n9184, B => n9186, S => n8445, Z => n8446);
   U15591 : NOR2_X1 port map( A1 => n329, A2 => n9200, ZN => n8451);
   U15592 : NAND2_X1 port map( A1 => n9199, A2 => n28862, ZN => n8450);
   U15593 : XNOR2_X1 port map( A => n10298, B => n10038, ZN => n8453);
   U15594 : XNOR2_X1 port map( A => n1902, B => n1184, ZN => n8452);
   U15595 : XNOR2_X1 port map( A => n8453, B => n8452, ZN => n8454);
   U15596 : INV_X1 port map( A => n10748, ZN => n11198);
   U15597 : AOI21_X1 port map( B1 => n8456, B2 => n8980, A => n8983, ZN => 
                           n9399);
   U15598 : INV_X1 port map( A => n9399, ZN => n8458);
   U15599 : NAND2_X1 port map( A1 => n8642, A2 => n8980, ZN => n9397);
   U15600 : OAI21_X1 port map( B1 => n436, B2 => n596, A => n9397, ZN => n9179)
                           ;
   U15601 : NAND2_X1 port map( A1 => n9179, A2 => n9396, ZN => n8457);
   U15602 : NAND2_X1 port map( A1 => n8458, A2 => n8457, ZN => n9656);
   U15603 : NAND2_X1 port map( A1 => n8681, A2 => n8809, ZN => n8459);
   U15604 : NAND2_X1 port map( A1 => n8810, A2 => n8809, ZN => n8460);
   U15605 : XNOR2_X1 port map( A => n9930, B => n9656, ZN => n8469);
   U15606 : INV_X1 port map( A => n8827, ZN => n8825);
   U15607 : XNOR2_X1 port map( A => n9964, B => n3386, ZN => n8468);
   U15608 : XNOR2_X1 port map( A => n8469, B => n8468, ZN => n8480);
   U15609 : AOI22_X1 port map( A1 => n8964, A2 => n9171, B1 => n8838, B2 => 
                           n8966, ZN => n9174);
   U15610 : AND2_X1 port map( A1 => n8836, A2 => n8838, ZN => n8967);
   U15611 : OAI21_X1 port map( B1 => n8967, B2 => n8837, A => n8961, ZN => 
                           n8470);
   U15612 : NAND2_X1 port map( A1 => n8954, A2 => n8956, ZN => n8805);
   U15613 : OAI21_X1 port map( B1 => n8472, B2 => n9161, A => n8471, ZN => 
                           n8474);
   U15614 : NAND3_X1 port map( A1 => n8801, A2 => n8802, A3 => n8956, ZN => 
                           n8473);
   U15615 : OAI211_X1 port map( C1 => n9164, C2 => n8805, A => n8474, B => 
                           n8473, ZN => n10008);
   U15616 : XNOR2_X1 port map( A => n28616, B => n10263, ZN => n10306);
   U15618 : INV_X1 port map( A => n10193, ZN => n8476);
   U15619 : XNOR2_X1 port map( A => n8476, B => n10302, ZN => n8477);
   U15621 : NAND2_X1 port map( A1 => n11198, A2 => n28157, ZN => n8623);
   U15622 : AOI22_X1 port map( A1 => n8481, A2 => n9013, B1 => n9018, B2 => 
                           n8662, ZN => n8484);
   U15623 : NAND2_X1 port map( A1 => n284, A2 => n29304, ZN => n8485);
   U15624 : OAI21_X1 port map( B1 => n8664, B2 => n8665, A => n8490, ZN => 
                           n8496);
   U15626 : OR2_X1 port map( A1 => n8500, A2 => n8499, ZN => n8654);
   U15627 : NAND2_X1 port map( A1 => n8634, A2 => n8653, ZN => n8503);
   U15628 : INV_X1 port map( A => n9430, ZN => n9976);
   U15629 : XNOR2_X1 port map( A => n9976, B => n9771, ZN => n9924);
   U15630 : NAND2_X1 port map( A1 => n8009, A2 => n8889, ZN => n8505);
   U15631 : AOI21_X1 port map( B1 => n8506, B2 => n8505, A => n8504, ZN => 
                           n8510);
   U15632 : OAI21_X1 port map( B1 => n8892, B2 => n8887, A => n8508, ZN => 
                           n8509);
   U15634 : NAND3_X1 port map( A1 => n8916, A2 => n8512, A3 => n8511, ZN => 
                           n8516);
   U15635 : NAND3_X1 port map( A1 => n9106, A2 => n8513, A3 => n8917, ZN => 
                           n8515);
   U15636 : NAND3_X2 port map( A1 => n8515, A2 => n8516, A3 => n8514, ZN => 
                           n10021);
   U15637 : XNOR2_X1 port map( A => n9678, B => n10021, ZN => n8518);
   U15638 : XNOR2_X1 port map( A => n9550, B => n3211, ZN => n8517);
   U15639 : XNOR2_X1 port map( A => n8518, B => n8517, ZN => n8519);
   U15641 : INV_X1 port map( A => n28638, ZN => n10751);
   U15642 : NAND2_X1 port map( A1 => n9224, A2 => n8687, ZN => n8527);
   U15643 : NAND2_X1 port map( A1 => n9228, A2 => n8687, ZN => n8528);
   U15644 : XNOR2_X1 port map( A => n9991, B => n9755, ZN => n9936);
   U15645 : INV_X1 port map( A => n9412, ZN => n8530);
   U15646 : INV_X1 port map( A => n9244, ZN => n8529);
   U15647 : OAI21_X1 port map( B1 => n8693, B2 => n8109, A => n8529, ZN => 
                           n9414);
   U15648 : NAND2_X1 port map( A1 => n9410, A2 => n8109, ZN => n9409);
   U15649 : OAI211_X1 port map( C1 => n8530, C2 => n8109, A => n9414, B => 
                           n9409, ZN => n8535);
   U15650 : AOI21_X1 port map( B1 => n8404, B2 => n8874, A => n8873, ZN => 
                           n8534);
   U15651 : AND2_X1 port map( A1 => n8873, A2 => n8881, ZN => n8878);
   U15652 : INV_X1 port map( A => n8874, ZN => n8531);
   U15653 : NAND3_X1 port map( A1 => n8532, A2 => n8403, A3 => n8531, ZN => 
                           n8533);
   U15654 : OAI21_X1 port map( B1 => n8534, B2 => n8878, A => n8533, ZN => 
                           n9717);
   U15655 : XNOR2_X1 port map( A => n8535, B => n9717, ZN => n10291);
   U15656 : XNOR2_X1 port map( A => n9936, B => n10291, ZN => n8548);
   U15657 : NOR2_X1 port map( A1 => n8537, A2 => n8734, ZN => n8540);
   U15659 : OAI211_X1 port map( C1 => n9045, C2 => n9047, A => n9237, B => 
                           n9233, ZN => n8543);
   U15660 : OAI211_X1 port map( C1 => n8544, C2 => n9045, A => n8543, B => 
                           n9238, ZN => n10029);
   U15661 : XNOR2_X1 port map( A => n9626, B => n10029, ZN => n8546);
   U15662 : XNOR2_X1 port map( A => n9447, B => n3336, ZN => n8545);
   U15663 : XNOR2_X1 port map( A => n8546, B => n8545, ZN => n8547);
   U15664 : XNOR2_X1 port map( A => n8548, B => n8547, ZN => n10747);
   U15665 : INV_X1 port map( A => n10747, ZN => n11197);
   U15666 : INV_X1 port map( A => n8550, ZN => n9137);
   U15667 : INV_X1 port map( A => n9340, ZN => n8924);
   U15668 : MUX2_X1 port map( A => n8550, B => n8549, S => n7410, Z => n8551);
   U15669 : XNOR2_X1 port map( A => n9851, B => n9504, ZN => n8559);
   U15670 : NAND2_X1 port map( A1 => n8553, A2 => n8941, ZN => n8554);
   U15671 : NAND3_X1 port map( A1 => n8557, A2 => n8765, A3 => n8554, ZN => 
                           n8556);
   U15672 : NAND3_X1 port map( A1 => n8945, A2 => n9562, A3 => n10401, ZN => 
                           n8555);
   U15673 : OAI211_X1 port map( C1 => n8557, C2 => n8945, A => n8556, B => 
                           n8555, ZN => n10434);
   U15674 : XNOR2_X1 port map( A => n10434, B => n3457, ZN => n8558);
   U15675 : XNOR2_X1 port map( A => n8559, B => n8558, ZN => n8573);
   U15676 : NAND3_X1 port map( A1 => n9144, A2 => n8563, A3 => n9139, ZN => 
                           n8566);
   U15677 : INV_X1 port map( A => n8185, ZN => n8564);
   U15678 : INV_X1 port map( A => n10436, ZN => n8572);
   U15679 : INV_X1 port map( A => n9149, ZN => n8931);
   U15680 : NAND2_X1 port map( A1 => n8760, A2 => n8931, ZN => n9152);
   U15681 : OAI211_X1 port map( C1 => n8570, C2 => n8760, A => n8930, B => 
                           n9152, ZN => n9378);
   U15682 : XNOR2_X1 port map( A => n8572, B => n10311, ZN => n9668);
   U15683 : AND2_X1 port map( A1 => n8574, A2 => n603, ZN => n9419);
   U15684 : INV_X1 port map( A => n9531, ZN => n8751);
   U15685 : XNOR2_X1 port map( A => n9763, B => n10359, ZN => n9940);
   U15686 : NAND2_X1 port map( A1 => n8580, A2 => n8579, ZN => n8583);
   U15687 : OAI21_X1 port map( B1 => n8828, B2 => n8826, A => n8824, ZN => 
                           n8585);
   U15688 : AOI22_X1 port map( A1 => n8585, A2 => n8584, B1 => n1839, B2 => 
                           n8828, ZN => n8588);
   U15689 : OR2_X1 port map( A1 => n8588, A2 => n8587, ZN => n9645);
   U15690 : XNOR2_X1 port map( A => n9645, B => n1878, ZN => n8602);
   U15691 : NAND2_X1 port map( A1 => n8977, A2 => n8589, ZN => n8973);
   U15692 : NAND2_X1 port map( A1 => n8594, A2 => n8978, ZN => n8590);
   U15694 : NAND2_X1 port map( A1 => n8591, A2 => n8817, ZN => n8595);
   U15695 : NAND2_X1 port map( A1 => n8593, A2 => n8592, ZN => n8818);
   U15696 : OAI21_X1 port map( B1 => n8595, B2 => n8594, A => n8818, ZN => 
                           n8596);
   U15697 : NAND3_X1 port map( A1 => n9064, A2 => n8872, A3 => n8865, ZN => 
                           n8599);
   U15698 : AND2_X1 port map( A1 => n8599, A2 => n8598, ZN => n8600);
   U15699 : XNOR2_X1 port map( A => n10285, B => n8602, ZN => n8621);
   U15700 : NOR2_X1 port map( A1 => n9080, A2 => n8603, ZN => n10234);
   U15701 : NAND2_X1 port map( A1 => n10234, A2 => n8724, ZN => n8604);
   U15702 : OAI21_X1 port map( B1 => n8724, B2 => n10240, A => n8604, ZN => 
                           n10245);
   U15703 : NAND2_X1 port map( A1 => n8848, A2 => n28500, ZN => n10237);
   U15704 : INV_X1 port map( A => n10237, ZN => n8607);
   U15705 : OR3_X2 port map( A1 => n10245, A2 => n8607, A3 => n8606, ZN => 
                           n9749);
   U15706 : NAND2_X1 port map( A1 => n8610, A2 => n9530, ZN => n8752);
   U15707 : NAND3_X1 port map( A1 => n9531, A2 => n8609, A3 => n9530, ZN => 
                           n8613);
   U15709 : INV_X1 port map( A => n8857, ZN => n8742);
   U15710 : NAND2_X1 port map( A1 => n9075, A2 => n9070, ZN => n8616);
   U15711 : NAND2_X1 port map( A1 => n9075, A2 => n8857, ZN => n8615);
   U15712 : NAND2_X1 port map( A1 => n9071, A2 => n8740, ZN => n8614);
   U15713 : NAND4_X1 port map( A1 => n8617, A2 => n8616, A3 => n8615, A4 => 
                           n8614, ZN => n8618);
   U15714 : XNOR2_X1 port map( A => n10043, B => n3662, ZN => n8619);
   U15715 : XNOR2_X1 port map( A => n9946, B => n8619, ZN => n8620);
   U15716 : NAND3_X1 port map( A1 => n3585, A2 => n10563, A3 => n28207, ZN => 
                           n8622);
   U15718 : NAND2_X1 port map( A1 => n8802, A2 => n8955, ZN => n8804);
   U15719 : XNOR2_X1 port map( A => n9306, B => n1246, ZN => n8626);
   U15720 : XNOR2_X1 port map( A => n8626, B => n1877, ZN => n8639);
   U15721 : INV_X1 port map( A => n9095, ZN => n8627);
   U15723 : NAND3_X1 port map( A1 => n9099, A2 => n8627, A3 => n8666, ZN => 
                           n8628);
   U15724 : NAND2_X1 port map( A1 => n8629, A2 => n8628, ZN => n8633);
   U15725 : AOI21_X1 port map( B1 => n8631, B2 => n9100, A => n8630, ZN => 
                           n8632);
   U15726 : NAND2_X1 port map( A1 => n8634, A2 => n8635, ZN => n8638);
   U15727 : NAND3_X1 port map( A1 => n8635, A2 => n8656, A3 => n8655, ZN => 
                           n8637);
   U15728 : NAND3_X1 port map( A1 => n8653, A2 => n8652, A3 => n8658, ZN => 
                           n8636);
   U15729 : XNOR2_X1 port map( A => n9986, B => n10160, ZN => n8904);
   U15730 : XNOR2_X1 port map( A => n8904, B => n8639, ZN => n8649);
   U15731 : NAND2_X1 port map( A1 => n8836, A2 => n8966, ZN => n8842);
   U15732 : NAND3_X1 port map( A1 => n8963, A2 => n8962, A3 => n8838, ZN => 
                           n8641);
   U15733 : NAND2_X1 port map( A1 => n8836, A2 => n9171, ZN => n8965);
   U15734 : NAND2_X1 port map( A1 => n8982, A2 => n8642, ZN => n8643);
   U15735 : AOI21_X1 port map( B1 => n9398, B2 => n8644, A => n8982, ZN => 
                           n8645);
   U15736 : XNOR2_X1 port map( A => n9746, B => n10184, ZN => n8648);
   U15737 : OAI21_X1 port map( B1 => n9566, B2 => n9561, A => n8943, ZN => 
                           n10403);
   U15738 : NAND2_X1 port map( A1 => n10403, A2 => n8944, ZN => n10407);
   U15741 : INV_X1 port map( A => n10283, ZN => n8647);
   U15742 : OAI211_X1 port map( C1 => n1966, C2 => n12202, A => n11438, B => 
                           n8650, ZN => n9259);
   U15743 : OAI21_X1 port map( B1 => n8656, B2 => n8655, A => n8654, ZN => 
                           n8657);
   U15744 : INV_X1 port map( A => n8657, ZN => n8659);
   U15745 : XNOR2_X1 port map( A => n9614, B => n9915, ZN => n9660);
   U15746 : XNOR2_X1 port map( A => n10134, B => n9696, ZN => n10255);
   U15747 : XNOR2_X1 port map( A => n9660, B => n10255, ZN => n8677);
   U15748 : NAND2_X1 port map( A1 => n8665, A2 => n8664, ZN => n9098);
   U15749 : OAI21_X1 port map( B1 => n9100, B2 => n8665, A => n9098, ZN => 
                           n8667);
   U15750 : MUX2_X1 port map( A => n8670, B => n8669, S => n8914, Z => n8674);
   U15751 : MUX2_X1 port map( A => n8672, B => n8671, S => n8914, Z => n8673);
   U15752 : XNOR2_X1 port map( A => n10133, B => n10257, ZN => n9831);
   U15753 : XNOR2_X1 port map( A => n9698, B => n3191, ZN => n8675);
   U15754 : XNOR2_X1 port map( A => n9831, B => n8675, ZN => n8676);
   U15755 : XNOR2_X1 port map( A => n8676, B => n8677, ZN => n10558);
   U15756 : NAND2_X1 port map( A1 => n8810, A2 => n8811, ZN => n8678);
   U15757 : AOI21_X1 port map( B1 => n8679, B2 => n8678, A => n8812, ZN => 
                           n8684);
   U15758 : NAND2_X1 port map( A1 => n8680, A2 => n8809, ZN => n8682);
   U15760 : OAI21_X1 port map( B1 => n8682, B2 => n8810, A => n8814, ZN => 
                           n8683);
   U15761 : XNOR2_X1 port map( A => n9645, B => n9949, ZN => n8692);
   U15762 : NAND3_X1 port map( A1 => n8685, A2 => n9221, A3 => n9222, ZN => 
                           n8690);
   U15763 : NAND3_X1 port map( A1 => n8688, A2 => n8687, A3 => n8686, ZN => 
                           n8689);
   U15764 : NAND3_X1 port map( A1 => n9230, A2 => n9233, A3 => n9229, ZN => 
                           n8691);
   U15765 : XNOR2_X1 port map( A => n8692, B => n9603, ZN => n8707);
   U15766 : NAND2_X1 port map( A1 => n9042, A2 => n8693, ZN => n8696);
   U15767 : NAND2_X1 port map( A1 => n9041, A2 => n9247, ZN => n8695);
   U15768 : XNOR2_X1 port map( A => n10330, B => n10232, ZN => n9304);
   U15769 : INV_X1 port map( A => n9304, ZN => n8705);
   U15770 : INV_X1 port map( A => n8877, ZN => n8698);
   U15771 : NAND2_X1 port map( A1 => n8878, A2 => n8698, ZN => n8703);
   U15772 : NAND2_X1 port map( A1 => n8404, A2 => n8699, ZN => n8702);
   U15773 : NAND3_X1 port map( A1 => n8403, A2 => n8698, A3 => n8874, ZN => 
                           n8701);
   U15774 : NAND3_X1 port map( A1 => n8873, A2 => n8699, A3 => n8877, ZN => 
                           n8700);
   U15775 : XNOR2_X1 port map( A => n10231, B => n3180, ZN => n8704);
   U15776 : XNOR2_X1 port map( A => n8705, B => n8704, ZN => n8706);
   U15777 : NAND3_X1 port map( A1 => n8404, A2 => n8874, A3 => n8877, ZN => 
                           n8711);
   U15778 : NAND2_X1 port map( A1 => n8712, A2 => n8711, ZN => n8713);
   U15780 : XNOR2_X1 port map( A => n9963, B => n8715, ZN => n9705);
   U15781 : NAND2_X1 port map( A1 => n8719, A2 => n8718, ZN => n8722);
   U15782 : AOI21_X1 port map( B1 => n8722, B2 => n4321, A => n8720, ZN => 
                           n8723);
   U15783 : NAND2_X1 port map( A1 => n8848, A2 => n8726, ZN => n8725);
   U15784 : AOI21_X1 port map( B1 => n8850, B2 => n8725, A => n8724, ZN => 
                           n8728);
   U15785 : NAND2_X1 port map( A1 => n28500, A2 => n8726, ZN => n9078);
   U15786 : AOI21_X1 port map( B1 => n9078, B2 => n8848, A => n29311, ZN => 
                           n8727);
   U15787 : XNOR2_X1 port map( A => n10264, B => n9877, ZN => n9817);
   U15788 : XNOR2_X1 port map( A => n9705, B => n9817, ZN => n8746);
   U15789 : NOR2_X1 port map( A1 => n8730, A2 => n8729, ZN => n8732);
   U15790 : OAI21_X1 port map( B1 => n8732, B2 => n8731, A => n8739, ZN => 
                           n8737);
   U15791 : AOI22_X1 port map( A1 => n8856, A2 => n9075, B1 => n8740, B2 => 
                           n8741, ZN => n8743);
   U15792 : XNOR2_X1 port map( A => n9931, B => n10265, ZN => n9742);
   U15793 : XNOR2_X1 port map( A => n9656, B => n3323, ZN => n8744);
   U15794 : XNOR2_X1 port map( A => n9742, B => n8744, ZN => n8745);
   U15795 : MUX2_X1 port map( A => n11345, B => n1898, S => n11334, Z => n8846)
                           ;
   U15796 : NAND3_X1 port map( A1 => n9529, A2 => n29395, A3 => n29662, ZN => 
                           n8750);
   U15797 : NAND2_X1 port map( A1 => n9133, A2 => n9340, ZN => n8754);
   U15798 : NOR2_X1 port map( A1 => n9341, A2 => n8756, ZN => n8757);
   U15799 : XNOR2_X1 port map( A => n10149, B => n8757, ZN => n9842);
   U15800 : NAND3_X1 port map( A1 => n9148, A2 => n6747, A3 => n11, ZN => n8758
                           );
   U15801 : MUX2_X1 port map( A => n8762, B => n8945, S => n8941, Z => n8766);
   U15802 : XNOR2_X1 port map( A => n9710, B => n10151, ZN => n10252);
   U15803 : XNOR2_X1 port map( A => n10252, B => n9842, ZN => n8775);
   U15805 : XNOR2_X1 port map( A => n9678, B => n9908, ZN => n8773);
   U15806 : INV_X1 port map( A => n1123, ZN => n26656);
   U15808 : XNOR2_X1 port map( A => n8773, B => n8772, ZN => n8774);
   U15809 : INV_X1 port map( A => n11337, ZN => n11174);
   U15810 : NOR2_X1 port map( A1 => n8995, A2 => n9210, ZN => n8776);
   U15814 : XNOR2_X1 port map( A => n9446, B => n10218, ZN => n9836);
   U15815 : NAND2_X1 port map( A1 => n9188, A2 => n8782, ZN => n9006);
   U15816 : NAND3_X1 port map( A1 => n9187, A2 => n9009, A3 => n9007, ZN => 
                           n8783);
   U15817 : XNOR2_X1 port map( A => n9992, B => n9716, ZN => n9310);
   U15818 : XNOR2_X1 port map( A => n9310, B => n9836, ZN => n8799);
   U15819 : OAI211_X1 port map( C1 => n8788, C2 => n8787, A => n8786, B => 
                           n8785, ZN => n8789);
   U15820 : XNOR2_X1 port map( A => n9626, B => n9934, ZN => n8797);
   U15821 : INV_X1 port map( A => n2353, ZN => n25378);
   U15822 : XNOR2_X1 port map( A => n301, B => n25378, ZN => n8796);
   U15823 : XNOR2_X1 port map( A => n8797, B => n8796, ZN => n8798);
   U15824 : XNOR2_X1 port map( A => n8799, B => n8798, ZN => n10830);
   U15825 : AND2_X1 port map( A1 => n8957, A2 => n8803, ZN => n8807);
   U15826 : MUX2_X1 port map( A => n8805, B => n8804, S => n8958, Z => n8806);
   U15827 : OAI21_X2 port map( B1 => n8807, B2 => n29096, A => n8806, ZN => 
                           n10275);
   U15829 : XNOR2_X1 port map( A => n9852, B => n10275, ZN => n9591);
   U15830 : INV_X1 port map( A => n8818, ZN => n8820);
   U15831 : NAND2_X1 port map( A1 => n8820, A2 => n8819, ZN => n8821);
   U15832 : NAND3_X1 port map( A1 => n1839, A2 => n8826, A3 => n8825, ZN => 
                           n8833);
   U15833 : NAND3_X1 port map( A1 => n8830, A2 => n8829, A3 => n8828, ZN => 
                           n8831);
   U15834 : XNOR2_X1 port map( A => n9591, B => n8835, ZN => n8845);
   U15835 : NOR2_X1 port map( A1 => n8837, A2 => n8836, ZN => n8840);
   U15836 : NOR2_X1 port map( A1 => n8966, A2 => n8838, ZN => n8839);
   U15837 : NAND3_X1 port map( A1 => n8964, A2 => n605, A3 => n9170, ZN => 
                           n8841);
   U15838 : INV_X1 port map( A => n2889, ZN => n27778);
   U15839 : XNOR2_X1 port map( A => n10436, B => n27778, ZN => n8843);
   U15840 : INV_X1 port map( A => n8847, ZN => n11702);
   U15841 : NAND2_X1 port map( A1 => n11702, A2 => n12202, ZN => n9058);
   U15842 : OAI21_X1 port map( B1 => n28500, B2 => n8848, A => n2320, ZN => 
                           n8849);
   U15843 : NAND3_X1 port map( A1 => n8852, A2 => n29311, A3 => n8851, ZN => 
                           n8853);
   U15846 : OAI21_X2 port map( B1 => n8862, B2 => n8861, A => n8860, ZN => 
                           n10385);
   U15847 : XNOR2_X1 port map( A => n10385, B => n9619, ZN => n10177);
   U15848 : XNOR2_X1 port map( A => n10321, B => n2350, ZN => n8863);
   U15849 : NAND3_X1 port map( A1 => n9062, A2 => n8864, A3 => n9064, ZN => 
                           n8870);
   U15850 : NAND2_X1 port map( A1 => n9062, A2 => n8865, ZN => n8867);
   U15851 : NAND3_X1 port map( A1 => n8868, A2 => n8867, A3 => n8866, ZN => 
                           n8869);
   U15852 : MUX2_X1 port map( A => n8403, B => n8876, S => n8874, Z => n8882);
   U15853 : NAND3_X1 port map( A1 => n8403, A2 => n8876, A3 => n8875, ZN => 
                           n8880);
   U15854 : NAND2_X1 port map( A1 => n8878, A2 => n8877, ZN => n8879);
   U15855 : XNOR2_X1 port map( A => n8884, B => n8885, ZN => n10473);
   U15856 : INV_X1 port map( A => n10473, ZN => n11323);
   U15857 : OAI22_X1 port map( A1 => n8888, A2 => n8887, B1 => n8886, B2 => 
                           n8890, ZN => n8895);
   U15858 : NAND2_X1 port map( A1 => n8890, A2 => n8889, ZN => n8893);
   U15859 : INV_X1 port map( A => n9824, ZN => n8896);
   U15860 : XNOR2_X1 port map( A => n10282, B => n8896, ZN => n8903);
   U15861 : INV_X1 port map( A => n9125, ZN => n8897);
   U15862 : NAND2_X1 port map( A1 => n8900, A2 => n8899, ZN => n8901);
   U15863 : XNOR2_X1 port map( A => n8902, B => n8903, ZN => n8923);
   U15864 : INV_X1 port map( A => n8904, ZN => n8921);
   U15865 : INV_X1 port map( A => n9012, ZN => n8905);
   U15866 : AND2_X1 port map( A1 => n8907, A2 => n8906, ZN => n8913);
   U15867 : NAND2_X1 port map( A1 => n8908, A2 => n9012, ZN => n8909);
   U15868 : OAI21_X1 port map( B1 => n608, B2 => n9012, A => n8909, ZN => n8911
                           );
   U15869 : NAND2_X1 port map( A1 => n8911, A2 => n8910, ZN => n8912);
   U15870 : NAND2_X1 port map( A1 => n8913, A2 => n8912, ZN => n10411);
   U15871 : NAND2_X1 port map( A1 => n8916, A2 => n8915, ZN => n8919);
   U15872 : AND2_X1 port map( A1 => n8917, A2 => n9107, ZN => n8918);
   U15873 : XNOR2_X1 port map( A => n10411, B => n9647, ZN => n9903);
   U15874 : XNOR2_X1 port map( A => n8921, B => n9903, ZN => n8922);
   U15876 : NAND2_X1 port map( A1 => n11323, A2 => n10810, ZN => n10859);
   U15877 : OAI21_X1 port map( B1 => n9133, B2 => n9134, A => n8924, ZN => 
                           n8927);
   U15879 : XNOR2_X1 port map( A => n10202, B => n3650, ZN => n8928);
   U15880 : XNOR2_X1 port map( A => n9779, B => n8928, ZN => n8940);
   U15881 : NAND2_X1 port map( A1 => n6747, A2 => n8929, ZN => n9147);
   U15882 : NAND2_X1 port map( A1 => n8931, A2 => n9148, ZN => n8934);
   U15883 : NAND2_X1 port map( A1 => n9374, A2 => n5958, ZN => n8932);
   U15884 : AOI21_X2 port map( B1 => n8935, B2 => n8934, A => n8933, ZN => 
                           n10396);
   U15885 : XNOR2_X1 port map( A => n10396, B => n1868, ZN => n9523);
   U15886 : XNOR2_X1 port map( A => n9996, B => n10289, ZN => n8951);
   U15887 : NOR2_X1 port map( A1 => n8941, A2 => n9561, ZN => n8942);
   U15888 : AOI21_X1 port map( B1 => n8947, B2 => n8943, A => n8942, ZN => 
                           n8949);
   U15889 : NAND2_X1 port map( A1 => n8945, A2 => n8944, ZN => n8946);
   U15890 : NOR2_X1 port map( A1 => n8947, A2 => n8946, ZN => n8948);
   U15891 : INV_X1 port map( A => n10371, ZN => n8950);
   U15892 : XNOR2_X1 port map( A => n8951, B => n8950, ZN => n8952);
   U15893 : INV_X1 port map( A => n10472, ZN => n11184);
   U15894 : INV_X1 port map( A => n8953, ZN => n8972);
   U15895 : MUX2_X1 port map( A => n8956, B => n8955, S => n29096, Z => n8960);
   U15896 : NOR2_X1 port map( A1 => n8962, A2 => n8961, ZN => n8971);
   U15897 : OAI21_X1 port map( B1 => n8964, B2 => n8963, A => n605, ZN => n8970
                           );
   U15898 : OAI21_X1 port map( B1 => n605, B2 => n8966, A => n8965, ZN => n8969
                           );
   U15899 : INV_X1 port map( A => n8967, ZN => n8968);
   U15900 : INV_X1 port map( A => n9540, ZN => n10419);
   U15901 : XNOR2_X1 port map( A => n10419, B => n9613, ZN => n9872);
   U15902 : XNOR2_X1 port map( A => n9872, B => n8972, ZN => n8991);
   U15903 : XNOR2_X1 port map( A => n10294, B => n2982, ZN => n8989);
   U15904 : INV_X1 port map( A => n8973, ZN => n8975);
   U15905 : NAND2_X1 port map( A1 => n607, A2 => n8978, ZN => n8979);
   U15906 : NAND3_X1 port map( A1 => n8982, A2 => n8981, A3 => n8980, ZN => 
                           n8986);
   U15908 : INV_X1 port map( A => n10258, ZN => n9528);
   U15909 : XNOR2_X1 port map( A => n9528, B => n10345, ZN => n9833);
   U15910 : XNOR2_X1 port map( A => n8989, B => n9833, ZN => n8990);
   U15911 : NAND3_X1 port map( A1 => n10859, A2 => n8992, A3 => n11322, ZN => 
                           n9056);
   U15912 : NAND3_X1 port map( A1 => n9434, A2 => n8996, A3 => n4305, ZN => 
                           n8997);
   U15913 : NAND2_X1 port map( A1 => n9196, A2 => n9206, ZN => n8999);
   U15914 : AND2_X1 port map( A1 => n8999, A2 => n9197, ZN => n9002);
   U15915 : XNOR2_X1 port map( A => n10189, B => n9003, ZN => n9022);
   U15916 : NAND2_X1 port map( A1 => n9009, A2 => n9007, ZN => n9005);
   U15917 : AOI21_X1 port map( B1 => n9006, B2 => n9005, A => n9004, ZN => 
                           n9011);
   U15918 : NAND2_X1 port map( A1 => n9184, A2 => n9007, ZN => n9008);
   U15919 : AOI21_X1 port map( B1 => n9009, B2 => n9008, A => n9188, ZN => 
                           n9010);
   U15920 : NAND3_X1 port map( A1 => n9013, A2 => n9012, A3 => n9014, ZN => 
                           n9017);
   U15921 : XNOR2_X1 port map( A => n9512, B => n10362, ZN => n9820);
   U15922 : XNOR2_X1 port map( A => n10304, B => n2598, ZN => n9020);
   U15923 : XNOR2_X1 port map( A => n9820, B => n9020, ZN => n9021);
   U15924 : NAND2_X1 port map( A1 => n9222, A2 => n9220, ZN => n9023);
   U15925 : NAND2_X1 port map( A1 => n597, A2 => n9023, ZN => n9025);
   U15927 : NOR2_X1 port map( A1 => n9035, A2 => n9034, ZN => n9036);
   U15928 : NAND2_X1 port map( A1 => n9037, A2 => n9036, ZN => n9038);
   U15929 : NOR2_X1 port map( A1 => n9039, A2 => n8109, ZN => n9040);
   U15931 : INV_X1 port map( A => n9849, ZN => n9044);
   U15932 : XNOR2_X1 port map( A => n9044, B => n9631, ZN => n9053);
   U15933 : XNOR2_X1 port map( A => n9592, B => n10071, ZN => n9051);
   U15934 : XNOR2_X1 port map( A => n10435, B => n3321, ZN => n9050);
   U15935 : XNOR2_X1 port map( A => n9051, B => n9050, ZN => n9052);
   U15936 : NAND3_X1 port map( A1 => n11187, A2 => n11181, A3 => n11321, ZN => 
                           n9054);
   U15937 : NAND2_X1 port map( A1 => n12205, A2 => n12200, ZN => n9057);
   U15939 : MUX2_X1 port map( A => n9059, B => n9060, S => n9062, Z => n9065);
   U15940 : XNOR2_X1 port map( A => n10258, B => n2509, ZN => n9066);
   U15941 : XNOR2_X1 port map( A => n9066, B => n1891, ZN => n9068);
   U15942 : XNOR2_X1 port map( A => n10297, B => n1902, ZN => n9067);
   U15943 : XNOR2_X1 port map( A => n9068, B => n9067, ZN => n9093);
   U15944 : OAI21_X1 port map( B1 => n9071, B2 => n9070, A => n9069, ZN => 
                           n9077);
   U15945 : OAI21_X1 port map( B1 => n9074, B2 => n9073, A => n9072, ZN => 
                           n9076);
   U15946 : OAI21_X1 port map( B1 => n9079, B2 => n28500, A => n9078, ZN => 
                           n9091);
   U15947 : NAND2_X1 port map( A1 => n28500, A2 => n29310, ZN => n9089);
   U15948 : INV_X1 port map( A => n9082, ZN => n9086);
   U15949 : INV_X1 port map( A => n9083, ZN => n9085);
   U15950 : OAI21_X1 port map( B1 => n9086, B2 => n9085, A => n9084, ZN => 
                           n9087);
   U15951 : NAND2_X1 port map( A1 => n9089, A2 => n9088, ZN => n9090);
   U15952 : XNOR2_X1 port map( A => n9695, B => n10344, ZN => n10057);
   U15953 : XNOR2_X1 port map( A => n1920, B => n10057, ZN => n9092);
   U15954 : INV_X1 port map( A => n9094, ZN => n9462);
   U15955 : OAI21_X1 port map( B1 => n9097, B2 => n9096, A => n9095, ZN => 
                           n9103);
   U15956 : INV_X1 port map( A => n9098, ZN => n9101);
   U15957 : OAI21_X1 port map( B1 => n9101, B2 => n9100, A => n9099, ZN => 
                           n9102);
   U15958 : NAND2_X1 port map( A1 => n9103, A2 => n9102, ZN => n10363);
   U15959 : INV_X1 port map( A => n9107, ZN => n9104);
   U15960 : NAND3_X1 port map( A1 => n9108, A2 => n9118, A3 => n9107, ZN => 
                           n9120);
   U15961 : INV_X1 port map( A => n9109, ZN => n9111);
   U15962 : NAND2_X1 port map( A1 => n9111, A2 => n28810, ZN => n9117);
   U15963 : INV_X1 port map( A => n9112, ZN => n9114);
   U15964 : NAND2_X1 port map( A1 => n9114, A2 => n29135, ZN => n9115);
   U15965 : NAND4_X1 port map( A1 => n9118, A2 => n9117, A3 => n9116, A4 => 
                           n9115, ZN => n9119);
   U15966 : XNOR2_X1 port map( A => n9462, B => n10086, ZN => n9130);
   U15967 : AOI22_X1 port map( A1 => n9125, A2 => n9124, B1 => n29304, B2 => 
                           n9122, ZN => n9126);
   U15968 : INV_X1 port map( A => n9512, ZN => n9881);
   U15969 : XNOR2_X1 port map( A => n9794, B => n9881, ZN => n9128);
   U15970 : XNOR2_X1 port map( A => n9964, B => n3232, ZN => n9127);
   U15971 : XNOR2_X1 port map( A => n9128, B => n9127, ZN => n9129);
   U15972 : AND2_X1 port map( A1 => n9132, A2 => n9133, ZN => n9135);
   U15973 : XNOR2_X1 port map( A => n1877, B => n10283, ZN => n9138);
   U15974 : XNOR2_X1 port map( A => n10332, B => n9138, ZN => n9159);
   U15975 : OAI21_X1 port map( B1 => n598, B2 => n9142, A => n9141, ZN => n9143
                           );
   U15976 : XNOR2_X1 port map( A => n10159, B => n9824, ZN => n9157);
   U15977 : INV_X1 port map( A => n9147, ZN => n9154);
   U15978 : AOI21_X1 port map( B1 => n6747, B2 => n9149, A => n9148, ZN => 
                           n9151);
   U15979 : NAND2_X1 port map( A1 => n9152, A2 => n9151, ZN => n9153);
   U15980 : XNOR2_X1 port map( A => n1918, B => n27452, ZN => n9156);
   U15981 : XNOR2_X1 port map( A => n9157, B => n9156, ZN => n9158);
   U15982 : OAI21_X1 port map( B1 => n9161, B2 => n9160, A => n9164, ZN => 
                           n9168);
   U15983 : INV_X1 port map( A => n9162, ZN => n9166);
   U15984 : NAND2_X1 port map( A1 => n9164, A2 => n9163, ZN => n9165);
   U15985 : INV_X1 port map( A => n9357, ZN => n9175);
   U15986 : XNOR2_X1 port map( A => n9175, B => n10373, ZN => n9182);
   U15987 : INV_X1 port map( A => n9176, ZN => n9178);
   U15988 : XNOR2_X1 port map( A => n9684, B => n10395, ZN => n9450);
   U15989 : XNOR2_X1 port map( A => n1868, B => n3035, ZN => n9180);
   U15990 : XNOR2_X1 port map( A => n9450, B => n9180, ZN => n9181);
   U15991 : NAND2_X1 port map( A1 => n10847, A2 => n11347, ZN => n9219);
   U15992 : XNOR2_X1 port map( A => n9504, B => n26909, ZN => n9183);
   U15993 : XNOR2_X1 port map( A => n9183, B => n10271, ZN => n9193);
   U15994 : MUX2_X1 port map( A => n9188, B => n9187, S => n9184, Z => n9192);
   U15997 : XNOR2_X1 port map( A => n10072, B => n10353, ZN => n9811);
   U15998 : XNOR2_X1 port map( A => n9811, B => n9193, ZN => n9217);
   U15999 : NAND2_X1 port map( A1 => n9195, A2 => n9194, ZN => n9205);
   U16000 : NOR2_X1 port map( A1 => n9196, A2 => n9200, ZN => n9198);
   U16001 : OAI21_X1 port map( B1 => n9199, B2 => n9198, A => n9197, ZN => 
                           n9204);
   U16002 : NAND3_X1 port map( A1 => n9202, A2 => n9201, A3 => n9200, ZN => 
                           n9203);
   U16003 : OAI211_X1 port map( C1 => n9206, C2 => n9205, A => n9204, B => 
                           n9203, ZN => n9629);
   U16004 : INV_X1 port map( A => n9207, ZN => n9215);
   U16005 : OAI21_X1 port map( B1 => n9209, B2 => n4305, A => n9208, ZN => 
                           n9214);
   U16006 : NAND3_X1 port map( A1 => n9211, A2 => n9210, A3 => n4305, ZN => 
                           n9213);
   U16007 : NAND3_X1 port map( A1 => n9434, A2 => n9436, A3 => n9438, ZN => 
                           n9212);
   U16009 : XNOR2_X1 port map( A => n10356, B => n9629, ZN => n10432);
   U16010 : XNOR2_X1 port map( A => n10432, B => n10359, ZN => n9216);
   U16012 : INV_X1 port map( A => n11349, ZN => n9218);
   U16013 : NAND3_X1 port map( A1 => n9224, A2 => n9223, A3 => n9228, ZN => 
                           n9225);
   U16014 : NOR2_X1 port map( A1 => n9229, A2 => n9233, ZN => n9231);
   U16015 : INV_X1 port map( A => n9232, ZN => n9234);
   U16016 : OAI21_X1 port map( B1 => n9238, B2 => n9237, A => n9236, ZN => 
                           n9239);
   U16018 : XNOR2_X1 port map( A => n10251, B => n10384, ZN => n9241);
   U16019 : NAND2_X1 port map( A1 => n9246, A2 => n9245, ZN => n9250);
   U16020 : XNOR2_X1 port map( A => n9677, B => n9976, ZN => n9253);
   U16021 : XNOR2_X1 port map( A => n9550, B => n3625, ZN => n9252);
   U16022 : XNOR2_X1 port map( A => n9253, B => n9252, ZN => n9254);
   U16023 : NAND2_X1 port map( A1 => n10476, A2 => n11347, ZN => n10477);
   U16024 : AOI21_X1 port map( B1 => n10477, B2 => n10847, A => n11192, ZN => 
                           n9256);
   U16025 : MUX2_X2 port map( A => n9259, B => n9258, S => n5825, Z => n12738);
   U16026 : XNOR2_X1 port map( A => n12738, B => n3015, ZN => n9478);
   U16027 : XNOR2_X1 port map( A => n9763, B => n9629, ZN => n9260);
   U16028 : XNOR2_X1 port map( A => n9849, B => n9260, ZN => n9264);
   U16029 : XNOR2_X1 port map( A => n9509, B => n9852, ZN => n10127);
   U16030 : INV_X1 port map( A => n10127, ZN => n9262);
   U16031 : XNOR2_X1 port map( A => n10071, B => n3722, ZN => n9261);
   U16032 : XNOR2_X1 port map( A => n9262, B => n9261, ZN => n9263);
   U16034 : INV_X1 port map( A => n9820, ZN => n9265);
   U16035 : XNOR2_X1 port map( A => n9929, B => n9877, ZN => n10119);
   U16036 : XNOR2_X1 port map( A => n9265, B => n10119, ZN => n9270);
   U16037 : XNOR2_X1 port map( A => n9930, B => n1923, ZN => n9267);
   U16038 : XNOR2_X1 port map( A => n9268, B => n9267, ZN => n9269);
   U16040 : INV_X1 port map( A => n10941, ZN => n10110);
   U16041 : XNOR2_X1 port map( A => n10371, B => n10391, ZN => n10079);
   U16042 : XNOR2_X1 port map( A => n9755, B => n9894, ZN => n10220);
   U16043 : XNOR2_X1 port map( A => n10145, B => n3196, ZN => n9271);
   U16044 : XNOR2_X1 port map( A => n10220, B => n9271, ZN => n9272);
   U16045 : INV_X1 port map( A => n10940, ZN => n10446);
   U16046 : XNOR2_X1 port map( A => n9824, B => n9948, ZN => n9520);
   U16047 : XNOR2_X1 port map( A => n10328, B => n10412, ZN => n10065);
   U16048 : INV_X1 port map( A => n10065, ZN => n9646);
   U16049 : XNOR2_X1 port map( A => n9646, B => n9520, ZN => n9276);
   U16050 : XNOR2_X1 port map( A => n9749, B => n9899, ZN => n9274);
   U16051 : XNOR2_X1 port map( A => n10160, B => n27956, ZN => n9273);
   U16052 : XNOR2_X1 port map( A => n9274, B => n9273, ZN => n9275);
   U16053 : NAND2_X1 port map( A1 => n10446, A2 => n10703, ZN => n9281);
   U16054 : XNOR2_X1 port map( A => n9918, B => n9833, ZN => n9280);
   U16055 : XNOR2_X1 port map( A => n9695, B => n10133, ZN => n9278);
   U16056 : XNOR2_X1 port map( A => n9799, B => n3369, ZN => n9277);
   U16057 : XNOR2_X1 port map( A => n9278, B => n9277, ZN => n9279);
   U16059 : XNOR2_X1 port map( A => n10251, B => n1884, ZN => n9283);
   U16060 : INV_X1 port map( A => n9352, ZN => n9711);
   U16061 : XNOR2_X1 port map( A => n10149, B => n9711, ZN => n9282);
   U16062 : XNOR2_X1 port map( A => n9282, B => n9283, ZN => n9288);
   U16063 : XNOR2_X1 port map( A => n1852, B => n27231, ZN => n9286);
   U16064 : XNOR2_X1 port map( A => n28488, B => n9771, ZN => n9285);
   U16065 : XNOR2_X1 port map( A => n9286, B => n9285, ZN => n9287);
   U16067 : NOR2_X1 port map( A1 => n10705, A2 => n10942, ZN => n10704);
   U16068 : INV_X1 port map( A => n10704, ZN => n9290);
   U16069 : AOI21_X1 port map( B1 => n10942, B2 => n10110, A => n10703, ZN => 
                           n9289);
   U16070 : NAND2_X1 port map( A1 => n9290, A2 => n9289, ZN => n9291);
   U16072 : XNOR2_X1 port map( A => n9710, B => n10335, ZN => n9293);
   U16073 : XNOR2_X1 port map( A => n10319, B => n9293, ZN => n9297);
   U16074 : INV_X1 port map( A => n3164, ZN => n9294);
   U16075 : XNOR2_X1 port map( A => n10178, B => n9294, ZN => n9296);
   U16076 : XNOR2_X1 port map( A => n10356, B => n2527, ZN => n9298);
   U16077 : XNOR2_X1 port map( A => n9956, B => n9298, ZN => n9300);
   U16078 : XNOR2_X1 port map( A => n9851, B => n9941, ZN => n10315);
   U16079 : XNOR2_X1 port map( A => n10315, B => n9590, ZN => n9299);
   U16080 : XNOR2_X1 port map( A => n10038, B => n9971, ZN => n9302);
   U16081 : XNOR2_X1 port map( A => n10183, B => n3422, ZN => n9303);
   U16082 : XNOR2_X1 port map( A => n9303, B => n10064, ZN => n9305);
   U16083 : XNOR2_X1 port map( A => n9305, B => n9304, ZN => n9308);
   U16084 : XNOR2_X1 port map( A => n9949, B => n10043, ZN => n9307);
   U16086 : XNOR2_X1 port map( A => n9307, B => n9725, ZN => n10286);
   U16087 : XNOR2_X1 port map( A => n9308, B => n10286, ZN => n10973);
   U16089 : XNOR2_X1 port map( A => n9818, B => n9705, ZN => n9309);
   U16090 : XNOR2_X1 port map( A => n9311, B => n9310, ZN => n9317);
   U16091 : XNOR2_X1 port map( A => n10143, B => n857, ZN => n9315);
   U16092 : XNOR2_X1 port map( A => n5412, B => n9997, ZN => n9314);
   U16093 : XNOR2_X1 port map( A => n9315, B => n9314, ZN => n9316);
   U16095 : XNOR2_X1 port map( A => n10088, B => n9930, ZN => n10268);
   U16096 : INV_X1 port map( A => n10268, ZN => n9319);
   U16097 : INV_X1 port map( A => n10264, ZN => n9318);
   U16098 : XNOR2_X1 port map( A => n9319, B => n9962, ZN => n9322);
   U16099 : XNOR2_X1 port map( A => n9878, B => n10304, ZN => n9741);
   U16100 : XNOR2_X1 port map( A => n10426, B => n1161, ZN => n9320);
   U16101 : XNOR2_X1 port map( A => n9741, B => n9320, ZN => n9321);
   U16102 : XNOR2_X1 port map( A => n9322, B => n9321, ZN => n9344);
   U16103 : INV_X1 port map( A => n9344, ZN => n10605);
   U16104 : XNOR2_X1 port map( A => n9735, B => n9323, ZN => n10256);
   U16105 : INV_X1 port map( A => n10256, ZN => n9324);
   U16106 : XNOR2_X1 port map( A => n9324, B => n9736, ZN => n9328);
   U16107 : XNOR2_X1 port map( A => n10257, B => n9971, ZN => n9326);
   U16108 : XNOR2_X1 port map( A => n10419, B => n2981, ZN => n9325);
   U16109 : XNOR2_X1 port map( A => n9325, B => n9326, ZN => n9327);
   U16110 : NAND2_X1 port map( A1 => n10605, A2 => n10913, ZN => n10732);
   U16111 : INV_X1 port map( A => n10732, ZN => n9333);
   U16112 : XNOR2_X1 port map( A => n10128, B => n9592, ZN => n9767);
   U16113 : XNOR2_X1 port map( A => n10277, B => n9767, ZN => n9332);
   U16114 : XNOR2_X1 port map( A => n10275, B => n10310, ZN => n9330);
   U16115 : XNOR2_X1 port map( A => n10435, B => n3752, ZN => n9329);
   U16116 : XNOR2_X1 port map( A => n9330, B => n9329, ZN => n9331);
   U16117 : XNOR2_X1 port map( A => n9332, B => n9331, ZN => n10735);
   U16118 : INV_X1 port map( A => n10735, ZN => n10914);
   U16119 : NAND2_X1 port map( A1 => n9333, A2 => n10914, ZN => n11526);
   U16120 : XNOR2_X1 port map( A => n9997, B => n9755, ZN => n9335);
   U16121 : XNOR2_X1 port map( A => n10289, B => n2274, ZN => n9334);
   U16122 : XNOR2_X1 port map( A => n9335, B => n9334, ZN => n9338);
   U16123 : XNOR2_X1 port map( A => n10396, B => n10218, ZN => n9780);
   U16124 : INV_X1 port map( A => n10912, ZN => n10689);
   U16125 : XNOR2_X1 port map( A => n10322, B => n28693, ZN => n9339);
   U16126 : XNOR2_X1 port map( A => n9771, B => n9979, ZN => n9342);
   U16127 : XNOR2_X1 port map( A => n9342, B => n10060, ZN => n10253);
   U16128 : XNOR2_X2 port map( A => n9343, B => n10253, ZN => n10911);
   U16129 : NAND2_X1 port map( A1 => n10689, A2 => n10911, ZN => n10733);
   U16130 : INV_X1 port map( A => n10913, ZN => n10609);
   U16131 : OAI211_X1 port map( C1 => n10605, C2 => n10689, A => n10733, B => 
                           n10609, ZN => n11525);
   U16132 : XNOR2_X1 port map( A => n9749, B => n9823, ZN => n9491);
   U16133 : XNOR2_X1 port map( A => n9748, B => n9491, ZN => n9347);
   U16134 : XNOR2_X1 port map( A => n10411, B => n3451, ZN => n9345);
   U16135 : XNOR2_X1 port map( A => n9306, B => n10227, ZN => n9984);
   U16136 : XNOR2_X1 port map( A => n9345, B => n9984, ZN => n9346);
   U16137 : NAND3_X1 port map( A1 => n10911, A2 => n10916, A3 => n9348, ZN => 
                           n11523);
   U16138 : NAND2_X1 port map( A1 => n13087, A2 => n11982, ZN => n9349);
   U16139 : OAI21_X1 port map( B1 => n11810, B2 => n13087, A => n9349, ZN => 
                           n9477);
   U16140 : XNOR2_X1 port map( A => n1917, B => n1247, ZN => n9350);
   U16141 : XNOR2_X1 port map( A => n9986, B => n9948, ZN => n9351);
   U16142 : XNOR2_X1 port map( A => n9647, B => n9517, ZN => n10188);
   U16143 : XNOR2_X1 port map( A => n10019, B => n9352, ZN => n10383);
   U16144 : INV_X1 port map( A => n10383, ZN => n9620);
   U16145 : XNOR2_X1 port map( A => n10250, B => n28488, ZN => n9353);
   U16146 : XNOR2_X1 port map( A => n9620, B => n9353, ZN => n9356);
   U16147 : INV_X1 port map( A => n2973, ZN => n24959);
   U16148 : XNOR2_X1 port map( A => n9619, B => n24959, ZN => n9354);
   U16149 : XNOR2_X1 port map( A => n10179, B => n9354, ZN => n9355);
   U16150 : XNOR2_X1 port map( A => n9356, B => n9355, ZN => n9863);
   U16151 : INV_X1 port map( A => n9863, ZN => n9362);
   U16152 : XNOR2_X1 port map( A => n10372, B => n9717, ZN => n10027);
   U16153 : XNOR2_X1 port map( A => n9357, B => n10027, ZN => n9361);
   U16154 : XNOR2_X1 port map( A => n9996, B => n28634, ZN => n9359);
   U16155 : XNOR2_X1 port map( A => n10202, B => n3015, ZN => n9358);
   U16156 : XNOR2_X1 port map( A => n9358, B => n9359, ZN => n9360);
   U16157 : NAND2_X1 port map( A1 => n9362, A2 => n10962, ZN => n10602);
   U16158 : OAI21_X1 port map( B1 => n10958, B2 => n28173, A => n10602, ZN => 
                           n9391);
   U16160 : XNOR2_X1 port map( A => n9368, B => n10352, ZN => n9369);
   U16161 : XNOR2_X1 port map( A => n9631, B => n9369, ZN => n9382);
   U16162 : INV_X1 port map( A => n9370, ZN => n9372);
   U16163 : NAND2_X1 port map( A1 => n9372, A2 => n11, ZN => n9377);
   U16164 : INV_X1 port map( A => n9373, ZN => n9375);
   U16165 : NAND2_X1 port map( A1 => n9375, A2 => n9374, ZN => n9376);
   U16166 : NAND3_X1 port map( A1 => n9378, A2 => n9377, A3 => n9376, ZN => 
                           n9379);
   U16167 : XNOR2_X1 port map( A => n9504, B => n1911, ZN => n9380);
   U16168 : XNOR2_X1 port map( A => n9721, B => n9380, ZN => n9381);
   U16169 : XNOR2_X1 port map( A => n9382, B => n9381, ZN => n10956);
   U16170 : INV_X1 port map( A => n9695, ZN => n9383);
   U16171 : XNOR2_X1 port map( A => n10138, B => n27462, ZN => n9384);
   U16172 : XNOR2_X1 port map( A => n10169, B => n9384, ZN => n9385);
   U16173 : XNOR2_X1 port map( A => n9386, B => n9385, ZN => n10963);
   U16174 : XNOR2_X1 port map( A => n10191, B => n10263, ZN => n10005);
   U16175 : XNOR2_X1 port map( A => n10005, B => n10424, ZN => n9389);
   U16176 : XNOR2_X1 port map( A => n9639, B => n9929, ZN => n9388);
   U16177 : XNOR2_X1 port map( A => n10193, B => n2446, ZN => n9387);
   U16178 : OAI21_X1 port map( B1 => n9858, B2 => n10780, A => n10687, ZN => 
                           n9390);
   U16179 : AOI22_X1 port map( A1 => n9391, A2 => n9390, B1 => n28173, B2 => 
                           n9858, ZN => n12226);
   U16180 : XNOR2_X1 port map( A => n10298, B => n10134, ZN => n9969);
   U16181 : XNOR2_X1 port map( A => n9732, B => n9613, ZN => n9453);
   U16182 : XNOR2_X1 port map( A => n9969, B => n9453, ZN => n9395);
   U16183 : XNOR2_X1 port map( A => n10344, B => n9392, ZN => n10418);
   U16184 : XNOR2_X1 port map( A => n1920, B => n3378, ZN => n9393);
   U16185 : XNOR2_X1 port map( A => n10418, B => n9393, ZN => n9394);
   U16186 : OAI22_X1 port map( A1 => n436, A2 => n9398, B1 => n9397, B2 => n609
                           , ZN => n9400);
   U16187 : NOR2_X1 port map( A1 => n9400, A2 => n9399, ZN => n9401);
   U16188 : XNOR2_X1 port map( A => n9961, B => n10425, ZN => n9405);
   U16189 : XNOR2_X1 port map( A => n9964, B => n1887, ZN => n9402);
   U16190 : XNOR2_X1 port map( A => n9403, B => n9402, ZN => n9404);
   U16191 : XNOR2_X1 port map( A => n9985, B => n10332, ZN => n9408);
   U16192 : XNOR2_X1 port map( A => n9647, B => n3483, ZN => n9406);
   U16193 : XNOR2_X1 port map( A => n9687, B => n9406, ZN => n9407);
   U16194 : INV_X1 port map( A => n9409, ZN => n9413);
   U16195 : OAI22_X1 port map( A1 => n9413, A2 => n9412, B1 => n28211, B2 => 
                           n9410, ZN => n9415);
   U16196 : XNOR2_X1 port map( A => n10202, B => n3256, ZN => n9416);
   U16197 : OAI21_X1 port map( B1 => n11004, B2 => n6779, A => n9417, ZN => 
                           n9694);
   U16198 : OAI21_X1 port map( B1 => n10997, B2 => n6779, A => n9694, ZN => 
                           n11528);
   U16199 : XNOR2_X1 port map( A => n10208, B => n10356, ZN => n9418);
   U16200 : XNOR2_X1 port map( A => n10272, B => n10434, ZN => n9958);
   U16201 : XNOR2_X1 port map( A => n9418, B => n9958, ZN => n9429);
   U16202 : INV_X1 port map( A => n9419, ZN => n9424);
   U16203 : INV_X1 port map( A => n9420, ZN => n9423);
   U16204 : OAI211_X1 port map( C1 => n9425, C2 => n9424, A => n9423, B => 
                           n9422, ZN => n9426);
   U16205 : XNOR2_X1 port map( A => n10436, B => n3686, ZN => n9427);
   U16206 : XNOR2_X1 port map( A => n9722, B => n9427, ZN => n9428);
   U16207 : XNOR2_X1 port map( A => n9428, B => n9429, ZN => n11000);
   U16208 : XNOR2_X1 port map( A => n9772, B => n9430, ZN => n10337);
   U16209 : INV_X1 port map( A => n10337, ZN => n9712);
   U16210 : XNOR2_X1 port map( A => n10151, B => n10386, ZN => n9981);
   U16211 : XNOR2_X1 port map( A => n9712, B => n9981, ZN => n9432);
   U16212 : XNOR2_X1 port map( A => n9431, B => n10335, ZN => n10382);
   U16213 : OAI211_X1 port map( C1 => n5573, C2 => n592, A => n10936, B => 
                           n10999, ZN => n11524);
   U16214 : NAND2_X1 port map( A1 => n11528, A2 => n11524, ZN => n11980);
   U16215 : NAND2_X1 port map( A1 => n9433, A2 => n12227, ZN => n13082);
   U16218 : INV_X1 port map( A => n10045, ZN => n9440);
   U16219 : XNOR2_X1 port map( A => n10283, B => n9440, ZN => n9442);
   U16220 : XNOR2_X1 port map( A => n9899, B => n3219, ZN => n9441);
   U16221 : XNOR2_X1 port map( A => n9442, B => n9441, ZN => n9445);
   U16222 : XNOR2_X1 port map( A => n10159, B => n9746, ZN => n9443);
   U16223 : XNOR2_X1 port map( A => n9443, B => n10188, ZN => n9444);
   U16224 : INV_X1 port map( A => n1879, ZN => n10458);
   U16225 : XNOR2_X1 port map( A => n9446, B => n10202, ZN => n9893);
   U16226 : INV_X1 port map( A => n9893, ZN => n9448);
   U16227 : XNOR2_X1 port map( A => n9447, B => n10028, ZN => n10199);
   U16228 : XNOR2_X1 port map( A => n10199, B => n9448, ZN => n9452);
   U16229 : XNOR2_X1 port map( A => n9754, B => n2411, ZN => n9449);
   U16230 : XNOR2_X1 port map( A => n9450, B => n9449, ZN => n9451);
   U16231 : XNOR2_X1 port map( A => n9452, B => n9451, ZN => n10924);
   U16232 : INV_X1 port map( A => n10924, ZN => n9475);
   U16233 : NAND2_X1 port map( A1 => n10458, A2 => n9475, ZN => n10108);
   U16234 : INV_X1 port map( A => n9453, ZN => n9455);
   U16235 : XNOR2_X1 port map( A => n10133, B => n1892, ZN => n9454);
   U16236 : XNOR2_X1 port map( A => n9455, B => n9454, ZN => n9459);
   U16237 : XNOR2_X1 port map( A => n10033, B => n10297, ZN => n9457);
   U16238 : XNOR2_X1 port map( A => n1902, B => n25992, ZN => n9456);
   U16239 : XNOR2_X1 port map( A => n9457, B => n9456, ZN => n9458);
   U16240 : XNOR2_X1 port map( A => n9639, B => n9877, ZN => n9461);
   U16241 : XNOR2_X1 port map( A => n10009, B => n891, ZN => n9460);
   U16242 : XNOR2_X1 port map( A => n9461, B => n9460, ZN => n9464);
   U16243 : XNOR2_X1 port map( A => n9462, B => n9658, ZN => n9463);
   U16246 : XNOR2_X1 port map( A => n9852, B => n10208, ZN => n9887);
   U16247 : XNOR2_X1 port map( A => n10357, B => n9504, ZN => n9466);
   U16248 : XNOR2_X1 port map( A => n10073, B => n3633, ZN => n9465);
   U16249 : XNOR2_X1 port map( A => n9772, B => n10384, ZN => n9470);
   U16252 : INV_X1 port map( A => n9906, ZN => n9469);
   U16253 : XNOR2_X1 port map( A => n9469, B => n9470, ZN => n9474);
   U16254 : XNOR2_X1 port map( A => n9677, B => n10059, ZN => n9472);
   U16255 : XNOR2_X1 port map( A => n9550, B => n5490, ZN => n9471);
   U16256 : XNOR2_X1 port map( A => n9472, B => n9471, ZN => n9473);
   U16257 : AOI21_X1 port map( B1 => n10459, B2 => n10458, A => n590, ZN => 
                           n9476);
   U16258 : XNOR2_X1 port map( A => n9478, B => n13051, ZN => n9869);
   U16259 : INV_X1 port map( A => n9771, ZN => n9479);
   U16260 : XNOR2_X1 port map( A => n9479, B => n10060, ZN => n9480);
   U16261 : XNOR2_X1 port map( A => n9981, B => n9480, ZN => n9483);
   U16262 : XNOR2_X1 port map( A => n10021, B => n3751, ZN => n9481);
   U16263 : XNOR2_X1 port map( A => n10338, B => n9481, ZN => n9482);
   U16264 : XNOR2_X1 port map( A => n9851, B => n10352, ZN => n10018);
   U16265 : XNOR2_X1 port map( A => n10277, B => n10018, ZN => n9486);
   U16266 : XNOR2_X1 port map( A => n9958, B => n9484, ZN => n9485);
   U16267 : INV_X1 port map( A => n11318, ZN => n11254);
   U16268 : XNOR2_X1 port map( A => n9969, B => n10256, ZN => n9490);
   U16269 : XNOR2_X1 port map( A => n28643, B => n10038, ZN => n9488);
   U16270 : XNOR2_X1 port map( A => n9698, B => n2385, ZN => n9487);
   U16271 : XNOR2_X1 port map( A => n9488, B => n9487, ZN => n9489);
   U16272 : XNOR2_X1 port map( A => n10043, B => n27225, ZN => n9492);
   U16273 : XNOR2_X1 port map( A => n10201, B => n10392, ZN => n9494);
   U16274 : INV_X1 port map( A => n3462, ZN => n27656);
   U16275 : XNOR2_X1 port map( A => n301, B => n27656, ZN => n9493);
   U16276 : XNOR2_X1 port map( A => n9494, B => n9493, ZN => n9497);
   U16277 : XNOR2_X1 port map( A => n10029, B => n10219, ZN => n9838);
   U16278 : XNOR2_X1 port map( A => n9992, B => n9755, ZN => n9495);
   U16279 : XNOR2_X1 port map( A => n10191, B => n9963, ZN => n10367);
   U16280 : INV_X1 port map( A => n9743, ZN => n9498);
   U16281 : XNOR2_X1 port map( A => n9498, B => n10367, ZN => n9501);
   U16282 : XNOR2_X1 port map( A => n10088, B => n2402, ZN => n9499);
   U16283 : XNOR2_X1 port map( A => n9961, B => n9499, ZN => n9500);
   U16284 : XNOR2_X1 port map( A => n9501, B => n9500, ZN => n10482);
   U16285 : MUX2_X2 port map( A => n9503, B => n9502, S => n4296, Z => n12211);
   U16286 : XNOR2_X1 port map( A => n9505, B => n9504, ZN => n9506);
   U16287 : XNOR2_X1 port map( A => n9506, B => n10271, ZN => n9508);
   U16288 : XNOR2_X1 port map( A => n10128, B => n3482, ZN => n9507);
   U16289 : XNOR2_X1 port map( A => n9508, B => n9507, ZN => n9510);
   U16290 : XNOR2_X1 port map( A => n10435, B => n10073, ZN => n10212);
   U16291 : XNOR2_X1 port map( A => n10212, B => n9509, ZN => n9812);
   U16292 : XNOR2_X1 port map( A => n10193, B => n1119, ZN => n9511);
   U16293 : XNOR2_X1 port map( A => n9511, B => n9878, ZN => n9513);
   U16294 : XNOR2_X1 port map( A => n9513, B => n1985, ZN => n9516);
   U16295 : INV_X1 port map( A => n9929, ZN => n9514);
   U16296 : XNOR2_X1 port map( A => n9515, B => n9516, ZN => n10522);
   U16297 : INV_X1 port map( A => n10522, ZN => n11274);
   U16298 : NAND2_X1 port map( A1 => n11038, A2 => n11274, ZN => n9548);
   U16299 : XNOR2_X1 port map( A => n9900, B => n1878, ZN => n9518);
   U16300 : XNOR2_X1 port map( A => n10232, B => n3223, ZN => n9519);
   U16301 : XNOR2_X1 port map( A => n9520, B => n9519, ZN => n9521);
   U16302 : XNOR2_X1 port map( A => n9522, B => n9521, ZN => n11269);
   U16303 : INV_X1 port map( A => n11269, ZN => n11034);
   U16304 : XNOR2_X1 port map( A => n9523, B => n10199, ZN => n9527);
   U16305 : XNOR2_X1 port map( A => n28634, B => n10144, ZN => n9525);
   U16306 : XNOR2_X1 port map( A => n9716, B => n5633, ZN => n9524);
   U16307 : XNOR2_X1 port map( A => n9525, B => n9524, ZN => n9526);
   U16308 : XNOR2_X1 port map( A => n9527, B => n9526, ZN => n11272);
   U16309 : NAND2_X1 port map( A1 => n11034, A2 => n28612, ZN => n9547);
   U16310 : XNOR2_X1 port map( A => n10137, B => n9528, ZN => n9873);
   U16311 : INV_X1 port map( A => n9873, ZN => n9541);
   U16312 : OAI21_X1 port map( B1 => n29662, B2 => n9533, A => n9532, ZN => 
                           n9535);
   U16313 : NAND2_X1 port map( A1 => n9536, A2 => n9535, ZN => n9538);
   U16314 : NAND2_X1 port map( A1 => n9538, A2 => n9537, ZN => n9539);
   U16315 : XNOR2_X1 port map( A => n9540, B => n9539, ZN => n10173);
   U16316 : XNOR2_X1 port map( A => n9541, B => n10173, ZN => n9546);
   U16317 : XNOR2_X1 port map( A => n9542, B => n9696, ZN => n9544);
   U16318 : XNOR2_X1 port map( A => n10138, B => n2523, ZN => n9543);
   U16319 : XNOR2_X1 port map( A => n9544, B => n9543, ZN => n9545);
   U16320 : MUX2_X1 port map( A => n9548, B => n9547, S => n279, Z => n9557);
   U16321 : XNOR2_X1 port map( A => n9907, B => n9549, ZN => n9554);
   U16322 : XNOR2_X1 port map( A => n9710, B => n10385, ZN => n9552);
   U16323 : XNOR2_X1 port map( A => n9550, B => n3660, ZN => n9551);
   U16324 : XNOR2_X1 port map( A => n9552, B => n9551, ZN => n9553);
   U16325 : NAND2_X1 port map( A1 => n9555, A2 => n11269, ZN => n9556);
   U16326 : XNOR2_X1 port map( A => n10386, B => n2984, ZN => n9559);
   U16327 : INV_X1 port map( A => n9786, ZN => n9558);
   U16328 : XNOR2_X1 port map( A => n9559, B => n9558, ZN => n9560);
   U16329 : XNOR2_X1 port map( A => n9560, B => n9842, ZN => n9571);
   U16330 : XNOR2_X1 port map( A => n10321, B => n10178, ZN => n9570);
   U16331 : NAND3_X1 port map( A1 => n9566, A2 => n9562, A3 => n9561, ZN => 
                           n9563);
   U16332 : OAI211_X1 port map( C1 => n9566, C2 => n9565, A => n9564, B => 
                           n9563, ZN => n9568);
   U16333 : NOR2_X1 port map( A1 => n9568, A2 => n9567, ZN => n9569);
   U16334 : XNOR2_X1 port map( A => n9570, B => n9569, ZN => n9926);
   U16335 : INV_X1 port map( A => n9817, ZN => n9574);
   U16336 : XNOR2_X1 port map( A => n9795, B => n3635, ZN => n9572);
   U16337 : XNOR2_X1 port map( A => n9572, B => n10302, ZN => n9573);
   U16338 : XNOR2_X1 port map( A => n9574, B => n9573, ZN => n9578);
   U16339 : XNOR2_X1 port map( A => n9575, B => n10304, ZN => n9576);
   U16342 : NAND2_X1 port map( A1 => n9579, A2 => n24906, ZN => n9585);
   U16343 : NAND4_X1 port map( A1 => n9581, A2 => n9582, A3 => n1196, A4 => 
                           n9580, ZN => n9584);
   U16344 : NAND3_X1 port map( A1 => n9585, A2 => n9584, A3 => n9583, ZN => 
                           n9586);
   U16345 : XNOR2_X1 port map( A => n9586, B => n10392, ZN => n9587);
   U16346 : XNOR2_X1 port map( A => n9587, B => n9836, ZN => n9589);
   U16347 : XNOR2_X1 port map( A => n10143, B => n9716, ZN => n9588);
   U16348 : XNOR2_X1 port map( A => n9757, B => n9588, ZN => n9938);
   U16349 : XNOR2_X1 port map( A => n9589, B => n9938, ZN => n11252);
   U16350 : XNOR2_X1 port map( A => n9592, B => n10434, ZN => n10314);
   U16351 : XNOR2_X1 port map( A => n10071, B => n3643, ZN => n9593);
   U16352 : XNOR2_X1 port map( A => n9593, B => n10314, ZN => n9594);
   U16353 : XNOR2_X1 port map( A => n9595, B => n9594, ZN => n10524);
   U16354 : INV_X1 port map( A => n10524, ZN => n10833);
   U16355 : XNOR2_X1 port map( A => n9596, B => n10294, ZN => n9919);
   U16356 : INV_X1 port map( A => n9919, ZN => n9600);
   U16357 : XNOR2_X1 port map( A => n9799, B => n3414, ZN => n9597);
   U16358 : XNOR2_X1 port map( A => n10298, B => n9597, ZN => n9598);
   U16359 : XNOR2_X1 port map( A => n9598, B => n9831, ZN => n9599);
   U16361 : XNOR2_X1 port map( A => n10160, B => n3317, ZN => n9602);
   U16362 : INV_X1 port map( A => n9601, ZN => n10409);
   U16363 : XNOR2_X1 port map( A => n9602, B => n10409, ZN => n9604);
   U16364 : XNOR2_X1 port map( A => n9604, B => n9603, ZN => n9607);
   U16365 : INV_X1 port map( A => n10282, ZN => n9605);
   U16366 : XNOR2_X1 port map( A => n9606, B => n9605, ZN => n9947);
   U16367 : XNOR2_X1 port map( A => n9607, B => n9947, ZN => n10834);
   U16369 : MUX2_X1 port map( A => n11355, B => n10476, S => n11349, Z => n9611
                           );
   U16370 : INV_X1 port map( A => n9608, ZN => n11351);
   U16371 : NAND2_X1 port map( A1 => n11351, A2 => n11347, ZN => n9609);
   U16372 : INV_X1 port map( A => n10847, ZN => n11352);
   U16373 : OAI22_X1 port map( A1 => n9609, A2 => n11349, B1 => n11352, B2 => 
                           n11351, ZN => n9610);
   U16374 : AOI21_X2 port map( B1 => n9611, B2 => n3161, A => n9610, ZN => 
                           n12110);
   U16376 : XNOR2_X1 port map( A => n9612, B => n9613, ZN => n10170);
   U16377 : INV_X1 port map( A => n10170, ZN => n9616);
   U16378 : XNOR2_X1 port map( A => n9614, B => n1892, ZN => n9615);
   U16379 : XNOR2_X1 port map( A => n9616, B => n9615, ZN => n9618);
   U16381 : XNOR2_X1 port map( A => n9677, B => n1853, ZN => n9622);
   U16382 : INV_X1 port map( A => Key(122), ZN => n15576);
   U16383 : XNOR2_X1 port map( A => n9622, B => n9621, ZN => n9623);
   U16384 : NAND2_X1 port map( A1 => n28204, A2 => n11045, ZN => n9644);
   U16385 : XNOR2_X1 port map( A => n9684, B => n10202, ZN => n9625);
   U16386 : XNOR2_X1 port map( A => n10144, B => n26531, ZN => n9624);
   U16387 : XNOR2_X1 port map( A => n9625, B => n9624, ZN => n9628);
   U16388 : XNOR2_X1 port map( A => n9626, B => n9996, ZN => n10393);
   U16389 : INV_X1 port map( A => n10393, ZN => n9627);
   U16390 : XNOR2_X1 port map( A => n10072, B => n9629, ZN => n9630);
   U16391 : XNOR2_X1 port map( A => n9631, B => n9630, ZN => n9635);
   U16392 : XNOR2_X1 port map( A => n10128, B => n10436, ZN => n9633);
   U16393 : INV_X1 port map( A => n3276, ZN => n28013);
   U16394 : XNOR2_X1 port map( A => n10350, B => n28013, ZN => n9632);
   U16395 : XNOR2_X1 port map( A => n9633, B => n9632, ZN => n9634);
   U16396 : XNOR2_X1 port map( A => n10362, B => n9878, ZN => n9638);
   U16397 : INV_X1 port map( A => n2996, ZN => n9636);
   U16398 : XNOR2_X1 port map( A => n9656, B => n9636, ZN => n9637);
   U16399 : XNOR2_X1 port map( A => n9638, B => n9637, ZN => n9643);
   U16400 : INV_X1 port map( A => n9639, ZN => n9640);
   U16401 : XNOR2_X1 port map( A => n9794, B => n9640, ZN => n9641);
   U16402 : XNOR2_X1 port map( A => n10424, B => n9641, ZN => n9642);
   U16403 : XNOR2_X1 port map( A => n9642, B => n9643, ZN => n10528);
   U16404 : OAI22_X1 port map( A1 => n9644, A2 => n11044, B1 => n11264, B2 => 
                           n28204, ZN => n9654);
   U16405 : XNOR2_X1 port map( A => n9645, B => n9986, ZN => n10048);
   U16406 : XNOR2_X1 port map( A => n9646, B => n10048, ZN => n9652);
   U16407 : XNOR2_X1 port map( A => n9647, B => n10159, ZN => n9650);
   U16408 : XNOR2_X1 port map( A => n9648, B => n1919, ZN => n9649);
   U16409 : XNOR2_X1 port map( A => n9650, B => n9649, ZN => n9651);
   U16410 : NAND2_X1 port map( A1 => n28204, A2 => n11267, ZN => n11043);
   U16411 : XNOR2_X1 port map( A => n9656, B => n1046, ZN => n9657);
   U16412 : XNOR2_X1 port map( A => n10303, B => n9657, ZN => n9659);
   U16413 : INV_X1 port map( A => n9660, ZN => n9664);
   U16416 : XNOR2_X1 port map( A => n9664, B => n9663, ZN => n9667);
   U16417 : XNOR2_X1 port map( A => n10295, B => n9971, ZN => n9665);
   U16418 : XNOR2_X1 port map( A => n9665, B => n9732, ZN => n9701);
   U16419 : XNOR2_X1 port map( A => n10072, B => n10352, ZN => n9670);
   U16420 : INV_X1 port map( A => n9668, ZN => n9669);
   U16421 : XNOR2_X1 port map( A => n9669, B => n9670, ZN => n9673);
   U16422 : XNOR2_X1 port map( A => n9941, B => n3537, ZN => n9671);
   U16423 : INV_X1 port map( A => n9908, ZN => n9922);
   U16424 : XNOR2_X1 port map( A => n9922, B => n9674, ZN => n9676);
   U16425 : XNOR2_X1 port map( A => n9676, B => n9675, ZN => n9682);
   U16426 : XNOR2_X1 port map( A => n9677, B => n9678, ZN => n9680);
   U16427 : XNOR2_X1 port map( A => n10022, B => n2577, ZN => n9679);
   U16428 : XNOR2_X1 port map( A => n9680, B => n9679, ZN => n9681);
   U16429 : XNOR2_X1 port map( A => n9681, B => n9682, ZN => n10855);
   U16430 : XNOR2_X1 port map( A => n9997, B => n2522, ZN => n9685);
   U16431 : XNOR2_X1 port map( A => n10046, B => n9687, ZN => n9691);
   U16432 : XNOR2_X1 port map( A => n10159, B => n9949, ZN => n9689);
   U16433 : XNOR2_X1 port map( A => n9725, B => n2946, ZN => n9688);
   U16434 : XNOR2_X1 port map( A => n9689, B => n9688, ZN => n9690);
   U16438 : XNOR2_X1 port map( A => n9695, B => n1175, ZN => n9697);
   U16439 : XNOR2_X1 port map( A => n9697, B => n9696, ZN => n9699);
   U16440 : XNOR2_X1 port map( A => n10342, B => n9699, ZN => n9700);
   U16441 : XNOR2_X1 port map( A => n9700, B => n9701, ZN => n10622);
   U16442 : INV_X1 port map( A => n10622, ZN => n9709);
   U16443 : INV_X1 port map( A => n9964, ZN => n9702);
   U16446 : XNOR2_X1 port map( A => n9705, B => n9706, ZN => n9707);
   U16447 : XNOR2_X2 port map( A => n9708, B => n9707, ZN => n10797);
   U16448 : NAND2_X1 port map( A1 => n9709, A2 => n10797, ZN => n10569);
   U16449 : XNOR2_X1 port map( A => n9710, B => n9711, ZN => n9713);
   U16450 : XNOR2_X1 port map( A => n9712, B => n9713, ZN => n9714);
   U16451 : XNOR2_X1 port map( A => n10391, B => n9991, ZN => n9715);
   U16452 : XNOR2_X1 port map( A => n10376, B => n9715, ZN => n9720);
   U16453 : XNOR2_X1 port map( A => n9313, B => n2381, ZN => n9718);
   U16454 : XNOR2_X1 port map( A => n9716, B => n9717, ZN => n10223);
   U16455 : XNOR2_X1 port map( A => n9718, B => n10223, ZN => n9719);
   U16456 : INV_X1 port map( A => n11227, ZN => n10795);
   U16457 : XNOR2_X1 port map( A => n10330, B => n9746, ZN => n9723);
   U16458 : XNOR2_X1 port map( A => n9723, B => n9724, ZN => n9729);
   U16459 : XNOR2_X1 port map( A => n1917, B => n9725, ZN => n9727);
   U16460 : INV_X1 port map( A => n21865, ZN => n27737);
   U16461 : XNOR2_X1 port map( A => n10232, B => n27737, ZN => n9726);
   U16462 : XNOR2_X1 port map( A => n9727, B => n9726, ZN => n9728);
   U16463 : XNOR2_X1 port map( A => n9729, B => n9728, ZN => n11225);
   U16464 : NAND2_X1 port map( A1 => n28568, A2 => n11225, ZN => n11231);
   U16465 : NAND2_X1 port map( A1 => n10797, A2 => n11227, ZN => n11898);
   U16466 : AOI21_X1 port map( B1 => n11231, B2 => n11898, A => n11099, ZN => 
                           n9730);
   U16467 : INV_X1 port map( A => n12198, ZN => n11818);
   U16468 : XNOR2_X1 port map( A => n10134, B => n9732, ZN => n9734);
   U16469 : XNOR2_X1 port map( A => n10038, B => n2441, ZN => n9733);
   U16470 : XNOR2_X1 port map( A => n9733, B => n9734, ZN => n9739);
   U16471 : XNOR2_X1 port map( A => n9915, B => n9735, ZN => n9737);
   U16472 : XNOR2_X1 port map( A => n9737, B => n9736, ZN => n9738);
   U16473 : INV_X1 port map( A => n11237, ZN => n10628);
   U16474 : XNOR2_X1 port map( A => n9741, B => n9740, ZN => n9745);
   U16475 : XNOR2_X1 port map( A => n9742, B => n9743, ZN => n9744);
   U16476 : XNOR2_X1 port map( A => n9949, B => n9746, ZN => n9747);
   U16477 : XNOR2_X1 port map( A => n9748, B => n9747, ZN => n9753);
   U16478 : INV_X1 port map( A => n10231, ZN => n10158);
   U16479 : XNOR2_X1 port map( A => n9749, B => n10158, ZN => n9751);
   U16481 : XNOR2_X1 port map( A => n9751, B => n9750, ZN => n9752);
   U16482 : XNOR2_X1 port map( A => n9753, B => n9752, ZN => n11013);
   U16483 : XNOR2_X1 port map( A => n9754, B => n9755, ZN => n9756);
   U16484 : XNOR2_X1 port map( A => n10287, B => n9756, ZN => n9761);
   U16485 : XNOR2_X1 port map( A => n9757, B => n301, ZN => n9759);
   U16486 : XNOR2_X1 port map( A => n10144, B => n2541, ZN => n9758);
   U16487 : XNOR2_X1 port map( A => n9759, B => n9758, ZN => n9760);
   U16488 : XNOR2_X1 port map( A => n9761, B => n9760, ZN => n11236);
   U16489 : NAND2_X1 port map( A1 => n11013, A2 => n11236, ZN => n11233);
   U16490 : INV_X1 port map( A => n11233, ZN => n9762);
   U16491 : NAND2_X1 port map( A1 => n9762, A2 => n5710, ZN => n9778);
   U16492 : XNOR2_X1 port map( A => n9763, B => n10272, ZN => n9765);
   U16493 : INV_X1 port map( A => n10315, ZN => n9764);
   U16494 : XNOR2_X1 port map( A => n9765, B => n9764, ZN => n9769);
   U16495 : XNOR2_X1 port map( A => n10357, B => n2476, ZN => n9766);
   U16496 : XNOR2_X1 port map( A => n9767, B => n9766, ZN => n9768);
   U16497 : XNOR2_X1 port map( A => n10319, B => n9770, ZN => n9776);
   U16498 : XNOR2_X1 port map( A => n9772, B => n9771, ZN => n9774);
   U16499 : INV_X1 port map( A => n22489, ZN => n28007);
   U16500 : XNOR2_X1 port map( A => n10151, B => n28007, ZN => n9773);
   U16501 : XNOR2_X1 port map( A => n9774, B => n9773, ZN => n9775);
   U16502 : INV_X1 port map( A => n11235, ZN => n11014);
   U16503 : INV_X1 port map( A => n11236, ZN => n10776);
   U16504 : OAI211_X1 port map( C1 => n3441, C2 => n1381, A => n11014, B => 
                           n10776, ZN => n9777);
   U16505 : XNOR2_X1 port map( A => n10080, B => n9780, ZN => n9784);
   U16506 : XNOR2_X1 port map( A => n10395, B => n28327, ZN => n9781);
   U16507 : XNOR2_X1 port map( A => n9782, B => n9781, ZN => n9783);
   U16508 : XNOR2_X1 port map( A => n9784, B => n9783, ZN => n10990);
   U16509 : XNOR2_X1 port map( A => n28488, B => n10385, ZN => n9787);
   U16510 : INV_X1 port map( A => n10059, ZN => n9788);
   U16511 : XNOR2_X1 port map( A => n9788, B => n10384, ZN => n9790);
   U16512 : XNOR2_X1 port map( A => n9979, B => n3644, ZN => n9789);
   U16513 : XNOR2_X1 port map( A => n9790, B => n9789, ZN => n9791);
   U16514 : INV_X1 port map( A => n10990, ZN => n10785);
   U16515 : XNOR2_X1 port map( A => n9794, B => n9795, ZN => n10120);
   U16516 : INV_X1 port map( A => n10120, ZN => n10085);
   U16517 : XNOR2_X1 port map( A => n10264, B => n28294, ZN => n9796);
   U16518 : XNOR2_X1 port map( A => n9796, B => n10364, ZN => n9797);
   U16519 : XNOR2_X1 port map( A => n10085, B => n9797, ZN => n9798);
   U16520 : XNOR2_X1 port map( A => n9799, B => n9661, ZN => n10135);
   U16521 : INV_X1 port map( A => n10135, ZN => n9801);
   U16522 : XNOR2_X1 port map( A => n10257, B => n10297, ZN => n9800);
   U16523 : XNOR2_X1 port map( A => n9801, B => n9800, ZN => n9804);
   U16524 : XNOR2_X1 port map( A => n10138, B => n27105, ZN => n9802);
   U16525 : XNOR2_X1 port map( A => n10173, B => n9802, ZN => n9803);
   U16526 : INV_X1 port map( A => n10992, ZN => n10791);
   U16527 : NAND3_X1 port map( A1 => n10693, A2 => n10691, A3 => n10791, ZN => 
                           n9816);
   U16528 : XNOR2_X1 port map( A => n10283, B => n10159, ZN => n9805);
   U16529 : XNOR2_X1 port map( A => n10227, B => n9948, ZN => n9807);
   U16530 : XNOR2_X1 port map( A => n10160, B => n3742, ZN => n9806);
   U16531 : XNOR2_X1 port map( A => n9807, B => n9806, ZN => n9808);
   U16532 : NAND3_X1 port map( A1 => n10995, A2 => n10993, A3 => n4538, ZN => 
                           n9815);
   U16533 : XNOR2_X1 port map( A => n10275, B => n3565, ZN => n9810);
   U16537 : MUX2_X1 port map( A => n11818, B => n12189, S => n12190, Z => n9868
                           );
   U16538 : XNOR2_X1 port map( A => n9818, B => n9817, ZN => n9822);
   U16539 : XNOR2_X1 port map( A => n10088, B => n26032, ZN => n9819);
   U16540 : XNOR2_X1 port map( A => n9820, B => n9819, ZN => n9821);
   U16541 : XNOR2_X1 port map( A => n9822, B => n9821, ZN => n10982);
   U16542 : XNOR2_X1 port map( A => n10229, B => n9825, ZN => n9829);
   U16543 : XNOR2_X1 port map( A => n10328, B => n10043, ZN => n9827);
   U16544 : XNOR2_X1 port map( A => n10183, B => n72, ZN => n9826);
   U16545 : XNOR2_X1 port map( A => n9827, B => n9826, ZN => n9828);
   U16546 : XNOR2_X1 port map( A => n9829, B => n9828, ZN => n10984);
   U16547 : NAND2_X1 port map( A1 => n10982, A2 => n10984, ZN => n10631);
   U16548 : XNOR2_X1 port map( A => n9870, B => n10038, ZN => n9830);
   U16549 : XNOR2_X1 port map( A => n9831, B => n9830, ZN => n9835);
   U16550 : XNOR2_X1 port map( A => n10171, B => n2404, ZN => n9832);
   U16551 : XNOR2_X1 port map( A => n9833, B => n9832, ZN => n9834);
   U16552 : NOR2_X1 port map( A1 => n10989, A2 => n10982, ZN => n10630);
   U16553 : XNOR2_X1 port map( A => n10371, B => n10143, ZN => n10200);
   U16554 : XNOR2_X1 port map( A => n10200, B => n9836, ZN => n9840);
   U16555 : XNOR2_X1 port map( A => n1868, B => n26665, ZN => n9837);
   U16556 : XNOR2_X1 port map( A => n9838, B => n9837, ZN => n9839);
   U16557 : XNOR2_X1 port map( A => n9840, B => n9839, ZN => n10981);
   U16558 : AND2_X1 port map( A1 => n10985, A2 => n10982, ZN => n9841);
   U16559 : NOR2_X1 port map( A1 => n10630, A2 => n9841, ZN => n9848);
   U16560 : XNOR2_X1 port map( A => n9843, B => n9842, ZN => n9847);
   U16561 : XNOR2_X1 port map( A => n10021, B => n3654, ZN => n9844);
   U16562 : XNOR2_X1 port map( A => n9845, B => n9844, ZN => n9846);
   U16563 : XNOR2_X1 port map( A => n9847, B => n9846, ZN => n10980);
   U16564 : XNOR2_X1 port map( A => n9849, B => n9850, ZN => n9856);
   U16565 : XNOR2_X1 port map( A => n9851, B => n10275, ZN => n9854);
   U16566 : XNOR2_X1 port map( A => n9852, B => n3380, ZN => n9853);
   U16567 : XNOR2_X1 port map( A => n9854, B => n9853, ZN => n9855);
   U16568 : INV_X1 port map( A => n10958, ZN => n10686);
   U16569 : NAND2_X1 port map( A1 => n10686, A2 => n10962, ZN => n9857);
   U16570 : NAND2_X1 port map( A1 => n9857, A2 => n10780, ZN => n9862);
   U16571 : INV_X1 port map( A => n10966, ZN => n9860);
   U16572 : NAND2_X1 port map( A1 => n9862, A2 => n9861, ZN => n12188);
   U16573 : MUX2_X1 port map( A => n10780, B => n10687, S => n10957, Z => n9864
                           );
   U16574 : NAND2_X1 port map( A1 => n9864, A2 => n10958, ZN => n12187);
   U16575 : NAND2_X1 port map( A1 => n11816, A2 => n12128, ZN => n12129);
   U16576 : NAND3_X1 port map( A1 => n9865, A2 => n12194, A3 => n12190, ZN => 
                           n9866);
   U16577 : NAND3_X1 port map( A1 => n12129, A2 => n12186, A3 => n9866, ZN => 
                           n9867);
   U16578 : XNOR2_X1 port map( A => n9869, B => n12454, ZN => n10444);
   U16579 : XNOR2_X1 port map( A => n9870, B => n9915, ZN => n9871);
   U16580 : XNOR2_X1 port map( A => n9872, B => n9871, ZN => n9876);
   U16581 : XNOR2_X1 port map( A => n10133, B => n26825, ZN => n9874);
   U16582 : XNOR2_X1 port map( A => n9873, B => n9874, ZN => n9875);
   U16583 : XNOR2_X1 port map( A => n9876, B => n9875, ZN => n9913);
   U16584 : INV_X1 port map( A => n9877, ZN => n9879);
   U16585 : XNOR2_X1 port map( A => n9879, B => n9878, ZN => n9880);
   U16586 : XNOR2_X1 port map( A => n10189, B => n9880, ZN => n9885);
   U16587 : XNOR2_X1 port map( A => n9931, B => n9881, ZN => n9883);
   U16588 : XNOR2_X1 port map( A => n10088, B => n730, ZN => n9882);
   U16589 : XNOR2_X1 port map( A => n9883, B => n9882, ZN => n9884);
   U16590 : NAND2_X1 port map( A1 => n11127, A2 => n11123, ZN => n10507);
   U16591 : XNOR2_X1 port map( A => n10074, B => n10271, ZN => n9886);
   U16592 : XNOR2_X1 port map( A => n9887, B => n9886, ZN => n9891);
   U16593 : INV_X1 port map( A => n3606, ZN => n25044);
   U16594 : XNOR2_X1 port map( A => n10128, B => n25044, ZN => n9889);
   U16595 : XNOR2_X1 port map( A => n9941, B => n10435, ZN => n9888);
   U16596 : XNOR2_X1 port map( A => n9888, B => n9889, ZN => n9890);
   U16597 : XNOR2_X1 port map( A => n9890, B => n9891, ZN => n11119);
   U16598 : INV_X1 port map( A => n11119, ZN => n10504);
   U16599 : XNOR2_X1 port map( A => n9892, B => n9893, ZN => n9898);
   U16600 : XNOR2_X1 port map( A => n10396, B => n9934, ZN => n9896);
   U16601 : XNOR2_X1 port map( A => n1868, B => n2987, ZN => n9895);
   U16602 : XNOR2_X1 port map( A => n9896, B => n9895, ZN => n9897);
   U16603 : XNOR2_X1 port map( A => n9949, B => n24897, ZN => n9902);
   U16605 : INV_X1 port map( A => n10156, ZN => n9901);
   U16606 : XNOR2_X1 port map( A => n9901, B => n9902, ZN => n9905);
   U16607 : XNOR2_X1 port map( A => n10229, B => n9903, ZN => n9904);
   U16608 : XNOR2_X1 port map( A => n9905, B => n9904, ZN => n10114);
   U16609 : XNOR2_X1 port map( A => n9906, B => n9907, ZN => n9912);
   U16610 : XNOR2_X1 port map( A => n9908, B => n10385, ZN => n9910);
   U16611 : XNOR2_X1 port map( A => n10060, B => n3586, ZN => n9909);
   U16612 : XNOR2_X1 port map( A => n9910, B => n9909, ZN => n9911);
   U16613 : INV_X1 port map( A => n11124, ZN => n11126);
   U16614 : INV_X1 port map( A => n11390, ZN => n11922);
   U16615 : XNOR2_X1 port map( A => n9915, B => n3154, ZN => n9917);
   U16616 : XNOR2_X1 port map( A => n9920, B => n9919, ZN => n10096);
   U16617 : XNOR2_X1 port map( A => n9921, B => n3527, ZN => n9923);
   U16618 : XNOR2_X1 port map( A => n9922, B => n9923, ZN => n9925);
   U16619 : XNOR2_X1 port map( A => n9924, B => n9925, ZN => n9927);
   U16620 : INV_X1 port map( A => n135, ZN => n26176);
   U16621 : XNOR2_X1 port map( A => n9964, B => n26176, ZN => n9928);
   U16622 : XNOR2_X1 port map( A => n9931, B => n9930, ZN => n9932);
   U16623 : XNOR2_X1 port map( A => n9935, B => n9934, ZN => n9937);
   U16624 : XNOR2_X1 port map( A => n9936, B => n9937, ZN => n9939);
   U16625 : XNOR2_X1 port map( A => n9939, B => n9938, ZN => n10490);
   U16626 : INV_X1 port map( A => n10490, ZN => n10492);
   U16627 : XNOR2_X1 port map( A => n9941, B => n1927, ZN => n9942);
   U16628 : XNOR2_X1 port map( A => n9943, B => n9942, ZN => n9944);
   U16629 : XNOR2_X1 port map( A => n9947, B => n9946, ZN => n9952);
   U16630 : XNOR2_X1 port map( A => n9948, B => n3491, ZN => n9950);
   U16631 : XNOR2_X1 port map( A => n9950, B => n9949, ZN => n9951);
   U16632 : INV_X1 port map( A => n10275, ZN => n9954);
   U16633 : XNOR2_X1 port map( A => n9955, B => n9954, ZN => n9957);
   U16634 : XNOR2_X1 port map( A => n9956, B => n9957, ZN => n9960);
   U16635 : XNOR2_X1 port map( A => n10359, B => n9958, ZN => n9959);
   U16636 : XNOR2_X1 port map( A => n9962, B => n9961, ZN => n9968);
   U16637 : XNOR2_X1 port map( A => n10007, B => n9963, ZN => n9966);
   U16638 : XNOR2_X1 port map( A => n9964, B => n2960, ZN => n9965);
   U16639 : XNOR2_X1 port map( A => n9966, B => n9965, ZN => n9967);
   U16640 : INV_X1 port map( A => n9969, ZN => n9970);
   U16641 : XNOR2_X1 port map( A => n9970, B => n10342, ZN => n9975);
   U16642 : XNOR2_X1 port map( A => n10037, B => n10257, ZN => n9973);
   U16643 : XNOR2_X1 port map( A => n9971, B => n2505, ZN => n9972);
   U16644 : XNOR2_X1 port map( A => n9973, B => n9972, ZN => n9974);
   U16645 : NAND2_X1 port map( A1 => n5672, A2 => n10713, ZN => n10457);
   U16647 : XNOR2_X1 port map( A => n9976, B => n26713, ZN => n9978);
   U16648 : XNOR2_X1 port map( A => n9978, B => n9977, ZN => n9983);
   U16649 : XNOR2_X1 port map( A => n10019, B => n9979, ZN => n9980);
   U16650 : XNOR2_X1 port map( A => n9981, B => n9980, ZN => n9982);
   U16651 : INV_X1 port map( A => n10498, ZN => n11132);
   U16652 : XNOR2_X1 port map( A => n9985, B => n9984, ZN => n9990);
   U16653 : XNOR2_X1 port map( A => n9986, B => n2477, ZN => n9987);
   U16654 : XNOR2_X1 port map( A => n9988, B => n9987, ZN => n9989);
   U16655 : XNOR2_X1 port map( A => n9989, B => n9990, ZN => n10715);
   U16656 : INV_X1 port map( A => n10715, ZN => n10500);
   U16657 : OAI21_X1 port map( B1 => n10498, B2 => n10500, A => n10502, ZN => 
                           n10003);
   U16658 : XNOR2_X1 port map( A => n10392, B => n9991, ZN => n9995);
   U16659 : INV_X1 port map( A => n9992, ZN => n9993);
   U16660 : XNOR2_X1 port map( A => n9993, B => n10218, ZN => n9994);
   U16661 : XNOR2_X1 port map( A => n9995, B => n9994, ZN => n10001);
   U16662 : XNOR2_X1 port map( A => n9996, B => n301, ZN => n9999);
   U16663 : XNOR2_X1 port map( A => n9997, B => n3374, ZN => n9998);
   U16664 : XNOR2_X1 port map( A => n9998, B => n9999, ZN => n10000);
   U16665 : XNOR2_X1 port map( A => n10000, B => n10001, ZN => n10711);
   U16666 : NAND2_X1 port map( A1 => n10711, A2 => n1834, ZN => n10714);
   U16667 : INV_X1 port map( A => n10714, ZN => n10002);
   U16668 : INV_X1 port map( A => n10005, ZN => n10006);
   U16669 : XNOR2_X1 port map( A => n10006, B => n10425, ZN => n10013);
   U16670 : XNOR2_X1 port map( A => n10007, B => n28616, ZN => n10011);
   U16671 : XNOR2_X1 port map( A => n10009, B => n3516, ZN => n10010);
   U16672 : XNOR2_X1 port map( A => n10010, B => n10011, ZN => n10012);
   U16673 : XNOR2_X2 port map( A => n10013, B => n10012, ZN => n11136);
   U16674 : INV_X1 port map( A => n11136, ZN => n10718);
   U16675 : XNOR2_X1 port map( A => n10436, B => n3372, ZN => n10014);
   U16676 : XNOR2_X1 port map( A => n10015, B => n10014, ZN => n10017);
   U16677 : XNOR2_X1 port map( A => n10311, B => n10073, ZN => n10016);
   U16678 : INV_X1 port map( A => n11142, ZN => n10920);
   U16679 : XNOR2_X1 port map( A => n10019, B => n10250, ZN => n10020);
   U16680 : XNOR2_X1 port map( A => n10382, B => n10020, ZN => n10026);
   U16681 : XNOR2_X1 port map( A => n10059, B => n10021, ZN => n10024);
   U16682 : XNOR2_X1 port map( A => n10022, B => n26680, ZN => n10023);
   U16683 : XNOR2_X1 port map( A => n10024, B => n10023, ZN => n10025);
   U16684 : XNOR2_X1 port map( A => n10026, B => n10025, ZN => n11140);
   U16685 : XNOR2_X1 port map( A => n5412, B => n10028, ZN => n10081);
   U16686 : XNOR2_X1 port map( A => n10029, B => n1179, ZN => n10030);
   U16687 : INV_X1 port map( A => n11135, ZN => n10031);
   U16690 : XNOR2_X1 port map( A => n10034, B => n10033, ZN => n10036);
   U16691 : INV_X1 port map( A => n10418, ZN => n10035);
   U16692 : XNOR2_X1 port map( A => n10036, B => n10035, ZN => n10042);
   U16693 : XNOR2_X1 port map( A => n28643, B => n10037, ZN => n10040);
   U16694 : XNOR2_X1 port map( A => n10038, B => n1062, ZN => n10039);
   U16695 : XNOR2_X1 port map( A => n10040, B => n10039, ZN => n10041);
   U16696 : XNOR2_X1 port map( A => n10043, B => n3695, ZN => n10044);
   U16697 : XNOR2_X1 port map( A => n10045, B => n10044, ZN => n10047);
   U16698 : XNOR2_X1 port map( A => n10047, B => n10046, ZN => n10049);
   U16699 : XNOR2_X1 port map( A => n10048, B => n10064, ZN => n10415);
   U16700 : OAI21_X1 port map( B1 => n10458, B2 => n10726, A => n10051, ZN => 
                           n10054);
   U16701 : OAI21_X1 port map( B1 => n10932, B2 => n10930, A => n10927, ZN => 
                           n10053);
   U16702 : NOR2_X1 port map( A1 => n588, A2 => n10928, ZN => n10052);
   U16704 : INV_X1 port map( A => n11853, ZN => n11924);
   U16705 : XNOR2_X1 port map( A => n10345, B => n1248, ZN => n10056);
   U16706 : XNOR2_X1 port map( A => n10057, B => n10056, ZN => n10058);
   U16707 : XNOR2_X1 port map( A => n10059, B => n1852, ZN => n10176);
   U16708 : XNOR2_X1 port map( A => n10060, B => n27894, ZN => n10061);
   U16709 : XNOR2_X1 port map( A => n10176, B => n10061, ZN => n10062);
   U16710 : XNOR2_X1 port map( A => n10159, B => n10064, ZN => n10066);
   U16711 : XNOR2_X1 port map( A => n10065, B => n10066, ZN => n10070);
   U16712 : XNOR2_X1 port map( A => n10160, B => n3622, ZN => n10067);
   U16713 : XNOR2_X1 port map( A => n10068, B => n10067, ZN => n10069);
   U16714 : XNOR2_X1 port map( A => n10072, B => n10071, ZN => n10126);
   U16715 : XNOR2_X1 port map( A => n10432, B => n10126, ZN => n10078);
   U16716 : XNOR2_X1 port map( A => n10074, B => n10073, ZN => n10076);
   U16717 : XNOR2_X1 port map( A => n10350, B => n22072, ZN => n10075);
   U16718 : XNOR2_X1 port map( A => n10076, B => n10075, ZN => n10077);
   U16719 : INV_X1 port map( A => n10556, ZN => n11153);
   U16720 : XNOR2_X1 port map( A => n10080, B => n10079, ZN => n10084);
   U16721 : XNOR2_X1 port map( A => n10219, B => n3423, ZN => n10082);
   U16722 : XNOR2_X1 port map( A => n10082, B => n10081, ZN => n10083);
   U16723 : XNOR2_X1 port map( A => n10087, B => n10362, ZN => n10190);
   U16724 : INV_X1 port map( A => n10190, ZN => n10090);
   U16725 : XNOR2_X1 port map( A => n10088, B => n2544, ZN => n10089);
   U16726 : MUX2_X1 port map( A => n4788, B => n593, S => n11154, Z => n10092);
   U16727 : INV_X1 port map( A => n10096, ZN => n11115);
   U16728 : INV_X1 port map( A => n10097, ZN => n10549);
   U16729 : MUX2_X1 port map( A => n10099, B => n10098, S => n29150, Z => 
                           n10100);
   U16730 : NOR2_X1 port map( A1 => n10502, A2 => n10715, ZN => n10101);
   U16731 : NOR2_X1 port map( A1 => n3862, A2 => n11136, ZN => n10103);
   U16732 : NAND3_X1 port map( A1 => n3862, A2 => n10919, A3 => n11136, ZN => 
                           n10104);
   U16733 : MUX2_X1 port map( A => n10108, B => n10932, S => n10927, Z => 
                           n10109);
   U16734 : INV_X1 port map( A => n10705, ZN => n10946);
   U16735 : INV_X1 port map( A => n10592, ZN => n10593);
   U16736 : NAND2_X1 port map( A1 => n10593, A2 => n28495, ZN => n10113);
   U16737 : NAND2_X1 port map( A1 => n10110, A2 => n10703, ZN => n10943);
   U16738 : OAI211_X1 port map( C1 => n28176, C2 => n10592, A => n10943, B => 
                           n10942, ZN => n10112);
   U16739 : INV_X1 port map( A => n10942, ZN => n10445);
   U16740 : NAND3_X1 port map( A1 => n1865, A2 => n10593, A3 => n10445, ZN => 
                           n10111);
   U16741 : INV_X1 port map( A => n10114, ZN => n11122);
   U16742 : AOI21_X1 port map( B1 => n11120, B2 => n11126, A => n11122, ZN => 
                           n10116);
   U16743 : NAND2_X1 port map( A1 => n10540, A2 => n11119, ZN => n10115);
   U16744 : XNOR2_X1 port map( A => n13219, B => n13167, ZN => n10442);
   U16745 : XNOR2_X1 port map( A => n10120, B => n10119, ZN => n10125);
   U16746 : INV_X1 port map( A => n2916, ZN => n10121);
   U16747 : XNOR2_X1 port map( A => n10265, B => n10121, ZN => n10122);
   U16748 : XNOR2_X1 port map( A => n10123, B => n10122, ZN => n10124);
   U16749 : XNOR2_X1 port map( A => n10126, B => n10127, ZN => n10132);
   U16750 : XNOR2_X1 port map( A => n10207, B => n10272, ZN => n10130);
   U16751 : XNOR2_X1 port map( A => n10128, B => n3081, ZN => n10129);
   U16752 : XNOR2_X1 port map( A => n10130, B => n10129, ZN => n10131);
   U16753 : XNOR2_X1 port map( A => n10132, B => n10131, ZN => n10882);
   U16754 : AND2_X1 port map( A1 => n10882, A2 => n11210, ZN => n10572);
   U16755 : XNOR2_X1 port map( A => n10134, B => n10133, ZN => n10136);
   U16756 : XNOR2_X1 port map( A => n10135, B => n10136, ZN => n10142);
   U16757 : XNOR2_X1 port map( A => n10137, B => n10171, ZN => n10140);
   U16758 : XNOR2_X1 port map( A => n10138, B => n3134, ZN => n10139);
   U16759 : XNOR2_X1 port map( A => n10140, B => n10139, ZN => n10141);
   U16760 : XNOR2_X1 port map( A => n10146, B => n28634, ZN => n10147);
   U16761 : XNOR2_X1 port map( A => n10149, B => n28488, ZN => n10150);
   U16762 : XNOR2_X1 port map( A => n10178, B => n3666, ZN => n10153);
   U16763 : XNOR2_X1 port map( A => n10152, B => n10153, ZN => n10154);
   U16764 : NAND3_X1 port map( A1 => n11084, A2 => n11209, A3 => n11086, ZN => 
                           n10166);
   U16765 : XNOR2_X1 port map( A => n10156, B => n10157, ZN => n10164);
   U16766 : XNOR2_X1 port map( A => n10159, B => n10158, ZN => n10162);
   U16767 : XNOR2_X1 port map( A => n10160, B => n2961, ZN => n10161);
   U16768 : XNOR2_X1 port map( A => n10162, B => n10161, ZN => n10163);
   U16769 : XNOR2_X1 port map( A => n10163, B => n10164, ZN => n11085);
   U16770 : NAND2_X1 port map( A1 => n11084, A2 => n28624, ZN => n11216);
   U16771 : NOR2_X1 port map( A1 => n11216, A2 => n11209, ZN => n10167);
   U16772 : XNOR2_X1 port map( A => n10169, B => n10170, ZN => n10175);
   U16773 : XNOR2_X1 port map( A => n10171, B => n2389, ZN => n10172);
   U16774 : XNOR2_X1 port map( A => n10173, B => n10172, ZN => n10174);
   U16775 : XNOR2_X1 port map( A => n10176, B => n10177, ZN => n10182);
   U16776 : XNOR2_X1 port map( A => n10178, B => n3109, ZN => n10180);
   U16777 : XNOR2_X1 port map( A => n10179, B => n10180, ZN => n10181);
   U16778 : XNOR2_X1 port map( A => n10183, B => n27298, ZN => n10186);
   U16779 : XNOR2_X1 port map( A => n10185, B => n10186, ZN => n10187);
   U16780 : INV_X1 port map( A => n11243, ZN => n10640);
   U16781 : XNOR2_X1 port map( A => n10190, B => n10189, ZN => n10197);
   U16782 : XNOR2_X1 port map( A => n10191, B => n10192, ZN => n10195);
   U16783 : XNOR2_X1 port map( A => n10193, B => n2510, ZN => n10194);
   U16784 : XNOR2_X1 port map( A => n10195, B => n10194, ZN => n10196);
   U16786 : OAI211_X1 port map( C1 => n1900, C2 => n11242, A => n10640, B => 
                           n10198, ZN => n10217);
   U16787 : XNOR2_X1 port map( A => n10200, B => n10199, ZN => n10206);
   U16788 : XNOR2_X1 port map( A => n10201, B => n10396, ZN => n10204);
   U16789 : XNOR2_X1 port map( A => n10202, B => n4029, ZN => n10203);
   U16790 : XNOR2_X1 port map( A => n10204, B => n10203, ZN => n10205);
   U16791 : NAND3_X1 port map( A1 => n1900, A2 => n11240, A3 => n11243, ZN => 
                           n10216);
   U16792 : XNOR2_X1 port map( A => n10208, B => n10207, ZN => n10210);
   U16793 : XNOR2_X1 port map( A => n10210, B => n10209, ZN => n10214);
   U16794 : INV_X1 port map( A => n21537, ZN => n27669);
   U16795 : XNOR2_X1 port map( A => n10350, B => n27669, ZN => n10211);
   U16796 : XNOR2_X1 port map( A => n10212, B => n10211, ZN => n10213);
   U16797 : NAND3_X1 port map( A1 => n10880, A2 => n11069, A3 => n11066, ZN => 
                           n10215);
   U16798 : XNOR2_X1 port map( A => n10219, B => n10218, ZN => n10221);
   U16799 : XNOR2_X1 port map( A => n10220, B => n10221, ZN => n10226);
   U16800 : INV_X1 port map( A => n2306, ZN => n27850);
   U16801 : XNOR2_X1 port map( A => n10222, B => n27850, ZN => n10224);
   U16802 : XNOR2_X1 port map( A => n10223, B => n10224, ZN => n10225);
   U16803 : XNOR2_X1 port map( A => n10225, B => n10226, ZN => n11218);
   U16804 : XNOR2_X1 port map( A => n10227, B => n10228, ZN => n10230);
   U16805 : XNOR2_X1 port map( A => n10229, B => n10230, ZN => n10249);
   U16806 : XNOR2_X1 port map( A => n10232, B => n10231, ZN => n10248);
   U16807 : INV_X1 port map( A => n10233, ZN => n10236);
   U16808 : INV_X1 port map( A => n10234, ZN => n10235);
   U16809 : NAND3_X1 port map( A1 => n10237, A2 => n10236, A3 => n10235, ZN => 
                           n10239);
   U16810 : INV_X1 port map( A => n3116, ZN => n27605);
   U16811 : NAND2_X1 port map( A1 => n10237, A2 => n10241, ZN => n10238);
   U16812 : NAND3_X1 port map( A1 => n10239, A2 => n27605, A3 => n10238, ZN => 
                           n10244);
   U16813 : INV_X1 port map( A => n10240, ZN => n10242);
   U16814 : NAND3_X1 port map( A1 => n10242, A2 => n10241, A3 => n27605, ZN => 
                           n10243);
   U16815 : OAI211_X1 port map( C1 => n10246, C2 => n10245, A => n10244, B => 
                           n10243, ZN => n10247);
   U16816 : XNOR2_X1 port map( A => n10254, B => n10253, ZN => n10657);
   U16817 : XNOR2_X1 port map( A => n10256, B => n10255, ZN => n10262);
   U16818 : XNOR2_X1 port map( A => n10295, B => n10257, ZN => n10260);
   U16819 : XNOR2_X1 port map( A => n10258, B => n1928, ZN => n10259);
   U16820 : XNOR2_X1 port map( A => n10260, B => n10259, ZN => n10261);
   U16821 : NOR2_X1 port map( A1 => n11222, A2 => n10876, ZN => n10269);
   U16822 : XNOR2_X1 port map( A => n10264, B => n10263, ZN => n10267);
   U16823 : XNOR2_X1 port map( A => n10265, B => n3036, ZN => n10266);
   U16825 : XNOR2_X1 port map( A => n10272, B => n3334, ZN => n10273);
   U16826 : XNOR2_X1 port map( A => n10274, B => n10273, ZN => n10279);
   U16827 : XNOR2_X1 port map( A => n10311, B => n10275, ZN => n10276);
   U16828 : XNOR2_X1 port map( A => n10277, B => n10276, ZN => n10278);
   U16830 : INV_X1 port map( A => n10876, ZN => n10871);
   U16833 : XNOR2_X1 port map( A => n10282, B => n2465, ZN => n10284);
   U16834 : XNOR2_X1 port map( A => n10288, B => n10287, ZN => n10293);
   U16835 : XNOR2_X1 port map( A => n10289, B => n1215, ZN => n10290);
   U16836 : XNOR2_X1 port map( A => n10291, B => n10290, ZN => n10292);
   U16837 : XNOR2_X1 port map( A => n10293, B => n10292, ZN => n11287);
   U16838 : XNOR2_X1 port map( A => n10294, B => n1079, ZN => n10296);
   U16839 : XNOR2_X1 port map( A => n10295, B => n10296, ZN => n10299);
   U16840 : XNOR2_X1 port map( A => n10298, B => n10297, ZN => n10417);
   U16841 : XNOR2_X1 port map( A => n10364, B => n10302, ZN => n10428);
   U16842 : XNOR2_X1 port map( A => n10303, B => n10428, ZN => n10308);
   U16843 : XNOR2_X1 port map( A => n10304, B => n2995, ZN => n10305);
   U16844 : XNOR2_X1 port map( A => n10306, B => n10305, ZN => n10307);
   U16845 : XNOR2_X1 port map( A => n10308, B => n10307, ZN => n10318);
   U16846 : OAI21_X1 port map( B1 => n11290, B2 => n11287, A => n10309, ZN => 
                           n11292);
   U16847 : XNOR2_X1 port map( A => n10310, B => n10311, ZN => n10313);
   U16848 : XNOR2_X1 port map( A => n10353, B => n1133, ZN => n10312);
   U16849 : XNOR2_X1 port map( A => n10313, B => n10312, ZN => n10317);
   U16850 : XNOR2_X1 port map( A => n10315, B => n10314, ZN => n10316);
   U16851 : XNOR2_X1 port map( A => n10316, B => n10317, ZN => n11075);
   U16852 : INV_X1 port map( A => n10318, ZN => n11072);
   U16853 : XNOR2_X1 port map( A => n10319, B => n10320, ZN => n10326);
   U16854 : XNOR2_X1 port map( A => n10321, B => n10384, ZN => n10324);
   U16855 : XNOR2_X1 port map( A => n10322, B => n2894, ZN => n10323);
   U16856 : XNOR2_X1 port map( A => n10324, B => n10323, ZN => n10325);
   U16857 : AND3_X1 port map( A1 => n10891, A2 => n11287, A3 => n29116, ZN => 
                           n10327);
   U16858 : XNOR2_X1 port map( A => n10328, B => n3049, ZN => n10329);
   U16859 : XNOR2_X1 port map( A => n10329, B => n10330, ZN => n10331);
   U16860 : XNOR2_X1 port map( A => n10331, B => n10332, ZN => n10333);
   U16861 : XNOR2_X1 port map( A => n10333, B => n10334, ZN => n10518);
   U16862 : XNOR2_X1 port map( A => n10335, B => n10384, ZN => n10336);
   U16863 : XNOR2_X1 port map( A => n10336, B => n10337, ZN => n10341);
   U16864 : XNOR2_X1 port map( A => n1852, B => n3728, ZN => n10339);
   U16865 : XNOR2_X1 port map( A => n10338, B => n10339, ZN => n10340);
   U16866 : NAND2_X1 port map( A1 => n11027, A2 => n11282, ZN => n11286);
   U16867 : XNOR2_X1 port map( A => n10342, B => n10343, ZN => n10349);
   U16868 : XNOR2_X1 port map( A => n10344, B => n10345, ZN => n10348);
   U16869 : XNOR2_X1 port map( A => n28643, B => n900, ZN => n10347);
   U16870 : INV_X1 port map( A => n2986, ZN => n24060);
   U16871 : XNOR2_X1 port map( A => n10350, B => n24060, ZN => n10351);
   U16872 : XNOR2_X1 port map( A => n10351, B => n10352, ZN => n10355);
   U16873 : XNOR2_X1 port map( A => n10355, B => n10354, ZN => n10361);
   U16874 : XNOR2_X1 port map( A => n10357, B => n10356, ZN => n10358);
   U16875 : XNOR2_X1 port map( A => n10359, B => n10358, ZN => n10360);
   U16876 : XNOR2_X1 port map( A => n10361, B => n10360, ZN => n10517);
   U16877 : XNOR2_X1 port map( A => n10363, B => n10362, ZN => n10366);
   U16878 : XNOR2_X1 port map( A => n10364, B => n3463, ZN => n10365);
   U16879 : XNOR2_X1 port map( A => n10366, B => n10365, ZN => n10370);
   U16880 : XNOR2_X1 port map( A => n10368, B => n10367, ZN => n10369);
   U16881 : NAND3_X1 port map( A1 => n585, A2 => n10517, A3 => n10884, ZN => 
                           n10381);
   U16882 : INV_X1 port map( A => n10517, ZN => n11283);
   U16884 : XNOR2_X1 port map( A => n10371, B => n10372, ZN => n10374);
   U16885 : XNOR2_X1 port map( A => n10373, B => n10374, ZN => n10378);
   U16886 : XNOR2_X1 port map( A => n10395, B => n3673, ZN => n10375);
   U16887 : XNOR2_X1 port map( A => n10376, B => n10375, ZN => n10377);
   U16888 : NAND3_X1 port map( A1 => n10517, A2 => n584, A3 => n11281, ZN => 
                           n10379);
   U16889 : XNOR2_X1 port map( A => n10383, B => n10382, ZN => n10390);
   U16890 : XNOR2_X1 port map( A => n10384, B => n3710, ZN => n10388);
   U16891 : XNOR2_X1 port map( A => n10386, B => n10385, ZN => n10387);
   U16892 : XNOR2_X1 port map( A => n10388, B => n10387, ZN => n10389);
   U16893 : XNOR2_X1 port map( A => n10391, B => n10392, ZN => n10394);
   U16894 : XNOR2_X1 port map( A => n10393, B => n10394, ZN => n10400);
   U16895 : XNOR2_X1 port map( A => n10396, B => n10395, ZN => n10398);
   U16896 : INV_X1 port map( A => n3508, ZN => n26899);
   U16897 : XNOR2_X1 port map( A => n5412, B => n26899, ZN => n10397);
   U16898 : XNOR2_X1 port map( A => n10398, B => n10397, ZN => n10399);
   U16899 : NOR2_X1 port map( A1 => n10401, A2 => n3787, ZN => n10402);
   U16900 : NAND3_X1 port map( A1 => n10407, A2 => n3787, A3 => n10406, ZN => 
                           n10408);
   U16902 : XNOR2_X1 port map( A => n10411, B => n1918, ZN => n10413);
   U16903 : XNOR2_X1 port map( A => n10414, B => n10413, ZN => n10416);
   U16904 : XNOR2_X1 port map( A => n10417, B => n10418, ZN => n10423);
   U16905 : XNOR2_X1 port map( A => n10419, B => n3062, ZN => n10420);
   U16906 : XNOR2_X1 port map( A => n10421, B => n10420, ZN => n10422);
   U16907 : XNOR2_X1 port map( A => n10422, B => n10423, ZN => n11204);
   U16908 : INV_X1 port map( A => n11204, ZN => n11090);
   U16909 : XNOR2_X1 port map( A => n10425, B => n10424, ZN => n10430);
   U16910 : XNOR2_X1 port map( A => n10426, B => n3598, ZN => n10427);
   U16911 : XNOR2_X1 port map( A => n10428, B => n10427, ZN => n10429);
   U16913 : NOR2_X1 port map( A1 => n11204, A2 => n11206, ZN => n10637);
   U16914 : XNOR2_X1 port map( A => n10432, B => n10433, ZN => n10440);
   U16915 : XNOR2_X1 port map( A => n10435, B => n10434, ZN => n10438);
   U16916 : XNOR2_X1 port map( A => n10436, B => n3554, ZN => n10437);
   U16917 : XNOR2_X1 port map( A => n10438, B => n10437, ZN => n10439);
   U16918 : XNOR2_X1 port map( A => n10440, B => n10439, ZN => n11093);
   U16919 : XNOR2_X1 port map( A => n13144, B => n10442, ZN => n10443);
   U16920 : INV_X1 port map( A => n13606, ZN => n14102);
   U16921 : NAND2_X1 port map( A1 => n10705, A2 => n28495, ZN => n10448);
   U16922 : NOR2_X1 port map( A1 => n10592, A2 => n28495, ZN => n10706);
   U16923 : NAND2_X1 port map( A1 => n10912, A2 => n10911, ZN => n10449);
   U16924 : NAND2_X1 port map( A1 => n10732, A2 => n10449, ZN => n10450);
   U16925 : NAND2_X1 port map( A1 => n10450, A2 => n10735, ZN => n10451);
   U16926 : NOR2_X1 port map( A1 => n10711, A2 => n10715, ZN => n10454);
   U16927 : NAND2_X1 port map( A1 => n10499, A2 => n10454, ZN => n10456);
   U16928 : OAI211_X1 port map( C1 => n10457, C2 => n2646, A => n10456, B => 
                           n10455, ZN => n10868);
   U16929 : NAND2_X1 port map( A1 => n10458, A2 => n10726, ZN => n10926);
   U16930 : NAND2_X1 port map( A1 => n10926, A2 => n10459, ZN => n10460);
   U16931 : AND3_X1 port map( A1 => n3862, A2 => n11138, A3 => n10718, ZN => 
                           n10767);
   U16932 : INV_X1 port map( A => n11876, ZN => n10464);
   U16933 : NAND2_X1 port map( A1 => n10464, A2 => n287, ZN => n10465);
   U16934 : NOR2_X1 port map( A1 => n10745, A2 => n11168, ZN => n10471);
   U16935 : INV_X1 port map( A => n11168, ZN => n11170);
   U16936 : NAND2_X1 port map( A1 => n11166, A2 => n11170, ZN => n10466);
   U16937 : NAND2_X1 port map( A1 => n10467, A2 => n11330, ZN => n11332);
   U16938 : NOR2_X1 port map( A1 => n10821, A2 => n11170, ZN => n10468);
   U16939 : AOI21_X1 port map( B1 => n10469, B2 => n11332, A => n10468, ZN => 
                           n10470);
   U16941 : NAND3_X1 port map( A1 => n11184, A2 => n11181, A3 => n10810, ZN => 
                           n10474);
   U16943 : OAI21_X1 port map( B1 => n11349, B2 => n11192, A => n10478, ZN => 
                           n10479);
   U16944 : NAND2_X1 port map( A1 => n11022, A2 => n11255, ZN => n10484);
   U16946 : NOR2_X1 port map( A1 => n10855, A2 => n11165, ZN => n10487);
   U16947 : INV_X1 port map( A => n10855, ZN => n11164);
   U16948 : NOR2_X1 port map( A1 => n11164, A2 => n11053, ZN => n10486);
   U16949 : INV_X1 port map( A => n12338, ZN => n11913);
   U16950 : OAI21_X1 port map( B1 => n12343, B2 => n11913, A => n12339, ZN => 
                           n10489);
   U16951 : XNOR2_X1 port map( A => n13097, B => n13227, ZN => n10539);
   U16953 : AOI21_X1 port map( B1 => n10554, B2 => n10494, A => n11154, ZN => 
                           n10495);
   U16954 : MUX2_X1 port map( A => n10499, B => n10498, S => n10497, Z => 
                           n10503);
   U16955 : MUX2_X1 port map( A => n10506, B => n10505, S => n4024, Z => n10509
                           );
   U16956 : OAI21_X1 port map( B1 => n11461, B2 => n1836, A => n11874, ZN => 
                           n10516);
   U16958 : NAND2_X1 port map( A1 => n11500, A2 => n11458, ZN => n11870);
   U16962 : INV_X1 port map( A => n10518, ZN => n11280);
   U16963 : MUX2_X1 port map( A => n10520, B => n10519, S => n11284, Z => 
                           n10521);
   U16964 : INV_X1 port map( A => n11449, ZN => n11888);
   U16966 : INV_X1 port map( A => n11037, ZN => n11273);
   U16967 : INV_X1 port map( A => n12328, ZN => n11884);
   U16968 : OAI21_X1 port map( B1 => n11888, B2 => n11884, A => n11747, ZN => 
                           n10531);
   U16969 : INV_X1 port map( A => n10528, ZN => n11266);
   U16970 : NOR2_X1 port map( A1 => n11261, A2 => n11047, ZN => n10530);
   U16971 : NAND2_X1 port map( A1 => n10530, A2 => n28204, ZN => n11886);
   U16972 : INV_X1 port map( A => n12327, ZN => n12333);
   U16973 : NAND2_X1 port map( A1 => n10665, A2 => n11076, ZN => n10894);
   U16974 : INV_X1 port map( A => n11287, ZN => n10893);
   U16975 : INV_X1 port map( A => n11075, ZN => n11291);
   U16976 : NAND2_X1 port map( A1 => n11291, A2 => n11072, ZN => n10532);
   U16977 : INV_X1 port map( A => n11223, ZN => n10878);
   U16978 : XNOR2_X1 port map( A => n10539, B => n10538, ZN => n10619);
   U16979 : NOR2_X1 port map( A1 => n11119, A2 => n11118, ZN => n10542);
   U16980 : INV_X1 port map( A => n11120, ZN => n11125);
   U16981 : NAND2_X1 port map( A1 => n11125, A2 => n11124, ZN => n10541);
   U16982 : OAI21_X1 port map( B1 => n10805, B2 => n11146, A => n10543, ZN => 
                           n10546);
   U16983 : NOR2_X2 port map( A1 => n10546, A2 => n10545, ZN => n11754);
   U16984 : OAI21_X1 port map( B1 => n10548, B2 => n10461, A => n10547, ZN => 
                           n10552);
   U16985 : NAND2_X1 port map( A1 => n29150, A2 => n11113, ZN => n10551);
   U16986 : OAI21_X1 port map( B1 => n11111, B2 => n11113, A => n10549, ZN => 
                           n10550);
   U16987 : NAND2_X1 port map( A1 => n10555, A2 => n11158, ZN => n10557);
   U16988 : AOI21_X1 port map( B1 => n11338, B2 => n11337, A => n10828, ZN => 
                           n10561);
   U16989 : NOR2_X1 port map( A1 => n10558, A2 => n11176, ZN => n10827);
   U16990 : NOR2_X1 port map( A1 => n10830, A2 => n1898, ZN => n10559);
   U16991 : OAI21_X1 port map( B1 => n10827, B2 => n10559, A => n11341, ZN => 
                           n10560);
   U16992 : OAI21_X1 port map( B1 => n11345, B2 => n10561, A => n10560, ZN => 
                           n11755);
   U16993 : NOR2_X1 port map( A1 => n10748, A2 => n10814, ZN => n10815);
   U16994 : NOR2_X1 port map( A1 => n11198, A2 => n10563, ZN => n10564);
   U16996 : NOR3_X1 port map( A1 => n5914, A2 => n5917, A3 => n28157, ZN => 
                           n10566);
   U16997 : XNOR2_X1 port map( A => n13226, B => n3752, ZN => n10617);
   U16998 : INV_X1 port map( A => n10797, ZN => n11232);
   U16999 : INV_X1 port map( A => n11225, ZN => n10794);
   U17000 : NAND3_X1 port map( A1 => n11099, A2 => n6814, A3 => n10794, ZN => 
                           n11899);
   U17001 : OAI211_X1 port map( C1 => n11066, C2 => n11244, A => n11240, B => 
                           n1851, ZN => n10571);
   U17002 : INV_X1 port map( A => n11240, ZN => n11063);
   U17003 : NAND3_X1 port map( A1 => n10640, A2 => n11063, A3 => n11069, ZN => 
                           n10570);
   U17004 : NAND2_X1 port map( A1 => n12352, A2 => n11901, ZN => n11468);
   U17005 : MUX2_X1 port map( A => n11212, B => n11213, S => n433, Z => n10575)
                           ;
   U17006 : NAND2_X1 port map( A1 => n433, A2 => n11211, ZN => n10573);
   U17007 : OAI21_X2 port map( B1 => n10575, B2 => n10574, A => n10573, ZN => 
                           n12350);
   U17008 : INV_X1 port map( A => n12350, ZN => n10586);
   U17009 : AND2_X1 port map( A1 => n11205, A2 => n10576, ZN => n10578);
   U17010 : NAND2_X1 port map( A1 => n10579, A2 => n11013, ZN => n10583);
   U17011 : NAND3_X1 port map( A1 => n10628, A2 => n5710, A3 => n3441, ZN => 
                           n10582);
   U17013 : NAND2_X1 port map( A1 => n29648, A2 => n11237, ZN => n11239);
   U17014 : INV_X1 port map( A => n11239, ZN => n10580);
   U17015 : NAND2_X1 port map( A1 => n10580, A2 => n10776, ZN => n10581);
   U17017 : AOI22_X1 port map( A1 => n10989, A2 => n3804, B1 => n10983, B2 => 
                           n10984, ZN => n10585);
   U17019 : MUX2_X1 port map( A => n28405, B => n10999, S => n11003, Z => 
                           n10589);
   U17020 : NOR2_X1 port map( A1 => n10589, A2 => n10936, ZN => n10590);
   U17021 : NAND2_X1 port map( A1 => n10592, A2 => n28495, ZN => n10944);
   U17023 : AOI21_X1 port map( B1 => n10702, B2 => n28176, A => n10946, ZN => 
                           n10595);
   U17024 : INV_X1 port map( A => n10995, ZN => n10787);
   U17025 : NAND2_X1 port map( A1 => n10693, A2 => n10597, ZN => n10601);
   U17026 : OAI21_X1 port map( B1 => n10992, B2 => n10991, A => n3454, ZN => 
                           n10600);
   U17027 : INV_X1 port map( A => n10991, ZN => n10598);
   U17028 : NOR2_X1 port map( A1 => n10598, A2 => n10787, ZN => n10599);
   U17029 : INV_X1 port map( A => n10602, ZN => n10964);
   U17030 : OAI21_X1 port map( B1 => n896, B2 => n9858, A => n10964, ZN => 
                           n10604);
   U17031 : INV_X1 port map( A => n10962, ZN => n10778);
   U17033 : NAND2_X1 port map( A1 => n11740, A2 => n12356, ZN => n10898);
   U17034 : INV_X1 port map( A => n10911, ZN => n10915);
   U17037 : INV_X1 port map( A => n12362, ZN => n11741);
   U17038 : AOI21_X1 port map( B1 => n10611, B2 => n10898, A => n11741, ZN => 
                           n10616);
   U17041 : NOR2_X1 port map( A1 => n10616, A2 => n10615, ZN => n12594);
   U17042 : INV_X1 port map( A => n12594, ZN => n13381);
   U17043 : XNOR2_X1 port map( A => n13381, B => n12593, ZN => n12654);
   U17044 : XNOR2_X1 port map( A => n12654, B => n10617, ZN => n10618);
   U17045 : XNOR2_X2 port map( A => n10619, B => n10618, ZN => n14593);
   U17046 : NAND2_X1 port map( A1 => n14102, A2 => n14593, ZN => n11372);
   U17048 : MUX2_X1 port map( A => n10624, B => n10623, S => n10797, Z => 
                           n10625);
   U17049 : NOR2_X2 port map( A1 => n10626, A2 => n10625, ZN => n12220);
   U17050 : NOR2_X1 port map( A1 => n6108, A2 => n11013, ZN => n10627);
   U17052 : INV_X1 port map( A => n10981, ZN => n10985);
   U17053 : INV_X1 port map( A => n10631, ZN => n10632);
   U17054 : NAND2_X1 port map( A1 => n10632, A2 => n10783, ZN => n10633);
   U17055 : MUX2_X1 port map( A => n12220, B => n28726, S => n12218, Z => 
                           n10645);
   U17056 : NAND2_X1 port map( A1 => n10785, A2 => n10786, ZN => n10635);
   U17057 : NAND2_X1 port map( A1 => n10995, A2 => n10786, ZN => n10994);
   U17058 : OAI211_X1 port map( C1 => n10785, C2 => n4538, A => n10992, B => 
                           n10994, ZN => n11693);
   U17059 : INV_X1 port map( A => n12218, ZN => n12041);
   U17060 : INV_X1 port map( A => n10637, ZN => n10638);
   U17061 : NOR2_X1 port map( A1 => n11069, A2 => n11066, ZN => n10639);
   U17062 : NAND3_X1 port map( A1 => n11066, A2 => n11242, A3 => n11244, ZN => 
                           n10642);
   U17063 : INV_X1 port map( A => n11066, ZN => n10641);
   U17064 : OAI22_X1 port map( A1 => n10643, A2 => n12224, B1 => n12042, B2 => 
                           n11962, ZN => n10644);
   U17065 : XNOR2_X1 port map( A => n13359, B => n3114, ZN => n10677);
   U17066 : NAND2_X1 port map( A1 => n431, A2 => n12337, ZN => n12027);
   U17067 : NAND2_X1 port map( A1 => n12343, A2 => n12338, ZN => n10646);
   U17069 : NAND2_X1 port map( A1 => n10647, A2 => n1291, ZN => n10651);
   U17071 : AOI22_X1 port map( A1 => n10649, A2 => n12026, B1 => n10648, B2 => 
                           n12339, ZN => n10650);
   U17073 : NOR2_X1 port map( A1 => n11280, A2 => n11282, ZN => n10652);
   U17074 : INV_X1 port map( A => n11281, ZN => n11029);
   U17075 : AOI22_X1 port map( A1 => n10883, A2 => n11086, B1 => n11211, B2 => 
                           n11212, ZN => n10656);
   U17076 : NAND2_X1 port map( A1 => n1986, A2 => n375, ZN => n11682);
   U17077 : MUX2_X1 port map( A => n11218, B => n10872, S => n10659, Z => 
                           n10658);
   U17078 : NAND2_X1 port map( A1 => n10659, A2 => n29593, ZN => n10661);
   U17079 : OAI22_X1 port map( A1 => n10872, A2 => n10661, B1 => n10660, B2 => 
                           n10876, ZN => n10662);
   U17080 : OAI21_X1 port map( B1 => n10893, B2 => n10665, A => n10664, ZN => 
                           n10667);
   U17081 : NAND3_X1 port map( A1 => n11290, A2 => n11072, A3 => n29116, ZN => 
                           n10666);
   U17082 : NAND2_X1 port map( A1 => n11048, A2 => n11261, ZN => n10670);
   U17083 : INV_X1 port map( A => n11047, ZN => n10888);
   U17084 : NAND3_X1 port map( A1 => n11979, A2 => n12232, A3 => n12233, ZN => 
                           n10675);
   U17085 : OAI21_X2 port map( B1 => n10673, B2 => n11274, A => n10672, ZN => 
                           n12234);
   U17086 : NAND4_X2 port map( A1 => n11977, A2 => n10676, A3 => n10674, A4 => 
                           n10675, ZN => n13337);
   U17087 : XNOR2_X1 port map( A => n12560, B => n13337, ZN => n13549);
   U17088 : XNOR2_X1 port map( A => n13549, B => n10677, ZN => n10773);
   U17089 : NAND2_X1 port map( A1 => n10973, A2 => n29577, ZN => n10679);
   U17090 : MUX2_X1 port map( A => n10679, B => n10678, S => n10681, Z => 
                           n11495);
   U17091 : MUX2_X1 port map( A => n10936, B => n6779, S => n10937, Z => n10685
                           );
   U17092 : INV_X1 port map( A => n12304, ZN => n10701);
   U17093 : OAI21_X1 port map( B1 => n10913, B2 => n10916, A => n10688, ZN => 
                           n10737);
   U17094 : NAND2_X1 port map( A1 => n10690, A2 => n10913, ZN => n11494);
   U17095 : NAND2_X1 port map( A1 => n10791, A2 => n3454, ZN => n10692);
   U17096 : NAND2_X1 port map( A1 => n12304, A2 => n12303, ZN => n10700);
   U17097 : INV_X1 port map( A => n10983, ZN => n10694);
   U17099 : MUX2_X1 port map( A => n10695, B => n589, S => n10783, Z => n10699)
                           ;
   U17101 : INV_X1 port map( A => n10982, ZN => n10988);
   U17102 : NAND2_X1 port map( A1 => n10701, A2 => n11491, ZN => n11363);
   U17104 : NAND2_X1 port map( A1 => n10706, A2 => n10705, ZN => n10707);
   U17105 : OAI211_X1 port map( C1 => n10710, C2 => n10110, A => n10708, B => 
                           n10707, ZN => n11794);
   U17106 : NAND2_X1 port map( A1 => n10711, A2 => n10715, ZN => n10712);
   U17107 : AOI21_X1 port map( B1 => n10715, B2 => n10714, A => n10713, ZN => 
                           n10716);
   U17108 : OAI21_X1 port map( B1 => n3862, B2 => n2968, A => n10919, ZN => 
                           n10720);
   U17109 : OAI21_X1 port map( B1 => n10721, B2 => n10720, A => n10719, ZN => 
                           n10722);
   U17110 : NAND2_X1 port map( A1 => n6482, A2 => n11486, ZN => n11718);
   U17111 : OAI21_X1 port map( B1 => n10976, B2 => n29577, A => n10970, ZN => 
                           n10724);
   U17112 : NAND2_X1 port map( A1 => n11718, A2 => n11430, ZN => n10731);
   U17113 : OAI21_X1 port map( B1 => n10924, B2 => n10927, A => n590, ZN => 
                           n10729);
   U17115 : NAND2_X1 port map( A1 => n10731, A2 => n28436, ZN => n10739);
   U17116 : NAND2_X1 port map( A1 => n10737, A2 => n10732, ZN => n10734);
   U17117 : NAND2_X1 port map( A1 => n10734, A2 => n10733, ZN => n11428);
   U17118 : NAND2_X1 port map( A1 => n10735, A2 => n10916, ZN => n10736);
   U17120 : INV_X1 port map( A => n11486, ZN => n11431);
   U17121 : NAND3_X1 port map( A1 => n11487, A2 => n11431, A3 => n2194, ZN => 
                           n10738);
   U17122 : XNOR2_X1 port map( A => n13036, B => n12919, ZN => n12065);
   U17123 : INV_X1 port map( A => n11166, ZN => n10819);
   U17124 : MUX2_X1 port map( A => n28638, B => n28157, S => n10563, Z => 
                           n10750);
   U17125 : OAI21_X1 port map( B1 => n11152, B2 => n10752, A => n28175, ZN => 
                           n10753);
   U17126 : NAND2_X1 port map( A1 => n10753, A2 => n10803, ZN => n10756);
   U17128 : NOR2_X1 port map( A1 => n11401, A2 => n11672, ZN => n10758);
   U17129 : INV_X1 port map( A => n10828, ZN => n11336);
   U17130 : NAND2_X1 port map( A1 => n11341, A2 => n11176, ZN => n10757);
   U17131 : OR2_X1 port map( A1 => n11340, A2 => n1898, ZN => n11634);
   U17132 : INV_X1 port map( A => n11515, ZN => n11845);
   U17133 : OAI21_X1 port map( B1 => n11677, B2 => n10758, A => n11845, ZN => 
                           n10765);
   U17134 : NOR2_X1 port map( A1 => n11640, A2 => n29139, ZN => n10763);
   U17135 : NAND2_X1 port map( A1 => n11120, A2 => n11124, ZN => n10759);
   U17136 : AOI21_X1 port map( B1 => n10760, B2 => n10759, A => n11119, ZN => 
                           n10762);
   U17137 : NOR2_X1 port map( A1 => n11124, A2 => n11123, ZN => n10761);
   U17138 : INV_X1 port map( A => n11848, ZN => n11641);
   U17139 : AOI22_X1 port map( A1 => n10763, A2 => n11515, B1 => n11641, B2 => 
                           n11401, ZN => n10764);
   U17140 : INV_X1 port map( A => n10868, ZN => n11583);
   U17141 : NAND2_X1 port map( A1 => n11877, A2 => n11583, ZN => n10771);
   U17142 : INV_X1 port map( A => n11881, ZN => n11582);
   U17143 : INV_X1 port map( A => n10766, ZN => n10769);
   U17144 : INV_X1 port map( A => n10767, ZN => n10768);
   U17145 : NAND4_X1 port map( A1 => n10769, A2 => n11583, A3 => n10768, A4 => 
                           n10453, ZN => n10770);
   U17146 : XNOR2_X1 port map( A => n13109, B => n13547, ZN => n13237);
   U17147 : XNOR2_X1 port map( A => n13237, B => n12065, ZN => n10772);
   U17148 : NOR2_X1 port map( A1 => n29648, A2 => n11235, ZN => n10775);
   U17149 : NOR2_X1 port map( A1 => n11012, A2 => n10776, ZN => n10777);
   U17151 : OAI21_X1 port map( B1 => n9362, B2 => n10962, A => n10958, ZN => 
                           n10781);
   U17154 : AND3_X1 port map( A1 => n10980, A2 => n10988, A3 => n589, ZN => 
                           n10784);
   U17155 : INV_X1 port map( A => n10784, ZN => n12094);
   U17156 : MUX2_X1 port map( A => n10785, B => n10787, S => n10786, Z => 
                           n10792);
   U17157 : NAND2_X1 port map( A1 => n10791, A2 => n10991, ZN => n10789);
   U17158 : NAND2_X1 port map( A1 => n10787, A2 => n10786, ZN => n10788);
   U17159 : MUX2_X1 port map( A => n10789, B => n10788, S => n3454, Z => n10790
                           );
   U17160 : OAI21_X1 port map( B1 => n10792, B2 => n10791, A => n10790, ZN => 
                           n11385);
   U17161 : INV_X1 port map( A => n11385, ZN => n12100);
   U17162 : AND2_X1 port map( A1 => n11099, A2 => n333, ZN => n11893);
   U17163 : NAND2_X1 port map( A1 => n6814, A2 => n10795, ZN => n10796);
   U17164 : NAND2_X1 port map( A1 => n11896, A2 => n10797, ZN => n10798);
   U17165 : AOI21_X1 port map( B1 => n12100, B2 => n12155, A => n12088, ZN => 
                           n10801);
   U17166 : NOR2_X1 port map( A1 => n10431, A2 => n11093, ZN => n10800);
   U17167 : OAI21_X1 port map( B1 => n11206, B2 => n587, A => n11207, ZN => 
                           n10799);
   U17168 : MUX2_X1 port map( A => n10800, B => n10799, S => n11094, Z => 
                           n12091);
   U17169 : NOR2_X1 port map( A1 => n11205, A2 => n29517, ZN => n12092);
   U17170 : OAI21_X1 port map( B1 => n11146, B2 => n10806, A => n10805, ZN => 
                           n10807);
   U17171 : OAI211_X1 port map( C1 => n10808, C2 => n11149, A => n11146, B => 
                           n28627, ZN => n10809);
   U17172 : AOI22_X1 port map( A1 => n11322, A2 => n11323, B1 => n11321, B2 => 
                           n10810, ZN => n10811);
   U17173 : NOR2_X1 port map( A1 => n10811, A2 => n11183, ZN => n10812);
   U17174 : NOR3_X1 port map( A1 => n581, A2 => n11198, A3 => n28157, ZN => 
                           n10817);
   U17175 : INV_X1 port map( A => n11646, ZN => n11645);
   U17176 : NAND2_X1 port map( A1 => n11645, A2 => n11715, ZN => n11414);
   U17177 : INV_X1 port map( A => n10821, ZN => n11329);
   U17178 : OR2_X1 port map( A1 => n10823, A2 => n11331, ZN => n10824);
   U17179 : NOR2_X1 port map( A1 => n11335, A2 => n11176, ZN => n10826);
   U17180 : NOR2_X1 port map( A1 => n11338, A2 => n434, ZN => n10825);
   U17181 : MUX2_X1 port map( A => n10826, B => n10825, S => n11345, Z => 
                           n10832);
   U17182 : INV_X1 port map( A => n10827, ZN => n11179);
   U17183 : NAND3_X1 port map( A1 => n11176, A2 => n11174, A3 => n1898, ZN => 
                           n10829);
   U17184 : OAI21_X1 port map( B1 => n11179, B2 => n10830, A => n10829, ZN => 
                           n10831);
   U17185 : XNOR2_X1 port map( A => n12723, B => n13386, ZN => n10867);
   U17186 : NAND2_X1 port map( A1 => n586, A2 => n10833, ZN => n10837);
   U17187 : AND2_X1 port map( A1 => n10834, A2 => n11252, ZN => n11250);
   U17188 : INV_X1 port map( A => n11250, ZN => n10835);
   U17189 : MUX2_X1 port map( A => n10837, B => n10836, S => n29148, Z => 
                           n10841);
   U17190 : INV_X1 port map( A => n10838, ZN => n10839);
   U17191 : NAND2_X1 port map( A1 => n10839, A2 => n11033, ZN => n10840);
   U17192 : NAND2_X1 port map( A1 => n11034, A2 => n279, ZN => n10843);
   U17193 : NAND3_X1 port map( A1 => n10847, A2 => n11350, A3 => n11347, ZN => 
                           n10848);
   U17194 : INV_X1 port map( A => n11347, ZN => n11191);
   U17195 : OAI21_X1 port map( B1 => n11349, B2 => n11348, A => n10849, ZN => 
                           n10850);
   U17196 : NOR2_X1 port map( A1 => n11308, A2 => n10851, ZN => n10854);
   U17197 : INV_X1 port map( A => n11053, ZN => n11312);
   U17198 : AOI22_X1 port map( A1 => n10854, A2 => n1933, B1 => n10852, B2 => 
                           n10851, ZN => n10857);
   U17199 : INV_X1 port map( A => n11321, ZN => n10858);
   U17200 : NAND3_X1 port map( A1 => n11184, A2 => n10858, A3 => n10473, ZN => 
                           n10860);
   U17201 : OAI21_X1 port map( B1 => n12037, B2 => n12241, A => n10861, ZN => 
                           n12239);
   U17203 : OAI211_X1 port map( C1 => n3653, C2 => n12507, A => n12512, B => 
                           n11990, ZN => n10865);
   U17204 : XNOR2_X1 port map( A => n11684, B => n10867, ZN => n10904);
   U17205 : NAND2_X1 port map( A1 => n11878, A2 => n11877, ZN => n10870);
   U17206 : INV_X1 port map( A => n13195, ZN => n12914);
   U17207 : NAND2_X1 port map( A1 => n10871, A2 => n435, ZN => n10874);
   U17209 : MUX2_X1 port map( A => n10874, B => n28329, S => n11220, Z => 
                           n11658);
   U17210 : INV_X1 port map( A => n11217, ZN => n10879);
   U17211 : NOR2_X1 port map( A1 => n10876, A2 => n435, ZN => n10877);
   U17212 : AOI22_X1 port map( A1 => n10879, A2 => n10878, B1 => n10877, B2 => 
                           n11222, ZN => n11657);
   U17213 : AOI21_X1 port map( B1 => n11063, B2 => n11242, A => n11243, ZN => 
                           n10881);
   U17214 : INV_X1 port map( A => n10882, ZN => n11083);
   U17215 : NAND2_X1 port map( A1 => n1854, A2 => n10884, ZN => n11028);
   U17216 : NAND3_X1 port map( A1 => n11027, A2 => n11284, A3 => n11281, ZN => 
                           n10886);
   U17217 : OAI211_X1 port map( C1 => n11283, C2 => n10884, A => n11029, B => 
                           n584, ZN => n10885);
   U17218 : INV_X1 port map( A => n12164, ZN => n10887);
   U17219 : OAI21_X1 port map( B1 => n1931, B2 => n12163, A => n10887, ZN => 
                           n10897);
   U17220 : AND2_X1 port map( A1 => n11264, A2 => n11267, ZN => n10890);
   U17221 : OAI21_X1 port map( B1 => n10890, B2 => n29510, A => n10889, ZN => 
                           n11656);
   U17223 : MUX2_X1 port map( A => n11294, B => n11290, S => n10318, Z => 
                           n11659);
   U17224 : AND2_X1 port map( A1 => n11659, A2 => n29116, ZN => n10895);
   U17225 : XNOR2_X1 port map( A => n12914, B => n13556, ZN => n10902);
   U17226 : NOR2_X1 port map( A1 => n12359, A2 => n12362, ZN => n10900);
   U17227 : INV_X1 port map( A => n12356, ZN => n11907);
   U17228 : XNOR2_X1 port map( A => n13101, B => n3742, ZN => n10901);
   U17229 : XNOR2_X1 port map( A => n10902, B => n10901, ZN => n10903);
   U17230 : XNOR2_X1 port map( A => n10904, B => n10903, ZN => n14105);
   U17231 : NAND2_X1 port map( A1 => n11547, A2 => n11855, ZN => n10907);
   U17232 : MUX2_X1 port map( A => n10907, B => n10906, S => n11549, Z => 
                           n10910);
   U17233 : NAND3_X1 port map( A1 => n11137, A2 => n10918, A3 => n10919, ZN => 
                           n10922);
   U17234 : NAND2_X1 port map( A1 => n1879, A2 => n10924, ZN => n10925);
   U17235 : AOI21_X1 port map( B1 => n10926, B2 => n10925, A => n590, ZN => 
                           n10935);
   U17236 : NAND2_X1 port map( A1 => n10930, A2 => n10929, ZN => n10931);
   U17237 : NAND2_X1 port map( A1 => n11951, A2 => n11861, ZN => n10955);
   U17238 : NOR2_X1 port map( A1 => n11002, A2 => n592, ZN => n10938);
   U17239 : INV_X1 port map( A => n11944, ZN => n11857);
   U17240 : OAI22_X1 port map( A1 => n10944, A2 => n10946, B1 => n10943, B2 => 
                           n10942, ZN => n10945);
   U17241 : NAND2_X1 port map( A1 => n10949, A2 => n28608, ZN => n10951);
   U17242 : NAND3_X1 port map( A1 => n11862, A2 => n11945, A3 => n11943, ZN => 
                           n10953);
   U17243 : INV_X1 port map( A => n11859, ZN => n11948);
   U17244 : NOR2_X1 port map( A1 => n10956, A2 => n10963, ZN => n10961);
   U17245 : NAND2_X1 port map( A1 => n10963, A2 => n10962, ZN => n10965);
   U17246 : NOR2_X1 port map( A1 => n29577, A2 => n10970, ZN => n10974);
   U17247 : OAI21_X1 port map( B1 => n10974, B2 => n10973, A => n10972, ZN => 
                           n10979);
   U17248 : OAI211_X1 port map( C1 => n10983, C2 => n10982, A => n10981, B => 
                           n10980, ZN => n10987);
   U17249 : NAND3_X1 port map( A1 => n10985, A2 => n10988, A3 => n10984, ZN => 
                           n10986);
   U17251 : AOI21_X1 port map( B1 => n10999, B2 => n10998, A => n10997, ZN => 
                           n11009);
   U17252 : NOR2_X1 port map( A1 => n5573, A2 => n11000, ZN => n11001);
   U17253 : NOR2_X1 port map( A1 => n11001, A2 => n28405, ZN => n11008);
   U17254 : NAND2_X1 port map( A1 => n11005, A2 => n28405, ZN => n11006);
   U17255 : NOR2_X1 port map( A1 => n3441, A2 => n11010, ZN => n11011);
   U17256 : NAND2_X1 port map( A1 => n11237, A2 => n11011, ZN => n11018);
   U17257 : NAND3_X1 port map( A1 => n5709, A2 => n11236, A3 => n11014, ZN => 
                           n11015);
   U17258 : NOR2_X1 port map( A1 => n12252, A2 => n12253, ZN => n11019);
   U17259 : AOI22_X1 port map( A1 => n11020, A2 => n12070, B1 => n11019, B2 => 
                           n349, ZN => n11021);
   U17260 : AND2_X1 port map( A1 => n11022, A2 => n11315, ZN => n11319);
   U17261 : NAND2_X1 port map( A1 => n11319, A2 => n11258, ZN => n11025);
   U17262 : NAND4_X1 port map( A1 => n11317, A2 => n11025, A3 => n11024, A4 => 
                           n11023, ZN => n12263);
   U17263 : INV_X1 port map( A => n12263, ZN => n12133);
   U17264 : NAND2_X1 port map( A1 => n11282, A2 => n11281, ZN => n11026);
   U17266 : INV_X1 port map( A => n11028, ZN => n11031);
   U17267 : NOR2_X1 port map( A1 => n11280, A2 => n11029, ZN => n11030);
   U17268 : OAI21_X1 port map( B1 => n12133, B2 => n11435, A => n12132, ZN => 
                           n11062);
   U17269 : NAND2_X1 port map( A1 => n11273, A2 => n28612, ZN => n11036);
   U17271 : MUX2_X1 port map( A => n11036, B => n11035, S => n28147, Z => 
                           n11042);
   U17272 : NAND2_X1 port map( A1 => n12133, A2 => n11574, ZN => n11928);
   U17273 : INV_X1 port map( A => n11928, ZN => n11061);
   U17274 : AOI21_X1 port map( B1 => n11045, B2 => n11266, A => n11267, ZN => 
                           n11046);
   U17275 : NAND2_X1 port map( A1 => n11262, A2 => n11046, ZN => n11050);
   U17276 : NAND3_X1 port map( A1 => n11048, A2 => n11047, A3 => n11266, ZN => 
                           n11049);
   U17277 : NAND2_X1 port map( A1 => n10855, A2 => n11165, ZN => n11052);
   U17278 : NAND2_X1 port map( A1 => n11164, A2 => n11053, ZN => n11054);
   U17279 : OAI211_X1 port map( C1 => n11057, C2 => n29637, A => n11055, B => 
                           n11054, ZN => n12264);
   U17280 : NAND3_X1 port map( A1 => n12134, A2 => n11574, A3 => n12267, ZN => 
                           n11059);
   U17281 : XNOR2_X1 port map( A => n12827, B => n13371, ZN => n12466);
   U17282 : XNOR2_X1 port map( A => n12087, B => n12466, ZN => n11203);
   U17283 : NOR2_X1 port map( A1 => n1900, A2 => n11063, ZN => n11065);
   U17284 : NAND2_X1 port map( A1 => n1900, A2 => n11066, ZN => n11241);
   U17285 : OAI22_X1 port map( A1 => n11069, A2 => n11241, B1 => n11068, B2 => 
                           n11240, ZN => n11070);
   U17286 : INV_X1 port map( A => n11290, ZN => n11071);
   U17287 : NAND2_X1 port map( A1 => n11071, A2 => n10665, ZN => n11080);
   U17288 : OAI21_X1 port map( B1 => n11075, B2 => n11072, A => n10665, ZN => 
                           n11074);
   U17289 : OAI21_X1 port map( B1 => n11291, B2 => n11287, A => n29116, ZN => 
                           n11073);
   U17290 : NAND2_X1 port map( A1 => n11074, A2 => n11073, ZN => n11079);
   U17291 : NAND3_X1 port map( A1 => n11077, A2 => n11076, A3 => n11075, ZN => 
                           n11078);
   U17292 : INV_X1 port map( A => n12270, ZN => n12576);
   U17293 : NAND2_X1 port map( A1 => n11213, A2 => n28624, ZN => n11081);
   U17294 : NOR2_X1 port map( A1 => n11084, A2 => n11083, ZN => n11088);
   U17295 : NOR2_X1 port map( A1 => n11086, A2 => n11085, ZN => n11087);
   U17296 : MUX2_X1 port map( A => n11088, B => n11087, S => n11210, Z => 
                           n11089);
   U17297 : NAND2_X1 port map( A1 => n11207, A2 => n10431, ZN => n11091);
   U17298 : AOI21_X1 port map( B1 => n11092, B2 => n11091, A => n11090, ZN => 
                           n11098);
   U17299 : NAND2_X1 port map( A1 => n29517, A2 => n11093, ZN => n11096);
   U17300 : OAI21_X1 port map( B1 => n5277, B2 => n11096, A => n11095, ZN => 
                           n11097);
   U17301 : NOR2_X1 port map( A1 => n12578, A2 => n12517, ZN => n12273);
   U17302 : OAI21_X1 port map( B1 => n11099, B2 => n333, A => n11225, ZN => 
                           n11100);
   U17303 : NAND2_X1 port map( A1 => n11100, A2 => n9709, ZN => n11102);
   U17304 : INV_X1 port map( A => n11898, ZN => n11101);
   U17305 : INV_X1 port map( A => n12516, ZN => n11940);
   U17306 : MUX2_X1 port map( A => n11103, B => n12273, S => n11940, Z => 
                           n11110);
   U17307 : NOR2_X1 port map( A1 => n11222, A2 => n435, ZN => n11107);
   U17308 : NAND2_X1 port map( A1 => n11104, A2 => n11220, ZN => n11105);
   U17309 : OAI21_X1 port map( B1 => n5974, B2 => n28202, A => n12578, ZN => 
                           n11108);
   U17310 : NOR2_X1 port map( A1 => n11121, A2 => n11120, ZN => n11130);
   U17311 : NAND3_X1 port map( A1 => n11124, A2 => n11123, A3 => n11122, ZN => 
                           n11129);
   U17312 : NAND3_X1 port map( A1 => n11127, A2 => n11126, A3 => n11125, ZN => 
                           n11128);
   U17313 : NAND2_X1 port map( A1 => n11774, A2 => n11131, ZN => n11134);
   U17314 : NAND3_X1 port map( A1 => n11133, A2 => n11132, A3 => n4555, ZN => 
                           n11775);
   U17315 : INV_X1 port map( A => n11551, ZN => n11422);
   U17316 : NAND2_X1 port map( A1 => n11422, A2 => n11782, ZN => n11151);
   U17317 : AOI22_X1 port map( A1 => n11137, A2 => n11136, B1 => n11135, B2 => 
                           n3862, ZN => n11143);
   U17319 : NAND2_X1 port map( A1 => n11421, A2 => n11553, ZN => n11150);
   U17320 : OAI21_X1 port map( B1 => n11146, B2 => n28627, A => n11144, ZN => 
                           n11147);
   U17321 : MUX2_X1 port map( A => n11151, B => n11150, S => n11785, Z => 
                           n11161);
   U17322 : NAND2_X1 port map( A1 => n28175, A2 => n11153, ZN => n11156);
   U17323 : INV_X1 port map( A => n11154, ZN => n11155);
   U17324 : XNOR2_X1 port map( A => n13249, B => n1905, ZN => n13532);
   U17325 : NAND2_X1 port map( A1 => n11166, A2 => n11168, ZN => n11167);
   U17326 : OAI211_X1 port map( C1 => n11169, C2 => n11168, A => n11167, B => 
                           n11330, ZN => n11172);
   U17327 : NAND3_X1 port map( A1 => n28208, A2 => n11331, A3 => n11170, ZN => 
                           n11171);
   U17331 : NAND3_X1 port map( A1 => n11349, A2 => n11192, A3 => n11350, ZN => 
                           n11193);
   U17332 : XNOR2_X1 port map( A => n13118, B => n3378, ZN => n11201);
   U17333 : XNOR2_X1 port map( A => n13532, B => n11201, ZN => n11202);
   U17334 : OAI211_X1 port map( C1 => n11211, C2 => n28624, A => n433, B => 
                           n11209, ZN => n11215);
   U17335 : OAI21_X1 port map( B1 => n11222, B2 => n11218, A => n11217, ZN => 
                           n11224);
   U17336 : OAI21_X1 port map( B1 => n11223, B2 => n11220, A => n11219, ZN => 
                           n11221);
   U17337 : OAI21_X1 port map( B1 => n333, B2 => n11225, A => n11231, ZN => 
                           n11229);
   U17338 : NAND2_X1 port map( A1 => n11232, A2 => n28270, ZN => n11228);
   U17342 : AND2_X1 port map( A1 => n12315, A2 => n12321, ZN => n11246);
   U17343 : NOR2_X1 port map( A1 => n11243, A2 => n11242, ZN => n11245);
   U17344 : NAND2_X1 port map( A1 => n11254, A2 => n11315, ZN => n11256);
   U17345 : MUX2_X1 port map( A => n11256, B => n11314, S => n11255, Z => 
                           n11257);
   U17346 : OAI21_X1 port map( B1 => n11259, B2 => n11258, A => n11257, ZN => 
                           n12081);
   U17347 : NOR2_X1 port map( A1 => n12080, A2 => n12081, ZN => n11297);
   U17348 : NAND2_X1 port map( A1 => n11264, A2 => n28204, ZN => n11265);
   U17349 : NAND3_X1 port map( A1 => n28174, A2 => n11267, A3 => n11266, ZN => 
                           n12290);
   U17350 : NAND2_X1 port map( A1 => n12289, A2 => n12081, ZN => n12062);
   U17351 : OAI21_X1 port map( B1 => n11271, B2 => n10523, A => n11270, ZN => 
                           n11279);
   U17352 : NAND2_X1 port map( A1 => n10523, A2 => n11272, ZN => n11277);
   U17353 : AOI21_X1 port map( B1 => n11277, B2 => n11276, A => n11275, ZN => 
                           n11278);
   U17354 : NOR2_X1 port map( A1 => n11288, A2 => n11287, ZN => n11289);
   U17355 : MUX2_X1 port map( A => n12062, B => n11295, S => n29324, Z => 
                           n11296);
   U17356 : XNOR2_X1 port map( A => n13539, B => n12841, ZN => n11307);
   U17357 : NAND2_X1 port map( A1 => n11782, A2 => n11785, ZN => n11301);
   U17358 : OR2_X1 port map( A1 => n11552, A2 => n11785, ZN => n11300);
   U17359 : INV_X1 port map( A => n11782, ZN => n11298);
   U17360 : OAI211_X1 port map( C1 => n11551, C2 => n29137, A => n11552, B => 
                           n11298, ZN => n11299);
   U17361 : OAI211_X1 port map( C1 => n11550, C2 => n11301, A => n11300, B => 
                           n11299, ZN => n12931);
   U17362 : NAND2_X1 port map( A1 => n11789, A2 => n28436, ZN => n11305);
   U17363 : NAND3_X1 port map( A1 => n10717, A2 => n2194, A3 => n2748, ZN => 
                           n11304);
   U17364 : NAND2_X1 port map( A1 => n10717, A2 => n11302, ZN => n11303);
   U17365 : XNOR2_X1 port map( A => n12931, B => n13075, ZN => n12136);
   U17366 : XNOR2_X1 port map( A => n11307, B => n12136, ZN => n11370);
   U17367 : NOR2_X1 port map( A1 => n11315, A2 => n11314, ZN => n11320);
   U17370 : NOR2_X1 port map( A1 => n11330, A2 => n11329, ZN => n11333);
   U17371 : INV_X1 port map( A => n12402, ZN => n11346);
   U17372 : NAND2_X1 port map( A1 => n11335, A2 => n11334, ZN => n11344);
   U17373 : NOR2_X1 port map( A1 => n11341, A2 => n11337, ZN => n11339);
   U17374 : AOI22_X1 port map( A1 => n11339, A2 => n11338, B1 => n11337, B2 => 
                           n11336, ZN => n11343);
   U17375 : OAI21_X1 port map( B1 => n11346, B2 => n12281, A => n12286, ZN => 
                           n11357);
   U17377 : NAND3_X1 port map( A1 => n11352, A2 => n11351, A3 => n11350, ZN => 
                           n11353);
   U17378 : OAI211_X2 port map( C1 => n11356, C2 => n11355, A => n11354, B => 
                           n11353, ZN => n12407);
   U17381 : OAI211_X1 port map( C1 => n11868, C2 => n11500, A => n11457, B => 
                           n578, ZN => n11361);
   U17382 : INV_X1 port map( A => n12303, ZN => n11769);
   U17385 : OAI21_X1 port map( B1 => n569, B2 => n12300, A => n12305, ZN => 
                           n11365);
   U17386 : INV_X1 port map( A => n11363, ZN => n11364);
   U17387 : AOI22_X2 port map( A1 => n11366, A2 => n11365, B1 => n11364, B2 => 
                           n12300, ZN => n13404);
   U17388 : XNOR2_X1 port map( A => n13404, B => n3164, ZN => n11367);
   U17389 : XNOR2_X1 port map( A => n11368, B => n11367, ZN => n11369);
   U17390 : NOR2_X1 port map( A1 => n12111, A2 => n12110, ZN => n11831);
   U17391 : OAI21_X1 port map( B1 => n12207, B2 => n12208, A => n28203, ZN => 
                           n11375);
   U17392 : NOR2_X1 port map( A1 => n12110, A2 => n9692, ZN => n11374);
   U17394 : INV_X1 port map( A => n12171, ZN => n11382);
   U17395 : INV_X1 port map( A => n11656, ZN => n12103);
   U17396 : NAND2_X1 port map( A1 => n12103, A2 => n12164, ZN => n11376);
   U17397 : INV_X1 port map( A => n12163, ZN => n11378);
   U17398 : XNOR2_X1 port map( A => n13297, B => n13401, ZN => n12490);
   U17399 : NOR2_X1 port map( A1 => n12151, A2 => n579, ZN => n11384);
   U17400 : NOR2_X1 port map( A1 => n11856, A2 => n12088, ZN => n11383);
   U17401 : NOR3_X1 port map( A1 => n11384, A2 => n12150, A3 => n11383, ZN => 
                           n11388);
   U17402 : AND2_X1 port map( A1 => n12151, A2 => n11856, ZN => n12152);
   U17403 : NAND2_X1 port map( A1 => n12152, A2 => n12990, ZN => n11386);
   U17404 : NAND2_X1 port map( A1 => n11927, A2 => n11851, ZN => n11394);
   U17405 : OAI21_X1 port map( B1 => n11853, B2 => n11855, A => n11852, ZN => 
                           n11392);
   U17407 : NAND3_X1 port map( A1 => n11944, A2 => n11858, A3 => n11945, ZN => 
                           n11397);
   U17408 : NAND2_X1 port map( A1 => n11952, A2 => n11947, ZN => n11395);
   U17409 : NAND2_X1 port map( A1 => n11397, A2 => n11396, ZN => n11400);
   U17410 : NAND2_X1 port map( A1 => n11857, A2 => n11948, ZN => n11398);
   U17411 : AOI21_X1 port map( B1 => n11665, B2 => n11398, A => n11862, ZN => 
                           n11399);
   U17412 : NOR2_X2 port map( A1 => n11400, A2 => n11399, ZN => n13208);
   U17413 : XNOR2_X1 port map( A => n13025, B => n13208, ZN => n12930);
   U17414 : NOR2_X1 port map( A1 => n11402, A2 => n11848, ZN => n11407);
   U17415 : INV_X1 port map( A => n11672, ZN => n11404);
   U17416 : NOR3_X1 port map( A1 => n11405, A2 => n11404, A3 => n11403, ZN => 
                           n11406);
   U17417 : XNOR2_X1 port map( A => n12747, B => n13405, ZN => n11409);
   U17418 : XNOR2_X1 port map( A => n12930, B => n11409, ZN => n11410);
   U17419 : INV_X1 port map( A => n12176, ZN => n12124);
   U17420 : INV_X1 port map( A => n11824, ZN => n12180);
   U17421 : AOI22_X1 port map( A1 => n11730, A2 => n12125, B1 => n12124, B2 => 
                           n12180, ZN => n11413);
   U17422 : MUX2_X1 port map( A => n11411, B => n12124, S => n11730, Z => 
                           n11412);
   U17423 : XNOR2_X1 port map( A => n12788, B => n12595, ZN => n11432);
   U17424 : INV_X1 port map( A => n11419, ZN => n11502);
   U17425 : AOI21_X1 port map( B1 => n11422, B2 => n11778, A => n11421, ZN => 
                           n11423);
   U17426 : INV_X1 port map( A => n11426, ZN => n11427);
   U17427 : NOR2_X1 port map( A1 => n11427, A2 => n11430, ZN => n11429);
   U17429 : NAND3_X1 port map( A1 => n12128, A2 => n12189, A3 => n11818, ZN => 
                           n11434);
   U17430 : INV_X1 port map( A => n12189, ZN => n11724);
   U17431 : OAI211_X2 port map( C1 => n11727, C2 => n11816, A => n11434, B => 
                           n11433, ZN => n13230);
   U17432 : AOI22_X1 port map( A1 => n12132, A2 => n11058, B1 => n12264, B2 => 
                           n12263, ZN => n11930);
   U17433 : NAND2_X1 port map( A1 => n575, A2 => n12263, ZN => n11436);
   U17434 : NAND2_X1 port map( A1 => n11436, A2 => n12264, ZN => n11437);
   U17435 : XNOR2_X1 port map( A => n13230, B => n13380, ZN => n11443);
   U17436 : NAND2_X1 port map( A1 => n12200, A2 => n12203, ZN => n11441);
   U17437 : OAI211_X1 port map( C1 => n12204, C2 => n11441, A => n11440, B => 
                           n11439, ZN => n12948);
   U17438 : XNOR2_X1 port map( A => n12948, B => n3334, ZN => n11442);
   U17439 : XNOR2_X1 port map( A => n11443, B => n11442, ZN => n11444);
   U17440 : XNOR2_X2 port map( A => n11445, B => n11444, ZN => n15194);
   U17441 : INV_X1 port map( A => n11740, ZN => n12357);
   U17442 : OAI21_X1 port map( B1 => n12363, B2 => n12362, A => n11446, ZN => 
                           n11447);
   U17443 : NAND3_X1 port map( A1 => n12327, A2 => n12018, A3 => n11449, ZN => 
                           n11452);
   U17444 : INV_X1 port map( A => n11747, ZN => n12329);
   U17445 : OAI211_X1 port map( C1 => n11888, C2 => n12328, A => n11450, B => 
                           n12332, ZN => n11451);
   U17447 : XNOR2_X1 port map( A => n13166, B => n13278, ZN => n11466);
   U17448 : NAND2_X1 port map( A1 => n11875, A2 => n11877, ZN => n11454);
   U17449 : AOI22_X1 port map( A1 => n130, A2 => n11454, B1 => n287, B2 => 
                           n11453, ZN => n11456);
   U17450 : NAND3_X1 port map( A1 => n11881, A2 => n11877, A3 => n11876, ZN => 
                           n11455);
   U17452 : NOR2_X1 port map( A1 => n4712, A2 => n11458, ZN => n11459);
   U17453 : OAI211_X1 port map( C1 => n1836, C2 => n11869, A => n11462, B => 
                           n11500, ZN => n11464);
   U17454 : XNOR2_X1 port map( A => n12894, B => n12817, ZN => n11465);
   U17455 : XNOR2_X1 port map( A => n11465, B => n11466, ZN => n11481);
   U17456 : INV_X1 port map( A => n12352, ZN => n11467);
   U17458 : NAND3_X1 port map( A1 => n29209, A2 => n12353, A3 => n29735, ZN => 
                           n11470);
   U17459 : NAND2_X1 port map( A1 => n12339, A2 => n12337, ZN => n11474);
   U17460 : XNOR2_X1 port map( A => n13018, B => n12514, ZN => n12681);
   U17461 : INV_X1 port map( A => n11755, ZN => n11996);
   U17462 : AND2_X1 port map( A1 => n11754, A2 => n12000, ZN => n11995);
   U17463 : NAND3_X1 port map( A1 => n11998, A2 => n11754, A3 => n11755, ZN => 
                           n11476);
   U17464 : OAI211_X1 port map( C1 => n11995, C2 => n11755, A => n11477, B => 
                           n11476, ZN => n11478);
   U17466 : XNOR2_X1 port map( A => n12763, B => n26531, ZN => n11479);
   U17467 : XNOR2_X1 port map( A => n12681, B => n11479, ZN => n11480);
   U17468 : INV_X1 port map( A => n12081, ZN => n12291);
   U17469 : NAND2_X1 port map( A1 => n29498, A2 => n11795, ZN => n12296);
   U17470 : NOR2_X1 port map( A1 => n12058, A2 => n29499, ZN => n11796);
   U17471 : INV_X1 port map( A => n12289, ZN => n11482);
   U17473 : NOR2_X1 port map( A1 => n12053, A2 => n12313, ZN => n12312);
   U17474 : INV_X1 port map( A => n12312, ZN => n11485);
   U17475 : NOR2_X1 port map( A1 => n12315, A2 => n12049, ZN => n11484);
   U17476 : INV_X1 port map( A => n12320, ZN => n12054);
   U17477 : NAND2_X1 port map( A1 => n12054, A2 => n12313, ZN => n11613);
   U17478 : OR2_X1 port map( A1 => n11613, A2 => n12049, ZN => n11483);
   U17480 : NAND3_X1 port map( A1 => n11793, A2 => n2194, A3 => n4046, ZN => 
                           n11488);
   U17481 : INV_X1 port map( A => n13263, ZN => n11498);
   U17482 : AND3_X1 port map( A1 => n11769, A2 => n12304, A3 => n11768, ZN => 
                           n11496);
   U17483 : NOR2_X2 port map( A1 => n11497, A2 => n11496, ZN => n13104);
   U17484 : XNOR2_X1 port map( A => n11498, B => n13104, ZN => n12912);
   U17485 : INV_X1 port map( A => n12912, ZN => n11499);
   U17486 : XNOR2_X1 port map( A => n11499, B => n12966, ZN => n11511);
   U17487 : OAI211_X1 port map( C1 => n3900, C2 => n11502, A => n11551, B => 
                           n11553, ZN => n11503);
   U17488 : INV_X1 port map( A => n12722, ZN => n11937);
   U17489 : XNOR2_X1 port map( A => n11937, B => n12965, ZN => n11509);
   U17490 : OR2_X1 port map( A1 => n12402, A2 => n12407, ZN => n11507);
   U17491 : NAND2_X1 port map( A1 => n11801, A2 => n12400, ZN => n12283);
   U17492 : NAND3_X1 port map( A1 => n12280, A2 => n12402, A3 => n12281, ZN => 
                           n11506);
   U17493 : XNOR2_X1 port map( A => n13150, B => n3223, ZN => n11508);
   U17494 : XNOR2_X1 port map( A => n11509, B => n11508, ZN => n11510);
   U17495 : INV_X1 port map( A => n14241, ZN => n14243);
   U17496 : NAND3_X1 port map( A1 => n11970, A2 => n12159, A3 => n12037, ZN => 
                           n11513);
   U17497 : INV_X1 port map( A => n11673, ZN => n11639);
   U17499 : NAND3_X1 port map( A1 => n11848, A2 => n29139, A3 => n11640, ZN => 
                           n11516);
   U17500 : XNOR2_X1 port map( A => n12780, B => n13137, ZN => n13375);
   U17501 : NOR2_X1 port map( A1 => n3653, A2 => n12508, ZN => n11836);
   U17502 : NAND3_X1 port map( A1 => n12512, A2 => n6374, A3 => n10863, ZN => 
                           n11520);
   U17503 : INV_X1 port map( A => n13081, ZN => n13084);
   U17504 : INV_X1 port map( A => n303, ZN => n11522);
   U17505 : NAND3_X1 port map( A1 => n13083, A2 => n13084, A3 => n11522, ZN => 
                           n11531);
   U17506 : AND2_X1 port map( A1 => n11524, A2 => n11523, ZN => n11527);
   U17507 : NAND4_X1 port map( A1 => n11528, A2 => n11527, A3 => n11526, A4 => 
                           n11525, ZN => n11529);
   U17508 : XNOR2_X1 port map( A => n13270, B => n13533, ZN => n12905);
   U17509 : XNOR2_X1 port map( A => n13375, B => n12905, ZN => n11546);
   U17510 : INV_X1 port map( A => n12220, ZN => n11963);
   U17511 : INV_X1 port map( A => n12219, ZN => n11965);
   U17512 : NAND2_X1 port map( A1 => n12043, A2 => n11965, ZN => n11534);
   U17513 : NAND2_X1 port map( A1 => n12044, A2 => n11963, ZN => n11533);
   U17514 : NAND3_X1 port map( A1 => n12220, A2 => n12219, A3 => n12218, ZN => 
                           n11532);
   U17515 : NAND4_X2 port map( A1 => n11535, A2 => n11533, A3 => n11534, A4 => 
                           n11532, ZN => n13420);
   U17516 : OAI21_X1 port map( B1 => n11754, B2 => n11536, A => n12000, ZN => 
                           n11537);
   U17517 : INV_X1 port map( A => n11998, ZN => n12001);
   U17518 : NAND3_X1 port map( A1 => n12001, A2 => n11754, A3 => n11996, ZN => 
                           n11539);
   U17519 : XNOR2_X1 port map( A => n12830, B => n13420, ZN => n11544);
   U17520 : NAND3_X1 port map( A1 => n1986, A2 => n12236, A3 => n375, ZN => 
                           n11542);
   U17521 : XNOR2_X1 port map( A => n11544, B => n11543, ZN => n11545);
   U17522 : INV_X1 port map( A => n14171, ZN => n14239);
   U17524 : INV_X1 port map( A => n11861, ZN => n11558);
   U17525 : NOR2_X1 port map( A1 => n11952, A2 => n11947, ZN => n11555);
   U17526 : AOI22_X1 port map( A1 => n11951, A2 => n11555, B1 => n11944, B2 => 
                           n11858, ZN => n11557);
   U17527 : INV_X1 port map( A => n11947, ZN => n11556);
   U17528 : AOI21_X1 port map( B1 => n349, B2 => n12249, A => n12070, ZN => 
                           n11559);
   U17529 : NAND2_X1 port map( A1 => n11559, A2 => n11934, ZN => n11562);
   U17530 : NAND2_X1 port map( A1 => n11594, A2 => n12070, ZN => n11561);
   U17531 : INV_X1 port map( A => n12253, ZN => n11932);
   U17532 : NOR2_X1 port map( A1 => n349, A2 => n11932, ZN => n11560);
   U17533 : XNOR2_X1 port map( A => n13364, B => n13190, ZN => n12920);
   U17534 : XNOR2_X1 port map( A => n11563, B => n12920, ZN => n11578);
   U17535 : NOR2_X1 port map( A1 => n12271, A2 => n12270, ZN => n12583);
   U17536 : INV_X1 port map( A => n12583, ZN => n11565);
   U17537 : INV_X1 port map( A => n28202, ZN => n11564);
   U17538 : NAND3_X1 port map( A1 => n12271, A2 => n12517, A3 => n11564, ZN => 
                           n12519);
   U17539 : AND2_X1 port map( A1 => n11565, A2 => n12519, ZN => n11566);
   U17540 : INV_X1 port map( A => n11622, ZN => n11953);
   U17541 : OAI21_X1 port map( B1 => n571, B2 => n11953, A => n6706, ZN => 
                           n11569);
   U17543 : AOI21_X1 port map( B1 => n11574, B2 => n12266, A => n12267, ZN => 
                           n11571);
   U17544 : OAI21_X1 port map( B1 => n12265, B2 => n12266, A => n11571, ZN => 
                           n11573);
   U17545 : NAND3_X1 port map( A1 => n11574, A2 => n568, A3 => n12263, ZN => 
                           n11572);
   U17546 : INV_X1 port map( A => n2402, ZN => n27678);
   U17547 : XNOR2_X1 port map( A => n13291, B => n27678, ZN => n11575);
   U17548 : XNOR2_X1 port map( A => n11578, B => n11577, ZN => n14238);
   U17549 : NAND3_X1 port map( A1 => n28172, A2 => n14239, A3 => n563, ZN => 
                           n11579);
   U17550 : NAND2_X1 port map( A1 => n14893, A2 => n15415, ZN => n15412);
   U17551 : INV_X1 port map( A => n15412, ZN => n12012);
   U17552 : XNOR2_X1 port map( A => n12881, B => n12841, ZN => n13540);
   U17553 : NOR2_X1 port map( A1 => n11881, A2 => n11877, ZN => n11589);
   U17554 : OAI21_X1 port map( B1 => n11878, B2 => n11582, A => n11876, ZN => 
                           n11588);
   U17555 : NOR2_X1 port map( A1 => n11877, A2 => n11583, ZN => n11584);
   U17556 : NOR2_X1 port map( A1 => n10453, A2 => n11876, ZN => n11585);
   U17557 : NAND2_X1 port map( A1 => n287, A2 => n11585, ZN => n11586);
   U17559 : XNOR2_X1 port map( A => n13540, B => n12349, ZN => n11606);
   U17560 : NAND2_X1 port map( A1 => n12583, A2 => n11940, ZN => n12581);
   U17561 : NAND2_X1 port map( A1 => n28202, A2 => n12270, ZN => n11590);
   U17562 : NAND2_X1 port map( A1 => n12575, A2 => n11590, ZN => n11591);
   U17563 : INV_X1 port map( A => n12251, ZN => n12256);
   U17564 : NOR2_X1 port map( A1 => n12253, A2 => n12249, ZN => n11593);
   U17565 : AOI21_X1 port map( B1 => n349, B2 => n12253, A => n11593, ZN => 
                           n11598);
   U17566 : NAND2_X1 port map( A1 => n11595, A2 => n12256, ZN => n11596);
   U17567 : XNOR2_X1 port map( A => n13504, B => n13458, ZN => n12933);
   U17568 : NAND2_X1 port map( A1 => n12204, A2 => n4844, ZN => n11600);
   U17569 : AOI21_X1 port map( B1 => n11601, B2 => n11600, A => n11702, ZN => 
                           n11603);
   U17570 : NOR2_X1 port map( A1 => n12205, A2 => n11807, ZN => n11602);
   U17571 : XNOR2_X1 port map( A => n12933, B => n11604, ZN => n11605);
   U17572 : XNOR2_X1 port map( A => n11606, B => n11605, ZN => n14157);
   U17573 : INV_X1 port map( A => n14157, ZN => n13935);
   U17574 : NOR2_X1 port map( A1 => n12303, A2 => n12302, ZN => n11607);
   U17575 : NOR2_X1 port map( A1 => n12305, A2 => n11607, ZN => n11611);
   U17576 : INV_X1 port map( A => n11608, ZN => n11609);
   U17577 : INV_X1 port map( A => n12548, ZN => n13473);
   U17578 : NAND2_X1 port map( A1 => n285, A2 => n12313, ZN => n11614);
   U17579 : AOI21_X1 port map( B1 => n11614, B2 => n12054, A => n12316, ZN => 
                           n11615);
   U17580 : XNOR2_X1 port map( A => n13473, B => n13450, ZN => n12899);
   U17581 : OAI21_X1 port map( B1 => n11617, B2 => n11616, A => n3653, ZN => 
                           n11620);
   U17582 : NOR2_X1 port map( A1 => n12512, A2 => n12508, ZN => n11618);
   U17583 : XNOR2_X1 port map( A => n13563, B => n13055, ZN => n11621);
   U17584 : XNOR2_X1 port map( A => n12899, B => n11621, ZN => n11631);
   U17585 : INV_X1 port map( A => n11800, ZN => n11623);
   U17586 : NAND2_X1 port map( A1 => n11623, A2 => n12286, ZN => n11624);
   U17587 : XNOR2_X1 port map( A => n13567, B => n3372, ZN => n11628);
   U17588 : XNOR2_X1 port map( A => n11629, B => n11628, ZN => n11630);
   U17589 : XNOR2_X2 port map( A => n11631, B => n11630, ZN => n14480);
   U17590 : INV_X1 port map( A => n11632, ZN => n11638);
   U17591 : INV_X1 port map( A => n11633, ZN => n11635);
   U17592 : NAND2_X1 port map( A1 => n11635, A2 => n11634, ZN => n11637);
   U17593 : NOR3_X1 port map( A1 => n11638, A2 => n11637, A3 => n11636, ZN => 
                           n11675);
   U17594 : MUX2_X1 port map( A => n11675, B => n11640, S => n11671, Z => 
                           n11644);
   U17595 : NOR2_X1 port map( A1 => n11640, A2 => n11672, ZN => n11849);
   U17596 : NOR2_X1 port map( A1 => n11849, A2 => n29139, ZN => n11643);
   U17597 : NAND3_X1 port map( A1 => n11641, A2 => n11640, A3 => n11639, ZN => 
                           n11642);
   U17599 : XNOR2_X1 port map( A => n29140, B => n13219, ZN => n11652);
   U17600 : XNOR2_X1 port map( A => n12867, B => n13523, ZN => n13168);
   U17601 : XNOR2_X1 port map( A => n11652, B => n13168, ZN => n11670);
   U17602 : NOR2_X1 port map( A1 => n12150, A2 => n12100, ZN => n11653);
   U17603 : NAND2_X1 port map( A1 => n1931, A2 => n12164, ZN => n11654);
   U17605 : AOI21_X1 port map( B1 => n11655, B2 => n11654, A => n28828, ZN => 
                           n11664);
   U17607 : INV_X1 port map( A => n11660, ZN => n11661);
   U17608 : MUX2_X1 port map( A => n11844, B => n11662, S => n12102, Z => 
                           n11663);
   U17609 : MUX2_X1 port map( A => n11951, B => n11948, S => n11945, Z => 
                           n11666);
   U17610 : XNOR2_X1 port map( A => n13048, B => n2274, ZN => n11669);
   U17612 : NOR2_X1 port map( A1 => n11676, A2 => n11675, ZN => n11679);
   U17613 : INV_X1 port map( A => n11680, ZN => n11683);
   U17614 : OAI21_X2 port map( B1 => n11682, B2 => n11683, A => n11681, ZN => 
                           n13245);
   U17615 : XNOR2_X1 port map( A => n13553, B => n13245, ZN => n12911);
   U17616 : XNOR2_X1 port map( A => n11684, B => n12911, ZN => n11701);
   U17617 : NOR2_X1 port map( A1 => n12000, A2 => n6661, ZN => n11757);
   U17619 : AND2_X1 port map( A1 => n13081, A2 => n12231, ZN => n11811);
   U17620 : INV_X1 port map( A => n11811, ZN => n11689);
   U17621 : AND2_X1 port map( A1 => n11980, A2 => n12226, ZN => n12228);
   U17622 : OAI211_X1 port map( C1 => n13081, C2 => n13086, A => n13083, B => 
                           n11809, ZN => n11690);
   U17623 : INV_X1 port map( A => n13043, ZN => n11692);
   U17624 : XNOR2_X1 port map( A => n12686, B => n11692, ZN => n11699);
   U17625 : OAI211_X1 port map( C1 => n12219, C2 => n12218, A => n12224, B => 
                           n12042, ZN => n11696);
   U17626 : NAND4_X1 port map( A1 => n2846, A2 => n12221, A3 => n11694, A4 => 
                           n11693, ZN => n11695);
   U17627 : XNOR2_X1 port map( A => n13484, B => n3422, ZN => n11698);
   U17628 : XNOR2_X1 port map( A => n11699, B => n11698, ZN => n11700);
   U17629 : XNOR2_X1 port map( A => n11701, B => n11700, ZN => n13755);
   U17630 : INV_X1 port map( A => n13755, ZN => n13934);
   U17631 : NOR2_X1 port map( A1 => n12202, A2 => n12201, ZN => n11706);
   U17632 : NAND2_X1 port map( A1 => n12204, A2 => n11706, ZN => n11707);
   U17633 : XNOR2_X1 port map( A => n12495, B => n12827, ZN => n13535);
   U17634 : INV_X1 port map( A => n13535, ZN => n11717);
   U17635 : OAI211_X1 port map( C1 => n11712, C2 => n11711, A => n11710, B => 
                           n11709, ZN => n11713);
   U17636 : XNOR2_X1 port map( A => n1857, B => n3369, ZN => n11716);
   U17637 : XNOR2_X1 port map( A => n11717, B => n11716, ZN => n11735);
   U17638 : INV_X1 port map( A => n11718, ZN => n11720);
   U17639 : NOR2_X1 port map( A1 => n11787, A2 => n2748, ZN => n11719);
   U17640 : XNOR2_X1 port map( A => n13249, B => n13067, ZN => n12298);
   U17641 : NAND3_X1 port map( A1 => n11819, A2 => n12198, A3 => n12186, ZN => 
                           n11722);
   U17642 : NOR2_X1 port map( A1 => n12186, A2 => n11724, ZN => n11725);
   U17643 : NAND2_X1 port map( A1 => n2483, A2 => n11725, ZN => n11726);
   U17644 : OAI211_X1 port map( C1 => n11727, C2 => n2483, A => n6917, B => 
                           n11726, ZN => n12554);
   U17645 : INV_X1 port map( A => n12554, ZN => n12826);
   U17646 : INV_X1 port map( A => n11730, ZN => n12179);
   U17647 : NOR2_X1 port map( A1 => n12179, A2 => n11824, ZN => n11729);
   U17648 : NOR2_X1 port map( A1 => n12125, A2 => n12124, ZN => n11728);
   U17649 : MUX2_X1 port map( A => n11729, B => n11728, S => n570, Z => n11733)
                           ;
   U17650 : NAND2_X1 port map( A1 => n1890, A2 => n12177, ZN => n12183);
   U17651 : NOR2_X1 port map( A1 => n13206, A2 => n11731, ZN => n11732);
   U17652 : NOR2_X2 port map( A1 => n11733, A2 => n11732, ZN => n13418);
   U17653 : XNOR2_X1 port map( A => n13418, B => n12826, ZN => n12904);
   U17654 : NAND2_X1 port map( A1 => n13934, A2 => n14158, ZN => n14163);
   U17655 : OAI21_X1 port map( B1 => n29735, B2 => n12022, A => n12354, ZN => 
                           n11738);
   U17656 : MUX2_X1 port map( A => n580, B => n12350, S => n12352, Z => n11737)
                           ;
   U17657 : NOR2_X1 port map( A1 => n12353, A2 => n12352, ZN => n11736);
   U17658 : INV_X1 port map( A => n13511, ZN => n11746);
   U17659 : INV_X1 port map( A => n12363, ZN => n12358);
   U17660 : NAND3_X1 port map( A1 => n12358, A2 => n11741, A3 => n12359, ZN => 
                           n11745);
   U17661 : NAND3_X1 port map( A1 => n11741, A2 => n11908, A3 => n12356, ZN => 
                           n11744);
   U17662 : NAND3_X1 port map( A1 => n12362, A2 => n11742, A3 => n12359, ZN => 
                           n11743);
   U17663 : XNOR2_X1 port map( A => n11746, B => n13039, ZN => n12809);
   U17665 : NAND2_X1 port map( A1 => n11449, A2 => n11747, ZN => n12330);
   U17666 : XNOR2_X1 port map( A => n13432, B => n13547, ZN => n11749);
   U17667 : XNOR2_X1 port map( A => n12809, B => n11749, ZN => n11764);
   U17668 : NOR2_X1 port map( A1 => n11751, A2 => n390, ZN => n11753);
   U17669 : NAND2_X1 port map( A1 => n4712, A2 => n11868, ZN => n11752);
   U17670 : XNOR2_X1 port map( A => n12560, B => n12699, ZN => n11762);
   U17672 : NAND2_X1 port map( A1 => n11998, A2 => n1831, ZN => n11758);
   U17673 : XNOR2_X1 port map( A => n13191, B => n2446, ZN => n11761);
   U17674 : XNOR2_X1 port map( A => n11762, B => n11761, ZN => n11763);
   U17675 : XNOR2_X1 port map( A => n11764, B => n11763, ZN => n13936);
   U17676 : INV_X1 port map( A => n13936, ZN => n13754);
   U17677 : NAND2_X1 port map( A1 => n14163, A2 => n13754, ZN => n11765);
   U17678 : NAND2_X1 port map( A1 => n14473, A2 => n13935, ZN => n11766);
   U17679 : INV_X1 port map( A => n11770, ZN => n11773);
   U17680 : OAI211_X2 port map( C1 => n11773, C2 => n285, A => n11772, B => 
                           n11771, ZN => n13170);
   U17681 : XNOR2_X1 port map( A => n13170, B => n13014, ZN => n13277);
   U17682 : INV_X1 port map( A => n11774, ZN => n11777);
   U17683 : INV_X1 port map( A => n11131, ZN => n11776);
   U17684 : OAI21_X1 port map( B1 => n11777, B2 => n11776, A => n11775, ZN => 
                           n11779);
   U17685 : MUX2_X1 port map( A => n11780, B => n11779, S => n11778, Z => 
                           n11781);
   U17686 : INV_X1 port map( A => n11781, ZN => n11786);
   U17687 : INV_X1 port map( A => n12542, ZN => n12866);
   U17688 : NAND2_X1 port map( A1 => n11789, A2 => n2194, ZN => n11790);
   U17690 : XNOR2_X1 port map( A => n13020, B => n12866, ZN => n12634);
   U17691 : XNOR2_X1 port map( A => n12634, B => n13277, ZN => n11805);
   U17692 : NAND3_X1 port map( A1 => n12289, A2 => n12080, A3 => n29499, ZN => 
                           n11798);
   U17693 : NAND2_X1 port map( A1 => n11796, A2 => n11795, ZN => n11797);
   U17694 : XNOR2_X1 port map( A => n12734, B => n12817, ZN => n11803);
   U17695 : INV_X1 port map( A => n12407, ZN => n12278);
   U17696 : INV_X1 port map( A => n3087, ZN => n27560);
   U17697 : XNOR2_X1 port map( A => n12760, B => n27560, ZN => n11802);
   U17698 : XNOR2_X1 port map( A => n11803, B => n11802, ZN => n11804);
   U17699 : NAND3_X1 port map( A1 => n12201, A2 => n12202, A3 => n12200, ZN => 
                           n11806);
   U17700 : NAND3_X1 port map( A1 => n8847, A2 => n11807, A3 => n12201, ZN => 
                           n11808);
   U17701 : XNOR2_X1 port map( A => n12776, B => n29247, ZN => n11815);
   U17702 : OAI21_X1 port map( B1 => n11812, B2 => n303, A => n11982, ZN => 
                           n11813);
   U17703 : XNOR2_X1 port map( A => n11815, B => n12985, ZN => n11829);
   U17704 : INV_X1 port map( A => n12128, ZN => n11820);
   U17705 : NOR2_X1 port map( A1 => n11819, A2 => n12186, ZN => n11817);
   U17706 : NAND2_X1 port map( A1 => n12128, A2 => n11817, ZN => n11822);
   U17707 : NAND3_X1 port map( A1 => n11820, A2 => n11819, A3 => n12189, ZN => 
                           n11821);
   U17708 : NAND4_X1 port map( A1 => n11823, A2 => n11822, A3 => n12127, A4 => 
                           n11821, ZN => n13436);
   U17709 : AOI21_X1 port map( B1 => n12179, B2 => n11824, A => n570, ZN => 
                           n11828);
   U17710 : NAND2_X1 port map( A1 => n12125, A2 => n12176, ZN => n11825);
   U17711 : AND2_X1 port map( A1 => n12183, A2 => n11825, ZN => n11827);
   U17712 : NAND2_X1 port map( A1 => n1890, A2 => n12180, ZN => n11826);
   U17713 : XNOR2_X1 port map( A => n13360, B => n13436, ZN => n13290);
   U17714 : XNOR2_X1 port map( A => n11829, B => n13290, ZN => n11839);
   U17717 : OAI21_X2 port map( B1 => n11833, B2 => n12109, A => n11832, ZN => 
                           n13035);
   U17718 : INV_X1 port map( A => n12512, ZN => n12510);
   U17719 : OAI21_X1 port map( B1 => n12512, B2 => n10863, A => n6374, ZN => 
                           n11834);
   U17720 : XNOR2_X1 port map( A => n11839, B => n11838, ZN => n13778);
   U17721 : INV_X1 port map( A => n13778, ZN => n14249);
   U17722 : NAND3_X1 port map( A1 => n12210, A2 => n12206, A3 => n12211, ZN => 
                           n11841);
   U17723 : OAI21_X1 port map( B1 => n11849, B2 => n11848, A => n5079, ZN => 
                           n11850);
   U17724 : AOI21_X1 port map( B1 => n11858, B2 => n11943, A => n11857, ZN => 
                           n11863);
   U17725 : XNOR2_X1 port map( A => n13566, B => n13175, ZN => n12792);
   U17726 : XNOR2_X1 port map( A => n12595, B => n3537, ZN => n11864);
   U17727 : XNOR2_X1 port map( A => n12792, B => n11864, ZN => n11865);
   U17728 : MUX2_X1 port map( A => n13744, B => n14249, S => n29312, Z => 
                           n12010);
   U17729 : OAI21_X1 port map( B1 => n578, B2 => n11869, A => n390, ZN => 
                           n11871);
   U17730 : OAI211_X1 port map( C1 => n390, C2 => n4712, A => n11871, B => 
                           n11870, ZN => n11873);
   U17731 : OAI21_X1 port map( B1 => n11875, B2 => n11877, A => n567, ZN => 
                           n11882);
   U17732 : NOR2_X1 port map( A1 => n11877, A2 => n11876, ZN => n11880);
   U17733 : XNOR2_X1 port map( A => n12849, B => n13478, ZN => n12638);
   U17734 : OAI21_X1 port map( B1 => n11884, B2 => n12332, A => n12327, ZN => 
                           n11891);
   U17735 : NAND3_X1 port map( A1 => n11888, A2 => n12018, A3 => n12329, ZN => 
                           n11889);
   U17736 : OAI211_X2 port map( C1 => n12014, C2 => n11891, A => n11890, B => 
                           n11889, ZN => n13136);
   U17737 : XNOR2_X1 port map( A => n12830, B => n13136, ZN => n11892);
   U17738 : XNOR2_X1 port map( A => n12638, B => n11892, ZN => n11920);
   U17740 : INV_X1 port map( A => n11893, ZN => n11895);
   U17741 : NAND2_X1 port map( A1 => n11895, A2 => n11894, ZN => n11897);
   U17742 : NAND2_X1 port map( A1 => n11900, A2 => n11899, ZN => n11903);
   U17743 : NOR2_X1 port map( A1 => n11903, A2 => n11901, ZN => n12427);
   U17744 : INV_X1 port map( A => n12427, ZN => n11902);
   U17745 : INV_X1 port map( A => n11903, ZN => n11904);
   U17746 : NAND3_X1 port map( A1 => n11904, A2 => n29209, A3 => n12350, ZN => 
                           n12430);
   U17748 : NAND2_X1 port map( A1 => n12362, A2 => n12359, ZN => n11911);
   U17749 : NAND3_X1 port map( A1 => n12361, A2 => n11908, A3 => n12357, ZN => 
                           n11909);
   U17752 : INV_X1 port map( A => n431, ZN => n12340);
   U17753 : NAND2_X1 port map( A1 => n11915, A2 => n12338, ZN => n11914);
   U17754 : INV_X1 port map( A => n12339, ZN => n12344);
   U17755 : NAND3_X1 port map( A1 => n12344, A2 => n12343, A3 => n11915, ZN => 
                           n11916);
   U17756 : XNOR2_X1 port map( A => n13482, B => n2982, ZN => n11918);
   U17757 : XNOR2_X1 port map( A => n13274, B => n11918, ZN => n11919);
   U17758 : XNOR2_X1 port map( A => n11919, B => n11920, ZN => n13775);
   U17759 : AOI21_X1 port map( B1 => n11922, B2 => n11927, A => n11921, ZN => 
                           n11926);
   U17760 : NOR2_X1 port map( A1 => n11924, A2 => n10905, ZN => n11925);
   U17761 : NOR2_X1 port map( A1 => n12132, A2 => n12267, ZN => n11929);
   U17762 : OAI21_X1 port map( B1 => n11930, B2 => n11929, A => n11928, ZN => 
                           n11931);
   U17763 : INV_X1 port map( A => n12249, ZN => n12072);
   U17764 : OAI22_X1 port map( A1 => n12251, A2 => n11933, B1 => n11932, B2 => 
                           n12072, ZN => n12071);
   U17765 : NAND2_X1 port map( A1 => n12071, A2 => n11934, ZN => n11936);
   U17766 : OAI211_X1 port map( C1 => n12070, C2 => n12252, A => n349, B => 
                           n12072, ZN => n11935);
   U17767 : XNOR2_X1 port map( A => n13265, B => n11937, ZN => n11938);
   U17768 : XNOR2_X1 port map( A => n11939, B => n11938, ZN => n11961);
   U17769 : XNOR2_X1 port map( A => n13008, B => n13262, ZN => n11959);
   U17770 : NAND3_X1 port map( A1 => n571, A2 => n6706, A3 => n11953, ZN => 
                           n11957);
   U17771 : XNOR2_X1 port map( A => n13488, B => n3180, ZN => n11958);
   U17772 : XNOR2_X1 port map( A => n11958, B => n11959, ZN => n11960);
   U17773 : XNOR2_X1 port map( A => n11961, B => n11960, ZN => n14078);
   U17774 : NAND2_X1 port map( A1 => n12224, A2 => n11962, ZN => n11968);
   U17775 : AOI21_X1 port map( B1 => n11963, B2 => n12042, A => n11962, ZN => 
                           n11964);
   U17777 : NAND3_X1 port map( A1 => n11963, A2 => n11965, A3 => n12218, ZN => 
                           n11966);
   U17778 : XNOR2_X1 port map( A => n13209, B => n3625, ZN => n11975);
   U17779 : NAND3_X1 port map( A1 => n5839, A2 => n12035, A3 => n12037, ZN => 
                           n11974);
   U17780 : INV_X1 port map( A => n11969, ZN => n11970);
   U17781 : NAND3_X1 port map( A1 => n11970, A2 => n12157, A3 => n12241, ZN => 
                           n11972);
   U17782 : NAND3_X1 port map( A1 => n11969, A2 => n12159, A3 => n12241, ZN => 
                           n11971);
   U17783 : NOR2_X1 port map( A1 => n776, A2 => n12234, ZN => n11976);
   U17784 : NOR2_X1 port map( A1 => n11976, A2 => n5009, ZN => n11978);
   U17785 : NAND3_X1 port map( A1 => n13081, A2 => n11982, A3 => n303, ZN => 
                           n11986);
   U17786 : NAND4_X1 port map( A1 => n11984, A2 => n13086, A3 => n13084, A4 => 
                           n11983, ZN => n11985);
   U17787 : XNOR2_X1 port map( A => n13133, B => n13543, ZN => n12492);
   U17788 : XNOR2_X1 port map( A => n11988, B => n12492, ZN => n12007);
   U17789 : INV_X1 port map( A => n12747, ZN => n12005);
   U17791 : NAND2_X1 port map( A1 => n11990, A2 => n11989, ZN => n11991);
   U17792 : NAND2_X1 port map( A1 => n12000, A2 => n11996, ZN => n12003);
   U17793 : INV_X1 port map( A => n11995, ZN => n11999);
   U17794 : NAND2_X1 port map( A1 => n11996, A2 => n1831, ZN => n11997);
   U17795 : NAND3_X1 port map( A1 => n6658, A2 => n572, A3 => n12001, ZN => 
                           n12002);
   U17796 : XNOR2_X1 port map( A => n13028, B => n12879, ZN => n12648);
   U17797 : XNOR2_X1 port map( A => n12005, B => n12648, ZN => n12006);
   U17798 : XNOR2_X1 port map( A => n12007, B => n12006, ZN => n13776);
   U17799 : NAND2_X1 port map( A1 => n13776, A2 => n14252, ZN => n13745);
   U17800 : INV_X1 port map( A => n13745, ZN => n12008);
   U17801 : NAND2_X1 port map( A1 => n12008, A2 => n14254, ZN => n12009);
   U17803 : AOI22_X1 port map( A1 => n12012, A2 => n15406, B1 => n12011, B2 => 
                           n3362, ZN => n12372);
   U17804 : AND2_X1 port map( A1 => n12013, A2 => n12018, ZN => n12021);
   U17805 : INV_X1 port map( A => n12014, ZN => n12020);
   U17806 : OAI21_X1 port map( B1 => n12021, B2 => n12020, A => n12019, ZN => 
                           n12388);
   U17807 : XNOR2_X1 port map( A => n12684, B => n3787, ZN => n12025);
   U17808 : OAI211_X1 port map( C1 => n12022, C2 => n12354, A => n11467, B => 
                           n580, ZN => n12023);
   U17809 : OAI211_X1 port map( C1 => n29735, C2 => n29209, A => n12024, B => 
                           n12023, ZN => n13348);
   U17810 : XNOR2_X1 port map( A => n13246, B => n12025, ZN => n12033);
   U17811 : XNOR2_X1 port map( A => n13195, B => n12965, ZN => n12797);
   U17812 : NOR2_X1 port map( A1 => n12026, A2 => n12337, ZN => n12031);
   U17813 : OAI21_X1 port map( B1 => n12028, B2 => n12337, A => n12027, ZN => 
                           n12029);
   U17814 : XNOR2_X1 port map( A => n12913, B => n12686, ZN => n13425);
   U17815 : XNOR2_X1 port map( A => n13425, B => n12797, ZN => n12032);
   U17816 : XNOR2_X1 port map( A => n12033, B => n12032, ZN => n14481);
   U17817 : XNOR2_X1 port map( A => n12954, B => n2381, ZN => n12034);
   U17818 : XNOR2_X1 port map( A => n12396, B => n13012, ZN => n13441);
   U17819 : MUX2_X1 port map( A => n12042, B => n12041, S => n12220, Z => 
                           n12046);
   U17820 : XNOR2_X1 port map( A => n13525, B => n13171, ZN => n13015);
   U17821 : XNOR2_X1 port map( A => n13051, B => n13015, ZN => n12047);
   U17822 : NOR2_X1 port map( A1 => n12053, A2 => n12051, ZN => n12052);
   U17823 : OAI21_X1 port map( B1 => n6920, B2 => n12052, A => n566, ZN => 
                           n12056);
   U17824 : NAND2_X1 port map( A1 => n12054, A2 => n285, ZN => n12055);
   U17825 : OAI211_X1 port map( C1 => n566, C2 => n12057, A => n12056, B => 
                           n12055, ZN => n13341);
   U17826 : INV_X1 port map( A => n12058, ZN => n12297);
   U17827 : NAND2_X1 port map( A1 => n12288, A2 => n12297, ZN => n12063);
   U17828 : XNOR2_X1 port map( A => n13341, B => n12697, ZN => n12410);
   U17829 : NAND2_X1 port map( A1 => n12279, A2 => n12401, ZN => n12068);
   U17830 : NAND3_X1 port map( A1 => n12408, A2 => n12278, A3 => n12402, ZN => 
                           n12066);
   U17831 : NAND4_X1 port map( A1 => n12068, A2 => n12067, A3 => n12404, A4 => 
                           n12066, ZN => n12069);
   U17832 : NAND2_X1 port map( A1 => n29306, A2 => n12120, ZN => n13766);
   U17833 : OAI21_X1 port map( B1 => n349, B2 => n12072, A => n12253, ZN => 
                           n12073);
   U17834 : NAND2_X1 port map( A1 => n12073, A2 => n12251, ZN => n12074);
   U17835 : OAI21_X1 port map( B1 => n12271, B2 => n28202, A => n12576, ZN => 
                           n12076);
   U17836 : XNOR2_X1 port map( A => n12677, B => n3565, ZN => n12078);
   U17837 : XNOR2_X1 port map( A => n13229, B => n12078, ZN => n12086);
   U17838 : XNOR2_X1 port map( A => n12948, B => n565, ZN => n12789);
   U17839 : NOR2_X1 port map( A1 => n12080, A2 => n3558, ZN => n12083);
   U17842 : XNOR2_X1 port map( A => n13451, B => n13447, ZN => n13283);
   U17843 : XNOR2_X1 port map( A => n13283, B => n12789, ZN => n12085);
   U17845 : NAND2_X1 port map( A1 => n12990, A2 => n12088, ZN => n12089);
   U17847 : INV_X1 port map( A => n12091, ZN => n12095);
   U17848 : INV_X1 port map( A => n12092, ZN => n12093);
   U17849 : NAND3_X1 port map( A1 => n12095, A2 => n12094, A3 => n12093, ZN => 
                           n12096);
   U17850 : NOR2_X1 port map( A1 => n12097, A2 => n12096, ZN => n12992);
   U17851 : NAND2_X1 port map( A1 => n12155, A2 => n12992, ZN => n12098);
   U17852 : MUX2_X1 port map( A => n28828, B => n12102, S => n12164, Z => 
                           n12107);
   U17854 : OAI21_X2 port map( B1 => n12107, B2 => n12167, A => n12106, ZN => 
                           n13370);
   U17855 : XNOR2_X1 port map( A => n13331, B => n13370, ZN => n12383);
   U17857 : OAI21_X1 port map( B1 => n12211, B2 => n12206, A => n12210, ZN => 
                           n12114);
   U17858 : NAND3_X1 port map( A1 => n12111, A2 => n12110, A3 => n12109, ZN => 
                           n12112);
   U17859 : XNOR2_X1 port map( A => n1857, B => n2441, ZN => n12116);
   U17860 : XNOR2_X1 port map( A => n12117, B => n12116, ZN => n12118);
   U17861 : INV_X1 port map( A => n29306, ZN => n14485);
   U17862 : NAND2_X1 port map( A1 => n570, A2 => n12180, ZN => n13205);
   U17863 : MUX2_X1 port map( A => n1890, B => n12177, S => n12176, Z => n13202
                           );
   U17864 : INV_X1 port map( A => n13202, ZN => n12123);
   U17865 : MUX2_X1 port map( A => n13205, B => n12123, S => n13206, Z => 
                           n12126);
   U17866 : NAND3_X1 port map( A1 => n12181, A2 => n12125, A3 => n12124, ZN => 
                           n13203);
   U17868 : NAND3_X1 port map( A1 => n12129, A2 => n12186, A3 => n12128, ZN => 
                           n12130);
   U17869 : INV_X1 port map( A => n13027, ZN => n12135);
   U17870 : XNOR2_X1 port map( A => n12135, B => n13296, ZN => n12139);
   U17871 : XNOR2_X1 port map( A => n13405, B => n3654, ZN => n12137);
   U17872 : XNOR2_X1 port map( A => n12136, B => n12137, ZN => n12138);
   U17873 : NAND3_X1 port map( A1 => n14485, A2 => n14484, A3 => n13947, ZN => 
                           n12140);
   U17874 : INV_X1 port map( A => n12142, ZN => n12143);
   U17875 : NOR2_X1 port map( A1 => n12146, A2 => n12145, ZN => n12147);
   U17876 : NOR3_X1 port map( A1 => n12151, A2 => n3961, A3 => n12991, ZN => 
                           n12153);
   U17877 : NOR2_X1 port map( A1 => n12153, A2 => n12152, ZN => n12154);
   U17878 : XNOR2_X1 port map( A => n13433, B => n12559, ZN => n12717);
   U17879 : INV_X1 port map( A => n12717, ZN => n12160);
   U17880 : XNOR2_X1 port map( A => n13236, B => n13039, ZN => n12609);
   U17881 : XNOR2_X1 port map( A => n12160, B => n12609, ZN => n12175);
   U17882 : XNOR2_X1 port map( A => n13547, B => n13338, ZN => n12173);
   U17883 : AND2_X1 port map( A1 => n12163, A2 => n1931, ZN => n12161);
   U17884 : NAND2_X1 port map( A1 => n12162, A2 => n12161, ZN => n12170);
   U17885 : NAND3_X1 port map( A1 => n28828, A2 => n11378, A3 => n12164, ZN => 
                           n12169);
   U17886 : NAND3_X1 port map( A1 => n12167, A2 => n11378, A3 => n1931, ZN => 
                           n12168);
   U17887 : XNOR2_X1 port map( A => n13113, B => n1923, ZN => n12172);
   U17888 : XNOR2_X1 port map( A => n12173, B => n12172, ZN => n12174);
   U17889 : NOR2_X1 port map( A1 => n12177, A2 => n12176, ZN => n12178);
   U17890 : MUX2_X1 port map( A => n12179, B => n12178, S => n570, Z => n12185)
                           ;
   U17891 : NOR2_X1 port map( A1 => n12181, A2 => n12180, ZN => n12182);
   U17892 : NOR2_X1 port map( A1 => n12183, A2 => n12182, ZN => n12184);
   U17894 : NAND2_X1 port map( A1 => n12186, A2 => n12189, ZN => n12197);
   U17895 : NAND2_X1 port map( A1 => n12187, A2 => n12186, ZN => n12193);
   U17896 : NOR2_X1 port map( A1 => n12190, A2 => n12189, ZN => n12191);
   U17897 : OAI21_X1 port map( B1 => n12193, B2 => n12192, A => n12191, ZN => 
                           n12196);
   U17898 : OAI211_X1 port map( C1 => n12198, C2 => n12197, A => n12196, B => 
                           n12195, ZN => n13428);
   U17899 : XNOR2_X1 port map( A => n13261, B => n13428, ZN => n12721);
   U17900 : XNOR2_X1 port map( A => n13552, B => n12854, ZN => n12199);
   U17901 : XNOR2_X1 port map( A => n12721, B => n12199, ZN => n12216);
   U17902 : OAI21_X1 port map( B1 => n12206, B2 => n12210, A => n12207, ZN => 
                           n12213);
   U17903 : AOI22_X1 port map( A1 => n12211, A2 => n12210, B1 => n12209, B2 => 
                           n12208, ZN => n12212);
   U17904 : OAI21_X1 port map( B1 => n6281, B2 => n12213, A => n12212, ZN => 
                           n12658);
   U17905 : XNOR2_X1 port map( A => n12658, B => n12799, ZN => n12484);
   U17906 : XNOR2_X1 port map( A => n13043, B => n3695, ZN => n12214);
   U17907 : XNOR2_X1 port map( A => n12484, B => n12214, ZN => n12215);
   U17908 : XNOR2_X1 port map( A => n12216, B => n12215, ZN => n14268);
   U17909 : AOI22_X1 port map( A1 => n28726, A2 => n12220, B1 => n12221, B2 => 
                           n12218, ZN => n12225);
   U17910 : MUX2_X1 port map( A => n12222, B => n12221, S => n12220, Z => 
                           n12223);
   U17911 : XNOR2_X1 port map( A => n12872, B => n13285, ZN => n12238);
   U17912 : NAND2_X1 port map( A1 => n12228, A2 => n13086, ZN => n12229);
   U17913 : XNOR2_X1 port map( A => n13448, B => n12472, ZN => n12423);
   U17914 : INV_X1 port map( A => n12423, ZN => n12237);
   U17915 : XNOR2_X1 port map( A => n12237, B => n12238, ZN => n12248);
   U17916 : XNOR2_X1 port map( A => n13055, B => n13226, ZN => n12246);
   U17917 : NAND2_X1 port map( A1 => n12242, A2 => n12241, ZN => n12243);
   U17918 : INV_X1 port map( A => n22072, ZN => n25361);
   U17919 : XNOR2_X1 port map( A => n12790, B => n25361, ZN => n12245);
   U17920 : XNOR2_X1 port map( A => n12245, B => n12246, ZN => n12247);
   U17921 : NAND2_X1 port map( A1 => n12252, A2 => n12249, ZN => n12250);
   U17922 : OAI21_X1 port map( B1 => n12251, B2 => n12252, A => n12250, ZN => 
                           n12255);
   U17923 : XNOR2_X1 port map( A => n12262, B => n12735, ZN => n12269);
   U17924 : XNOR2_X1 port map( A => n12866, B => n12632, ZN => n12268);
   U17925 : XNOR2_X1 port map( A => n12269, B => n12268, ZN => n12277);
   U17926 : MUX2_X1 port map( A => n28202, B => n12270, S => n12271, Z => 
                           n12274);
   U17927 : INV_X1 port map( A => n12271, ZN => n12272);
   U17928 : XNOR2_X1 port map( A => n13080, B => n13048, ZN => n12275);
   U17929 : XNOR2_X1 port map( A => n13219, B => n12275, ZN => n12276);
   U17930 : XNOR2_X1 port map( A => n12277, B => n12276, ZN => n13749);
   U17931 : INV_X1 port map( A => n13749, ZN => n14099);
   U17932 : MUX2_X1 port map( A => n12278, B => n12280, S => n12402, Z => 
                           n12287);
   U17933 : OAI21_X1 port map( B1 => n12407, B2 => n12281, A => n12280, ZN => 
                           n12282);
   U17934 : NAND3_X1 port map( A1 => n12284, A2 => n12283, A3 => n12282, ZN => 
                           n12285);
   U17935 : OAI21_X1 port map( B1 => n12287, B2 => n12286, A => n12285, ZN => 
                           n12752);
   U17936 : NAND4_X1 port map( A1 => n12061, A2 => n29324, A3 => n12291, A4 => 
                           n12290, ZN => n12294);
   U17937 : XNOR2_X1 port map( A => n12783, B => n13121, ZN => n12465);
   U17938 : XNOR2_X1 port map( A => n12465, B => n12298, ZN => n12326);
   U17940 : OAI21_X1 port map( B1 => n12305, B2 => n28807, A => n12300, ZN => 
                           n12310);
   U17941 : AND2_X1 port map( A1 => n12302, A2 => n12304, ZN => n12308);
   U17942 : NOR2_X1 port map( A1 => n12304, A2 => n12303, ZN => n12306);
   U17943 : AOI22_X1 port map( A1 => n12308, A2 => n4197, B1 => n12306, B2 => 
                           n12305, ZN => n12309);
   U17945 : NAND2_X1 port map( A1 => n12312, A2 => n12316, ZN => n12319);
   U17946 : NAND2_X1 port map( A1 => n12321, A2 => n12313, ZN => n12314);
   U17947 : OAI21_X1 port map( B1 => n12316, B2 => n12315, A => n12314, ZN => 
                           n12317);
   U17948 : INV_X1 port map( A => n12317, ZN => n12318);
   U17949 : NAND3_X1 port map( A1 => n12322, A2 => n12321, A3 => n12320, ZN => 
                           n12323);
   U17950 : XNOR2_X1 port map( A => n13419, B => n13272, ZN => n13140);
   U17951 : XNOR2_X1 port map( A => n12849, B => n3154, ZN => n12324);
   U17952 : XNOR2_X1 port map( A => n13140, B => n12324, ZN => n12325);
   U17953 : XNOR2_X2 port map( A => n12326, B => n12325, ZN => n14262);
   U17954 : NOR2_X1 port map( A1 => n14262, A2 => n1743, ZN => n12367);
   U17955 : AOI21_X1 port map( B1 => n12329, B2 => n12328, A => n12327, ZN => 
                           n12331);
   U17956 : MUX2_X1 port map( A => n12332, B => n12331, S => n12330, Z => 
                           n12336);
   U17957 : NOR2_X1 port map( A1 => n12334, A2 => n12333, ZN => n12335);
   U17958 : OAI22_X1 port map( A1 => n1291, A2 => n12341, B1 => n6919, B2 => 
                           n12340, ZN => n12348);
   U17960 : AOI21_X1 port map( B1 => n12346, B2 => n12345, A => n12344, ZN => 
                           n12347);
   U17961 : NOR2_X1 port map( A1 => n12348, A2 => n12347, ZN => n12572);
   U17962 : INV_X1 port map( A => n12572, ZN => n12768);
   U17963 : XNOR2_X1 port map( A => n12768, B => n12644, ZN => n12460);
   U17964 : XNOR2_X1 port map( A => n12460, B => n12349, ZN => n12366);
   U17965 : MUX2_X1 port map( A => n11467, B => n580, S => n12350, Z => n12351)
                           ;
   U17966 : NAND2_X1 port map( A1 => n12351, A2 => n29735, ZN => n12355);
   U17967 : XNOR2_X1 port map( A => n13298, B => n13461, ZN => n12749);
   U17968 : XNOR2_X1 port map( A => n12879, B => n3586, ZN => n12364);
   U17969 : XNOR2_X1 port map( A => n12749, B => n12364, ZN => n12365);
   U17970 : XNOR2_X1 port map( A => n12365, B => n12366, ZN => n14264);
   U17971 : OAI21_X1 port map( B1 => n13613, B2 => n12367, A => n13762, ZN => 
                           n12368);
   U17972 : XNOR2_X1 port map( A => n16310, B => n27105, ZN => n12631);
   U17973 : XNOR2_X1 port map( A => n13297, B => n29064, ZN => n12374);
   U17974 : XNOR2_X1 port map( A => n13459, B => n2511, ZN => n12373);
   U17975 : XNOR2_X1 port map( A => n12374, B => n12373, ZN => n12376);
   U17976 : XNOR2_X1 port map( A => n13027, B => n13542, ZN => n12375);
   U17977 : XNOR2_X1 port map( A => n12677, B => n3457, ZN => n12378);
   U17978 : XNOR2_X1 port map( A => n12379, B => n12378, ZN => n12382);
   U17979 : XNOR2_X1 port map( A => n13179, B => n13226, ZN => n13565);
   U17982 : INV_X1 port map( A => n14331, ZN => n14336);
   U17983 : XNOR2_X1 port map( A => n13249, B => n13533, ZN => n12691);
   U17984 : XNOR2_X1 port map( A => n12383, B => n12691, ZN => n12387);
   U17985 : XNOR2_X1 port map( A => n12385, B => n12384, ZN => n12386);
   U17986 : INV_X1 port map( A => n12388, ZN => n13005);
   U17987 : XNOR2_X1 port map( A => n12913, B => n12723, ZN => n12391);
   U17988 : XNOR2_X1 port map( A => n13348, B => n3491, ZN => n12390);
   U17989 : XNOR2_X1 port map( A => n12391, B => n12390, ZN => n12392);
   U17991 : INV_X1 port map( A => n14406, ZN => n13878);
   U17992 : NAND2_X1 port map( A1 => n14332, A2 => n13878, ZN => n12399);
   U17993 : INV_X1 port map( A => n13015, ZN => n12395);
   U17994 : XNOR2_X1 port map( A => n13278, B => n2987, ZN => n12394);
   U17995 : XNOR2_X1 port map( A => n12395, B => n12394, ZN => n12398);
   U17996 : XNOR2_X1 port map( A => n12738, B => n12868, ZN => n12815);
   U17997 : XNOR2_X1 port map( A => n13522, B => n12815, ZN => n12397);
   U17998 : INV_X1 port map( A => n14407, ZN => n13879);
   U17999 : NAND2_X1 port map( A1 => n12402, A2 => n12278, ZN => n12403);
   U18000 : NAND3_X1 port map( A1 => n12405, A2 => n12404, A3 => n12403, ZN => 
                           n12406);
   U18001 : OAI21_X1 port map( B1 => n12408, B2 => n12407, A => n12406, ZN => 
                           n12860);
   U18002 : XNOR2_X1 port map( A => n13109, B => n12860, ZN => n12807);
   U18003 : XNOR2_X1 port map( A => n13547, B => n13190, ZN => n12698);
   U18004 : XNOR2_X1 port map( A => n12698, B => n12807, ZN => n12412);
   U18005 : XNOR2_X1 port map( A => n13291, B => n3516, ZN => n12409);
   U18006 : XNOR2_X1 port map( A => n12410, B => n12409, ZN => n12411);
   U18007 : XNOR2_X1 port map( A => n12411, B => n12412, ZN => n14330);
   U18008 : INV_X1 port map( A => n14330, ZN => n14405);
   U18009 : NAND3_X1 port map( A1 => n13879, A2 => n14405, A3 => n29607, ZN => 
                           n12415);
   U18010 : NOR2_X1 port map( A1 => n29607, A2 => n13878, ZN => n12413);
   U18011 : NAND2_X1 port map( A1 => n14411, A2 => n12413, ZN => n12414);
   U18012 : NAND2_X1 port map( A1 => n14904, A2 => n14906, ZN => n14903);
   U18013 : INV_X1 port map( A => n14903, ZN => n13993);
   U18014 : XNOR2_X1 port map( A => n13402, B => n12588, ZN => n12419);
   U18015 : XNOR2_X1 port map( A => n13461, B => n22489, ZN => n12416);
   U18016 : XNOR2_X1 port map( A => n12417, B => n12416, ZN => n12418);
   U18017 : INV_X1 port map( A => n13287, ZN => n13378);
   U18018 : XNOR2_X1 port map( A => n12421, B => n13378, ZN => n12425);
   U18019 : XNOR2_X1 port map( A => n13451, B => n3380, ZN => n12422);
   U18020 : XNOR2_X1 port map( A => n12423, B => n12422, ZN => n12424);
   U18021 : NOR2_X1 port map( A1 => n30, A2 => n29628, ZN => n12452);
   U18022 : XNOR2_X1 port map( A => n13121, B => n13482, ZN => n12616);
   U18023 : INV_X1 port map( A => n12616, ZN => n12426);
   U18024 : XNOR2_X1 port map( A => n13419, B => n13270, ZN => n13374);
   U18025 : XNOR2_X1 port map( A => n12426, B => n13374, ZN => n12434);
   U18026 : XNOR2_X1 port map( A => n13269, B => n13136, ZN => n12433);
   U18027 : AND2_X1 port map( A1 => n12427, A2 => n12428, ZN => n12431);
   U18028 : XNOR2_X1 port map( A => n13369, B => n1175, ZN => n12432);
   U18029 : XNOR2_X1 port map( A => n12658, B => n13488, ZN => n12620);
   U18030 : XNOR2_X1 port map( A => n12620, B => n12435, ZN => n12439);
   U18031 : XNOR2_X1 port map( A => n13262, B => n12686, ZN => n12437);
   U18032 : XNOR2_X1 port map( A => n13428, B => n27298, ZN => n12436);
   U18033 : XNOR2_X1 port map( A => n12437, B => n12436, ZN => n12438);
   U18034 : NAND2_X1 port map( A1 => n13877, A2 => n14399, ZN => n12451);
   U18035 : XNOR2_X1 port map( A => n12776, B => n3036, ZN => n12440);
   U18036 : XNOR2_X1 port map( A => n13433, B => n12440, ZN => n12443);
   U18037 : INV_X1 port map( A => n13360, ZN => n12441);
   U18038 : XNOR2_X1 port map( A => n13236, B => n12441, ZN => n12442);
   U18039 : XNOR2_X1 port map( A => n12443, B => n12442, ZN => n12446);
   U18040 : INV_X1 port map( A => n13035, ZN => n12444);
   U18041 : XNOR2_X1 port map( A => n13364, B => n12699, ZN => n12987);
   U18042 : XNOR2_X1 port map( A => n12444, B => n12987, ZN => n12445);
   U18043 : NOR2_X1 port map( A1 => n14402, A2 => n14399, ZN => n13963);
   U18044 : XNOR2_X1 port map( A => n12894, B => n12632, ZN => n12449);
   U18045 : XNOR2_X1 port map( A => n12760, B => n3508, ZN => n12447);
   U18046 : XNOR2_X1 port map( A => n12447, B => n13445, ZN => n12448);
   U18047 : XNOR2_X1 port map( A => n13170, B => n12734, ZN => n12450);
   U18048 : INV_X1 port map( A => n15097, ZN => n14901);
   U18049 : XNOR2_X1 port map( A => n13020, B => n12453, ZN => n13147);
   U18050 : INV_X1 port map( A => n13147, ZN => n13497);
   U18051 : XNOR2_X1 port map( A => n13497, B => n12454, ZN => n12458);
   U18052 : XNOR2_X1 port map( A => n12763, B => n12632, ZN => n12456);
   U18053 : XNOR2_X1 port map( A => n12735, B => n5633, ZN => n12455);
   U18054 : XOR2_X1 port map( A => n12455, B => n12456, Z => n12457);
   U18055 : XNOR2_X1 port map( A => n12841, B => n13405, ZN => n12459);
   U18056 : XNOR2_X1 port map( A => n12460, B => n12459, ZN => n12464);
   U18057 : XNOR2_X1 port map( A => n13404, B => n3728, ZN => n12462);
   U18058 : XNOR2_X1 port map( A => n13028, B => n12461, ZN => n13505);
   U18059 : XNOR2_X1 port map( A => n12462, B => n13505, ZN => n12463);
   U18061 : XNOR2_X1 port map( A => n13478, B => n12780, ZN => n13141);
   U18062 : XNOR2_X1 port map( A => n13141, B => n12465, ZN => n12469);
   U18063 : XNOR2_X1 port map( A => n13272, B => n2912, ZN => n12467);
   U18064 : XNOR2_X1 port map( A => n12467, B => n12466, ZN => n12468);
   U18065 : XNOR2_X1 port map( A => n12469, B => n12468, ZN => n13686);
   U18066 : INV_X1 port map( A => n13686, ZN => n12481);
   U18067 : NAND2_X1 port map( A1 => n14417, A2 => n12470, ZN => n12475);
   U18068 : XNOR2_X1 port map( A => n13285, B => n12978, ZN => n13474);
   U18069 : XNOR2_X1 port map( A => n13054, B => n13563, ZN => n12471);
   U18070 : XNOR2_X1 port map( A => n12948, B => n13231, ZN => n12474);
   U18071 : INV_X1 port map( A => n1133, ZN => n28073);
   U18072 : XNOR2_X1 port map( A => n13381, B => n28073, ZN => n12473);
   U18073 : NAND2_X1 port map( A1 => n12475, A2 => n14414, ZN => n12489);
   U18074 : XNOR2_X1 port map( A => n13236, B => n13359, ZN => n12477);
   U18076 : XNOR2_X1 port map( A => n13113, B => n12985, ZN => n13509);
   U18077 : XNOR2_X1 port map( A => n12560, B => n1046, ZN => n12478);
   U18078 : XNOR2_X1 port map( A => n13509, B => n12478, ZN => n12479);
   U18079 : XNOR2_X1 port map( A => n13261, B => n13008, ZN => n13487);
   U18080 : XNOR2_X1 port map( A => n12965, B => n13386, ZN => n12482);
   U18081 : XNOR2_X1 port map( A => n13487, B => n12482, ZN => n12486);
   U18082 : XNOR2_X1 port map( A => n12566, B => n3317, ZN => n12483);
   U18083 : XNOR2_X1 port map( A => n12484, B => n12483, ZN => n12485);
   U18084 : XNOR2_X1 port map( A => n12486, B => n12485, ZN => n14215);
   U18085 : INV_X1 port map( A => n14215, ZN => n13891);
   U18086 : NAND3_X1 port map( A1 => n13891, A2 => n14415, A3 => n14217, ZN => 
                           n12487);
   U18087 : AND2_X1 port map( A1 => n14413, A2 => n12487, ZN => n12488);
   U18088 : NAND2_X1 port map( A1 => n12489, A2 => n12488, ZN => n14902);
   U18089 : INV_X1 port map( A => n14902, ZN => n14578);
   U18091 : XNOR2_X1 port map( A => n13457, B => n12490, ZN => n12494);
   U18092 : XNOR2_X1 port map( A => n12881, B => n27231, ZN => n12491);
   U18093 : XNOR2_X1 port map( A => n12492, B => n12491, ZN => n12493);
   U18095 : XNOR2_X1 port map( A => n13414, B => n13136, ZN => n12498);
   U18096 : INV_X1 port map( A => n12495, ZN => n12496);
   U18097 : XNOR2_X1 port map( A => n12496, B => n13137, ZN => n12847);
   U18098 : INV_X1 port map( A => n12847, ZN => n12497);
   U18099 : XNOR2_X1 port map( A => n12497, B => n12498, ZN => n12502);
   U18100 : XNOR2_X1 port map( A => n13413, B => n13420, ZN => n12500);
   U18101 : XNOR2_X1 port map( A => n12500, B => n12499, ZN => n12501);
   U18102 : INV_X1 port map( A => n857, ZN => n12503);
   U18103 : XNOR2_X1 port map( A => n12504, B => n12503, ZN => n12505);
   U18104 : XNOR2_X1 port map( A => n12505, B => n13278, ZN => n12506);
   U18105 : XNOR2_X1 port map( A => n13018, B => n12734, ZN => n13146);
   U18106 : XNOR2_X1 port map( A => n12506, B => n13146, ZN => n12515);
   U18107 : NOR2_X1 port map( A1 => n12508, A2 => n12507, ZN => n12509);
   U18108 : AOI22_X1 port map( A1 => n12511, A2 => n12510, B1 => n12509, B2 => 
                           n3653, ZN => n12513);
   U18109 : XNOR2_X1 port map( A => n12515, B => n13442, ZN => n13703);
   U18111 : XNOR2_X1 port map( A => n12696, B => n13035, ZN => n13155);
   U18112 : INV_X1 port map( A => n13155, ZN => n12522);
   U18113 : AOI21_X1 port map( B1 => n5947, B2 => n12578, A => n12516, ZN => 
                           n12518);
   U18114 : OAI22_X1 port map( A1 => n12518, A2 => n12583, B1 => n5947, B2 => 
                           n12272, ZN => n12520);
   U18115 : NAND2_X1 port map( A1 => n12520, A2 => n12519, ZN => n12521);
   U18117 : XNOR2_X1 port map( A => n13191, B => n13436, ZN => n12524);
   U18118 : XNOR2_X1 port map( A => n13291, B => n28294, ZN => n12523);
   U18119 : XNOR2_X1 port map( A => n12524, B => n12523, ZN => n12525);
   U18121 : INV_X1 port map( A => n3633, ZN => n12527);
   U18122 : XNOR2_X1 port map( A => n13159, B => n12527, ZN => n12528);
   U18123 : XNOR2_X1 port map( A => n13380, B => n13567, ZN => n12876);
   U18124 : XNOR2_X1 port map( A => n12528, B => n12876, ZN => n12531);
   U18125 : XNOR2_X1 port map( A => n13566, B => n12788, ZN => n13284);
   U18126 : XNOR2_X1 port map( A => n13230, B => n12529, ZN => n13180);
   U18128 : NAND2_X1 port map( A1 => n13872, A2 => n12534, ZN => n14425);
   U18129 : INV_X1 port map( A => n14425, ZN => n14306);
   U18130 : XNOR2_X1 port map( A => n13150, B => n3483, ZN => n12535);
   U18131 : XNOR2_X1 port map( A => n12535, B => n13260, ZN => n12537);
   U18132 : INV_X1 port map( A => n13265, ZN => n12536);
   U18133 : XNOR2_X1 port map( A => n12914, B => n12536, ZN => n13426);
   U18134 : XNOR2_X1 port map( A => n13426, B => n12537, ZN => n12540);
   U18135 : INV_X1 port map( A => n13553, ZN => n12657);
   U18136 : XNOR2_X1 port map( A => n12657, B => n12538, ZN => n12539);
   U18137 : NAND2_X1 port map( A1 => n14306, A2 => n14426, ZN => n14905);
   U18140 : INV_X1 port map( A => n15098, ZN => n15095);
   U18141 : XNOR2_X1 port map( A => n12762, B => n3035, ZN => n12543);
   U18142 : XNOR2_X1 port map( A => n12543, B => n13051, ZN => n12544);
   U18143 : XNOR2_X1 port map( A => n12544, B => n13315, ZN => n12547);
   U18144 : XNOR2_X1 port map( A => n13171, B => n12600, ZN => n12545);
   U18145 : XNOR2_X1 port map( A => n12816, B => n12545, ZN => n12546);
   U18146 : XNOR2_X1 port map( A => n12547, B => n12546, ZN => n14319);
   U18147 : INV_X1 port map( A => n14319, ZN => n14310);
   U18148 : XNOR2_X1 port map( A => n12548, B => n12872, ZN => n13095);
   U18149 : XNOR2_X1 port map( A => n13097, B => n13563, ZN => n12549);
   U18150 : XNOR2_X1 port map( A => n12549, B => n13095, ZN => n12553);
   U18151 : XNOR2_X1 port map( A => n12677, B => n3643, ZN => n12550);
   U18152 : XNOR2_X1 port map( A => n12550, B => n12551, ZN => n12552);
   U18153 : XNOR2_X1 port map( A => n13418, B => n13069, ZN => n12851);
   U18154 : XNOR2_X1 port map( A => n12851, B => n13332, ZN => n12558);
   U18155 : XNOR2_X1 port map( A => n13370, B => n12783, ZN => n12556);
   U18156 : XNOR2_X1 port map( A => n12827, B => n3501, ZN => n12555);
   U18157 : XNOR2_X1 port map( A => n12556, B => n12555, ZN => n12557);
   U18158 : XNOR2_X1 port map( A => n12558, B => n12557, ZN => n13257);
   U18159 : MUX2_X1 port map( A => n14310, B => n14313, S => n14320, Z => 
                           n12587);
   U18160 : XNOR2_X1 port map( A => n13432, B => n13034, ZN => n12562);
   U18161 : XNOR2_X1 port map( A => n12560, B => n12697, ZN => n13192);
   U18162 : INV_X1 port map( A => n13192, ZN => n12561);
   U18163 : XNOR2_X1 port map( A => n12561, B => n12562, ZN => n12565);
   U18164 : XNOR2_X1 port map( A => n13511, B => n13036, ZN => n13112);
   U18165 : XNOR2_X1 port map( A => n13338, B => n3323, ZN => n12563);
   U18166 : XNOR2_X1 port map( A => n13112, B => n12563, ZN => n12564);
   U18168 : INV_X1 port map( A => n14318, ZN => n13711);
   U18169 : XNOR2_X1 port map( A => n13005, B => n12566, ZN => n13197);
   U18170 : INV_X1 port map( A => n13197, ZN => n12567);
   U18171 : XNOR2_X1 port map( A => n12567, B => n13347, ZN => n12571);
   U18172 : XNOR2_X1 port map( A => n12568, B => n13245, ZN => n12570);
   U18173 : XNOR2_X1 port map( A => n13101, B => n3528, ZN => n12569);
   U18175 : NAND3_X1 port map( A1 => n14319, A2 => n13711, A3 => n13884, ZN => 
                           n12586);
   U18176 : XNOR2_X1 port map( A => n13406, B => n12841, ZN => n12574);
   U18177 : XNOR2_X1 port map( A => n12572, B => n13075, ZN => n12573);
   U18178 : XNOR2_X1 port map( A => n12574, B => n12573, ZN => n12584);
   U18179 : OAI21_X1 port map( B1 => n28202, B2 => n12576, A => n12575, ZN => 
                           n12582);
   U18180 : NAND2_X1 port map( A1 => n12579, A2 => n12578, ZN => n12580);
   U18181 : OAI211_X1 port map( C1 => n12583, C2 => n12582, A => n12581, B => 
                           n12580, ZN => n12883);
   U18182 : XNOR2_X1 port map( A => n13504, B => n12879, ZN => n13322);
   U18183 : XNOR2_X1 port map( A => n12747, B => n13404, ZN => n13503);
   U18184 : XNOR2_X1 port map( A => n12588, B => n13503, ZN => n12592);
   U18185 : XNOR2_X1 port map( A => n13458, B => n3666, ZN => n12590);
   U18186 : XNOR2_X1 port map( A => n13061, B => n12589, ZN => n13324);
   U18187 : XNOR2_X1 port map( A => n12590, B => n13324, ZN => n12591);
   U18188 : INV_X1 port map( A => n13803, ZN => n14297);
   U18189 : XNOR2_X1 port map( A => n12594, B => n12595, ZN => n13471);
   U18190 : XNOR2_X1 port map( A => n12833, B => n13471, ZN => n12599);
   U18191 : XNOR2_X1 port map( A => n12787, B => n13231, ZN => n12597);
   U18192 : XNOR2_X1 port map( A => n13450, B => n21537, ZN => n12596);
   U18193 : XNOR2_X1 port map( A => n12597, B => n12596, ZN => n12598);
   U18194 : XNOR2_X1 port map( A => n12599, B => n12598, ZN => n12607);
   U18195 : XNOR2_X1 port map( A => n12760, B => n1215, ZN => n12601);
   U18196 : XNOR2_X1 port map( A => n12601, B => n12600, ZN => n12602);
   U18197 : XNOR2_X1 port map( A => n12817, B => n13396, ZN => n13494);
   U18198 : XNOR2_X1 port map( A => n12602, B => n13494, ZN => n12606);
   U18199 : XNOR2_X1 port map( A => n12603, B => n13048, ZN => n12604);
   U18200 : XNOR2_X1 port map( A => n12604, B => n12813, ZN => n12605);
   U18201 : XNOR2_X1 port map( A => n13038, B => n12609, ZN => n12613);
   U18202 : XNOR2_X1 port map( A => n13432, B => n13337, ZN => n12611);
   U18203 : XNOR2_X1 port map( A => n12776, B => n1119, ZN => n12610);
   U18204 : XNOR2_X1 port map( A => n12611, B => n12610, ZN => n12612);
   U18205 : XNOR2_X1 port map( A => n12613, B => n12612, ZN => n14293);
   U18206 : AOI22_X1 port map( A1 => n12614, A2 => n14298, B1 => n14292, B2 => 
                           n14293, ZN => n12625);
   U18207 : XNOR2_X1 port map( A => n13418, B => n1928, ZN => n12615);
   U18208 : XNOR2_X1 port map( A => n13067, B => n1906, ZN => n13329);
   U18209 : XNOR2_X1 port map( A => n13329, B => n12615, ZN => n12618);
   U18210 : XNOR2_X1 port map( A => n13479, B => n12616, ZN => n12617);
   U18212 : INV_X1 port map( A => n14292, ZN => n13697);
   U18213 : OAI22_X1 port map( A1 => n14297, A2 => n14293, B1 => n14295, B2 => 
                           n13697, ZN => n12623);
   U18214 : XNOR2_X1 port map( A => n12722, B => n13386, ZN => n13490);
   U18215 : XNOR2_X1 port map( A => n13556, B => n13043, ZN => n13350);
   U18216 : XNOR2_X1 port map( A => n13490, B => n13350, ZN => n12622);
   U18217 : XNOR2_X1 port map( A => n13245, B => n3049, ZN => n12619);
   U18218 : XNOR2_X1 port map( A => n12620, B => n12619, ZN => n12621);
   U18219 : XNOR2_X1 port map( A => n12622, B => n12621, ZN => n13306);
   U18220 : NAND2_X1 port map( A1 => n12623, A2 => n14291, ZN => n12624);
   U18221 : AND2_X1 port map( A1 => n3315, A2 => n15094, ZN => n12627);
   U18222 : NOR2_X1 port map( A1 => n14578, A2 => n3315, ZN => n12626);
   U18223 : AOI22_X1 port map( A1 => n15095, A2 => n12627, B1 => n12626, B2 => 
                           n14903, ZN => n12628);
   U18224 : NAND2_X1 port map( A1 => n12629, A2 => n12628, ZN => n16527);
   U18225 : INV_X1 port map( A => n16527, ZN => n12630);
   U18226 : XNOR2_X1 port map( A => n12631, B => n12630, ZN => n13130);
   U18227 : XNOR2_X1 port map( A => n1885, B => n3423, ZN => n12633);
   U18228 : XNOR2_X1 port map( A => n13220, B => n12633, ZN => n12636);
   U18229 : XNOR2_X1 port map( A => n12637, B => n13121, ZN => n13247);
   U18230 : XNOR2_X1 port map( A => n13247, B => n12638, ZN => n12643);
   U18231 : INV_X1 port map( A => n13371, ZN => n12639);
   U18232 : XNOR2_X1 port map( A => n1905, B => n12639, ZN => n12641);
   U18233 : XNOR2_X1 port map( A => n12495, B => n26214, ZN => n12640);
   U18234 : XNOR2_X1 port map( A => n12641, B => n12640, ZN => n12642);
   U18235 : XNOR2_X1 port map( A => n12746, B => n12644, ZN => n13224);
   U18236 : INV_X1 port map( A => n13224, ZN => n12647);
   U18237 : INV_X1 port map( A => n12881, ZN => n12645);
   U18238 : XNOR2_X1 port map( A => n13539, B => n12645, ZN => n12646);
   U18239 : XNOR2_X1 port map( A => n12647, B => n12646, ZN => n12651);
   U18240 : XNOR2_X1 port map( A => n13404, B => n3211, ZN => n12649);
   U18241 : XNOR2_X1 port map( A => n12649, B => n12648, ZN => n12650);
   U18242 : XNOR2_X1 port map( A => n12651, B => n12650, ZN => n13851);
   U18243 : INV_X1 port map( A => n13851, ZN => n14176);
   U18244 : MUX2_X1 port map( A => n14177, B => n14181, S => n14176, Z => 
                           n12673);
   U18245 : INV_X1 port map( A => n13227, ZN => n12729);
   U18246 : XNOR2_X1 port map( A => n12729, B => n13231, ZN => n13096);
   U18247 : XNOR2_X1 port map( A => n12652, B => n13096, ZN => n12656);
   U18248 : XNOR2_X1 port map( A => n13567, B => n2889, ZN => n12653);
   U18249 : XNOR2_X1 port map( A => n12654, B => n12653, ZN => n12655);
   U18250 : XNOR2_X1 port map( A => n12657, B => n12854, ZN => n12659);
   U18251 : XNOR2_X1 port map( A => n12659, B => n13243, ZN => n12663);
   U18252 : XNOR2_X1 port map( A => n13386, B => n13556, ZN => n12661);
   U18253 : XNOR2_X1 port map( A => n4670, B => n24897, ZN => n12660);
   U18254 : XNOR2_X1 port map( A => n12661, B => n12660, ZN => n12662);
   U18255 : XNOR2_X1 port map( A => n12663, B => n12662, ZN => n13753);
   U18256 : NAND2_X1 port map( A1 => n5693, A2 => n14451, ZN => n12671);
   U18257 : INV_X1 port map( A => n12985, ZN => n12664);
   U18258 : XNOR2_X1 port map( A => n13236, B => n12664, ZN => n12666);
   U18259 : XNOR2_X1 port map( A => n13338, B => n13109, ZN => n12665);
   U18260 : XNOR2_X1 port map( A => n12665, B => n12666, ZN => n12670);
   U18261 : XNOR2_X1 port map( A => n13359, B => n13337, ZN => n12668);
   U18262 : XNOR2_X1 port map( A => n13191, B => n2960, ZN => n12667);
   U18263 : XNOR2_X1 port map( A => n12668, B => n12667, ZN => n12669);
   U18264 : XNOR2_X1 port map( A => n12670, B => n12669, ZN => n14178);
   U18265 : OAI21_X1 port map( B1 => n12671, B2 => n14176, A => n13932, ZN => 
                           n12672);
   U18266 : XNOR2_X1 port map( A => n13230, B => n2527, ZN => n12675);
   U18267 : INV_X1 port map( A => n12787, ZN => n12674);
   U18268 : XNOR2_X1 port map( A => n12675, B => n12674, ZN => n12676);
   U18269 : XNOR2_X1 port map( A => n12676, B => n13565, ZN => n12679);
   U18270 : XNOR2_X1 port map( A => n13451, B => n12677, ZN => n12678);
   U18271 : XNOR2_X1 port map( A => n12678, B => n13380, ZN => n12983);
   U18272 : XNOR2_X1 port map( A => n12679, B => n12983, ZN => n12711);
   U18273 : XNOR2_X1 port map( A => n12760, B => n28327, ZN => n12680);
   U18274 : XNOR2_X1 port map( A => n29140, B => n12681, ZN => n12682);
   U18275 : XNOR2_X1 port map( A => n12683, B => n12682, ZN => n12712);
   U18276 : XNOR2_X1 port map( A => n13150, B => n12684, ZN => n13388);
   U18277 : XNOR2_X1 port map( A => n12685, B => n13388, ZN => n12690);
   U18278 : XNOR2_X1 port map( A => n13488, B => n72, ZN => n12687);
   U18279 : XNOR2_X1 port map( A => n12688, B => n12687, ZN => n12689);
   U18280 : XNOR2_X1 port map( A => n12690, B => n12689, ZN => n13967);
   U18282 : XNOR2_X1 port map( A => n13370, B => n13137, ZN => n13000);
   U18283 : XNOR2_X1 port map( A => n13000, B => n12691, ZN => n12695);
   U18284 : XNOR2_X1 port map( A => n1857, B => n13420, ZN => n12693);
   U18285 : XNOR2_X1 port map( A => n13482, B => n27462, ZN => n12692);
   U18286 : XNOR2_X1 port map( A => n12693, B => n12692, ZN => n12694);
   U18287 : XNOR2_X1 port map( A => n12696, B => n12697, ZN => n13363);
   U18288 : XNOR2_X1 port map( A => n12698, B => n13363, ZN => n12703);
   U18289 : XNOR2_X1 port map( A => n12776, B => n2325, ZN => n12700);
   U18290 : XNOR2_X1 port map( A => n12701, B => n12700, ZN => n12702);
   U18291 : OAI21_X1 port map( B1 => n14463, B2 => n13967, A => n12704, ZN => 
                           n12715);
   U18292 : INV_X1 port map( A => n13967, ZN => n14456);
   U18293 : NOR2_X1 port map( A1 => n14455, A2 => n14456, ZN => n12714);
   U18294 : XNOR2_X1 port map( A => n13406, B => n13401, ZN => n12706);
   U18295 : XNOR2_X1 port map( A => n12705, B => n12706, ZN => n12710);
   U18296 : XNOR2_X1 port map( A => n13208, B => n3697, ZN => n12708);
   U18297 : XNOR2_X1 port map( A => n12707, B => n12708, ZN => n12709);
   U18298 : NOR2_X1 port map( A1 => n12711, A2 => n427, ZN => n12713);
   U18299 : XNOR2_X1 port map( A => n13035, B => n13109, ZN => n12716);
   U18300 : XNOR2_X1 port map( A => n12717, B => n12716, ZN => n12720);
   U18301 : XNOR2_X1 port map( A => n13113, B => n13364, ZN => n13293);
   U18302 : XNOR2_X1 port map( A => n12808, B => n2602, ZN => n12718);
   U18303 : XNOR2_X1 port map( A => n12718, B => n13293, ZN => n12719);
   U18304 : INV_X1 port map( A => n13933, ZN => n14465);
   U18305 : XNOR2_X1 port map( A => n13346, B => n12721, ZN => n12726);
   U18306 : XNOR2_X1 port map( A => n12722, B => n12723, ZN => n12822);
   U18307 : XNOR2_X1 port map( A => n13263, B => n27452, ZN => n12724);
   U18308 : XNOR2_X1 port map( A => n12822, B => n12724, ZN => n12725);
   U18309 : INV_X1 port map( A => n14469, ZN => n14185);
   U18310 : XNOR2_X1 port map( A => n12595, B => n13159, ZN => n12728);
   U18311 : XNOR2_X1 port map( A => n12980, B => n13285, ZN => n12727);
   U18312 : XNOR2_X1 port map( A => n12727, B => n12728, ZN => n12733);
   U18313 : XNOR2_X1 port map( A => n12790, B => n12729, ZN => n12731);
   U18314 : XNOR2_X1 port map( A => n13448, B => n3482, ZN => n12730);
   U18315 : XNOR2_X1 port map( A => n12731, B => n12730, ZN => n12732);
   U18316 : XNOR2_X1 port map( A => n12732, B => n12733, ZN => n12743);
   U18317 : NAND2_X1 port map( A1 => n14185, A2 => n12743, ZN => n12744);
   U18318 : XNOR2_X1 port map( A => n12894, B => n13080, ZN => n13280);
   U18319 : INV_X1 port map( A => n13280, ZN => n12737);
   U18320 : INV_X1 port map( A => n12734, ZN => n12736);
   U18321 : XNOR2_X1 port map( A => n12736, B => n12762, ZN => n13318);
   U18322 : XNOR2_X1 port map( A => n12737, B => n13318, ZN => n12742);
   U18323 : XNOR2_X1 port map( A => n12738, B => n2522, ZN => n12740);
   U18324 : XNOR2_X1 port map( A => n13445, B => n12817, ZN => n12739);
   U18325 : XNOR2_X1 port map( A => n12740, B => n12739, ZN => n12741);
   U18326 : XNOR2_X1 port map( A => n12742, B => n12741, ZN => n13677);
   U18327 : INV_X1 port map( A => n13677, ZN => n14184);
   U18330 : XNOR2_X1 port map( A => n13025, B => n2984, ZN => n12748);
   U18331 : XNOR2_X1 port map( A => n12747, B => n29064, ZN => n12839);
   U18332 : XNOR2_X1 port map( A => n12839, B => n12748, ZN => n12751);
   U18333 : XNOR2_X1 port map( A => n13325, B => n12749, ZN => n12750);
   U18334 : XNOR2_X1 port map( A => n12750, B => n12751, ZN => n13678);
   U18335 : INV_X1 port map( A => n12752, ZN => n12753);
   U18336 : XNOR2_X1 port map( A => n13374, B => n13328, ZN => n12757);
   U18337 : XNOR2_X1 port map( A => n12830, B => n13272, ZN => n12755);
   U18338 : XNOR2_X1 port map( A => n13118, B => n2385, ZN => n12754);
   U18339 : XNOR2_X1 port map( A => n12755, B => n12754, ZN => n12756);
   U18340 : NAND3_X1 port map( A1 => n14182, A2 => n14469, A3 => n14464, ZN => 
                           n12758);
   U18341 : XNOR2_X1 port map( A => n12760, B => n13278, ZN => n13496);
   U18342 : INV_X1 port map( A => n13496, ZN => n12761);
   U18343 : XNOR2_X1 port map( A => n12761, B => n13277, ZN => n12767);
   U18344 : XNOR2_X1 port map( A => n12762, B => n2306, ZN => n12764);
   U18345 : XNOR2_X1 port map( A => n12764, B => n12763, ZN => n12765);
   U18346 : XNOR2_X1 port map( A => n12765, B => n13167, ZN => n12766);
   U18348 : XNOR2_X1 port map( A => n12768, B => n13405, ZN => n12769);
   U18349 : XNOR2_X1 port map( A => n13501, B => n12769, ZN => n12773);
   U18350 : XNOR2_X1 port map( A => n13543, B => n12931, ZN => n12771);
   U18351 : XNOR2_X1 port map( A => n13209, B => n3109, ZN => n12770);
   U18352 : XNOR2_X1 port map( A => n12771, B => n12770, ZN => n12772);
   U18353 : XNOR2_X1 port map( A => n12773, B => n12772, ZN => n14497);
   U18355 : XNOR2_X1 port map( A => n13290, B => n12775, ZN => n12779);
   U18356 : XNOR2_X1 port map( A => n12919, B => n2996, ZN => n12777);
   U18357 : XNOR2_X1 port map( A => n12777, B => n13513, ZN => n12778);
   U18358 : XNOR2_X1 port map( A => n12780, B => n13414, ZN => n12782);
   U18359 : INV_X1 port map( A => n12944, ZN => n12781);
   U18360 : XNOR2_X1 port map( A => n12781, B => n12782, ZN => n12786);
   U18361 : INV_X1 port map( A => n3134, ZN => n27643);
   U18362 : XNOR2_X1 port map( A => n12783, B => n27643, ZN => n12784);
   U18363 : XNOR2_X1 port map( A => n12784, B => n13274, ZN => n12785);
   U18364 : XNOR2_X1 port map( A => n12786, B => n12785, ZN => n13672);
   U18365 : INV_X1 port map( A => n13672, ZN => n14491);
   U18366 : NAND2_X1 port map( A1 => n14154, A2 => n14491, ZN => n12795);
   U18367 : INV_X1 port map( A => n12949, ZN => n13472);
   U18368 : XNOR2_X1 port map( A => n13472, B => n12789, ZN => n12794);
   U18369 : XNOR2_X1 port map( A => n12790, B => n3554, ZN => n12791);
   U18370 : XNOR2_X1 port map( A => n12791, B => n12792, ZN => n12793);
   U18371 : MUX2_X1 port map( A => n12796, B => n12795, S => n14492, Z => 
                           n12805);
   U18372 : XNOR2_X1 port map( A => n13265, B => n13485, ZN => n12798);
   U18373 : XNOR2_X1 port map( A => n12798, B => n12797, ZN => n12803);
   U18374 : XNOR2_X1 port map( A => n12799, B => n13262, ZN => n12801);
   U18375 : XNOR2_X1 port map( A => n13488, B => n2465, ZN => n12800);
   U18376 : XNOR2_X1 port map( A => n12801, B => n12800, ZN => n12802);
   U18377 : XNOR2_X1 port map( A => n12803, B => n12802, ZN => n13855);
   U18378 : INV_X1 port map( A => n13855, ZN => n14493);
   U18379 : OAI21_X1 port map( B1 => n4549, B2 => n15101, A => n549, ZN => 
                           n12891);
   U18380 : INV_X1 port map( A => n13549, ZN => n12806);
   U18381 : XNOR2_X1 port map( A => n12806, B => n12807, ZN => n12812);
   U18382 : XNOR2_X1 port map( A => n12808, B => n2544, ZN => n12810);
   U18383 : INV_X1 port map( A => n12809, ZN => n13342);
   U18384 : XNOR2_X1 port map( A => n13342, B => n12810, ZN => n12811);
   U18385 : INV_X1 port map( A => n13048, ZN => n12814);
   U18386 : XNOR2_X1 port map( A => n12814, B => n12813, ZN => n13314);
   U18387 : XNOR2_X1 port map( A => n13314, B => n12815, ZN => n12821);
   U18388 : XNOR2_X1 port map( A => n12816, B => n13493, ZN => n12819);
   U18389 : XNOR2_X1 port map( A => n12817, B => n2353, ZN => n12818);
   U18390 : XNOR2_X1 port map( A => n12819, B => n12818, ZN => n12820);
   U18391 : XNOR2_X1 port map( A => n13557, B => n12913, ZN => n12824);
   U18392 : XNOR2_X1 port map( A => n13484, B => n3662, ZN => n12823);
   U18393 : XNOR2_X1 port map( A => n12824, B => n12823, ZN => n12825);
   U18394 : XNOR2_X1 port map( A => n12827, B => n5059, ZN => n12828);
   U18395 : XNOR2_X1 port map( A => n13118, B => n12830, ZN => n12831);
   U18396 : INV_X1 port map( A => n13329, ZN => n12832);
   U18397 : XNOR2_X1 port map( A => n13563, B => n12595, ZN => n12836);
   U18398 : XNOR2_X1 port map( A => n13473, B => n26909, ZN => n12835);
   U18399 : XNOR2_X1 port map( A => n12836, B => n12835, ZN => n12837);
   U18400 : INV_X1 port map( A => n12839, ZN => n12840);
   U18401 : XNOR2_X1 port map( A => n12840, B => n13324, ZN => n12845);
   U18402 : XNOR2_X1 port map( A => n12841, B => n13459, ZN => n12843);
   U18403 : XNOR2_X1 port map( A => n13504, B => n2350, ZN => n12842);
   U18404 : XNOR2_X1 port map( A => n12843, B => n12842, ZN => n12844);
   U18405 : NAND3_X1 port map( A1 => n4549, A2 => n15422, A3 => n14575, ZN => 
                           n12890);
   U18406 : XNOR2_X1 port map( A => n13331, B => n12849, ZN => n12850);
   U18407 : INV_X1 port map( A => n12851, ZN => n13248);
   U18408 : XNOR2_X1 port map( A => n13150, B => n3219, ZN => n12852);
   U18409 : XNOR2_X1 port map( A => n13553, B => n12852, ZN => n12853);
   U18410 : XNOR2_X1 port map( A => n13246, B => n12853, ZN => n12857);
   U18411 : XNOR2_X1 port map( A => n12913, B => n13245, ZN => n12855);
   U18412 : XNOR2_X1 port map( A => n12855, B => n12854, ZN => n12856);
   U18413 : XNOR2_X1 port map( A => n12857, B => n12856, ZN => n14207);
   U18414 : INV_X1 port map( A => n13036, ZN => n12858);
   U18415 : XNOR2_X1 port map( A => n13341, B => n12858, ZN => n13240);
   U18416 : XNOR2_X1 port map( A => n13338, B => n13432, ZN => n12859);
   U18417 : XNOR2_X1 port map( A => n13240, B => n12859, ZN => n12864);
   U18418 : XNOR2_X1 port map( A => n12860, B => n13191, ZN => n12924);
   U18419 : INV_X1 port map( A => n1161, ZN => n27730);
   U18420 : XNOR2_X1 port map( A => n12861, B => n27730, ZN => n12862);
   U18421 : XNOR2_X1 port map( A => n12924, B => n12862, ZN => n12863);
   U18422 : XNOR2_X1 port map( A => n12864, B => n12863, ZN => n14433);
   U18423 : MUX2_X1 port map( A => n1841, B => n14207, S => n14433, Z => n12888
                           );
   U18424 : XNOR2_X1 port map( A => n13018, B => n1179, ZN => n12865);
   U18425 : XNOR2_X1 port map( A => n12868, B => n12867, ZN => n12892);
   U18426 : XNOR2_X1 port map( A => n13444, B => n13525, ZN => n12869);
   U18427 : XNOR2_X1 port map( A => n12869, B => n13051, ZN => n13221);
   U18428 : INV_X1 port map( A => n13221, ZN => n12870);
   U18429 : XNOR2_X2 port map( A => n12871, B => n12870, ZN => n14438);
   U18430 : XNOR2_X1 port map( A => n12872, B => n13447, ZN => n12874);
   U18431 : INV_X1 port map( A => n13229, ZN => n12873);
   U18432 : XNOR2_X1 port map( A => n13450, B => n25044, ZN => n12875);
   U18433 : XNOR2_X1 port map( A => n12876, B => n12875, ZN => n12877);
   U18434 : XNOR2_X1 port map( A => n12879, B => n3527, ZN => n12880);
   U18435 : XNOR2_X1 port map( A => n12880, B => n29494, ZN => n12882);
   U18436 : XNOR2_X1 port map( A => n12881, B => n13459, ZN => n12929);
   U18437 : XNOR2_X1 port map( A => n12883, B => n13075, ZN => n12884);
   U18439 : INV_X1 port map( A => n15423, ZN => n14577);
   U18440 : NAND3_X1 port map( A1 => n15102, A2 => n15105, A3 => n14577, ZN => 
                           n12889);
   U18441 : XNOR2_X1 port map( A => n13167, B => n13493, ZN => n12893);
   U18442 : XNOR2_X1 port map( A => n12892, B => n12893, ZN => n12898);
   U18443 : XNOR2_X1 port map( A => n13166, B => n1225, ZN => n12896);
   U18444 : XNOR2_X1 port map( A => n12894, B => n13444, ZN => n12895);
   U18445 : XNOR2_X1 port map( A => n12895, B => n12896, ZN => n12897);
   U18446 : XNOR2_X1 port map( A => n13179, B => n13447, ZN => n12900);
   U18447 : XNOR2_X1 port map( A => n12899, B => n12900, ZN => n12903);
   U18448 : XNOR2_X1 port map( A => n13567, B => n3083, ZN => n12901);
   U18449 : XNOR2_X1 port map( A => n12904, B => n12905, ZN => n12910);
   U18450 : XNOR2_X1 port map( A => n12495, B => n2389, ZN => n12907);
   U18451 : XNOR2_X1 port map( A => n12908, B => n12907, ZN => n12909);
   U18452 : MUX2_X1 port map( A => n14082, B => n14084, S => n14287, Z => 
                           n12928);
   U18453 : INV_X1 port map( A => n12913, ZN => n12915);
   U18454 : XNOR2_X1 port map( A => n12914, B => n12915, ZN => n12917);
   U18455 : XNOR2_X1 port map( A => n13484, B => n3116, ZN => n12916);
   U18456 : XNOR2_X1 port map( A => n12917, B => n12916, ZN => n12918);
   U18457 : NOR2_X1 port map( A1 => n28625, A2 => n14282, ZN => n12927);
   U18459 : XNOR2_X1 port map( A => n12921, B => n12920, ZN => n12926);
   U18460 : INV_X1 port map( A => n3463, ZN => n12922);
   U18461 : XNOR2_X1 port map( A => n13511, B => n12922, ZN => n12923);
   U18462 : XNOR2_X1 port map( A => n12924, B => n12923, ZN => n12925);
   U18463 : XNOR2_X1 port map( A => n12926, B => n12925, ZN => n14083);
   U18464 : XNOR2_X1 port map( A => n12929, B => n12930, ZN => n12935);
   U18465 : XNOR2_X1 port map( A => n12931, B => n3710, ZN => n12932);
   U18466 : XNOR2_X1 port map( A => n12933, B => n12932, ZN => n12934);
   U18467 : XNOR2_X1 port map( A => n12935, B => n12934, ZN => n14286);
   U18468 : INV_X1 port map( A => n14084, ZN => n14281);
   U18471 : AND2_X1 port map( A1 => n14106, A2 => n14105, ZN => n14234);
   U18472 : NAND2_X1 port map( A1 => n14234, A2 => n14102, ZN => n12941);
   U18473 : BUF_X2 port map( A => n13606, Z => n14230);
   U18474 : NAND2_X1 port map( A1 => n12938, A2 => n14230, ZN => n12940);
   U18475 : NAND2_X1 port map( A1 => n14102, A2 => n14107, ZN => n12939);
   U18478 : XNOR2_X1 port map( A => n13141, B => n12943, ZN => n12947);
   U18479 : XNOR2_X1 port map( A => n13419, B => n1184, ZN => n12945);
   U18480 : XNOR2_X1 port map( A => n12944, B => n12945, ZN => n12946);
   U18481 : XNOR2_X1 port map( A => n13448, B => n12948, ZN => n13379);
   U18482 : XNOR2_X1 port map( A => n12949, B => n13379, ZN => n12953);
   U18483 : XNOR2_X1 port map( A => n13230, B => n3493, ZN => n12951);
   U18484 : XNOR2_X1 port map( A => n12978, B => n13055, ZN => n12950);
   U18485 : XNOR2_X1 port map( A => n12951, B => n12950, ZN => n12952);
   U18486 : XNOR2_X1 port map( A => n12954, B => n13445, ZN => n13394);
   U18487 : XNOR2_X1 port map( A => n13394, B => n13496, ZN => n12959);
   U18488 : XNOR2_X1 port map( A => n13020, B => n13048, ZN => n12957);
   U18489 : XNOR2_X1 port map( A => n12955, B => n3212, ZN => n12956);
   U18490 : XNOR2_X1 port map( A => n12956, B => n12957, ZN => n12958);
   U18491 : INV_X1 port map( A => n13061, ZN => n12960);
   U18492 : XNOR2_X1 port map( A => n13028, B => n1123, ZN => n12961);
   U18493 : XNOR2_X1 port map( A => n12962, B => n12961, ZN => n12964);
   U18494 : XNOR2_X1 port map( A => n13428, B => n12965, ZN => n13389);
   U18495 : XNOR2_X1 port map( A => n12966, B => n13389, ZN => n12970);
   U18496 : XNOR2_X1 port map( A => n13008, B => n13043, ZN => n12968);
   U18497 : XNOR2_X1 port map( A => n13488, B => n3622, ZN => n12967);
   U18498 : XNOR2_X1 port map( A => n12968, B => n12967, ZN => n12969);
   U18499 : XNOR2_X1 port map( A => n13039, B => n135, ZN => n12971);
   U18500 : XNOR2_X1 port map( A => n12985, B => n12971, ZN => n12973);
   U18501 : XNOR2_X1 port map( A => n12973, B => n12972, ZN => n12975);
   U18502 : XNOR2_X1 port map( A => n13513, B => n13433, ZN => n12974);
   U18503 : NAND2_X1 port map( A1 => n12976, A2 => n14365, ZN => n14370);
   U18504 : XNOR2_X1 port map( A => n12978, B => n3276, ZN => n12979);
   U18505 : XNOR2_X1 port map( A => n12979, B => n28587, ZN => n12982);
   U18506 : XNOR2_X1 port map( A => n12980, B => n13562, ZN => n12981);
   U18507 : XNOR2_X1 port map( A => n12982, B => n12981, ZN => n12984);
   U18508 : XNOR2_X1 port map( A => n12985, B => n2598, ZN => n12986);
   U18509 : XNOR2_X1 port map( A => n13341, B => n13436, ZN => n13545);
   U18510 : XNOR2_X1 port map( A => n12986, B => n13545, ZN => n12989);
   U18511 : XNOR2_X1 port map( A => n13363, B => n12987, ZN => n12988);
   U18512 : XNOR2_X1 port map( A => n12989, B => n12988, ZN => n13832);
   U18513 : MUX2_X1 port map( A => n12992, B => n12991, S => n12990, Z => 
                           n12993);
   U18514 : NAND2_X1 port map( A1 => n12994, A2 => n12993, ZN => n12997);
   U18515 : INV_X1 port map( A => n12995, ZN => n12996);
   U18516 : NAND2_X1 port map( A1 => n12997, A2 => n12996, ZN => n12999);
   U18517 : INV_X1 port map( A => n13413, ZN => n12998);
   U18518 : XNOR2_X1 port map( A => n12998, B => n12999, ZN => n13530);
   U18519 : XNOR2_X1 port map( A => n13000, B => n13530, ZN => n13004);
   U18520 : XNOR2_X1 port map( A => n1857, B => n13478, ZN => n13002);
   U18521 : XNOR2_X1 port map( A => n13270, B => n3414, ZN => n13001);
   U18522 : XNOR2_X1 port map( A => n13002, B => n13001, ZN => n13003);
   U18523 : NAND3_X1 port map( A1 => n13829, A2 => n13832, A3 => n14278, ZN => 
                           n13024);
   U18524 : XNOR2_X1 port map( A => n13005, B => n13263, ZN => n13007);
   U18525 : INV_X1 port map( A => n13348, ZN => n13006);
   U18526 : XNOR2_X1 port map( A => n13006, B => n13265, ZN => n13554);
   U18527 : XNOR2_X1 port map( A => n13150, B => n2946, ZN => n13009);
   U18528 : XNOR2_X1 port map( A => n13010, B => n13009, ZN => n13011);
   U18529 : XNOR2_X1 port map( A => n13013, B => n13014, ZN => n13016);
   U18530 : XNOR2_X1 port map( A => n13016, B => n13015, ZN => n13023);
   U18531 : INV_X1 port map( A => n13017, ZN => n13019);
   U18532 : XNOR2_X1 port map( A => n13018, B => n13019, ZN => n13393);
   U18533 : XNOR2_X1 port map( A => n13020, B => n3462, ZN => n13021);
   U18534 : XNOR2_X1 port map( A => n13393, B => n13021, ZN => n13022);
   U18535 : NAND2_X1 port map( A1 => n14362, A2 => n14358, ZN => n14275);
   U18536 : XNOR2_X1 port map( A => n13025, B => n29495, ZN => n13026);
   U18537 : XNOR2_X1 port map( A => n13027, B => n13026, ZN => n13031);
   U18538 : XNOR2_X1 port map( A => n13028, B => n3660, ZN => n13029);
   U18539 : XNOR2_X1 port map( A => n13456, B => n13029, ZN => n13030);
   U18540 : XNOR2_X1 port map( A => n13031, B => n13030, ZN => n14360);
   U18541 : OAI21_X1 port map( B1 => n14275, B2 => n14360, A => n13032, ZN => 
                           n13033);
   U18542 : XNOR2_X1 port map( A => n13035, B => n13034, ZN => n13340);
   U18543 : XNOR2_X1 port map( A => n13036, B => n13360, ZN => n13037);
   U18544 : XNOR2_X1 port map( A => n13340, B => n13037, ZN => n13041);
   U18545 : XNOR2_X1 port map( A => n13039, B => n1887, ZN => n13040);
   U18546 : INV_X1 port map( A => n13490, ZN => n13042);
   U18547 : XNOR2_X1 port map( A => n13346, B => n13042, ZN => n13047);
   U18548 : XNOR2_X1 port map( A => n13043, B => n13262, ZN => n13045);
   U18549 : XNOR2_X1 port map( A => n13101, B => n3451, ZN => n13044);
   U18550 : XNOR2_X1 port map( A => n13045, B => n13044, ZN => n13046);
   U18551 : XNOR2_X1 port map( A => n13170, B => n3196, ZN => n13049);
   U18552 : XNOR2_X1 port map( A => n13049, B => n13048, ZN => n13050);
   U18553 : XNOR2_X1 port map( A => n13050, B => n13318, ZN => n13053);
   U18554 : XNOR2_X1 port map( A => n13494, B => n13051, ZN => n13052);
   U18555 : XNOR2_X1 port map( A => n13353, B => n13471, ZN => n13059);
   U18556 : XNOR2_X1 port map( A => n13097, B => n13175, ZN => n13057);
   U18557 : XNOR2_X1 port map( A => n13055, B => n3385, ZN => n13056);
   U18558 : XNOR2_X1 port map( A => n13057, B => n13056, ZN => n13058);
   U18559 : XNOR2_X1 port map( A => n13059, B => n13058, ZN => n13824);
   U18560 : XNOR2_X1 port map( A => n13325, B => n13503, ZN => n13065);
   U18561 : XNOR2_X1 port map( A => n13061, B => n13075, ZN => n13063);
   U18562 : XNOR2_X1 port map( A => n13209, B => n26680, ZN => n13062);
   U18563 : XNOR2_X1 port map( A => n13063, B => n13062, ZN => n13064);
   U18564 : INV_X1 port map( A => n13369, ZN => n13066);
   U18565 : XNOR2_X1 port map( A => n13066, B => n13067, ZN => n13068);
   U18566 : XNOR2_X1 port map( A => n13328, B => n13068, ZN => n13072);
   U18567 : XNOR2_X1 port map( A => n429, B => n25992, ZN => n13070);
   U18568 : XNOR2_X1 port map( A => n13479, B => n13070, ZN => n13071);
   U18569 : OAI211_X1 port map( C1 => n14351, C2 => n13826, A => n4893, B => 
                           n14354, ZN => n13073);
   U18570 : INV_X1 port map( A => n13073, ZN => n13074);
   U18571 : AOI21_X2 port map( B1 => n14015, B2 => n14350, A => n13074, ZN => 
                           n15077);
   U18572 : XNOR2_X1 port map( A => n13298, B => n13075, ZN => n13077);
   U18573 : XNOR2_X1 port map( A => n13208, B => n3644, ZN => n13076);
   U18574 : XNOR2_X1 port map( A => n13077, B => n13076, ZN => n13079);
   U18575 : XNOR2_X1 port map( A => n13224, B => n13322, ZN => n13078);
   U18576 : XNOR2_X1 port map( A => n13078, B => n13079, ZN => n14342);
   U18577 : XNOR2_X1 port map( A => n13166, B => n13080, ZN => n13092);
   U18578 : NAND2_X1 port map( A1 => n13082, A2 => n13081, ZN => n13089);
   U18579 : NAND2_X1 port map( A1 => n13087, A2 => n13083, ZN => n13085);
   U18580 : OAI211_X1 port map( C1 => n13087, C2 => n13086, A => n13085, B => 
                           n13084, ZN => n13088);
   U18581 : NAND2_X1 port map( A1 => n13089, A2 => n13088, ZN => n13090);
   U18582 : XNOR2_X1 port map( A => n13090, B => n2541, ZN => n13091);
   U18583 : XNOR2_X1 port map( A => n13092, B => n13091, ZN => n13093);
   U18584 : INV_X1 port map( A => n13095, ZN => n13354);
   U18585 : XNOR2_X1 port map( A => n13354, B => n13096, ZN => n13100);
   U18586 : XNOR2_X1 port map( A => n13179, B => n13285, ZN => n13099);
   U18587 : XNOR2_X1 port map( A => n13097, B => n1911, ZN => n13098);
   U18589 : INV_X1 port map( A => n13101, ZN => n13102);
   U18590 : XNOR2_X1 port map( A => n28603, B => n13102, ZN => n13103);
   U18591 : XNOR2_X1 port map( A => n13103, B => n13347, ZN => n13107);
   U18592 : XNOR2_X1 port map( A => n13104, B => n21865, ZN => n13105);
   U18593 : XNOR2_X1 port map( A => n13243, B => n13105, ZN => n13106);
   U18594 : XNOR2_X1 port map( A => n13107, B => n13106, ZN => n13842);
   U18595 : XNOR2_X1 port map( A => n13338, B => n13236, ZN => n13111);
   U18596 : INV_X1 port map( A => n13190, ZN => n13108);
   U18597 : XNOR2_X1 port map( A => n13108, B => n13109, ZN => n13110);
   U18598 : XNOR2_X1 port map( A => n13111, B => n13110, ZN => n13117);
   U18599 : INV_X1 port map( A => n13112, ZN => n13115);
   U18600 : XNOR2_X1 port map( A => n13113, B => n2510, ZN => n13114);
   U18601 : XNOR2_X1 port map( A => n13115, B => n13114, ZN => n13116);
   U18602 : XNOR2_X1 port map( A => n13116, B => n13117, ZN => n14010);
   U18603 : XNOR2_X1 port map( A => n429, B => n13533, ZN => n13120);
   U18604 : XNOR2_X1 port map( A => n13118, B => n2404, ZN => n13119);
   U18605 : XNOR2_X1 port map( A => n13120, B => n13119, ZN => n13124);
   U18606 : XNOR2_X1 port map( A => n13272, B => n13121, ZN => n13122);
   U18607 : XNOR2_X1 port map( A => n13122, B => n13332, ZN => n13123);
   U18608 : INV_X1 port map( A => n14342, ZN => n14135);
   U18609 : INV_X1 port map( A => n14131, ZN => n14343);
   U18610 : NAND2_X1 port map( A1 => n14135, A2 => n14343, ZN => n13125);
   U18611 : MUX2_X1 port map( A => n14948, B => n15077, S => n15073, Z => 
                           n13126);
   U18612 : INV_X1 port map( A => n14874, ZN => n14572);
   U18613 : NAND2_X1 port map( A1 => n13126, A2 => n14572, ZN => n13127);
   U18614 : INV_X1 port map( A => n14948, ZN => n15072);
   U18615 : XNOR2_X1 port map( A => n16606, B => n16476, ZN => n13129);
   U18616 : XNOR2_X1 port map( A => n13130, B => n13129, ZN => n13605);
   U18617 : XNOR2_X1 port map( A => n13539, B => n29494, ZN => n13132);
   U18618 : XNOR2_X1 port map( A => n13131, B => n13132, ZN => n13135);
   U18619 : XNOR2_X1 port map( A => n13133, B => n2973, ZN => n13134);
   U18620 : XNOR2_X1 port map( A => n1906, B => n13136, ZN => n13139);
   U18621 : XNOR2_X1 port map( A => n13137, B => n27105, ZN => n13138);
   U18622 : XNOR2_X1 port map( A => n13139, B => n13138, ZN => n13143);
   U18623 : XNOR2_X1 port map( A => n13140, B => n13141, ZN => n13142);
   U18624 : XNOR2_X1 port map( A => n13143, B => n13142, ZN => n14061);
   U18625 : XNOR2_X1 port map( A => n13144, B => n26665, ZN => n13145);
   U18626 : XNOR2_X1 port map( A => n13145, B => n13394, ZN => n13149);
   U18627 : XNOR2_X1 port map( A => n13147, B => n13146, ZN => n13148);
   U18628 : MUX2_X1 port map( A => n14325, B => n14064, S => n14327, Z => 
                           n13165);
   U18629 : XNOR2_X1 port map( A => n13487, B => n13389, ZN => n13154);
   U18630 : XNOR2_X1 port map( A => n13150, B => n27422, ZN => n13151);
   U18631 : XNOR2_X1 port map( A => n13152, B => n13151, ZN => n13153);
   U18632 : XNOR2_X1 port map( A => n13154, B => n13153, ZN => n13653);
   U18633 : XNOR2_X1 port map( A => n13362, B => n13155, ZN => n13158);
   U18634 : XNOR2_X1 port map( A => n13337, B => n3598, ZN => n13156);
   U18635 : XNOR2_X1 port map( A => n13509, B => n13156, ZN => n13157);
   U18636 : XNOR2_X1 port map( A => n13157, B => n13158, ZN => n13652);
   U18637 : XNOR2_X1 port map( A => n13474, B => n13379, ZN => n13163);
   U18638 : XNOR2_X1 port map( A => n13159, B => n13380, ZN => n13161);
   U18639 : XNOR2_X1 port map( A => n12593, B => n3686, ZN => n13160);
   U18640 : XNOR2_X1 port map( A => n13161, B => n13160, ZN => n13162);
   U18641 : XNOR2_X2 port map( A => n13163, B => n13162, ZN => n14328);
   U18642 : INV_X1 port map( A => n15692, ZN => n15084);
   U18643 : XNOR2_X1 port map( A => n13166, B => n13167, ZN => n13169);
   U18644 : XNOR2_X1 port map( A => n13169, B => n13168, ZN => n13174);
   U18645 : XNOR2_X1 port map( A => n13170, B => n13171, ZN => n13398);
   U18646 : XNOR2_X1 port map( A => n13218, B => n3336, ZN => n13172);
   U18647 : XNOR2_X1 port map( A => n13172, B => n13398, ZN => n13173);
   U18648 : XNOR2_X1 port map( A => n13174, B => n13173, ZN => n14029);
   U18649 : XNOR2_X1 port map( A => n13567, B => n3321, ZN => n13176);
   U18650 : XNOR2_X1 port map( A => n13177, B => n13176, ZN => n13183);
   U18651 : XNOR2_X1 port map( A => n13178, B => n13179, ZN => n13181);
   U18652 : XNOR2_X1 port map( A => n13181, B => n13180, ZN => n13182);
   U18653 : XNOR2_X1 port map( A => n13370, B => n13414, ZN => n13184);
   U18654 : XNOR2_X1 port map( A => n13535, B => n13184, ZN => n13188);
   U18655 : XNOR2_X1 port map( A => n13369, B => n13420, ZN => n13186);
   U18656 : XNOR2_X1 port map( A => n13533, B => n3191, ZN => n13185);
   U18657 : XNOR2_X1 port map( A => n13186, B => n13185, ZN => n13187);
   U18659 : MUX2_X1 port map( A => n14029, B => n29107, S => n14031, Z => 
                           n13217);
   U18660 : XNOR2_X1 port map( A => n13360, B => n730, ZN => n13189);
   U18661 : XNOR2_X1 port map( A => n13189, B => n13434, ZN => n13194);
   U18662 : XNOR2_X1 port map( A => n13190, B => n13191, ZN => n13546);
   U18663 : XNOR2_X1 port map( A => n13192, B => n13546, ZN => n13193);
   U18664 : XNOR2_X1 port map( A => n13553, B => n13195, ZN => n13196);
   U18665 : XNOR2_X1 port map( A => n13197, B => n13196, ZN => n13201);
   U18666 : XNOR2_X1 port map( A => n13104, B => n1246, ZN => n13199);
   U18667 : XNOR2_X1 port map( A => n13244, B => n13262, ZN => n13198);
   U18668 : XNOR2_X1 port map( A => n13199, B => n13198, ZN => n13200);
   U18669 : XNOR2_X1 port map( A => n13201, B => n13200, ZN => n13917);
   U18670 : NAND2_X1 port map( A1 => n13917, A2 => n13793, ZN => n13215);
   U18671 : XNOR2_X1 port map( A => n13540, B => n13457, ZN => n13213);
   U18672 : NAND2_X1 port map( A1 => n13206, A2 => n13202, ZN => n13204);
   U18673 : OAI211_X1 port map( C1 => n13206, C2 => n13205, A => n13204, B => 
                           n13203, ZN => n13207);
   U18674 : XNOR2_X1 port map( A => n13208, B => n13207, ZN => n13211);
   U18675 : XNOR2_X1 port map( A => n13209, B => n3770, ZN => n13210);
   U18676 : XNOR2_X1 port map( A => n13211, B => n13210, ZN => n13212);
   U18677 : XNOR2_X2 port map( A => n13213, B => n13212, ZN => n14030);
   U18678 : NAND2_X1 port map( A1 => n14030, A2 => n29107, ZN => n13214);
   U18679 : MUX2_X1 port map( A => n13215, B => n13214, S => n14029, Z => 
                           n13216);
   U18680 : XNOR2_X1 port map( A => n13223, B => n13224, ZN => n13225);
   U18681 : NAND2_X1 port map( A1 => n14045, A2 => n14043, ZN => n13578);
   U18682 : INV_X1 port map( A => n13578, ZN => n13256);
   U18683 : XNOR2_X1 port map( A => n13227, B => n13226, ZN => n13228);
   U18684 : XNOR2_X1 port map( A => n13229, B => n13228, ZN => n13235);
   U18685 : XNOR2_X1 port map( A => n13230, B => n13231, ZN => n13233);
   U18686 : XNOR2_X1 port map( A => n13450, B => n2986, ZN => n13232);
   U18687 : XNOR2_X1 port map( A => n13233, B => n13232, ZN => n13234);
   U18688 : XNOR2_X2 port map( A => n13235, B => n13234, ZN => n14051);
   U18689 : NAND2_X1 port map( A1 => n14045, A2 => n14051, ZN => n13909);
   U18690 : XNOR2_X1 port map( A => n13432, B => n13236, ZN => n13238);
   U18691 : XNOR2_X1 port map( A => n13238, B => n13237, ZN => n13242);
   U18692 : XNOR2_X1 port map( A => n13240, B => n13239, ZN => n13241);
   U18693 : XNOR2_X1 port map( A => n13244, B => n13245, ZN => n13430);
   U18694 : NOR2_X1 port map( A1 => n14046, A2 => n14044, ZN => n13255);
   U18695 : XNOR2_X1 port map( A => n13248, B => n13247, ZN => n13253);
   U18696 : XNOR2_X1 port map( A => n13249, B => n13331, ZN => n13251);
   U18697 : XNOR2_X1 port map( A => n13420, B => n2523, ZN => n13250);
   U18698 : XNOR2_X1 port map( A => n13251, B => n13250, ZN => n13252);
   U18699 : NAND2_X1 port map( A1 => n1896, A2 => n14043, ZN => n13254);
   U18700 : AOI21_X1 port map( B1 => n14309, B2 => n14317, A => n14318, ZN => 
                           n13259);
   U18701 : NOR2_X1 port map( A1 => n14320, A2 => n13884, ZN => n13258);
   U18702 : XNOR2_X1 port map( A => n28603, B => n13260, ZN => n13264);
   U18703 : XNOR2_X1 port map( A => n13263, B => n13262, ZN => n13390);
   U18704 : XNOR2_X1 port map( A => n13390, B => n13264, ZN => n13268);
   U18705 : XNOR2_X1 port map( A => n13265, B => n27956, ZN => n13266);
   U18706 : XNOR2_X1 port map( A => n13425, B => n13266, ZN => n13267);
   U18707 : XNOR2_X1 port map( A => n13270, B => n1062, ZN => n13271);
   U18708 : XNOR2_X1 port map( A => n13412, B => n13271, ZN => n13276);
   U18709 : XNOR2_X1 port map( A => n13272, B => n13273, ZN => n13481);
   U18710 : XNOR2_X1 port map( A => n13481, B => n13274, ZN => n13275);
   U18711 : XNOR2_X1 port map( A => n13441, B => n13277, ZN => n13282);
   U18712 : XNOR2_X1 port map( A => n13278, B => n2411, ZN => n13279);
   U18713 : XNOR2_X1 port map( A => n13280, B => n13279, ZN => n13281);
   U18714 : XNOR2_X1 port map( A => n13283, B => n13284, ZN => n13289);
   U18715 : XNOR2_X1 port map( A => n13285, B => n1927, ZN => n13286);
   U18716 : XNOR2_X1 port map( A => n13287, B => n13286, ZN => n13288);
   U18718 : XNOR2_X1 port map( A => n13438, B => n13290, ZN => n13295);
   U18719 : XNOR2_X1 port map( A => n13291, B => n3244, ZN => n13292);
   U18720 : XNOR2_X1 port map( A => n13293, B => n13292, ZN => n13294);
   U18721 : XNOR2_X1 port map( A => n13294, B => n13295, ZN => n13646);
   U18722 : INV_X1 port map( A => n14053, ZN => n14303);
   U18723 : NAND3_X1 port map( A1 => n29611, A2 => n13646, A3 => n14303, ZN => 
                           n13304);
   U18724 : INV_X1 port map( A => n14301, ZN => n14054);
   U18725 : XNOR2_X1 port map( A => n13402, B => n13296, ZN => n13302);
   U18726 : XNOR2_X1 port map( A => n13297, B => n13298, ZN => n13300);
   U18727 : XNOR2_X1 port map( A => n13543, B => n1193, ZN => n13299);
   U18728 : XNOR2_X1 port map( A => n13300, B => n13299, ZN => n13301);
   U18729 : XNOR2_X1 port map( A => n13302, B => n13301, ZN => n14302);
   U18730 : NAND3_X1 port map( A1 => n14054, A2 => n14302, A3 => n14304, ZN => 
                           n13303);
   U18731 : NAND3_X1 port map( A1 => n14563, A2 => n15690, A3 => n15691, ZN => 
                           n13305);
   U18732 : INV_X1 port map( A => n15690, ZN => n15087);
   U18733 : INV_X1 port map( A => n14563, ZN => n15088);
   U18734 : NOR2_X1 port map( A1 => n13803, A2 => n13699, ZN => n13310);
   U18736 : OAI21_X1 port map( B1 => n14293, B2 => n13306, A => n14294, ZN => 
                           n13307);
   U18737 : NAND2_X1 port map( A1 => n14298, A2 => n13307, ZN => n13308);
   U18738 : INV_X1 port map( A => n15083, ZN => n15689);
   U18739 : NAND2_X1 port map( A1 => n15088, A2 => n15689, ZN => n13311);
   U18740 : AOI21_X1 port map( B1 => n14878, B2 => n13311, A => n15692, ZN => 
                           n13312);
   U18741 : INV_X1 port map( A => n13314, ZN => n13317);
   U18742 : INV_X1 port map( A => n13315, ZN => n13316);
   U18743 : XNOR2_X1 port map( A => n13317, B => n13316, ZN => n13321);
   U18744 : XNOR2_X1 port map( A => n13525, B => n4029, ZN => n13319);
   U18745 : XNOR2_X1 port map( A => n13319, B => n13318, ZN => n13320);
   U18746 : XNOR2_X1 port map( A => n13538, B => n3003, ZN => n13323);
   U18747 : XNOR2_X1 port map( A => n13322, B => n13323, ZN => n13327);
   U18748 : XNOR2_X1 port map( A => n13325, B => n13324, ZN => n13326);
   U18750 : INV_X1 port map( A => n13328, ZN => n13330);
   U18751 : XNOR2_X1 port map( A => n13329, B => n13330, ZN => n13335);
   U18752 : XNOR2_X1 port map( A => n13331, B => n3062, ZN => n13333);
   U18753 : XNOR2_X1 port map( A => n13332, B => n13333, ZN => n13334);
   U18754 : XNOR2_X1 port map( A => n13335, B => n13334, ZN => n13913);
   U18755 : INV_X1 port map( A => n13913, ZN => n13729);
   U18756 : NOR2_X1 port map( A1 => n6351, A2 => n13729, ZN => n13336);
   U18757 : XNOR2_X1 port map( A => n13338, B => n13337, ZN => n13339);
   U18758 : XNOR2_X1 port map( A => n13340, B => n13339, ZN => n13345);
   U18759 : XNOR2_X1 port map( A => n13341, B => n2995, ZN => n13343);
   U18760 : XNOR2_X1 port map( A => n13343, B => n13342, ZN => n13344);
   U18762 : XNOR2_X1 port map( A => n13346, B => n13347, ZN => n13352);
   U18763 : XNOR2_X1 port map( A => n13348, B => n2961, ZN => n13349);
   U18764 : XNOR2_X1 port map( A => n13350, B => n13349, ZN => n13351);
   U18765 : XNOR2_X1 port map( A => n13352, B => n13351, ZN => n13583);
   U18766 : MUX2_X1 port map( A => n13912, B => n13583, S => n13729, Z => 
                           n13358);
   U18767 : XNOR2_X1 port map( A => n13354, B => n13353, ZN => n13357);
   U18768 : XNOR2_X1 port map( A => n13562, B => n2476, ZN => n13355);
   U18769 : XNOR2_X1 port map( A => n13360, B => n13359, ZN => n13361);
   U18770 : XNOR2_X1 port map( A => n13362, B => n13361, ZN => n13368);
   U18771 : INV_X1 port map( A => n13363, ZN => n13366);
   U18772 : XNOR2_X1 port map( A => n13364, B => n891, ZN => n13365);
   U18773 : XNOR2_X1 port map( A => n13366, B => n13365, ZN => n13367);
   U18774 : XNOR2_X1 port map( A => n13369, B => n13370, ZN => n13373);
   U18775 : XNOR2_X1 port map( A => n13371, B => n26825, ZN => n13372);
   U18776 : XNOR2_X1 port map( A => n13373, B => n13372, ZN => n13377);
   U18777 : XNOR2_X1 port map( A => n13374, B => n13375, ZN => n13376);
   U18778 : NAND2_X1 port map( A1 => n13716, A2 => n14016, ZN => n14142);
   U18779 : XNOR2_X1 port map( A => n13378, B => n13379, ZN => n13385);
   U18780 : XNOR2_X1 port map( A => n13381, B => n1172, ZN => n13382);
   U18781 : XNOR2_X1 port map( A => n13383, B => n13382, ZN => n13384);
   U18782 : XNOR2_X2 port map( A => n13385, B => n13384, ZN => n14144);
   U18783 : INV_X1 port map( A => n14144, ZN => n13900);
   U18784 : XNOR2_X1 port map( A => n13386, B => n2477, ZN => n13387);
   U18785 : XNOR2_X1 port map( A => n13388, B => n13387, ZN => n13392);
   U18786 : XNOR2_X1 port map( A => n13390, B => n13389, ZN => n13391);
   U18787 : XNOR2_X1 port map( A => n13391, B => n13392, ZN => n13902);
   U18788 : INV_X1 port map( A => n13393, ZN => n13395);
   U18789 : XNOR2_X1 port map( A => n13395, B => n13394, ZN => n13399);
   U18790 : XNOR2_X1 port map( A => n13396, B => n2403, ZN => n13397);
   U18791 : XNOR2_X1 port map( A => n13461, B => n27894, ZN => n13400);
   U18792 : XNOR2_X1 port map( A => n13400, B => n29495, ZN => n13403);
   U18793 : XNOR2_X1 port map( A => n13403, B => n13402, ZN => n13409);
   U18794 : XNOR2_X1 port map( A => n13405, B => n13404, ZN => n13407);
   U18795 : XNOR2_X1 port map( A => n13406, B => n13407, ZN => n13408);
   U18796 : INV_X1 port map( A => n13412, ZN => n13417);
   U18797 : XNOR2_X1 port map( A => n13413, B => n2509, ZN => n13415);
   U18798 : XNOR2_X1 port map( A => n13415, B => n13414, ZN => n13416);
   U18799 : XNOR2_X1 port map( A => n13417, B => n13416, ZN => n13424);
   U18800 : INV_X1 port map( A => n13418, ZN => n13422);
   U18801 : XNOR2_X1 port map( A => n13419, B => n13420, ZN => n13421);
   U18802 : XNOR2_X1 port map( A => n13422, B => n13421, ZN => n13423);
   U18803 : INV_X1 port map( A => n13425, ZN => n13427);
   U18804 : XNOR2_X1 port map( A => n13428, B => n3607, ZN => n13429);
   U18805 : XNOR2_X1 port map( A => n13430, B => n13429, ZN => n13431);
   U18806 : XNOR2_X1 port map( A => n13432, B => n13433, ZN => n13435);
   U18807 : XNOR2_X1 port map( A => n13434, B => n13435, ZN => n13439);
   U18808 : INV_X1 port map( A => n3386, ZN => n19658);
   U18809 : XNOR2_X1 port map( A => n13436, B => n19658, ZN => n13437);
   U18810 : NOR2_X1 port map( A1 => n13440, A2 => n13726, ZN => n13464);
   U18811 : INV_X1 port map( A => n13441, ZN => n13443);
   U18812 : XNOR2_X1 port map( A => n13444, B => n3650, ZN => n13446);
   U18813 : XNOR2_X1 port map( A => n13448, B => n13447, ZN => n13449);
   U18814 : XNOR2_X1 port map( A => n28587, B => n13450, ZN => n13453);
   U18815 : INV_X1 port map( A => n1187, ZN => n27534);
   U18816 : XNOR2_X1 port map( A => n13451, B => n27534, ZN => n13452);
   U18817 : XNOR2_X1 port map( A => n13453, B => n13452, ZN => n13454);
   U18818 : XNOR2_X1 port map( A => n13455, B => n13454, ZN => n13595);
   U18819 : XNOR2_X1 port map( A => n13461, B => n2577, ZN => n13462);
   U18821 : NAND2_X1 port map( A1 => n14881, A2 => n388, ZN => n13519);
   U18822 : NAND2_X1 port map( A1 => n14030, A2 => n14031, ZN => n13465);
   U18823 : OAI21_X1 port map( B1 => n14029, B2 => n14030, A => n13465, ZN => 
                           n13467);
   U18824 : INV_X1 port map( A => n14030, ZN => n13796);
   U18825 : INV_X1 port map( A => n14031, ZN => n13916);
   U18826 : INV_X1 port map( A => n13793, ZN => n14032);
   U18827 : NAND2_X1 port map( A1 => n14031, A2 => n14032, ZN => n13466);
   U18828 : INV_X1 port map( A => n14046, ZN => n13662);
   U18829 : NAND3_X1 port map( A1 => n13662, A2 => n14051, A3 => n13661, ZN => 
                           n13468);
   U18830 : NAND3_X1 port map( A1 => n14043, A2 => n14044, A3 => n14051, ZN => 
                           n13469);
   U18831 : INV_X1 port map( A => n14045, ZN => n13907);
   U18832 : XNOR2_X1 port map( A => n13472, B => n13471, ZN => n13477);
   U18833 : XNOR2_X1 port map( A => n13473, B => n3722, ZN => n13475);
   U18834 : XNOR2_X1 port map( A => n13474, B => n13475, ZN => n13476);
   U18836 : XNOR2_X1 port map( A => n29640, B => n13478, ZN => n13480);
   U18837 : XNOR2_X1 port map( A => n13479, B => n13480, ZN => n13483);
   U18838 : INV_X1 port map( A => n3067, ZN => n27515);
   U18839 : XNOR2_X1 port map( A => n13485, B => n13484, ZN => n13486);
   U18840 : XNOR2_X1 port map( A => n13487, B => n13486, ZN => n13492);
   U18841 : XNOR2_X1 port map( A => n13488, B => n1247, ZN => n13489);
   U18842 : XNOR2_X1 port map( A => n13490, B => n13489, ZN => n13491);
   U18843 : XNOR2_X1 port map( A => n13493, B => n3256, ZN => n13495);
   U18844 : XNOR2_X1 port map( A => n13495, B => n13494, ZN => n13499);
   U18845 : XNOR2_X1 port map( A => n13496, B => n13497, ZN => n13498);
   U18846 : NAND2_X1 port map( A1 => n13589, A2 => n13719, ZN => n14000);
   U18847 : INV_X1 port map( A => n13501, ZN => n13502);
   U18848 : XNOR2_X1 port map( A => n13502, B => n13503, ZN => n13508);
   U18849 : XNOR2_X1 port map( A => n13504, B => n28693, ZN => n13506);
   U18850 : XNOR2_X1 port map( A => n13505, B => n13506, ZN => n13507);
   U18851 : XNOR2_X1 port map( A => n13509, B => n13510, ZN => n13515);
   U18852 : XNOR2_X1 port map( A => n13511, B => n26032, ZN => n13512);
   U18853 : XNOR2_X1 port map( A => n13513, B => n13512, ZN => n13514);
   U18855 : INV_X1 port map( A => n14974, ZN => n13517);
   U18856 : NAND2_X1 port map( A1 => n13517, A2 => n14972, ZN => n13518);
   U18857 : XNOR2_X1 port map( A => n16346, B => n16312, ZN => n13603);
   U18858 : XNOR2_X1 port map( A => n13522, B => n13521, ZN => n13529);
   U18859 : XNOR2_X1 port map( A => n13524, B => n13523, ZN => n13527);
   U18860 : XNOR2_X1 port map( A => n13525, B => n3673, ZN => n13526);
   U18861 : XNOR2_X1 port map( A => n13527, B => n13526, ZN => n13528);
   U18862 : INV_X1 port map( A => n14007, ZN => n14386);
   U18863 : INV_X1 port map( A => n13530, ZN => n13531);
   U18864 : XNOR2_X1 port map( A => n13531, B => n13532, ZN => n13537);
   U18865 : XNOR2_X1 port map( A => n13533, B => n1079, ZN => n13534);
   U18866 : XNOR2_X1 port map( A => n13535, B => n13534, ZN => n13536);
   U18867 : XNOR2_X1 port map( A => n13537, B => n13536, ZN => n13837);
   U18868 : XNOR2_X1 port map( A => n13538, B => n13539, ZN => n13541);
   U18869 : XNOR2_X1 port map( A => n13540, B => n13541, ZN => n13544);
   U18870 : XNOR2_X1 port map( A => n13546, B => n13545, ZN => n13551);
   U18871 : XNOR2_X1 port map( A => n13547, B => n3635, ZN => n13548);
   U18872 : XNOR2_X1 port map( A => n13549, B => n13548, ZN => n13550);
   U18873 : XNOR2_X1 port map( A => n13551, B => n13550, ZN => n14381);
   U18874 : AOI22_X1 port map( A1 => n14386, A2 => n14150, B1 => n13572, B2 => 
                           n14381, ZN => n13575);
   U18875 : XNOR2_X1 port map( A => n13552, B => n13553, ZN => n13555);
   U18876 : XNOR2_X1 port map( A => n13554, B => n13555, ZN => n13561);
   U18877 : XNOR2_X1 port map( A => n13104, B => n1919, ZN => n13559);
   U18878 : XNOR2_X1 port map( A => n13557, B => n13556, ZN => n13558);
   U18879 : XNOR2_X1 port map( A => n13559, B => n13558, ZN => n13560);
   U18880 : XNOR2_X1 port map( A => n13563, B => n13562, ZN => n13564);
   U18881 : XNOR2_X1 port map( A => n13565, B => n13564, ZN => n13571);
   U18882 : XNOR2_X1 port map( A => n13567, B => n3081, ZN => n13568);
   U18883 : XNOR2_X1 port map( A => n13569, B => n13568, ZN => n13570);
   U18884 : NOR2_X1 port map( A1 => n14007, A2 => n14381, ZN => n13734);
   U18885 : NOR2_X1 port map( A1 => n13573, A2 => n13734, ZN => n13574);
   U18886 : NAND2_X1 port map( A1 => n14043, A2 => n13661, ZN => n13576);
   U18887 : INV_X1 port map( A => n14043, ZN => n13906);
   U18888 : NAND2_X1 port map( A1 => n14047, A2 => n13906, ZN => n13577);
   U18889 : NAND3_X1 port map( A1 => n13578, A2 => n5731, A3 => n13577, ZN => 
                           n13579);
   U18890 : NOR2_X1 port map( A1 => n13716, A2 => n29589, ZN => n13581);
   U18891 : NAND2_X1 port map( A1 => n13912, A2 => n13583, ZN => n13582);
   U18892 : NAND2_X1 port map( A1 => n6351, A2 => n13914, ZN => n13585);
   U18893 : INV_X1 port map( A => n13583, ZN => n13910);
   U18894 : OAI211_X1 port map( C1 => n13730, C2 => n13914, A => n5847, B => 
                           n13910, ZN => n13584);
   U18895 : MUX2_X1 port map( A => n13589, B => n13587, S => n13719, Z => 
                           n13588);
   U18896 : NOR2_X1 port map( A1 => n13588, A2 => n14039, ZN => n13590);
   U18897 : NAND2_X1 port map( A1 => n13719, A2 => n28569, ZN => n13999);
   U18898 : NAND2_X1 port map( A1 => n13592, A2 => n28196, ZN => n13600);
   U18899 : NOR2_X1 port map( A1 => n13593, A2 => n13726, ZN => n13597);
   U18900 : NOR2_X1 port map( A1 => n28518, A2 => n13638, ZN => n14895);
   U18901 : INV_X1 port map( A => n14895, ZN => n13598);
   U18902 : NAND2_X1 port map( A1 => n13598, A2 => n15400, ZN => n13599);
   U18903 : NAND2_X1 port map( A1 => n13600, A2 => n13599, ZN => n13601);
   U18904 : XNOR2_X1 port map( A => n13603, B => n15777, ZN => n13604);
   U18905 : NOR2_X1 port map( A1 => n14231, A2 => n14107, ZN => n13607);
   U18906 : MUX2_X1 port map( A => n6956, B => n13607, S => n14593, Z => n13610
                           );
   U18907 : AOI21_X1 port map( B1 => n14235, B2 => n13608, A => n14230, ZN => 
                           n13609);
   U18908 : NOR2_X2 port map( A1 => n13610, A2 => n13609, ZN => n15004);
   U18909 : NAND2_X1 port map( A1 => n1743, A2 => n14262, ZN => n13763);
   U18910 : INV_X1 port map( A => n13763, ZN => n13612);
   U18912 : NAND2_X1 port map( A1 => n14362, A2 => n28507, ZN => n13617);
   U18913 : INV_X1 port map( A => n13832, ZN => n14271);
   U18914 : NAND3_X1 port map( A1 => n14272, A2 => n14271, A3 => n14278, ZN => 
                           n13616);
   U18916 : NAND2_X1 port map( A1 => n15001, A2 => n15127, ZN => n14688);
   U18917 : INV_X1 port map( A => n13770, ZN => n13620);
   U18920 : INV_X1 port map( A => n14091, ZN => n14369);
   U18921 : NAND2_X1 port map( A1 => n14091, A2 => n14365, ZN => n14118);
   U18922 : NOR2_X1 port map( A1 => n14118, A2 => n14366, ZN => n13624);
   U18923 : AOI21_X2 port map( B1 => n13625, B2 => n1960, A => n13624, ZN => 
                           n15000);
   U18924 : NAND2_X1 port map( A1 => n14351, A2 => n4893, ZN => n13626);
   U18925 : NAND3_X1 port map( A1 => n13627, A2 => n13626, A3 => n13826, ZN => 
                           n13631);
   U18926 : INV_X1 port map( A => n14354, ZN => n14353);
   U18927 : NAND3_X1 port map( A1 => n13825, A2 => n4893, A3 => n14353, ZN => 
                           n13629);
   U18928 : NAND2_X1 port map( A1 => n14126, A2 => n14355, ZN => n13628);
   U18929 : NAND2_X1 port map( A1 => n13631, A2 => n13630, ZN => n15123);
   U18930 : INV_X1 port map( A => n15004, ZN => n15125);
   U18931 : NOR2_X1 port map( A1 => n15127, A2 => n15123, ZN => n13633);
   U18932 : AOI21_X1 port map( B1 => n14686, B2 => n15125, A => n13633, ZN => 
                           n13634);
   U18933 : OAI21_X1 port map( B1 => n14944, B2 => n13637, A => n13636, ZN => 
                           n14945);
   U18934 : INV_X1 port map( A => n13638, ZN => n15401);
   U18935 : NAND2_X1 port map( A1 => n14945, A2 => n15401, ZN => n13642);
   U18936 : OAI21_X1 port map( B1 => n14944, B2 => n14943, A => n13639, ZN => 
                           n13640);
   U18937 : NAND2_X1 port map( A1 => n13640, A2 => n28196, ZN => n13641);
   U18938 : NAND2_X1 port map( A1 => n5887, A2 => n13583, ZN => n13643);
   U18939 : AOI21_X2 port map( B1 => n13645, B2 => n13730, A => n13644, ZN => 
                           n15115);
   U18940 : NAND2_X1 port map( A1 => n14301, A2 => n14304, ZN => n13651);
   U18941 : INV_X1 port map( A => n13647, ZN => n13648);
   U18942 : NAND2_X1 port map( A1 => n13648, A2 => n14054, ZN => n13649);
   U18943 : INV_X1 port map( A => n13652, ZN => n14324);
   U18944 : INV_X1 port map( A => n13653, ZN => n14065);
   U18945 : INV_X1 port map( A => n14328, ZN => n13654);
   U18946 : NOR2_X1 port map( A1 => n14327, A2 => n13654, ZN => n13656);
   U18947 : OAI211_X1 port map( C1 => n29626, C2 => n14328, A => n13653, B => 
                           n14064, ZN => n13655);
   U18948 : NAND2_X1 port map( A1 => n13808, A2 => n13803, ZN => n13659);
   U18949 : INV_X1 port map( A => n14295, ZN => n13806);
   U18950 : NAND3_X1 port map( A1 => n14295, A2 => n14291, A3 => n14297, ZN => 
                           n13657);
   U18951 : OAI21_X1 port map( B1 => n15115, B2 => n1001, A => n13660, ZN => 
                           n14114);
   U18952 : NOR2_X1 port map( A1 => n14045, A2 => n13661, ZN => n13664);
   U18953 : NOR2_X1 port map( A1 => n1896, A2 => n14051, ZN => n13663);
   U18954 : MUX2_X1 port map( A => n13664, B => n13663, S => n13662, Z => 
                           n13665);
   U18955 : INV_X1 port map( A => n14514, ZN => n15116);
   U18956 : INV_X1 port map( A => n14029, ZN => n13921);
   U18957 : NAND2_X1 port map( A1 => n13916, A2 => n29107, ZN => n13666);
   U18958 : OR2_X1 port map( A1 => n13666, A2 => n14032, ZN => n13667);
   U18960 : XNOR2_X1 port map( A => n29319, B => n28557, ZN => n13669);
   U18961 : XNOR2_X1 port map( A => n13669, B => n13670, ZN => n13760);
   U18962 : INV_X1 port map( A => n14207, ZN => n14439);
   U18963 : NOR2_X1 port map( A1 => n14207, A2 => n1876, ZN => n13671);
   U18964 : INV_X1 port map( A => n13672, ZN => n13673);
   U18965 : OAI21_X1 port map( B1 => n14492, B2 => n14497, A => n13856, ZN => 
                           n13676);
   U18967 : NAND2_X1 port map( A1 => n14492, A2 => n29036, ZN => n13675);
   U18968 : NAND2_X1 port map( A1 => n15389, A2 => n15388, ZN => n14723);
   U18969 : INV_X1 port map( A => n14464, ZN => n13852);
   U18970 : INV_X1 port map( A => n13678, ZN => n14467);
   U18971 : NAND3_X1 port map( A1 => n14467, A2 => n13852, A3 => n4840, ZN => 
                           n13681);
   U18972 : NAND3_X1 port map( A1 => n14185, A2 => n13678, A3 => n14464, ZN => 
                           n13679);
   U18973 : NOR2_X1 port map( A1 => n12711, A2 => n14456, ZN => n13682);
   U18977 : NAND2_X1 port map( A1 => n14416, A2 => n14414, ZN => n13893);
   U18978 : INV_X1 port map( A => n14193, ZN => n13867);
   U18979 : NAND3_X1 port map( A1 => n28805, A2 => n14192, A3 => n13867, ZN => 
                           n13688);
   U18982 : INV_X1 port map( A => n14992, ZN => n15391);
   U18985 : MUX2_X1 port map( A => n29133, B => n14406, S => n14407, Z => 
                           n13693);
   U18986 : INV_X1 port map( A => n14333, ZN => n13692);
   U18987 : OAI21_X1 port map( B1 => n13653, B2 => n14061, A => n14324, ZN => 
                           n13694);
   U18989 : AOI21_X1 port map( B1 => n14291, B2 => n14293, A => n13697, ZN => 
                           n13698);
   U18990 : NAND2_X1 port map( A1 => n13698, A2 => n13702, ZN => n13701);
   U18991 : NOR2_X1 port map( A1 => n14292, A2 => n13699, ZN => n13807);
   U18992 : NAND2_X1 port map( A1 => n13807, A2 => n13803, ZN => n13700);
   U18993 : OAI211_X1 port map( C1 => n13702, C2 => n14294, A => n13701, B => 
                           n13700, ZN => n15137);
   U18994 : NAND2_X1 port map( A1 => n15248, A2 => n15137, ZN => n15247);
   U18995 : NOR2_X1 port map( A1 => n13872, A2 => n14429, ZN => n13706);
   U18996 : INV_X1 port map( A => n14426, ZN => n13873);
   U18998 : NAND2_X1 port map( A1 => n15250, A2 => n15137, ZN => n13710);
   U19000 : OAI21_X1 port map( B1 => n14398, B2 => n28804, A => n14402, ZN => 
                           n13707);
   U19001 : MUX2_X1 port map( A => n13710, B => n14733, S => n15246, Z => 
                           n13715);
   U19002 : NAND3_X1 port map( A1 => n14312, A2 => n13711, A3 => n14313, ZN => 
                           n13713);
   U19003 : NAND3_X1 port map( A1 => n15249, A2 => n15135, A3 => n15250, ZN => 
                           n13714);
   U19004 : XNOR2_X1 port map( A => n16160, B => n16126, ZN => n16418);
   U19005 : INV_X1 port map( A => n15372, ZN => n15374);
   U19006 : NAND3_X1 port map( A1 => n13726, A2 => n5404, A3 => n14146, ZN => 
                           n13727);
   U19008 : INV_X1 port map( A => n14010, ZN => n14344);
   U19009 : NAND2_X1 port map( A1 => n14346, A2 => n14132, ZN => n14134);
   U19011 : NOR2_X1 port map( A1 => n14344, A2 => n14345, ZN => n13728);
   U19012 : INV_X1 port map( A => n14380, ZN => n14385);
   U19013 : MUX2_X1 port map( A => n14007, B => n14385, S => n14150, Z => 
                           n13736);
   U19014 : INV_X1 port map( A => n13572, ZN => n13836);
   U19015 : NOR2_X1 port map( A1 => n13836, A2 => n14380, ZN => n13733);
   U19016 : AOI22_X1 port map( A1 => n13734, A2 => n14004, B1 => n13733, B2 => 
                           n14007, ZN => n13735);
   U19017 : NAND2_X1 port map( A1 => n28172, A2 => n14241, ZN => n13769);
   U19018 : NOR2_X1 port map( A1 => n15194, A2 => n14241, ZN => n15192);
   U19019 : NAND2_X1 port map( A1 => n15192, A2 => n29097, ZN => n13741);
   U19020 : OAI211_X1 port map( C1 => n29097, C2 => n14238, A => n15194, B => 
                           n13739, ZN => n13740);
   U19021 : INV_X1 port map( A => n15379, ZN => n15152);
   U19022 : NOR2_X1 port map( A1 => n14166, A2 => n14484, ZN => n13742);
   U19023 : INV_X1 port map( A => n14481, ZN => n14164);
   U19024 : INV_X1 port map( A => n15382, ZN => n13752);
   U19025 : OAI22_X1 port map( A1 => n13744, A2 => n14252, B1 => n14078, B2 => 
                           n13778, ZN => n14076);
   U19026 : INV_X1 port map( A => n14078, ZN => n14251);
   U19027 : NOR2_X1 port map( A1 => n14251, A2 => n14250, ZN => n13746);
   U19028 : INV_X1 port map( A => n15383, ZN => n15150);
   U19029 : NOR2_X1 port map( A1 => n14268, A2 => n14262, ZN => n13748);
   U19030 : MUX2_X1 port map( A => n13748, B => n13747, S => n14264, Z => 
                           n13751);
   U19031 : NAND2_X1 port map( A1 => n14261, A2 => n14259, ZN => n14266);
   U19032 : OAI21_X1 port map( B1 => n14264, B2 => n14266, A => n14098, ZN => 
                           n13750);
   U19033 : AOI21_X1 port map( B1 => n13752, B2 => n15150, A => n15151, ZN => 
                           n13758);
   U19034 : OAI22_X1 port map( A1 => n14177, A2 => n14452, B1 => n13753, B2 => 
                           n14178, ZN => n13850);
   U19035 : OAI22_X1 port map( A1 => n15155, A2 => n15379, B1 => n15151, B2 => 
                           n15383, ZN => n15381);
   U19036 : NAND2_X1 port map( A1 => n14475, A2 => n13936, ZN => n13756);
   U19037 : NOR2_X1 port map( A1 => n14480, A2 => n13936, ZN => n13757);
   U19038 : INV_X1 port map( A => n14986, ZN => n15384);
   U19039 : XNOR2_X1 port map( A => n16456, B => n16318, ZN => n16162);
   U19040 : XNOR2_X1 port map( A => n16162, B => n16418, ZN => n13759);
   U19041 : XNOR2_X1 port map( A => n13760, B => n13759, ZN => n17716);
   U19042 : INV_X1 port map( A => n17716, ZN => n17720);
   U19043 : MUX2_X1 port map( A => n13762, B => n13761, S => n14099, Z => 
                           n13764);
   U19045 : NAND3_X1 port map( A1 => n29306, A2 => n14481, A3 => n14486, ZN => 
                           n13765);
   U19046 : NAND2_X1 port map( A1 => n15201, A2 => n15207, ZN => n14968);
   U19047 : MUX2_X1 port map( A => n15195, B => n13943, S => n28172, Z => 
                           n13768);
   U19048 : AND3_X1 port map( A1 => n13767, A2 => n14174, A3 => n14241, ZN => 
                           n15193);
   U19049 : MUX2_X1 port map( A => n14285, B => n14083, S => n14287, Z => 
                           n13774);
   U19050 : NAND2_X1 port map( A1 => n14082, A2 => n14084, ZN => n13771);
   U19051 : AND2_X1 port map( A1 => n13771, A2 => n13770, ZN => n13773);
   U19052 : INV_X1 port map( A => n14286, ZN => n14081);
   U19053 : NOR2_X1 port map( A1 => n14287, A2 => n14081, ZN => n13772);
   U19054 : INV_X1 port map( A => n14963, ZN => n15209);
   U19055 : INV_X1 port map( A => n13775, ZN => n14077);
   U19056 : MUX2_X1 port map( A => n14252, B => n14077, S => n14078, Z => 
                           n13781);
   U19057 : INV_X1 port map( A => n13776, ZN => n14253);
   U19058 : NAND3_X1 port map( A1 => n13778, A2 => n14252, A3 => n14077, ZN => 
                           n13779);
   U19060 : INV_X1 port map( A => n15208, ZN => n13782);
   U19061 : INV_X1 port map( A => n15207, ZN => n15204);
   U19062 : NAND3_X1 port map( A1 => n15209, A2 => n13782, A3 => n15204, ZN => 
                           n13787);
   U19063 : NAND2_X1 port map( A1 => n14230, A2 => n14593, ZN => n13784);
   U19064 : OAI211_X1 port map( C1 => n14960, C2 => n15207, A => n13785, B => 
                           n15202, ZN => n13786);
   U19066 : INV_X1 port map( A => n14881, ZN => n14976);
   U19067 : NAND2_X1 port map( A1 => n14882, A2 => n13789, ZN => n14970);
   U19068 : OAI21_X1 port map( B1 => n14976, B2 => n14970, A => n13788, ZN => 
                           n13792);
   U19069 : NOR2_X1 port map( A1 => n13789, A2 => n14972, ZN => n13790);
   U19070 : XNOR2_X1 port map( A => n15070, B => n16284, ZN => n16171);
   U19071 : NAND2_X1 port map( A1 => n6066, A2 => n14032, ZN => n13797);
   U19072 : AOI21_X1 port map( B1 => n6066, B2 => n14031, A => n13793, ZN => 
                           n13795);
   U19074 : NOR2_X1 port map( A1 => n14324, A2 => n14328, ZN => n13798);
   U19075 : NAND2_X1 port map( A1 => n14314, A2 => n14318, ZN => n13886);
   U19076 : NAND2_X1 port map( A1 => n13886, A2 => n14313, ZN => n13801);
   U19077 : AOI21_X1 port map( B1 => n14313, B2 => n560, A => n14314, ZN => 
                           n13800);
   U19078 : MUX2_X1 port map( A => n13805, B => n13804, S => n14294, Z => 
                           n13810);
   U19079 : AOI22_X1 port map( A1 => n13808, A2 => n14291, B1 => n13807, B2 => 
                           n13806, ZN => n13809);
   U19080 : NAND2_X1 port map( A1 => n14332, A2 => n14405, ZN => n13812);
   U19081 : OAI21_X1 port map( B1 => n14408, B2 => n13878, A => n13879, ZN => 
                           n13811);
   U19082 : OAI21_X1 port map( B1 => n13813, B2 => n13812, A => n13811, ZN => 
                           n13814);
   U19083 : NOR2_X1 port map( A1 => n15184, A2 => n14784, ZN => n15187);
   U19084 : NAND2_X1 port map( A1 => n28625, A2 => n14084, ZN => n14284);
   U19085 : OAI21_X1 port map( B1 => n14085, B2 => n14285, A => n561, ZN => 
                           n13821);
   U19086 : NAND2_X1 port map( A1 => n13821, A2 => n14082, ZN => n13823);
   U19087 : NAND3_X1 port map( A1 => n14286, A2 => n561, A3 => n14282, ZN => 
                           n13822);
   U19088 : NAND2_X1 port map( A1 => n14362, A2 => n13832, ZN => n14363);
   U19089 : INV_X1 port map( A => n14363, ZN => n13828);
   U19090 : NAND2_X1 port map( A1 => n13828, A2 => n13827, ZN => n13831);
   U19091 : INV_X1 port map( A => n14360, ZN => n14273);
   U19092 : NAND3_X1 port map( A1 => n14359, A2 => n14273, A3 => n28507, ZN => 
                           n13830);
   U19093 : NOR2_X1 port map( A1 => n308, A2 => n14091, ZN => n13834);
   U19095 : NAND2_X1 port map( A1 => n13836, A2 => n14380, ZN => n13840);
   U19096 : NAND3_X1 port map( A1 => n14006, A2 => n557, A3 => n14150, ZN => 
                           n13839);
   U19097 : OAI21_X1 port map( B1 => n13572, B2 => n14004, A => n556, ZN => 
                           n13838);
   U19098 : OAI21_X1 port map( B1 => n14797, B2 => n15460, A => n13841, ZN => 
                           n13846);
   U19099 : OAI21_X1 port map( B1 => n14135, B2 => n14346, A => n14343, ZN => 
                           n13843);
   U19100 : MUX2_X1 port map( A => n28803, B => n15180, S => n15175, Z => 
                           n13844);
   U19101 : XNOR2_X1 port map( A => n15738, B => n16366, ZN => n16044);
   U19102 : XNOR2_X1 port map( A => n16171, B => n16044, ZN => n13927);
   U19103 : AOI21_X1 port map( B1 => n14435, B2 => n14439, A => n14433, ZN => 
                           n13849);
   U19104 : OAI22_X1 port map( A1 => n14438, A2 => n14434, B1 => n14207, B2 => 
                           n14433, ZN => n14206);
   U19105 : NAND2_X1 port map( A1 => n14206, A2 => n14432, ZN => n13848);
   U19106 : NOR2_X1 port map( A1 => n15476, A2 => n15168, ZN => n13861);
   U19107 : NAND2_X1 port map( A1 => n13851, A2 => n14452, ZN => n14453);
   U19108 : NAND3_X1 port map( A1 => n14453, A2 => n13753, A3 => n14451, ZN => 
                           n14548);
   U19109 : OAI21_X1 port map( B1 => n14466, B2 => n4840, A => n14182, ZN => 
                           n14183);
   U19110 : NAND2_X1 port map( A1 => n13933, A2 => n14464, ZN => n13854);
   U19111 : NAND2_X1 port map( A1 => n14492, A2 => n14497, ZN => n14155);
   U19112 : NAND2_X1 port map( A1 => n14493, A2 => n13674, ZN => n13858);
   U19114 : NAND3_X1 port map( A1 => n14498, A2 => n14491, A3 => n14494, ZN => 
                           n13859);
   U19115 : OAI211_X1 port map( C1 => n29037, C2 => n14155, A => n13860, B => 
                           n13859, ZN => n15167);
   U19116 : INV_X1 port map( A => n15168, ZN => n14551);
   U19117 : NAND2_X1 port map( A1 => n13967, A2 => n14459, ZN => n13862);
   U19119 : INV_X1 port map( A => n15166, ZN => n15471);
   U19120 : NAND3_X1 port map( A1 => n14193, A2 => n14393, A3 => n14194, ZN => 
                           n13869);
   U19121 : OAI211_X1 port map( C1 => n13873, C2 => n13872, A => n13871, B => 
                           n28199, ZN => n13876);
   U19122 : NOR2_X1 port map( A1 => n15466, A2 => n4515, ZN => n13890);
   U19123 : MUX2_X1 port map( A => n13879, B => n13878, S => n14405, Z => 
                           n13880);
   U19124 : NAND3_X1 port map( A1 => n14332, A2 => n1830, A3 => n29133, ZN => 
                           n13881);
   U19125 : OAI21_X1 port map( B1 => n13884, B2 => n14312, A => n14318, ZN => 
                           n13885);
   U19126 : OR2_X1 port map( A1 => n560, A2 => n13886, ZN => n13887);
   U19129 : NAND3_X1 port map( A1 => n13891, A2 => n14216, A3 => n28647, ZN => 
                           n13892);
   U19130 : XNOR2_X1 port map( A => n16192, B => n16634, ZN => n16397);
   U19132 : INV_X1 port map( A => n14773, ZN => n14808);
   U19133 : NAND2_X1 port map( A1 => n14020, A2 => n13901, ZN => n13905);
   U19134 : NOR2_X1 port map( A1 => n14808, A2 => n14807, ZN => n14712);
   U19135 : OAI211_X1 port map( C1 => n14030, C2 => n14033, A => n13917, B => 
                           n13916, ZN => n13919);
   U19136 : NAND3_X1 port map( A1 => n6066, A2 => n14032, A3 => n29107, ZN => 
                           n13918);
   U19137 : OAI211_X1 port map( C1 => n13921, C2 => n29107, A => n13919, B => 
                           n13918, ZN => n14806);
   U19138 : INV_X1 port map( A => n14806, ZN => n14767);
   U19139 : NAND2_X1 port map( A1 => n14807, A2 => n28493, ZN => n13923);
   U19140 : INV_X1 port map( A => n14302, ZN => n14059);
   U19141 : AOI21_X1 port map( B1 => n14059, B2 => n5956, A => n29611, ZN => 
                           n14771);
   U19142 : MUX2_X1 port map( A => n14300, B => n14299, S => n28478, Z => 
                           n14770);
   U19143 : NAND2_X1 port map( A1 => n14302, A2 => n14303, ZN => n14769);
   U19144 : NAND3_X1 port map( A1 => n14810, A2 => n14807, A3 => n14713, ZN => 
                           n13925);
   U19145 : NAND2_X1 port map( A1 => n14176, A2 => n14452, ZN => n13928);
   U19146 : NAND2_X1 port map( A1 => n1320, A2 => n13928, ZN => n13929);
   U19147 : OAI21_X1 port map( B1 => n13930, B2 => n1320, A => n13929, ZN => 
                           n13931);
   U19149 : NAND2_X1 port map( A1 => n14249, A2 => n14250, ZN => n14237);
   U19150 : NAND2_X1 port map( A1 => n14251, A2 => n14077, ZN => n13938);
   U19151 : NAND2_X1 port map( A1 => n15438, A2 => n15300, ZN => n13941);
   U19152 : INV_X1 port map( A => n15438, ZN => n15302);
   U19153 : INV_X1 port map( A => n15018, ZN => n15437);
   U19154 : NOR2_X1 port map( A1 => n15444, A2 => n15437, ZN => n14667);
   U19155 : NAND2_X1 port map( A1 => n15303, A2 => n15302, ZN => n13949);
   U19156 : NOR2_X1 port map( A1 => n14193, A2 => n14192, ZN => n13952);
   U19158 : NAND2_X1 port map( A1 => n13956, A2 => n13955, ZN => n15015);
   U19159 : INV_X1 port map( A => n13957, ZN => n13958);
   U19160 : AOI21_X1 port map( B1 => n14438, B2 => n14432, A => n14437, ZN => 
                           n13960);
   U19161 : OAI21_X1 port map( B1 => n13963, B2 => n13962, A => n30, ZN => 
                           n13964);
   U19162 : OAI21_X2 port map( B1 => n13965, B2 => n14400, A => n13964, ZN => 
                           n15014);
   U19163 : INV_X1 port map( A => n14459, ZN => n13966);
   U19164 : NAND3_X1 port map( A1 => n14204, A2 => n14456, A3 => n13966, ZN => 
                           n13971);
   U19165 : AND2_X1 port map( A1 => n14455, A2 => n13967, ZN => n13968);
   U19166 : NAND2_X1 port map( A1 => n13968, A2 => n14200, ZN => n13970);
   U19167 : NAND4_X1 port map( A1 => n14463, A2 => n13971, A3 => n13970, A4 => 
                           n13969, ZN => n15013);
   U19168 : AOI21_X1 port map( B1 => n14155, B2 => n14494, A => n14491, ZN => 
                           n13975);
   U19169 : NAND2_X1 port map( A1 => n14493, A2 => n14491, ZN => n13972);
   U19170 : AOI21_X1 port map( B1 => n13973, B2 => n13972, A => n14497, ZN => 
                           n13974);
   U19171 : NAND2_X1 port map( A1 => n15447, A2 => n15321, ZN => n13976);
   U19172 : XNOR2_X1 port map( A => n16564, B => n16146, ZN => n16424);
   U19173 : NOR2_X1 port map( A1 => n15115, A2 => n15117, ZN => n14112);
   U19174 : INV_X1 port map( A => n14112, ZN => n13982);
   U19175 : INV_X1 port map( A => n14743, ZN => n15114);
   U19176 : OAI21_X1 port map( B1 => n15113, B2 => n1904, A => n14744, ZN => 
                           n13981);
   U19177 : NOR2_X1 port map( A1 => n14514, A2 => n14740, ZN => n13980);
   U19178 : AOI21_X1 port map( B1 => n13982, B2 => n13981, A => n13980, ZN => 
                           n13984);
   U19179 : NOR2_X1 port map( A1 => n15115, A2 => n15113, ZN => n15120);
   U19180 : AND2_X1 port map( A1 => n15120, A2 => n15116, ZN => n13983);
   U19181 : NOR2_X1 port map( A1 => n15125, A2 => n15000, ZN => n13987);
   U19182 : AOI22_X1 port map( A1 => n15132, A2 => n13987, B1 => n15004, B2 => 
                           n13986, ZN => n13988);
   U19183 : XNOR2_X1 port map( A => n28579, B => n15788, ZN => n16183);
   U19184 : XNOR2_X1 port map( A => n16183, B => n16424, ZN => n14028);
   U19185 : INV_X1 port map( A => n15085, ZN => n13989);
   U19186 : NAND2_X1 port map( A1 => n13989, A2 => n15691, ZN => n13992);
   U19187 : NAND2_X1 port map( A1 => n15691, A2 => n323, ZN => n14566);
   U19188 : OAI21_X1 port map( B1 => n1886, B2 => n14563, A => n15690, ZN => 
                           n13991);
   U19190 : OAI21_X1 port map( B1 => n15098, B2 => n15094, A => n15099, ZN => 
                           n13996);
   U19191 : OAI21_X1 port map( B1 => n13993, B2 => n14902, A => n14679, ZN => 
                           n13995);
   U19192 : AND2_X1 port map( A1 => n13993, A2 => n15094, ZN => n13994);
   U19193 : XNOR2_X1 port map( A => n16062, B => n16295, ZN => n14026);
   U19194 : MUX2_X1 port map( A => n13999, B => n13998, S => n14036, Z => 
                           n14003);
   U19195 : INV_X1 port map( A => n14000, ZN => n14001);
   U19196 : AOI22_X1 port map( A1 => n14001, A2 => n14036, B1 => n13587, B2 => 
                           n28569, ZN => n14002);
   U19197 : NAND2_X1 port map( A1 => n14003, A2 => n14002, ZN => n14824);
   U19198 : INV_X1 port map( A => n14004, ZN => n14382);
   U19199 : AND2_X1 port map( A1 => n14824, A2 => n15431, ZN => n14823);
   U19200 : INV_X1 port map( A => n14823, ZN => n14024);
   U19202 : NAND3_X1 port map( A1 => n14341, A2 => n14344, A3 => n14345, ZN => 
                           n14012);
   U19203 : NAND3_X1 port map( A1 => n14132, A2 => n14135, A3 => n14136, ZN => 
                           n14011);
   U19204 : INV_X1 port map( A => n14821, ZN => n15432);
   U19205 : NAND2_X1 port map( A1 => n2974, A2 => n14144, ZN => n14019);
   U19206 : NOR2_X1 port map( A1 => n29589, A2 => n4425, ZN => n14017);
   U19207 : AOI22_X1 port map( A1 => n14020, A2 => n14019, B1 => n14018, B2 => 
                           n14017, ZN => n14825);
   U19208 : INV_X1 port map( A => n14825, ZN => n15027);
   U19209 : NAND3_X1 port map( A1 => n15031, A2 => n14821, A3 => n15027, ZN => 
                           n14021);
   U19210 : XNOR2_X1 port map( A => n16059, B => n3380, ZN => n14025);
   U19211 : XNOR2_X1 port map( A => n14026, B => n14025, ZN => n14027);
   U19213 : INV_X1 port map( A => n17428, ZN => n17005);
   U19215 : MUX2_X1 port map( A => n14030, B => n14031, S => n14029, Z => 
                           n14035);
   U19216 : MUX2_X1 port map( A => n14032, B => n6066, S => n14031, Z => n14034
                           );
   U19218 : NAND2_X1 port map( A1 => n14046, A2 => n14051, ZN => n14048);
   U19219 : MUX2_X1 port map( A => n14049, B => n14048, S => n14047, Z => 
                           n14050);
   U19220 : NOR2_X1 port map( A1 => n14300, A2 => n28478, ZN => n14055);
   U19221 : INV_X1 port map( A => n14055, ZN => n14058);
   U19222 : OAI21_X1 port map( B1 => n14055, B2 => n5956, A => n14054, ZN => 
                           n14057);
   U19223 : NAND3_X1 port map( A1 => n29611, A2 => n14300, A3 => n14299, ZN => 
                           n14056);
   U19224 : OAI211_X2 port map( C1 => n14058, C2 => n14059, A => n14057, B => 
                           n14056, ZN => n14842);
   U19225 : NOR2_X1 port map( A1 => n28842, A2 => n14060, ZN => n14074);
   U19226 : INV_X1 port map( A => n14061, ZN => n14063);
   U19227 : MUX2_X1 port map( A => n14323, B => n14063, S => n29626, Z => 
                           n14067);
   U19228 : NAND2_X1 port map( A1 => n15286, A2 => n14601, ZN => n14073);
   U19229 : NAND2_X1 port map( A1 => n14068, A2 => n13583, ZN => n14069);
   U19230 : NOR2_X1 port map( A1 => n14696, A2 => n14071, ZN => n14072);
   U19231 : AOI21_X2 port map( B1 => n14074, B2 => n14073, A => n14072, ZN => 
                           n15801);
   U19232 : INV_X1 port map( A => n15292, ZN => n15289);
   U19233 : OAI21_X1 port map( B1 => n14078, B2 => n14077, A => n14249, ZN => 
                           n14079);
   U19234 : NOR2_X1 port map( A1 => n14080, A2 => n14082, ZN => n14090);
   U19236 : NAND3_X1 port map( A1 => n14085, A2 => n14083, A3 => n14084, ZN => 
                           n14087);
   U19237 : INV_X1 port map( A => n14365, ZN => n14368);
   U19238 : OAI21_X1 port map( B1 => n14094, B2 => n564, A => n14368, ZN => 
                           n14095);
   U19239 : MUX2_X1 port map( A => n1743, B => n14262, S => n14260, Z => n14100
                           );
   U19240 : INV_X1 port map( A => n14101, ZN => n14232);
   U19241 : NOR2_X1 port map( A1 => n14106, A2 => n14593, ZN => n14108);
   U19242 : INV_X1 port map( A => n14517, ZN => n15293);
   U19243 : XNOR2_X1 port map( A => n15801, B => n29516, ZN => n16179);
   U19244 : NAND2_X1 port map( A1 => n15115, A2 => n14514, ZN => n14111);
   U19245 : NAND2_X1 port map( A1 => n14112, A2 => n14744, ZN => n14113);
   U19246 : NAND2_X1 port map( A1 => n15138, A2 => n15250, ZN => n14730);
   U19247 : INV_X1 port map( A => n15137, ZN => n15251);
   U19248 : XNOR2_X1 port map( A => n16329, B => n16377, ZN => n14117);
   U19249 : XNOR2_X1 port map( A => n16179, B => n14117, ZN => n14225);
   U19250 : NAND2_X1 port map( A1 => n14119, A2 => n14118, ZN => n14124);
   U19251 : NAND2_X1 port map( A1 => n14120, A2 => n14365, ZN => n14121);
   U19253 : INV_X1 port map( A => n14153, ZN => n15355);
   U19255 : OAI211_X1 port map( C1 => n14127, C2 => n14355, A => n14126, B => 
                           n14125, ZN => n14130);
   U19256 : INV_X1 port map( A => n14752, ZN => n15243);
   U19257 : NAND2_X1 port map( A1 => n14132, A2 => n14131, ZN => n14133);
   U19258 : MUX2_X1 port map( A => n14134, B => n14133, S => n14345, Z => 
                           n14140);
   U19259 : NAND2_X1 port map( A1 => n14135, A2 => n14341, ZN => n14138);
   U19260 : NAND2_X1 port map( A1 => n14344, A2 => n14343, ZN => n14137);
   U19261 : MUX2_X1 port map( A => n14138, B => n14137, S => n14136, Z => 
                           n14139);
   U19262 : AOI21_X2 port map( B1 => n14144, B2 => n14145, A => n14143, ZN => 
                           n15060);
   U19263 : NOR2_X1 port map( A1 => n15060, A2 => n15355, ZN => n14149);
   U19264 : NAND2_X1 port map( A1 => n13594, A2 => n2849, ZN => n14147);
   U19265 : MUX2_X1 port map( A => n14150, B => n13572, S => n14386, Z => 
                           n14152);
   U19266 : NOR2_X1 port map( A1 => n15359, A2 => n14153, ZN => n14751);
   U19267 : XNOR2_X1 port map( A => n16467, B => n3516, ZN => n14223);
   U19268 : OAI22_X1 port map( A1 => n29036, A2 => n14491, B1 => n28601, B2 => 
                           n14494, ZN => n14156);
   U19269 : NAND2_X1 port map( A1 => n14156, A2 => n14493, ZN => n15344);
   U19270 : NAND2_X1 port map( A1 => n14157, A2 => n14480, ZN => n14476);
   U19271 : OAI21_X1 port map( B1 => n293, B2 => n14161, A => n14476, ZN => 
                           n14160);
   U19272 : AND2_X1 port map( A1 => n15222, A2 => n15343, ZN => n15228);
   U19273 : NAND2_X1 port map( A1 => n29565, A2 => n14164, ZN => n14168);
   U19274 : NOR2_X1 port map( A1 => n14757, A2 => n15222, ZN => n14191);
   U19275 : INV_X1 port map( A => n15342, ZN => n15225);
   U19276 : NAND2_X1 port map( A1 => n14178, A2 => n14451, ZN => n14179);
   U19277 : NAND2_X1 port map( A1 => n14183, A2 => n14182, ZN => n14190);
   U19278 : AOI21_X1 port map( B1 => n14465, B2 => n14185, A => n14184, ZN => 
                           n14186);
   U19279 : NAND2_X1 port map( A1 => n14187, A2 => n14186, ZN => n14188);
   U19280 : AOI21_X1 port map( B1 => n12534, B2 => n14426, A => n29558, ZN => 
                           n14197);
   U19281 : NAND2_X1 port map( A1 => n14199, A2 => n14198, ZN => n15238);
   U19282 : NAND2_X1 port map( A1 => n427, A2 => n14456, ZN => n14202);
   U19283 : MUX2_X1 port map( A => n14202, B => n14459, S => n28806, Z => 
                           n14203);
   U19285 : INV_X1 port map( A => n15238, ZN => n15233);
   U19286 : INV_X1 port map( A => n14206, ZN => n14209);
   U19287 : OAI211_X1 port map( C1 => n14432, C2 => n14437, A => n1841, B => 
                           n14207, ZN => n14208);
   U19288 : NAND3_X1 port map( A1 => n15338, A2 => n15233, A3 => n15334, ZN => 
                           n14222);
   U19289 : NAND2_X1 port map( A1 => n14402, A2 => n14399, ZN => n14211);
   U19290 : MUX2_X1 port map( A => n14211, B => n14210, S => n14400, Z => 
                           n14212);
   U19292 : INV_X1 port map( A => n15334, ZN => n15339);
   U19293 : OAI211_X1 port map( C1 => n14216, C2 => n14215, A => n14214, B => 
                           n29638, ZN => n14219);
   U19294 : NAND3_X1 port map( A1 => n14220, A2 => n15339, A3 => n15333, ZN => 
                           n14221);
   U19295 : XNOR2_X1 port map( A => n14225, B => n14224, ZN => n17426);
   U19296 : MUX2_X1 port map( A => n14227, B => n14226, S => n17426, Z => 
                           n14507);
   U19297 : MUX2_X1 port map( A => n14767, B => n14713, S => n14810, Z => 
                           n14228);
   U19298 : INV_X1 port map( A => n14595, ZN => n14233);
   U19299 : INV_X1 port map( A => n14234, ZN => n14236);
   U19300 : AND2_X1 port map( A1 => n14235, A2 => n14236, ZN => n14594);
   U19301 : OR2_X1 port map( A1 => n14237, A2 => n14252, ZN => n14596);
   U19302 : INV_X1 port map( A => n14596, ZN => n14248);
   U19303 : OAI21_X1 port map( B1 => n14240, B2 => n14239, A => n14238, ZN => 
                           n14242);
   U19304 : NAND2_X1 port map( A1 => n14242, A2 => n14241, ZN => n14247);
   U19305 : NAND3_X1 port map( A1 => n13943, A2 => n14243, A3 => n15194, ZN => 
                           n14246);
   U19306 : MUX2_X1 port map( A => n14251, B => n14250, S => n14249, Z => 
                           n14257);
   U19307 : NAND2_X1 port map( A1 => n14253, A2 => n14252, ZN => n14256);
   U19308 : INV_X1 port map( A => n14254, ZN => n14255);
   U19309 : NOR2_X1 port map( A1 => n14260, A2 => n14259, ZN => n14263);
   U19310 : INV_X1 port map( A => n14264, ZN => n14265);
   U19311 : OAI22_X1 port map( A1 => n14268, A2 => n14267, B1 => n14266, B2 => 
                           n14265, ZN => n14269);
   U19313 : NAND2_X1 port map( A1 => n14275, A2 => n14274, ZN => n14276);
   U19314 : NAND2_X1 port map( A1 => n14276, A2 => n14360, ZN => n14277);
   U19315 : NAND2_X1 port map( A1 => n14286, A2 => n14285, ZN => n14288);
   U19316 : INV_X1 port map( A => n15054, ZN => n15259);
   U19318 : OAI21_X1 port map( B1 => n14298, B2 => n14297, A => n14296, ZN => 
                           n14606);
   U19319 : NAND2_X1 port map( A1 => n15309, A2 => n14851, ZN => n14340);
   U19320 : AND2_X1 port map( A1 => n12534, A2 => n4522, ZN => n14607);
   U19321 : NOR2_X2 port map( A1 => n14610, A2 => n14607, ZN => n15319);
   U19322 : INV_X1 port map( A => n15319, ZN => n14854);
   U19323 : NAND2_X1 port map( A1 => n14311, A2 => n14313, ZN => n14316);
   U19324 : NOR2_X1 port map( A1 => n14314, A2 => n14313, ZN => n14315);
   U19325 : MUX2_X1 port map( A => n14319, B => n14318, S => n14317, Z => 
                           n14321);
   U19326 : NOR2_X1 port map( A1 => n14325, A2 => n14328, ZN => n14326);
   U19327 : NAND2_X1 port map( A1 => n14327, A2 => n14326, ZN => n14329);
   U19328 : AND2_X1 port map( A1 => n14406, A2 => n29133, ZN => n14409);
   U19329 : INV_X1 port map( A => n14409, ZN => n14337);
   U19330 : NOR2_X1 port map( A1 => n14332, A2 => n14406, ZN => n14334);
   U19331 : OAI21_X1 port map( B1 => n14337, B2 => n1830, A => n14335, ZN => 
                           n15307);
   U19332 : OAI21_X1 port map( B1 => n15309, B2 => n15307, A => n14851, ZN => 
                           n14338);
   U19333 : OAI21_X1 port map( B1 => n14340, B2 => n14854, A => n14339, ZN => 
                           n16339);
   U19334 : INV_X1 port map( A => n16339, ZN => n16130);
   U19335 : MUX2_X1 port map( A => n14343, B => n14342, S => n14341, Z => 
                           n14348);
   U19336 : MUX2_X1 port map( A => n14345, B => n14344, S => n14343, Z => 
                           n14347);
   U19337 : MUX2_X2 port map( A => n14348, B => n14347, S => n14346, Z => 
                           n15514);
   U19339 : NOR2_X1 port map( A1 => n15274, A2 => n15515, ZN => n14364);
   U19340 : NAND2_X1 port map( A1 => n15510, A2 => n15276, ZN => n14388);
   U19341 : AOI22_X1 port map( A1 => n13725, A2 => n14373, B1 => n14376, B2 => 
                           n14372, ZN => n14375);
   U19342 : INV_X1 port map( A => n15511, ZN => n14918);
   U19344 : OAI211_X1 port map( C1 => n14918, C2 => n15274, A => n14920, B => 
                           n15515, ZN => n14387);
   U19345 : XNOR2_X1 port map( A => n16130, B => n16443, ZN => n16028);
   U19346 : XNOR2_X1 port map( A => n16028, B => n16154, ZN => n14506);
   U19347 : NOR2_X1 port map( A1 => n15285, A2 => n14695, ZN => n14844);
   U19348 : INV_X1 port map( A => n14844, ZN => n14390);
   U19349 : OAI21_X1 port map( B1 => n6048, B2 => n14842, A => n14695, ZN => 
                           n14392);
   U19350 : XNOR2_X1 port map( A => n15452, B => n3528, ZN => n14504);
   U19352 : AOI21_X1 port map( B1 => n14332, B2 => n14406, A => n14405, ZN => 
                           n14412);
   U19354 : INV_X1 port map( A => n14413, ZN => n14423);
   U19355 : NAND2_X1 port map( A1 => n28648, A2 => n14414, ZN => n14422);
   U19356 : AOI21_X1 port map( B1 => n29638, B2 => n14415, A => n14414, ZN => 
                           n14418);
   U19357 : INV_X1 port map( A => n14621, ZN => n14705);
   U19358 : NAND2_X1 port map( A1 => n14436, A2 => n14435, ZN => n14443);
   U19359 : NAND3_X1 port map( A1 => n14438, A2 => n14440, A3 => n14437, ZN => 
                           n14442);
   U19360 : NAND3_X1 port map( A1 => n1841, A2 => n14440, A3 => n14439, ZN => 
                           n14441);
   U19361 : INV_X1 port map( A => n28647, ZN => n14445);
   U19362 : OR2_X1 port map( A1 => n14446, A2 => n14445, ZN => n14447);
   U19363 : NOR2_X1 port map( A1 => n427, A2 => n14459, ZN => n14457);
   U19364 : OAI21_X1 port map( B1 => n14458, B2 => n14457, A => n14456, ZN => 
                           n14462);
   U19365 : NAND2_X1 port map( A1 => n14460, A2 => n14459, ZN => n14461);
   U19366 : OAI211_X1 port map( C1 => n427, C2 => n14463, A => n14462, B => 
                           n14461, ZN => n15490);
   U19367 : INV_X1 port map( A => n15490, ZN => n14702);
   U19368 : NAND2_X1 port map( A1 => n14465, A2 => n14464, ZN => n14468);
   U19369 : MUX2_X1 port map( A => n14471, B => n14470, S => n14469, Z => 
                           n14472);
   U19370 : NAND2_X1 port map( A1 => n14473, A2 => n14480, ZN => n14478);
   U19371 : NAND3_X1 port map( A1 => n14476, A2 => n14475, A3 => n14474, ZN => 
                           n14477);
   U19373 : NAND2_X1 port map( A1 => n15491, A2 => n15485, ZN => n14917);
   U19374 : NAND2_X1 port map( A1 => n29565, A2 => n14481, ZN => n14482);
   U19375 : MUX2_X1 port map( A => n14483, B => n14482, S => n14166, Z => 
                           n14490);
   U19376 : NOR2_X1 port map( A1 => n14485, A2 => n14484, ZN => n14488);
   U19377 : AOI22_X1 port map( A1 => n14488, A2 => n14166, B1 => n14487, B2 => 
                           n14486, ZN => n14489);
   U19378 : NOR2_X1 port map( A1 => n29037, A2 => n14493, ZN => n14495);
   U19379 : AND3_X1 port map( A1 => n29036, A2 => n14498, A3 => n14497, ZN => 
                           n14616);
   U19380 : NOR2_X1 port map( A1 => n15490, A2 => n14616, ZN => n14500);
   U19381 : XNOR2_X1 port map( A => n16653, B => n16558, ZN => n16406);
   U19382 : XNOR2_X1 port map( A => n16406, B => n14504, ZN => n14505);
   U19383 : XNOR2_X1 port map( A => n14505, B => n14506, ZN => n17424);
   U19385 : OAI21_X1 port map( B1 => n15138, B2 => n15246, A => n15252, ZN => 
                           n14511);
   U19387 : INV_X1 port map( A => n15250, ZN => n15136);
   U19388 : NAND3_X1 port map( A1 => n15135, A2 => n15136, A3 => n15248, ZN => 
                           n14509);
   U19390 : NOR2_X1 port map( A1 => n14514, A2 => n15117, ZN => n14742);
   U19391 : NAND2_X1 port map( A1 => n14742, A2 => n15115, ZN => n14515);
   U19392 : OR2_X1 port map( A1 => n15215, A2 => n15292, ZN => n14522);
   U19393 : NAND3_X1 port map( A1 => n15036, A2 => n15290, A3 => n14517, ZN => 
                           n14519);
   U19394 : NAND4_X2 port map( A1 => n14522, A2 => n14521, A3 => n14520, A4 => 
                           n14519, ZN => n16262);
   U19395 : XNOR2_X1 port map( A => n16262, B => n72, ZN => n14523);
   U19396 : INV_X1 port map( A => n15224, ZN => n15348);
   U19397 : MUX2_X1 port map( A => n15225, B => n15348, S => n15046, Z => 
                           n14525);
   U19399 : NAND2_X1 port map( A1 => n15338, A2 => n15333, ZN => n14526);
   U19400 : AND3_X1 port map( A1 => n15238, A2 => n14526, A3 => n14781, ZN => 
                           n14527);
   U19401 : INV_X1 port map( A => n16024, ZN => n14529);
   U19402 : XNOR2_X1 port map( A => n14529, B => n16405, ZN => n15893);
   U19403 : NAND3_X1 port map( A1 => n15183, A2 => n552, A3 => n14785, ZN => 
                           n14530);
   U19404 : NAND3_X1 port map( A1 => n553, A2 => n15457, A3 => n15174, ZN => 
                           n14538);
   U19405 : NOR2_X1 port map( A1 => n15456, A2 => n15174, ZN => n15458);
   U19406 : NAND3_X1 port map( A1 => n15180, A2 => n15174, A3 => n28803, ZN => 
                           n14536);
   U19407 : NAND3_X1 port map( A1 => n14534, A2 => n5635, A3 => n15456, ZN => 
                           n14535);
   U19408 : XNOR2_X1 port map( A => n16052, B => n15927, ZN => n16311);
   U19409 : NAND3_X1 port map( A1 => n15202, A2 => n15204, A3 => n14967, ZN => 
                           n14543);
   U19410 : NOR2_X1 port map( A1 => n15202, A2 => n15208, ZN => n14539);
   U19411 : AND2_X1 port map( A1 => n15207, A2 => n15208, ZN => n14964);
   U19412 : NAND2_X1 port map( A1 => n15209, A2 => n14960, ZN => n14540);
   U19413 : NAND3_X2 port map( A1 => n14542, A2 => n14543, A3 => n14541, ZN => 
                           n16247);
   U19414 : XNOR2_X1 port map( A => n16247, B => n5059, ZN => n14544);
   U19415 : XNOR2_X1 port map( A => n16311, B => n14544, ZN => n14562);
   U19416 : INV_X1 port map( A => n15466, ZN => n15159);
   U19417 : NAND2_X1 port map( A1 => n15159, A2 => n15463, ZN => n14546);
   U19418 : NOR3_X1 port map( A1 => n15462, A2 => n14652, A3 => n29153, ZN => 
                           n14545);
   U19420 : NAND2_X1 port map( A1 => n15168, A2 => n15474, ZN => n15170);
   U19421 : INV_X1 port map( A => n15167, ZN => n14958);
   U19422 : NAND3_X1 port map( A1 => n15166, A2 => n14551, A3 => n1848, ZN => 
                           n14552);
   U19423 : OAI211_X1 port map( C1 => n1809, C2 => n15170, A => n14553, B => 
                           n14552, ZN => n16435);
   U19424 : INV_X1 port map( A => n16435, ZN => n14554);
   U19425 : XNOR2_X1 port map( A => n14554, B => n16603, ZN => n16343);
   U19426 : NOR2_X1 port map( A1 => n14810, A2 => n14713, ZN => n14559);
   U19427 : INV_X1 port map( A => n14713, ZN => n14766);
   U19428 : OAI21_X1 port map( B1 => n14767, B2 => n14766, A => n13922, ZN => 
                           n14558);
   U19429 : NAND2_X1 port map( A1 => n14559, A2 => n14715, ZN => n14557);
   U19430 : NAND2_X1 port map( A1 => n14775, A2 => n14555, ZN => n14556);
   U19431 : XNOR2_X1 port map( A => n16618, B => n16312, ZN => n14560);
   U19432 : XNOR2_X1 port map( A => n16343, B => n14560, ZN => n14561);
   U19433 : NAND2_X1 port map( A1 => n15690, A2 => n15083, ZN => n14877);
   U19434 : AND2_X1 port map( A1 => n14877, A2 => n14563, ZN => n14565);
   U19435 : NAND2_X1 port map( A1 => n14670, A2 => n323, ZN => n14564);
   U19436 : OAI21_X1 port map( B1 => n15692, B2 => n14565, A => n14564, ZN => 
                           n14568);
   U19437 : NOR2_X1 port map( A1 => n15084, A2 => n14566, ZN => n14567);
   U19438 : NOR2_X1 port map( A1 => n14568, A2 => n14567, ZN => n14921);
   U19439 : INV_X1 port map( A => n15082, ZN => n14574);
   U19441 : INV_X1 port map( A => n15077, ZN => n15075);
   U19442 : OR2_X1 port map( A1 => n14948, A2 => n15077, ZN => n14872);
   U19443 : NAND2_X1 port map( A1 => n14872, A2 => n14571, ZN => n14573);
   U19445 : INV_X1 port map( A => n16320, ZN => n14581);
   U19446 : OAI21_X1 port map( B1 => n15420, B2 => n15101, A => n4549, ZN => 
                           n14576);
   U19447 : AOI21_X1 port map( B1 => n14903, B2 => n15097, A => n14578, ZN => 
                           n14580);
   U19448 : XNOR2_X1 port map( A => n14581, B => n15903, ZN => n14592);
   U19449 : NAND2_X1 port map( A1 => n14881, A2 => n13789, ZN => n14585);
   U19450 : XNOR2_X1 port map( A => n29319, B => n16256, ZN => n14590);
   U19451 : NAND2_X1 port map( A1 => n15406, A2 => n14894, ZN => n14939);
   U19452 : INV_X1 port map( A => n15407, ZN => n15416);
   U19453 : AOI21_X1 port map( B1 => n14940, B2 => n14939, A => n15416, ZN => 
                           n14588);
   U19454 : NAND2_X1 port map( A1 => n15415, A2 => n15409, ZN => n14586);
   U19455 : AOI21_X1 port map( B1 => n14586, B2 => n14893, A => n14894, ZN => 
                           n14587);
   U19456 : XNOR2_X1 port map( A => n16257, B => n3728, ZN => n14589);
   U19457 : XNOR2_X1 port map( A => n14590, B => n14589, ZN => n14591);
   U19459 : INV_X1 port map( A => n29297, ZN => n16996);
   U19460 : INV_X1 port map( A => n14762, ZN => n15056);
   U19461 : NAND2_X1 port map( A1 => n14597, A2 => n14596, ZN => n15053);
   U19462 : NAND2_X1 port map( A1 => n15053, A2 => n14761, ZN => n14598);
   U19463 : NAND3_X1 port map( A1 => n15055, A2 => n15261, A3 => n14763, ZN => 
                           n14599);
   U19464 : INV_X1 port map( A => n15366, ZN => n14603);
   U19466 : NOR2_X1 port map( A1 => n15274, A2 => n15511, ZN => n14605);
   U19467 : NOR2_X1 port map( A1 => n15514, A2 => n14697, ZN => n14604);
   U19468 : INV_X1 port map( A => n15307, ZN => n15308);
   U19469 : INV_X1 port map( A => n15306, ZN => n15312);
   U19470 : OAI21_X1 port map( B1 => n15312, B2 => n15310, A => n14851, ZN => 
                           n14613);
   U19471 : INV_X1 port map( A => n14606, ZN => n14609);
   U19472 : INV_X1 port map( A => n14607, ZN => n14608);
   U19473 : NAND3_X1 port map( A1 => n1096, A2 => n14609, A3 => n14608, ZN => 
                           n14611);
   U19474 : OAI21_X1 port map( B1 => n14611, B2 => n14610, A => n15311, ZN => 
                           n14612);
   U19476 : NAND2_X1 port map( A1 => n14702, A2 => n15485, ZN => n14617);
   U19478 : INV_X1 port map( A => n15489, ZN => n15486);
   U19479 : NAND3_X1 port map( A1 => n15486, A2 => n14702, A3 => n14703, ZN => 
                           n14619);
   U19480 : NOR2_X1 port map( A1 => n15503, A2 => n15265, ZN => n14623);
   U19481 : AOI22_X1 port map( A1 => n14623, A2 => n15502, B1 => n14622, B2 => 
                           n15500, ZN => n14627);
   U19482 : INV_X1 port map( A => n15506, ZN => n14625);
   U19483 : INV_X1 port map( A => n14623, ZN => n14624);
   U19484 : OAI211_X1 port map( C1 => n14625, C2 => n15497, A => n14624, B => 
                           n14922, ZN => n14626);
   U19485 : XNOR2_X1 port map( A => n16399, B => n16043, ZN => n16367);
   U19486 : XNOR2_X1 port map( A => n16278, B => n16367, ZN => n14628);
   U19487 : NOR2_X1 port map( A1 => n14992, A2 => n15394, ZN => n14632);
   U19488 : AOI22_X1 port map( A1 => n15395, A2 => n14632, B1 => n15391, B2 => 
                           n14631, ZN => n14635);
   U19491 : MUX2_X1 port map( A => n15382, B => n15152, S => n14986, Z => 
                           n14638);
   U19492 : OR2_X1 port map( A1 => n15382, A2 => n15151, ZN => n15154);
   U19493 : NAND3_X1 port map( A1 => n15382, A2 => n14986, A3 => n15150, ZN => 
                           n14636);
   U19494 : AND2_X1 port map( A1 => n15154, A2 => n14636, ZN => n14637);
   U19495 : OAI21_X1 port map( B1 => n14638, B2 => n15155, A => n14637, ZN => 
                           n16426);
   U19496 : XNOR2_X1 port map( A => n16426, B => n16567, ZN => n16362);
   U19497 : INV_X1 port map( A => n16362, ZN => n14643);
   U19498 : OAI21_X1 port map( B1 => n15077, B2 => n15072, A => n15081, ZN => 
                           n14640);
   U19499 : XNOR2_X1 port map( A => n16272, B => n16295, ZN => n15426);
   U19500 : INV_X1 port map( A => n15426, ZN => n14642);
   U19501 : XNOR2_X1 port map( A => n14643, B => n14642, ZN => n14656);
   U19502 : NAND3_X1 port map( A1 => n15184, A2 => n15183, A3 => n15190, ZN => 
                           n14648);
   U19503 : INV_X1 port map( A => n15183, ZN => n14644);
   U19504 : NAND3_X1 port map( A1 => n15186, A2 => n14644, A3 => n15185, ZN => 
                           n14647);
   U19505 : NAND2_X1 port map( A1 => n14645, A2 => n14644, ZN => n14646);
   U19507 : NAND3_X1 port map( A1 => n3784, A2 => n6879, A3 => n15370, ZN => 
                           n14651);
   U19508 : NOR2_X1 port map( A1 => n15372, A2 => n14863, ZN => n14650);
   U19509 : XNOR2_X1 port map( A => n15817, B => n16294, ZN => n14654);
   U19510 : XNOR2_X1 port map( A => n321, B => n2889, ZN => n14653);
   U19511 : XNOR2_X1 port map( A => n14654, B => n14653, ZN => n14655);
   U19512 : OAI21_X1 port map( B1 => n16863, B2 => n16996, A => n16991, ZN => 
                           n14694);
   U19513 : NOR2_X1 port map( A1 => n16992, A2 => n17269, ZN => n14693);
   U19514 : NOR2_X1 port map( A1 => n15438, A2 => n15436, ZN => n15020);
   U19515 : INV_X1 port map( A => n14658, ZN => n14663);
   U19516 : INV_X1 port map( A => n14659, ZN => n14662);
   U19518 : NAND2_X1 port map( A1 => n14670, A2 => n28666, ZN => n14672);
   U19519 : OAI211_X1 port map( C1 => n323, C2 => n15691, A => n15087, B => 
                           n15689, ZN => n14671);
   U19520 : XNOR2_X1 port map( A => n28597, B => n16641, ZN => n14676);
   U19521 : NAND2_X1 port map( A1 => n15321, A2 => n15013, ZN => n15326);
   U19522 : INV_X1 port map( A => n15013, ZN => n15445);
   U19523 : OAI211_X1 port map( C1 => n15014, C2 => n15015, A => n15322, B => 
                           n15445, ZN => n14674);
   U19524 : NAND2_X1 port map( A1 => n1926, A2 => n15014, ZN => n14673);
   U19525 : XNOR2_X1 port map( A => n14676, B => n14675, ZN => n14692);
   U19526 : INV_X1 port map( A => n15094, ZN => n14680);
   U19527 : AOI21_X1 port map( B1 => n3315, B2 => n14680, A => n14679, ZN => 
                           n14681);
   U19528 : INV_X1 port map( A => n14824, ZN => n15032);
   U19529 : INV_X1 port map( A => n15029, ZN => n14684);
   U19530 : XNOR2_X1 port map( A => n15909, B => n15802, ZN => n16331);
   U19531 : NAND2_X1 port map( A1 => n14685, A2 => n15000, ZN => n14690);
   U19532 : INV_X1 port map( A => n15132, ZN => n14689);
   U19533 : XNOR2_X1 port map( A => n16329, B => n16238, ZN => n16082);
   U19534 : XNOR2_X1 port map( A => n16082, B => n16331, ZN => n14691);
   U19535 : XNOR2_X1 port map( A => n14692, B => n14691, ZN => n16995);
   U19536 : XNOR2_X1 port map( A => n16563, B => n1911, ZN => n14701);
   U19537 : NAND2_X1 port map( A1 => n14698, A2 => n15512, ZN => n14699);
   U19538 : NAND3_X1 port map( A1 => n15309, A2 => n15312, A3 => n15307, ZN => 
                           n14700);
   U19539 : XNOR2_X1 port map( A => n16216, B => n16421, ZN => n16536);
   U19540 : XNOR2_X1 port map( A => n16536, B => n14701, ZN => n14721);
   U19541 : INV_X1 port map( A => n15494, ZN => n15269);
   U19542 : AND2_X1 port map( A1 => n14922, A2 => n15503, ZN => n14707);
   U19544 : INV_X1 port map( A => n16185, ZN => n14709);
   U19545 : INV_X1 port map( A => n16270, ZN => n15878);
   U19546 : INV_X1 port map( A => n15053, ZN => n15262);
   U19547 : NOR2_X1 port map( A1 => n15262, A2 => n15260, ZN => n14710);
   U19549 : INV_X1 port map( A => n16568, ZN => n14719);
   U19550 : INV_X1 port map( A => n14712, ZN => n14714);
   U19551 : AOI21_X1 port map( B1 => n14714, B2 => n14713, A => n14810, ZN => 
                           n14718);
   U19552 : NAND2_X1 port map( A1 => n14810, A2 => n28493, ZN => n14716);
   U19553 : AOI21_X1 port map( B1 => n14811, B2 => n14716, A => n14773, ZN => 
                           n14717);
   U19554 : XNOR2_X1 port map( A => n15878, B => n16145, ZN => n14720);
   U19555 : NAND2_X1 port map( A1 => n15387, A2 => n15388, ZN => n14728);
   U19556 : NAND2_X1 port map( A1 => n15395, A2 => n14722, ZN => n14727);
   U19557 : NAND2_X1 port map( A1 => n15389, A2 => n3210, ZN => n14725);
   U19558 : INV_X1 port map( A => n15389, ZN => n15145);
   U19559 : OAI21_X1 port map( B1 => n15387, B2 => n15144, A => n15145, ZN => 
                           n14724);
   U19560 : OAI211_X1 port map( C1 => n14990, C2 => n14725, A => n14724, B => 
                           n14723, ZN => n14726);
   U19561 : NAND3_X1 port map( A1 => n15252, A2 => n15138, A3 => n15246, ZN => 
                           n14731);
   U19562 : XNOR2_X1 port map( A => n16280, B => n543, ZN => n15863);
   U19563 : INV_X1 port map( A => n15863, ZN => n14736);
   U19564 : NAND2_X1 port map( A1 => n28196, A2 => n28518, ZN => n15399);
   U19565 : XNOR2_X1 port map( A => n16365, B => n1225, ZN => n14735);
   U19566 : XNOR2_X1 port map( A => n14736, B => n14735, ZN => n14749);
   U19567 : MUX2_X1 port map( A => n15155, B => n15382, S => n15383, Z => 
                           n14739);
   U19568 : NOR2_X1 port map( A1 => n14740, A2 => n1904, ZN => n14741);
   U19569 : NAND2_X1 port map( A1 => n15115, A2 => n14743, ZN => n14745);
   U19570 : NAND2_X1 port map( A1 => n15000, A2 => n15127, ZN => n14747);
   U19571 : XNOR2_X1 port map( A => n16116, B => n16506, ZN => n14748);
   U19573 : OAI21_X1 port map( B1 => n15060, B2 => n14753, A => n15359, ZN => 
                           n14754);
   U19575 : AND2_X1 port map( A1 => n15343, A2 => n15342, ZN => n14756);
   U19576 : NAND2_X1 port map( A1 => n15226, A2 => n14756, ZN => n14759);
   U19577 : AOI22_X1 port map( A1 => n14757, A2 => n15223, B1 => n15348, B2 => 
                           n15343, ZN => n14758);
   U19578 : INV_X1 port map( A => n16578, ZN => n14760);
   U19579 : XNOR2_X1 port map( A => n14760, B => n16495, ZN => n16124);
   U19580 : OAI21_X1 port map( B1 => n14810, B2 => n14767, A => n14766, ZN => 
                           n14768);
   U19581 : NAND2_X1 port map( A1 => n14768, A2 => n13922, ZN => n14777);
   U19582 : INV_X1 port map( A => n14772, ZN => n14774);
   U19583 : XNOR2_X1 port map( A => n16416, B => n16012, ZN => n16497);
   U19584 : INV_X1 port map( A => n16497, ZN => n14778);
   U19585 : XNOR2_X1 port map( A => n14778, B => n16124, ZN => n14791);
   U19586 : XNOR2_X1 port map( A => n16579, B => n3586, ZN => n14789);
   U19587 : INV_X1 port map( A => n15239, ZN => n15235);
   U19588 : NAND3_X1 port map( A1 => n15234, A2 => n15338, A3 => n15334, ZN => 
                           n14782);
   U19589 : INV_X1 port map( A => n14784, ZN => n14783);
   U19590 : AOI21_X1 port map( B1 => n15184, B2 => n15185, A => n14783, ZN => 
                           n14788);
   U19591 : OAI21_X1 port map( B1 => n14785, B2 => n15182, A => n14799, ZN => 
                           n14786);
   U19592 : NAND2_X1 port map( A1 => n14786, A2 => n15183, ZN => n14787);
   U19593 : XNOR2_X1 port map( A => n16321, B => n16077, ZN => n16253);
   U19594 : XNOR2_X1 port map( A => n14789, B => n16253, ZN => n14790);
   U19595 : XNOR2_X1 port map( A => n14791, B => n14790, ZN => n14871);
   U19596 : OAI211_X1 port map( C1 => n14881, C2 => n13789, A => n14793, B => 
                           n5813, ZN => n14794);
   U19597 : AOI22_X1 port map( A1 => n15459, A2 => n15174, B1 => n15456, B2 => 
                           n28803, ZN => n15461);
   U19598 : OAI211_X1 port map( C1 => n14534, C2 => n28803, A => n28462, B => 
                           n15457, ZN => n14798);
   U19599 : XNOR2_X1 port map( A => n28585, B => n15760, ZN => n16514);
   U19600 : XNOR2_X1 port map( A => n16119, B => n16514, ZN => n14815);
   U19601 : INV_X1 port map( A => n15171, ZN => n15475);
   U19602 : NAND2_X1 port map( A1 => n15475, A2 => n15476, ZN => n15473);
   U19603 : OAI211_X1 port map( C1 => n15166, C2 => n15168, A => n15171, B => 
                           n14958, ZN => n14801);
   U19604 : NAND2_X1 port map( A1 => n545, A2 => n15462, ZN => n15164);
   U19605 : INV_X1 port map( A => n15164, ZN => n14804);
   U19606 : NAND2_X1 port map( A1 => n14802, A2 => n15161, ZN => n14803);
   U19607 : AOI21_X1 port map( B1 => n14808, B2 => n14807, A => n28493, ZN => 
                           n14809);
   U19608 : XNOR2_X1 port map( A => n16586, B => n135, ZN => n14813);
   U19609 : XNOR2_X1 port map( A => n16243, B => n14813, ZN => n14814);
   U19610 : XNOR2_X1 port map( A => n14815, B => n14814, ZN => n16999);
   U19611 : MUX2_X1 port map( A => n29572, B => n14871, S => n16999, Z => 
                           n14915);
   U19612 : AND3_X1 port map( A1 => n15437, A2 => n15438, A3 => n15300, ZN => 
                           n14816);
   U19613 : AOI21_X1 port map( B1 => n15444, B2 => n15302, A => n14816, ZN => 
                           n14820);
   U19614 : INV_X1 port map( A => n15300, ZN => n15440);
   U19615 : OAI21_X1 port map( B1 => n15444, B2 => n15436, A => n15440, ZN => 
                           n14819);
   U19616 : INV_X1 port map( A => n15303, ZN => n14817);
   U19617 : NOR2_X1 port map( A1 => n14817, A2 => n15022, ZN => n14818);
   U19618 : NOR2_X1 port map( A1 => n14821, A2 => n14826, ZN => n14822);
   U19619 : NAND2_X1 port map( A1 => n15032, A2 => n14825, ZN => n14827);
   U19620 : AOI21_X1 port map( B1 => n15433, B2 => n14827, A => n15430, ZN => 
                           n14828);
   U19621 : NOR2_X1 port map( A1 => n14832, A2 => n14831, ZN => n14835);
   U19622 : OAI21_X1 port map( B1 => n14837, B2 => n15294, A => n14836, ZN => 
                           n14840);
   U19623 : INV_X1 port map( A => n15291, ZN => n15037);
   U19624 : OAI21_X1 port map( B1 => n15215, B2 => n15037, A => n14838, ZN => 
                           n14839);
   U19625 : INV_X1 port map( A => n15284, ZN => n14841);
   U19626 : NOR2_X1 port map( A1 => n28996, A2 => n14842, ZN => n14843);
   U19627 : XNOR2_X1 port map( A => n16017, B => n15887, ZN => n16524);
   U19628 : INV_X1 port map( A => n16524, ZN => n14850);
   U19629 : INV_X1 port map( A => n15309, ZN => n14852);
   U19630 : NAND3_X1 port map( A1 => n14854, A2 => n14851, A3 => n14852, ZN => 
                           n14858);
   U19631 : NOR2_X1 port map( A1 => n14852, A2 => n15310, ZN => n14853);
   U19632 : NAND2_X1 port map( A1 => n14854, A2 => n14853, ZN => n14857);
   U19633 : NAND3_X1 port map( A1 => n15310, A2 => n15311, A3 => n15306, ZN => 
                           n14856);
   U19634 : NAND3_X1 port map( A1 => n15322, A2 => n546, A3 => n15321, ZN => 
                           n14862);
   U19635 : NAND3_X1 port map( A1 => n15447, A2 => n15321, A3 => n15014, ZN => 
                           n14861);
   U19636 : INV_X1 port map( A => n15321, ZN => n15446);
   U19637 : NAND3_X1 port map( A1 => n15446, A2 => n546, A3 => n15445, ZN => 
                           n14860);
   U19638 : INV_X1 port map( A => n15014, ZN => n15448);
   U19639 : NAND3_X1 port map( A1 => n1926, A2 => n15448, A3 => n15015, ZN => 
                           n14859);
   U19640 : XNOR2_X1 port map( A => n16165, B => n16313, ZN => n16249);
   U19641 : NOR2_X1 port map( A1 => n15009, A2 => n14863, ZN => n14864);
   U19642 : OAI21_X1 port map( B1 => n14865, B2 => n14864, A => n15373, ZN => 
                           n14866);
   U19643 : XNOR2_X1 port map( A => n16249, B => n14868, ZN => n14869);
   U19644 : XNOR2_X1 port map( A => n14870, B => n14869, ZN => n17396);
   U19645 : OAI21_X1 port map( B1 => n15073, B2 => n15072, A => n14872, ZN => 
                           n14873);
   U19646 : NAND2_X1 port map( A1 => n14873, A2 => n15071, ZN => n14875);
   U19647 : AND2_X1 port map( A1 => n15072, A2 => n14874, ZN => n15078);
   U19648 : MUX2_X1 port map( A => n323, B => n15690, S => n15692, Z => n14880)
                           ;
   U19649 : NAND2_X1 port map( A1 => n14878, A2 => n14877, ZN => n14879);
   U19650 : XNOR2_X1 port map( A => n15849, B => n15982, ZN => n16518);
   U19651 : INV_X1 port map( A => n16518, ZN => n14892);
   U19652 : NAND2_X1 port map( A1 => n14882, A2 => n14881, ZN => n14883);
   U19653 : NAND2_X1 port map( A1 => n14883, A2 => n388, ZN => n14889);
   U19654 : NOR2_X1 port map( A1 => n14884, A2 => n5813, ZN => n14888);
   U19655 : NAND3_X1 port map( A1 => n14886, A2 => n13789, A3 => n14885, ZN => 
                           n14887);
   U19656 : XNOR2_X1 port map( A => n16131, B => n14890, ZN => n14891);
   U19657 : XNOR2_X1 port map( A => n14892, B => n14891, ZN => n14914);
   U19658 : NAND2_X1 port map( A1 => n14895, A2 => n28196, ZN => n14899);
   U19659 : NAND2_X1 port map( A1 => n14944, A2 => n15402, ZN => n14897);
   U19660 : OAI211_X1 port map( C1 => n28196, C2 => n15398, A => n14899, B => 
                           n14898, ZN => n16409);
   U19661 : XNOR2_X1 port map( A => n16409, B => n16556, ZN => n16134);
   U19662 : NAND2_X1 port map( A1 => n14903, A2 => n14901, ZN => n15096);
   U19663 : NAND3_X1 port map( A1 => n15096, A2 => n15099, A3 => n15100, ZN => 
                           n14911);
   U19664 : NAND2_X1 port map( A1 => n14908, A2 => n14907, ZN => n14909);
   U19665 : OAI211_X1 port map( C1 => n15095, C2 => n15094, A => n3315, B => 
                           n14909, ZN => n14910);
   U19666 : XNOR2_X1 port map( A => n16070, B => n2946, ZN => n14912);
   U19667 : XNOR2_X1 port map( A => n16134, B => n14912, ZN => n14913);
   U19668 : INV_X1 port map( A => n17397, ZN => n17402);
   U19669 : INV_X1 port map( A => n16498, ZN => n15855);
   U19670 : NAND2_X1 port map( A1 => n15510, A2 => n14918, ZN => n14919);
   U19673 : XNOR2_X1 port map( A => n16455, B => n16038, ZN => n14931);
   U19674 : NAND2_X1 port map( A1 => n14927, A2 => n14967, ZN => n14929);
   U19675 : XNOR2_X1 port map( A => n15654, B => n3109, ZN => n14930);
   U19676 : XNOR2_X1 port map( A => n14931, B => n14930, ZN => n14932);
   U19677 : INV_X1 port map( A => n15802, ZN => n14933);
   U19678 : XNOR2_X1 port map( A => n14933, B => n16509, ZN => n14941);
   U19679 : INV_X1 port map( A => n15101, ZN => n15417);
   U19680 : OAI211_X1 port map( C1 => n15407, C2 => n15406, A => n14937, B => 
                           n15410, ZN => n14938);
   U19681 : XNOR2_X1 port map( A => n15583, B => n16241, ZN => n15948);
   U19682 : XNOR2_X1 port map( A => n15948, B => n14941, ZN => n14955);
   U19683 : XNOR2_X1 port map( A => n16641, B => n2916, ZN => n14953);
   U19684 : NOR2_X1 port map( A1 => n15401, A2 => n28518, ZN => n14947);
   U19685 : NAND2_X1 port map( A1 => n14945, A2 => n15399, ZN => n14946);
   U19686 : AOI21_X1 port map( B1 => n14949, B2 => n15071, A => n15076, ZN => 
                           n14951);
   U19688 : XNOR2_X1 port map( A => n15949, B => n15999, ZN => n16639);
   U19689 : XNOR2_X1 port map( A => n16639, B => n14953, ZN => n14954);
   U19690 : AOI22_X1 port map( A1 => n15475, A2 => n14958, B1 => n1850, B2 => 
                           n15168, ZN => n14956);
   U19691 : MUX2_X1 port map( A => n14956, B => n15170, S => n15166, Z => 
                           n14957);
   U19693 : NOR2_X1 port map( A1 => n15208, A2 => n14960, ZN => n14962);
   U19694 : AOI22_X1 port map( A1 => n14963, A2 => n15208, B1 => n14962, B2 => 
                           n14961, ZN => n14966);
   U19696 : XNOR2_X1 port map( A => n16296, B => n16534, ZN => n15944);
   U19697 : XNOR2_X1 port map( A => n321, B => n3537, ZN => n14978);
   U19698 : NAND2_X1 port map( A1 => n14972, A2 => n14971, ZN => n14973);
   U19700 : AOI21_X2 port map( B1 => n14977, B2 => n14976, A => n14975, ZN => 
                           n16211);
   U19701 : XNOR2_X1 port map( A => n14978, B => n16211, ZN => n14979);
   U19702 : XNOR2_X1 port map( A => n14979, B => n15944, ZN => n14985);
   U19703 : NAND2_X1 port map( A1 => n15180, A2 => n15174, ZN => n14982);
   U19704 : INV_X1 port map( A => n16422, ZN => n14983);
   U19705 : MUX2_X1 port map( A => n15383, B => n15151, S => n15382, Z => 
                           n14988);
   U19706 : MUX2_X1 port map( A => n15382, B => n14986, S => n15379, Z => 
                           n14987);
   U19707 : NOR2_X1 port map( A1 => n15394, A2 => n15388, ZN => n14991);
   U19708 : XNOR2_X1 port map( A => n16023, B => n3422, ZN => n14996);
   U19709 : INV_X1 port map( A => n16409, ZN => n14995);
   U19710 : XNOR2_X1 port map( A => n14996, B => n14995, ZN => n14997);
   U19711 : INV_X1 port map( A => n14999, ZN => n15005);
   U19712 : NAND2_X1 port map( A1 => n15001, A2 => n15000, ZN => n15002);
   U19713 : NOR2_X1 port map( A1 => n15002, A2 => n15132, ZN => n15003);
   U19714 : AOI21_X1 port map( B1 => n15005, B2 => n15004, A => n15003, ZN => 
                           n15006);
   U19715 : XNOR2_X1 port map( A => n15007, B => n15772, ZN => n15986);
   U19716 : XNOR2_X1 port map( A => n15986, B => n2206, ZN => n16658);
   U19717 : XNOR2_X1 port map( A => n16393, B => n15011, ZN => n15026);
   U19718 : AND2_X1 port map( A1 => n15447, A2 => n15445, ZN => n15012);
   U19719 : NAND2_X1 port map( A1 => n15320, A2 => n546, ZN => n15017);
   U19720 : NOR2_X1 port map( A1 => n15022, A2 => n15301, ZN => n15019);
   U19721 : NOR2_X1 port map( A1 => n15020, A2 => n15019, ZN => n15021);
   U19722 : NAND2_X1 port map( A1 => n15021, A2 => n15444, ZN => n15024);
   U19723 : NOR2_X1 port map( A1 => n15438, A2 => n15022, ZN => n15435);
   U19724 : NAND2_X1 port map( A1 => n15435, A2 => n15440, ZN => n15023);
   U19725 : XNOR2_X1 port map( A => n15026, B => n15965, ZN => n15044);
   U19727 : NAND3_X1 port map( A1 => n15037, A2 => n15036, A3 => n15293, ZN => 
                           n15038);
   U19729 : XNOR2_X1 port map( A => n15042, B => n16232, ZN => n16633);
   U19730 : INV_X1 port map( A => n16633, ZN => n15043);
   U19731 : INV_X1 port map( A => n15338, ZN => n15052);
   U19736 : XNOR2_X1 port map( A => n15780, B => n16618, ZN => n15057);
   U19737 : XNOR2_X1 port map( A => n15973, B => n15057, ZN => n15068);
   U19738 : INV_X1 port map( A => n15359, ZN => n15245);
   U19740 : NOR3_X1 port map( A1 => n15245, A2 => n15361, A3 => n28197, ZN => 
                           n15059);
   U19741 : NOR3_X1 port map( A1 => n15359, A2 => n14752, A3 => n15355, ZN => 
                           n15058);
   U19742 : NOR2_X1 port map( A1 => n15059, A2 => n15058, ZN => n15064);
   U19743 : NOR2_X1 port map( A1 => n15060, A2 => n15360, ZN => n15061);
   U19745 : XNOR2_X1 port map( A => n16619, B => n2385, ZN => n15066);
   U19746 : XNOR2_X1 port map( A => n16526, B => n16052, ZN => n15065);
   U19747 : XNOR2_X1 port map( A => n15066, B => n15065, ZN => n15067);
   U19748 : NAND3_X1 port map( A1 => n17435, A2 => n17438, A3 => n17440, ZN => 
                           n15069);
   U19749 : INV_X1 port map( A => n18304, ZN => n18475);
   U19750 : XNOR2_X1 port map( A => n15070, B => n2403, ZN => n15093);
   U19751 : NOR2_X1 port map( A1 => n15072, A2 => n15071, ZN => n15074);
   U19752 : NAND2_X1 port map( A1 => n15078, A2 => n15077, ZN => n15079);
   U19753 : NOR2_X1 port map( A1 => n15084, A2 => n15083, ZN => n15091);
   U19754 : OAI21_X1 port map( B1 => n15692, B2 => n323, A => n15691, ZN => 
                           n15090);
   U19756 : XNOR2_X1 port map( A => n16598, B => n15093, ZN => n15112);
   U19757 : NAND2_X1 port map( A1 => n15102, A2 => n15101, ZN => n15104);
   U19758 : INV_X1 port map( A => n16191, ZN => n15110);
   U19759 : NAND2_X1 port map( A1 => n15410, A2 => n15107, ZN => n15109);
   U19760 : XNOR2_X1 port map( A => n16365, B => n16398, ZN => n15741);
   U19761 : XNOR2_X1 port map( A => n15110, B => n15741, ZN => n15111);
   U19762 : INV_X1 port map( A => n17304, ZN => n17305);
   U19763 : XNOR2_X1 port map( A => n16477, B => n2509, ZN => n15133);
   U19764 : AND2_X1 port map( A1 => n15116, A2 => n15115, ZN => n15118);
   U19766 : NOR2_X1 port map( A1 => n13632, A2 => n15123, ZN => n15124);
   U19767 : AOI22_X1 port map( A1 => n15126, A2 => n15125, B1 => n15124, B2 => 
                           n1744, ZN => n15130);
   U19768 : NOR2_X1 port map( A1 => n551, A2 => n15127, ZN => n15128);
   U19769 : NAND2_X1 port map( A1 => n15132, A2 => n15128, ZN => n15129);
   U19770 : XNOR2_X1 port map( A => n15133, B => n16140, ZN => n15158);
   U19771 : INV_X1 port map( A => n15246, ZN => n15134);
   U19772 : OAI21_X1 port map( B1 => n15249, B2 => n15135, A => n15134, ZN => 
                           n15143);
   U19773 : AND2_X1 port map( A1 => n15135, A2 => n15138, ZN => n15142);
   U19774 : NAND2_X1 port map( A1 => n15246, A2 => n15136, ZN => n15140);
   U19775 : NAND2_X1 port map( A1 => n15138, A2 => n15137, ZN => n15139);
   U19776 : MUX2_X1 port map( A => n15140, B => n15139, S => n14733, Z => 
                           n15141);
   U19777 : OAI21_X1 port map( B1 => n15143, B2 => n15142, A => n15141, ZN => 
                           n16620);
   U19778 : MUX2_X1 port map( A => n15388, B => n15389, S => n15144, Z => 
                           n15146);
   U19779 : NOR3_X1 port map( A1 => n15395, A2 => n15391, A3 => n15387, ZN => 
                           n15148);
   U19780 : INV_X1 port map( A => n16196, ZN => n15156);
   U19781 : NAND3_X1 port map( A1 => n15155, A2 => n15152, A3 => n15384, ZN => 
                           n15153);
   U19782 : XNOR2_X1 port map( A => n15156, B => n16050, ZN => n15157);
   U19783 : AND2_X1 port map( A1 => n15161, A2 => n29153, ZN => n15162);
   U19784 : NOR2_X1 port map( A1 => n15171, A2 => n15170, ZN => n15172);
   U19785 : XNOR2_X1 port map( A => n16449, B => n1247, ZN => n15173);
   U19786 : XNOR2_X1 port map( A => n16203, B => n15173, ZN => n15214);
   U19787 : NAND2_X1 port map( A1 => n28462, A2 => n15180, ZN => n15178);
   U19788 : MUX2_X1 port map( A => n15178, B => n15177, S => n5635, Z => n15179
                           );
   U19789 : MUX2_X1 port map( A => n15184, B => n15183, S => n15182, Z => 
                           n15191);
   U19790 : NOR2_X1 port map( A1 => n15186, A2 => n15185, ZN => n15188);
   U19791 : OAI21_X1 port map( B1 => n15188, B2 => n15187, A => n15190, ZN => 
                           n15189);
   U19793 : XNOR2_X1 port map( A => n15850, B => n16407, ZN => n16554);
   U19794 : INV_X1 port map( A => n15192, ZN => n15198);
   U19795 : INV_X1 port map( A => n15193, ZN => n15197);
   U19796 : NAND2_X1 port map( A1 => n15195, A2 => n15194, ZN => n15196);
   U19797 : OAI211_X1 port map( C1 => n15199, C2 => n15198, A => n15197, B => 
                           n15196, ZN => n15200);
   U19798 : NAND2_X1 port map( A1 => n15201, A2 => n15200, ZN => n15205);
   U19799 : NAND2_X1 port map( A1 => n15202, A2 => n15208, ZN => n15203);
   U19801 : OAI211_X1 port map( C1 => n15209, C2 => n15208, A => n15207, B => 
                           n15206, ZN => n15210);
   U19802 : INV_X1 port map( A => n16404, ZN => n15212);
   U19803 : XNOR2_X1 port map( A => n16554, B => n15745, ZN => n15213);
   U19804 : XNOR2_X1 port map( A => n15213, B => n15214, ZN => n17012);
   U19806 : MUX2_X1 port map( A => n15216, B => n15215, S => n15217, Z => 
                           n15221);
   U19807 : INV_X1 port map( A => n15217, ZN => n15297);
   U19808 : NAND2_X1 port map( A1 => n15291, A2 => n14517, ZN => n15218);
   U19809 : AND2_X1 port map( A1 => n15219, A2 => n15218, ZN => n15220);
   U19810 : XNOR2_X1 port map( A => n16563, B => n15642, ZN => n16058);
   U19811 : NOR2_X1 port map( A1 => n15222, A2 => n15224, ZN => n15232);
   U19813 : OAI21_X1 port map( B1 => n15229, B2 => n15228, A => n15227, ZN => 
                           n15230);
   U19814 : NOR2_X1 port map( A1 => n15234, A2 => n15233, ZN => n15237);
   U19815 : AND2_X1 port map( A1 => n15334, A2 => n15333, ZN => n15236);
   U19816 : AND2_X1 port map( A1 => n15238, A2 => n15239, ZN => n15335);
   U19817 : INV_X1 port map( A => n16105, ZN => n15241);
   U19818 : XNOR2_X1 port map( A => n15241, B => n16271, ZN => n16218);
   U19819 : INV_X1 port map( A => n16218, ZN => n15242);
   U19820 : XNOR2_X1 port map( A => n16058, B => n15242, ZN => n15258);
   U19821 : XNOR2_X1 port map( A => n15788, B => n3321, ZN => n15256);
   U19822 : NAND2_X1 port map( A1 => n15355, A2 => n14752, ZN => n15244);
   U19823 : AOI21_X1 port map( B1 => n15247, B2 => n15246, A => n15252, ZN => 
                           n15255);
   U19824 : XNOR2_X1 port map( A => n15727, B => n16360, ZN => n16566);
   U19825 : INV_X1 port map( A => n16566, ZN => n16147);
   U19827 : NOR2_X1 port map( A1 => n15260, A2 => n15259, ZN => n15263);
   U19828 : XNOR2_X1 port map( A => n16388, B => n16586, ZN => n16031);
   U19829 : XNOR2_X1 port map( A => n16084, B => n16242, ZN => n15834);
   U19830 : XNOR2_X1 port map( A => n16031, B => n15834, ZN => n15281);
   U19831 : NAND2_X1 port map( A1 => n15312, A2 => n15311, ZN => n15955);
   U19832 : NAND2_X1 port map( A1 => n15956, A2 => n15955, ZN => n15273);
   U19833 : OR2_X1 port map( A1 => n15319, A2 => n15272, ZN => n15954);
   U19834 : OR3_X1 port map( A1 => n15276, A2 => n15275, A3 => n15274, ZN => 
                           n15278);
   U19836 : XNOR2_X1 port map( A => n16387, B => n15545, ZN => n16588);
   U19837 : NAND2_X1 port map( A1 => n17013, A2 => n16788, ZN => n15331);
   U19838 : OAI21_X1 port map( B1 => n15293, B2 => n15292, A => n15291, ZN => 
                           n15295);
   U19839 : NAND2_X1 port map( A1 => n15295, A2 => n15294, ZN => n15296);
   U19841 : INV_X1 port map( A => n16580, ZN => n15299);
   U19842 : XNOR2_X1 port map( A => n15299, B => n16575, ZN => n16123);
   U19843 : OAI21_X1 port map( B1 => n15302, B2 => n15301, A => n15300, ZN => 
                           n15305);
   U19844 : AOI22_X2 port map( A1 => n15305, A2 => n548, B1 => n15304, B2 => 
                           n15303, ZN => n16414);
   U19845 : XNOR2_X1 port map( A => n16414, B => n16579, ZN => n15762);
   U19846 : XNOR2_X1 port map( A => n16123, B => n15762, ZN => n15330);
   U19847 : NAND2_X1 port map( A1 => n15307, A2 => n15306, ZN => n15318);
   U19848 : OAI21_X1 port map( B1 => n15309, B2 => n15308, A => n15315, ZN => 
                           n15314);
   U19849 : OAI21_X1 port map( B1 => n15312, B2 => n15311, A => n15310, ZN => 
                           n15313);
   U19850 : NAND2_X1 port map( A1 => n15314, A2 => n15313, ZN => n15317);
   U19851 : OAI21_X1 port map( B1 => n15322, B2 => n15445, A => n15321, ZN => 
                           n15324);
   U19852 : NAND2_X1 port map( A1 => n15324, A2 => n546, ZN => n15325);
   U19853 : XNOR2_X1 port map( A => n16625, B => n16255, ZN => n16223);
   U19854 : XNOR2_X1 port map( A => n16456, B => n3029, ZN => n15328);
   U19855 : XNOR2_X1 port map( A => n16223, B => n15328, ZN => n15329);
   U19857 : MUX2_X2 port map( A => n15332, B => n15331, S => n29152, Z => 
                           n18011);
   U19858 : MUX2_X1 port map( A => n18476, B => n18475, S => n18011, Z => 
                           n15523);
   U19859 : NOR2_X1 port map( A1 => n15334, A2 => n15333, ZN => n15336);
   U19860 : XNOR2_X1 port map( A => n16170, B => n16366, ZN => n16484);
   U19861 : AOI21_X1 port map( B1 => n550, B2 => n15342, A => n15343, ZN => 
                           n15354);
   U19862 : AND2_X1 port map( A1 => n15345, A2 => n15344, ZN => n15347);
   U19863 : NAND4_X1 port map( A1 => n15349, A2 => n15348, A3 => n15347, A4 => 
                           n15346, ZN => n15350);
   U19864 : OAI21_X1 port map( B1 => n15351, B2 => n425, A => n15350, ZN => 
                           n15352);
   U19865 : AOI21_X1 port map( B1 => n15361, B2 => n15360, A => n15359, ZN => 
                           n15362);
   U19867 : XNOR2_X1 port map( A => n16279, B => n16230, ZN => n15994);
   U19868 : XNOR2_X1 port map( A => n16484, B => n15994, ZN => n15368);
   U19869 : XNOR2_X1 port map( A => n29084, B => n3508, ZN => n15365);
   U19870 : XNOR2_X1 port map( A => n15366, B => n15365, ZN => n15367);
   U19872 : NAND2_X1 port map( A1 => n15373, A2 => n426, ZN => n15375);
   U19873 : NAND2_X1 port map( A1 => n15375, A2 => n15374, ZN => n15377);
   U19874 : NAND2_X1 port map( A1 => n15381, A2 => n15380, ZN => n15386);
   U19875 : NAND2_X1 port map( A1 => n15386, A2 => n15385, ZN => n16373);
   U19876 : XNOR2_X1 port map( A => n16081, B => n16373, ZN => n15997);
   U19877 : XNOR2_X1 port map( A => n16082, B => n15997, ZN => n15397);
   U19878 : XNOR2_X1 port map( A => n15949, B => n2544, ZN => n15396);
   U19879 : OAI22_X1 port map( A1 => n15389, A2 => n15388, B1 => n15387, B2 => 
                           n15390, ZN => n15393);
   U19880 : NAND3_X1 port map( A1 => n15391, A2 => n15394, A3 => n15390, ZN => 
                           n15392);
   U19881 : XNOR2_X1 port map( A => n16589, B => n16377, ZN => n16468);
   U19882 : NAND2_X1 port map( A1 => n17298, A2 => n29072, ZN => n16831);
   U19883 : NAND2_X1 port map( A1 => n15402, A2 => n15400, ZN => n15403);
   U19884 : MUX2_X1 port map( A => n15403, B => n15402, S => n15401, Z => 
                           n15405);
   U19885 : OAI21_X1 port map( B1 => n3362, B2 => n15407, A => n15406, ZN => 
                           n15413);
   U19886 : NAND2_X1 port map( A1 => n15410, A2 => n15409, ZN => n15411);
   U19887 : NAND3_X1 port map( A1 => n15413, A2 => n15412, A3 => n15411, ZN => 
                           n15414);
   U19889 : XNOR2_X1 port map( A => n15914, B => n16649, ZN => n15789);
   U19890 : NAND3_X1 port map( A1 => n15420, A2 => n15423, A3 => n15417, ZN => 
                           n15418);
   U19891 : OAI211_X1 port map( C1 => n15423, C2 => n15422, A => n15421, B => 
                           n14575, ZN => n15424);
   U19892 : XNOR2_X1 port map( A => n16062, B => n16569, ZN => n16461);
   U19893 : INV_X1 port map( A => n16461, ZN => n15425);
   U19894 : XNOR2_X1 port map( A => n15425, B => n15789, ZN => n15429);
   U19895 : XNOR2_X1 port map( A => n16211, B => n2527, ZN => n15427);
   U19896 : XNOR2_X1 port map( A => n15426, B => n15427, ZN => n15428);
   U19898 : NAND2_X1 port map( A1 => n16831, A2 => n17411, ZN => n15522);
   U19899 : NAND2_X1 port map( A1 => n15444, A2 => n15435, ZN => n15443);
   U19900 : NOR2_X1 port map( A1 => n15438, A2 => n15437, ZN => n15441);
   U19901 : NOR2_X1 port map( A1 => n15437, A2 => n15436, ZN => n15439);
   U19902 : AOI22_X1 port map( A1 => n15441, A2 => n15440, B1 => n15439, B2 => 
                           n15438, ZN => n15442);
   U19903 : XNOR2_X1 port map( A => n16071, B => n16303, ZN => n15769);
   U19904 : MUX2_X1 port map( A => n15446, B => n15445, S => n15447, Z => 
                           n15450);
   U19905 : XNOR2_X1 port map( A => n16557, B => n16339, ZN => n16450);
   U19906 : INV_X1 port map( A => n16450, ZN => n15451);
   U19907 : XNOR2_X1 port map( A => n15769, B => n15451, ZN => n15455);
   U19908 : XNOR2_X1 port map( A => n16262, B => n3317, ZN => n15453);
   U19909 : XNOR2_X1 port map( A => n15852, B => n15453, ZN => n15454);
   U19910 : XNOR2_X1 port map( A => n16252, B => n29319, ZN => n15470);
   U19914 : INV_X1 port map( A => n16453, ZN => n15469);
   U19915 : XNOR2_X1 port map( A => n15469, B => n15470, ZN => n15483);
   U19916 : AOI21_X1 port map( B1 => n15473, B2 => n15472, A => n15471, ZN => 
                           n15479);
   U19917 : NAND2_X1 port map( A1 => n15475, A2 => n15474, ZN => n15477);
   U19918 : AOI21_X1 port map( B1 => n15477, B2 => n15476, A => n1848, ZN => 
                           n15478);
   U19919 : XNOR2_X1 port map( A => n16319, B => n15977, ZN => n15481);
   U19920 : XNOR2_X1 port map( A => n16257, B => n2511, ZN => n15480);
   U19921 : XNOR2_X1 port map( A => n15481, B => n15480, ZN => n15482);
   U19922 : XNOR2_X2 port map( A => n15483, B => n15482, ZN => n17413);
   U19923 : NAND2_X1 port map( A1 => n17411, A2 => n29072, ZN => n15484);
   U19924 : NAND2_X1 port map( A1 => n15486, A2 => n15485, ZN => n15488);
   U19925 : NAND2_X1 port map( A1 => n15491, A2 => n15489, ZN => n15487);
   U19926 : NAND3_X1 port map( A1 => n15491, A2 => n3748, A3 => n15489, ZN => 
                           n15492);
   U19928 : XNOR2_X1 port map( A => n16309, B => n2981, ZN => n15496);
   U19929 : XNOR2_X1 port map( A => n15496, B => n16619, ZN => n15508);
   U19930 : NAND2_X1 port map( A1 => n15497, A2 => n15500, ZN => n15507);
   U19931 : NAND3_X1 port map( A1 => n15503, A2 => n15499, A3 => n15498, ZN => 
                           n15505);
   U19932 : NAND2_X1 port map( A1 => n15500, A2 => n15502, ZN => n15501);
   U19933 : OAI211_X1 port map( C1 => n15503, C2 => n15502, A => n15501, B => 
                           n14923, ZN => n15504);
   U19934 : XNOR2_X1 port map( A => n16346, B => n16607, ZN => n16481);
   U19935 : INV_X1 port map( A => n16481, ZN => n15648);
   U19936 : XNOR2_X1 port map( A => n15648, B => n15508, ZN => n15521);
   U19937 : XNOR2_X1 port map( A => n16312, B => n16247, ZN => n15520);
   U19938 : INV_X1 port map( A => n15509, ZN => n15519);
   U19939 : OAI21_X1 port map( B1 => n5049, B2 => n15511, A => n15510, ZN => 
                           n15518);
   U19940 : NAND2_X1 port map( A1 => n15519, A2 => n15515, ZN => n15516);
   U19941 : XNOR2_X1 port map( A => n15928, B => n15520, ZN => n16098);
   U19943 : XNOR2_X1 port map( A => n16229, B => n16634, ZN => n16503);
   U19944 : XNOR2_X1 port map( A => n29084, B => n15992, ZN => n16190);
   U19945 : INV_X1 port map( A => n16190, ZN => n15525);
   U19946 : XNOR2_X1 port map( A => n15525, B => n16503, ZN => n15528);
   U19947 : XNOR2_X1 port map( A => n15865, B => n16284, ZN => n16369);
   U19948 : XNOR2_X1 port map( A => n16398, B => n2274, ZN => n15526);
   U19949 : XNOR2_X1 port map( A => n16369, B => n15526, ZN => n15527);
   U19950 : XNOR2_X1 port map( A => n15528, B => n15527, ZN => n15551);
   U19951 : XNOR2_X1 port map( A => n16619, B => n16434, ZN => n15530);
   U19952 : XNOR2_X1 port map( A => n16310, B => n26214, ZN => n15529);
   U19953 : XNOR2_X1 port map( A => n15530, B => n15529, ZN => n15534);
   U19954 : XNOR2_X1 port map( A => n16051, B => n16527, ZN => n15532);
   U19955 : XNOR2_X1 port map( A => n16017, B => n3661, ZN => n15531);
   U19956 : XNOR2_X1 port map( A => n15532, B => n15531, ZN => n15533);
   U19957 : XNOR2_X1 port map( A => n15533, B => n15534, ZN => n17349);
   U19958 : XNOR2_X1 port map( A => n16264, B => n15535, ZN => n16517);
   U19959 : INV_X1 port map( A => n16517, ZN => n15536);
   U19960 : INV_X1 port map( A => n16305, ZN => n15537);
   U19961 : XNOR2_X1 port map( A => n15537, B => n15850, ZN => n16340);
   U19962 : XNOR2_X1 port map( A => n16404, B => n3787, ZN => n15538);
   U19963 : XNOR2_X1 port map( A => n16340, B => n15538, ZN => n15539);
   U19964 : XNOR2_X1 port map( A => n16360, B => n16211, ZN => n15877);
   U19965 : XNOR2_X1 port map( A => n16271, B => n16146, ZN => n16532);
   U19966 : XNOR2_X1 port map( A => n16532, B => n15877, ZN => n15544);
   U19967 : XNOR2_X1 port map( A => n28579, B => n15642, ZN => n15542);
   U19968 : XNOR2_X1 port map( A => n16216, B => n22072, ZN => n15541);
   U19969 : XNOR2_X1 port map( A => n15542, B => n15541, ZN => n15543);
   U19970 : XNOR2_X1 port map( A => n15544, B => n15543, ZN => n17346);
   U19971 : INV_X1 port map( A => n17346, ZN => n17029);
   U19972 : XNOR2_X1 port map( A => n16510, B => n2402, ZN => n15546);
   U19973 : XNOR2_X1 port map( A => n16376, B => n15546, ZN => n15550);
   U19974 : XNOR2_X1 port map( A => n15949, B => n15760, ZN => n16208);
   U19975 : INV_X1 port map( A => n16208, ZN => n15548);
   U19976 : XNOR2_X1 port map( A => n16388, B => n16242, ZN => n15547);
   U19977 : XNOR2_X1 port map( A => n15548, B => n15547, ZN => n15549);
   U19978 : INV_X1 port map( A => n15551, ZN => n17192);
   U19979 : MUX2_X1 port map( A => n17029, B => n17347, S => n17192, Z => 
                           n15557);
   U19980 : INV_X1 port map( A => n16318, ZN => n15552);
   U19981 : XNOR2_X1 port map( A => n16414, B => n15552, ZN => n15553);
   U19982 : XNOR2_X1 port map( A => n16224, B => n15553, ZN => n15556);
   U19984 : XNOR2_X1 port map( A => n29151, B => n2984, ZN => n15554);
   U19985 : XNOR2_X1 port map( A => n16499, B => n15554, ZN => n15555);
   U19986 : XNOR2_X1 port map( A => n16568, B => n15790, ZN => n16214);
   U19987 : XNOR2_X1 port map( A => n15944, B => n16214, ZN => n15560);
   U19988 : XNOR2_X1 port map( A => n16185, B => n16295, ZN => n16102);
   U19989 : XNOR2_X1 port map( A => n16102, B => n15558, ZN => n15559);
   U19990 : XNOR2_X1 port map( A => n15561, B => n15965, ZN => n15564);
   U19991 : XNOR2_X1 port map( A => n16090, B => n15668, ZN => n15563);
   U19992 : XNOR2_X1 port map( A => n29571, B => n2411, ZN => n15562);
   U19993 : NOR2_X1 port map( A1 => n17338, A2 => n17340, ZN => n15582);
   U19994 : XNOR2_X1 port map( A => n16444, B => n15565, ZN => n16300);
   U19995 : XNOR2_X1 port map( A => n15900, B => n16519, ZN => n15566);
   U19996 : XNOR2_X1 port map( A => n16300, B => n15566, ZN => n15570);
   U19997 : XNOR2_X1 port map( A => n15772, B => n16070, ZN => n15567);
   U19998 : XNOR2_X1 port map( A => n15568, B => n15567, ZN => n15569);
   U19999 : XNOR2_X1 port map( A => n16165, B => n16312, ZN => n15572);
   U20000 : XNOR2_X1 port map( A => n15927, B => n3191, ZN => n15571);
   U20001 : XNOR2_X1 port map( A => n15572, B => n15571, ZN => n15574);
   U20002 : XNOR2_X1 port map( A => n15780, B => n16605, ZN => n16197);
   U20003 : XNOR2_X1 port map( A => n15973, B => n16197, ZN => n15573);
   U20004 : INV_X1 port map( A => n17155, ZN => n17200);
   U20005 : XNOR2_X1 port map( A => n16322, B => n16077, ZN => n15858);
   U20006 : XNOR2_X1 port map( A => n16578, B => n15654, ZN => n16221);
   U20007 : XNOR2_X1 port map( A => n15858, B => n16221, ZN => n15580);
   U20008 : XNOR2_X1 port map( A => n6454, B => n16498, ZN => n15578);
   U20009 : XNOR2_X1 port map( A => n15578, B => n15577, ZN => n15579);
   U20010 : INV_X1 port map( A => n17204, ZN => n17339);
   U20012 : XNOR2_X1 port map( A => n16085, B => n16329, ZN => n15872);
   U20013 : XNOR2_X1 port map( A => n15999, B => n16585, ZN => n16207);
   U20014 : XNOR2_X1 port map( A => n15872, B => n16207, ZN => n15587);
   U20015 : XNOR2_X1 port map( A => n15583, B => n15909, ZN => n15585);
   U20016 : XNOR2_X1 port map( A => n16241, B => n1119, ZN => n15584);
   U20017 : XNOR2_X1 port map( A => n15585, B => n15584, ZN => n15586);
   U20018 : MUX2_X1 port map( A => n28564, B => n17335, S => n17338, Z => 
                           n15588);
   U20019 : NOR2_X1 port map( A1 => n17336, A2 => n15588, ZN => n15589);
   U20020 : XNOR2_X1 port map( A => n16449, B => n16023, ZN => n15770);
   U20021 : XNOR2_X1 port map( A => n16557, B => n16519, ZN => n15591);
   U20022 : XNOR2_X1 port map( A => n15770, B => n15591, ZN => n15594);
   U20023 : XNOR2_X1 port map( A => n16303, B => n3607, ZN => n15592);
   U20024 : XNOR2_X1 port map( A => n15594, B => n15593, ZN => n17389);
   U20025 : XNOR2_X1 port map( A => n16456, B => n16038, ZN => n15782);
   U20026 : XNOR2_X1 port map( A => n16319, B => n16498, ZN => n15595);
   U20027 : XNOR2_X1 port map( A => n15782, B => n15595, ZN => n15599);
   U20028 : XNOR2_X1 port map( A => n16257, B => n26680, ZN => n15596);
   U20029 : XNOR2_X1 port map( A => n15597, B => n15596, ZN => n15598);
   U20030 : XNOR2_X1 port map( A => n15598, B => n15599, ZN => n16700);
   U20031 : NAND2_X1 port map( A1 => n17389, A2 => n29045, ZN => n17162);
   U20032 : XNOR2_X1 port map( A => n15802, B => n16467, ZN => n16032);
   U20033 : INV_X1 port map( A => n16238, ZN => n15711);
   U20034 : XNOR2_X1 port map( A => n15801, B => n15711, ZN => n15600);
   U20035 : XNOR2_X1 port map( A => n15600, B => n16032, ZN => n15604);
   U20036 : XNOR2_X1 port map( A => n16373, B => n16589, ZN => n15602);
   U20037 : XNOR2_X1 port map( A => n16241, B => n891, ZN => n15601);
   U20038 : XNOR2_X1 port map( A => n15602, B => n15601, ZN => n15603);
   U20039 : XNOR2_X1 port map( A => n15788, B => n16272, ZN => n15606);
   U20040 : XNOR2_X1 port map( A => n16569, B => n16534, ZN => n15605);
   U20041 : XNOR2_X1 port map( A => n15605, B => n15606, ZN => n15610);
   U20042 : INV_X1 port map( A => n2476, ZN => n24356);
   U20043 : XNOR2_X1 port map( A => n321, B => n24356, ZN => n15607);
   U20044 : XNOR2_X1 port map( A => n15608, B => n15607, ZN => n15609);
   U20045 : NAND2_X1 port map( A1 => n17386, A2 => n17385, ZN => n15611);
   U20046 : NAND2_X1 port map( A1 => n17162, A2 => n15611, ZN => n15616);
   U20047 : XNOR2_X1 port map( A => n16247, B => n2404, ZN => n15612);
   U20048 : XNOR2_X1 port map( A => n16309, B => n16607, ZN => n15613);
   U20049 : XNOR2_X1 port map( A => n15777, B => n15613, ZN => n15614);
   U20050 : XNOR2_X1 port map( A => n16483, B => n16233, ZN => n15698);
   U20052 : OAI21_X1 port map( B1 => n17382, B2 => n28497, A => n17385, ZN => 
                           n15615);
   U20054 : OAI21_X1 port map( B1 => n18493, B2 => n18292, A => n28633, ZN => 
                           n15737);
   U20057 : XNOR2_X1 port map( A => n16280, B => n16636, ZN => n15620);
   U20058 : XNOR2_X1 port map( A => n15620, B => n15619, ZN => n15624);
   U20059 : XNOR2_X1 port map( A => n16596, B => n16230, ZN => n15622);
   U20060 : XNOR2_X1 port map( A => n16398, B => n5633, ZN => n15621);
   U20061 : XNOR2_X1 port map( A => n15622, B => n15621, ZN => n15623);
   U20062 : XNOR2_X1 port map( A => n15624, B => n15623, ZN => n17355);
   U20064 : XNOR2_X1 port map( A => n16321, B => n16416, ZN => n15859);
   U20065 : XNOR2_X1 port map( A => n15625, B => n15859, ZN => n15628);
   U20066 : XNOR2_X1 port map( A => n16256, B => n16625, ZN => n15822);
   U20067 : XNOR2_X1 port map( A => n16578, B => n27231, ZN => n15626);
   U20068 : XNOR2_X1 port map( A => n15822, B => n15626, ZN => n15627);
   U20069 : XNOR2_X1 port map( A => n16081, B => n16641, ZN => n16240);
   U20070 : XNOR2_X1 port map( A => n28585, B => n16471, ZN => n15629);
   U20071 : XNOR2_X1 port map( A => n16240, B => n15629, ZN => n15633);
   U20072 : XNOR2_X1 port map( A => n15631, B => n15630, ZN => n15632);
   U20073 : XNOR2_X1 port map( A => n15633, B => n15632, ZN => n17357);
   U20074 : MUX2_X1 port map( A => n17355, B => n17359, S => n17357, Z => 
                           n15647);
   U20075 : XNOR2_X1 port map( A => n16404, B => n3662, ZN => n15634);
   U20076 : INV_X1 port map( A => n15849, ZN => n16408);
   U20077 : XNOR2_X1 port map( A => n16408, B => n16556, ZN => n15636);
   U20078 : XNOR2_X1 port map( A => n15636, B => n16654, ZN => n15637);
   U20080 : NOR2_X1 port map( A1 => n17354, A2 => n17359, ZN => n17198);
   U20081 : XNOR2_X1 port map( A => n16605, B => n16434, ZN => n15639);
   U20082 : XNOR2_X1 port map( A => n15928, B => n16618, ZN => n16246);
   U20083 : INV_X1 port map( A => n16620, ZN => n16095);
   U20084 : XNOR2_X1 port map( A => n16436, B => n16095, ZN => n15975);
   U20085 : INV_X1 port map( A => n17356, ZN => n17196);
   U20086 : NAND2_X1 port map( A1 => n17198, A2 => n17196, ZN => n15646);
   U20087 : XNOR2_X1 port map( A => n15914, B => n15817, ZN => n16269);
   U20088 : INV_X1 port map( A => n16269, ZN => n15641);
   U20089 : XNOR2_X1 port map( A => n16291, B => n16568, ZN => n15640);
   U20090 : XNOR2_X1 port map( A => n16105, B => n3554, ZN => n15643);
   U20091 : XNOR2_X1 port map( A => n15644, B => n15643, ZN => n15645);
   U20092 : INV_X1 port map( A => n17030, ZN => n16953);
   U20093 : INV_X1 port map( A => n18489, ZN => n17674);
   U20094 : NOR2_X1 port map( A1 => n18487, A2 => n17674, ZN => n15736);
   U20095 : XNOR2_X1 port map( A => n15649, B => n15648, ZN => n15653);
   U20096 : XNOR2_X1 port map( A => n29525, B => n15927, ZN => n15651);
   U20097 : XNOR2_X1 port map( A => n16247, B => n26825, ZN => n15650);
   U20098 : XNOR2_X1 port map( A => n15651, B => n15650, ZN => n15652);
   U20099 : XNOR2_X1 port map( A => n28557, B => n6449, ZN => n15656);
   U20100 : XNOR2_X1 port map( A => n16574, B => n15654, ZN => n15655);
   U20101 : XNOR2_X1 port map( A => n15656, B => n15655, ZN => n15660);
   U20102 : INV_X1 port map( A => n2577, ZN => n25902);
   U20103 : XNOR2_X1 port map( A => n16257, B => n25902, ZN => n15657);
   U20104 : XNOR2_X1 port map( A => n15658, B => n15657, ZN => n15659);
   U20105 : XNOR2_X1 port map( A => n16426, B => n16272, ZN => n16107);
   U20106 : INV_X1 port map( A => n16107, ZN => n15661);
   U20107 : INV_X1 port map( A => n16062, ZN => n16143);
   U20108 : XNOR2_X1 port map( A => n16143, B => n16563, ZN => n16359);
   U20109 : XNOR2_X1 port map( A => n16359, B => n15661, ZN => n15665);
   U20110 : XNOR2_X1 port map( A => n16294, B => n15790, ZN => n15663);
   U20111 : XNOR2_X1 port map( A => n16569, B => n1927, ZN => n15662);
   U20112 : XNOR2_X1 port map( A => n15663, B => n15662, ZN => n15664);
   U20113 : XNOR2_X1 port map( A => n15665, B => n15664, ZN => n16762);
   U20115 : INV_X1 port map( A => n16484, ZN => n15667);
   U20116 : XNOR2_X1 port map( A => n16233, B => n16365, ZN => n15666);
   U20117 : XNOR2_X1 port map( A => n15667, B => n15666, ZN => n15672);
   U20118 : XNOR2_X1 port map( A => n16399, B => n15668, ZN => n15670);
   U20119 : XNOR2_X1 port map( A => n15989, B => n3256, ZN => n15669);
   U20120 : XNOR2_X1 port map( A => n15670, B => n15669, ZN => n15671);
   U20121 : INV_X1 port map( A => n15772, ZN => n16199);
   U20122 : XNOR2_X1 port map( A => n15900, B => n15673, ZN => n15677);
   U20123 : XNOR2_X1 port map( A => n16262, B => n2961, ZN => n15674);
   U20124 : XNOR2_X1 port map( A => n15674, B => n16405, ZN => n15675);
   U20125 : XNOR2_X1 port map( A => n15675, B => n16450, ZN => n15676);
   U20126 : XNOR2_X1 port map( A => n15676, B => n15677, ZN => n16943);
   U20128 : NAND2_X1 port map( A1 => n17549, A2 => n16944, ZN => n16947);
   U20129 : INV_X1 port map( A => n16947, ZN => n15686);
   U20130 : XNOR2_X1 port map( A => n16238, B => n28597, ZN => n15680);
   U20131 : INV_X1 port map( A => n15999, ZN => n15678);
   U20132 : XNOR2_X1 port map( A => n15678, B => n16586, ZN => n15679);
   U20133 : XNOR2_X1 port map( A => n15679, B => n15680, ZN => n15684);
   U20134 : XNOR2_X1 port map( A => n16589, B => n3232, ZN => n15681);
   U20135 : XNOR2_X1 port map( A => n15682, B => n15681, ZN => n15683);
   U20136 : INV_X1 port map( A => n17548, ZN => n17239);
   U20137 : OAI21_X1 port map( B1 => n15686, B2 => n15685, A => n17552, ZN => 
                           n15687);
   U20138 : INV_X1 port map( A => n18490, ZN => n18015);
   U20141 : XNOR2_X1 port map( A => n16395, B => n1849, ZN => n15696);
   U20142 : XNOR2_X1 port map( A => n16043, B => n16393, ZN => n16504);
   U20143 : XNOR2_X1 port map( A => n15696, B => n16504, ZN => n15700);
   U20144 : XNOR2_X1 port map( A => n16284, B => n3462, ZN => n15697);
   U20145 : XNOR2_X1 port map( A => n15698, B => n15697, ZN => n15699);
   U20147 : INV_X1 port map( A => n17368, ZN => n17366);
   U20148 : XNOR2_X1 port map( A => n16495, B => n15701, ZN => n16415);
   U20149 : XNOR2_X1 port map( A => n16160, B => n16494, ZN => n16577);
   U20150 : XNOR2_X1 port map( A => n16577, B => n16415, ZN => n15705);
   U20151 : XNOR2_X1 port map( A => n16257, B => n3164, ZN => n15702);
   U20152 : XNOR2_X1 port map( A => n15703, B => n15702, ZN => n15704);
   U20153 : XNOR2_X1 port map( A => n15705, B => n15704, ZN => n17361);
   U20154 : XNOR2_X1 port map( A => n15706, B => n15971, ZN => n16433);
   U20155 : INV_X1 port map( A => n16433, ZN => n15707);
   U20156 : XNOR2_X1 port map( A => n15707, B => n259, ZN => n15710);
   U20157 : XNOR2_X1 port map( A => n16606, B => n16310, ZN => n16166);
   U20158 : XNOR2_X1 port map( A => n16247, B => n2389, ZN => n15708);
   U20159 : XNOR2_X1 port map( A => n16166, B => n15708, ZN => n15709);
   U20160 : INV_X1 port map( A => n17365, ZN => n17369);
   U20161 : XNOR2_X1 port map( A => n15711, B => n16509, ZN => n15712);
   U20162 : XNOR2_X1 port map( A => n15712, B => n16591, ZN => n15716);
   U20163 : XNOR2_X1 port map( A => n16387, B => n16467, ZN => n15714);
   U20164 : XNOR2_X1 port map( A => n16332, B => n1887, ZN => n15713);
   U20165 : XNOR2_X1 port map( A => n15714, B => n15713, ZN => n15715);
   U20166 : XNOR2_X1 port map( A => n15716, B => n15715, ZN => n15731);
   U20167 : XNOR2_X1 port map( A => n16558, B => n16407, ZN => n15718);
   U20168 : XNOR2_X1 port map( A => n16024, B => n16409, ZN => n16521);
   U20169 : XNOR2_X1 port map( A => n15718, B => n16521, ZN => n15722);
   U20170 : XNOR2_X1 port map( A => n16305, B => n3622, ZN => n15719);
   U20171 : XNOR2_X1 port map( A => n15720, B => n15719, ZN => n15721);
   U20173 : XNOR2_X1 port map( A => n16422, B => n15723, ZN => n16533);
   U20174 : INV_X1 port map( A => n16533, ZN => n15726);
   U20175 : XNOR2_X1 port map( A => n16059, B => n3081, ZN => n15724);
   U20176 : XNOR2_X1 port map( A => n15724, B => n16272, ZN => n15725);
   U20177 : XNOR2_X1 port map( A => n15725, B => n15726, ZN => n15730);
   U20178 : XNOR2_X1 port map( A => n28579, B => n16427, ZN => n15728);
   U20179 : INV_X1 port map( A => n16564, ZN => n16213);
   U20180 : XNOR2_X1 port map( A => n16213, B => n15728, ZN => n15729);
   U20181 : XNOR2_X1 port map( A => n15730, B => n15729, ZN => n17234);
   U20182 : INV_X1 port map( A => n28632, ZN => n18486);
   U20183 : OAI211_X1 port map( C1 => n18015, C2 => n18489, A => n15734, B => 
                           n18486, ZN => n15735);
   U20184 : XNOR2_X1 port map( A => n19495, B => n19103, ZN => n19650);
   U20185 : XNOR2_X1 port map( A => n15668, B => n2541, ZN => n15740);
   U20186 : XNOR2_X1 port map( A => n15738, B => n15992, ZN => n15739);
   U20187 : XNOR2_X1 port map( A => n15740, B => n15739, ZN => n15743);
   U20188 : XNOR2_X1 port map( A => n16397, B => n15741, ZN => n15742);
   U20189 : XNOR2_X1 port map( A => n16443, B => n1919, ZN => n15744);
   U20190 : XNOR2_X1 port map( A => n15744, B => n15982, ZN => n15747);
   U20191 : INV_X1 port map( A => n15745, ZN => n15746);
   U20192 : XNOR2_X1 port map( A => n15747, B => n15746, ZN => n15749);
   U20193 : XNOR2_X1 port map( A => n16406, B => n15900, ZN => n15748);
   U20194 : XNOR2_X1 port map( A => n16527, B => n16606, ZN => n16432);
   U20195 : XNOR2_X1 port map( A => n16432, B => n16050, ZN => n15753);
   U20196 : XNOR2_X1 port map( A => n16017, B => n16476, ZN => n15751);
   U20197 : XNOR2_X1 port map( A => n15927, B => n25992, ZN => n15750);
   U20198 : XNOR2_X1 port map( A => n15751, B => n15750, ZN => n15752);
   U20199 : XNOR2_X1 port map( A => n15753, B => n15752, ZN => n16918);
   U20200 : NOR2_X1 port map( A1 => n17317, A2 => n16918, ZN => n15754);
   U20201 : AOI21_X1 port map( B1 => n17316, B2 => n17317, A => n15754, ZN => 
                           n15768);
   U20202 : INV_X1 port map( A => n16058, ZN => n15755);
   U20203 : XNOR2_X1 port map( A => n15755, B => n16424, ZN => n15759);
   U20204 : XNOR2_X1 port map( A => n16294, B => n16216, ZN => n15757);
   U20205 : XNOR2_X1 port map( A => n16059, B => n3722, ZN => n15756);
   U20206 : XNOR2_X1 port map( A => n15757, B => n15756, ZN => n15758);
   U20207 : XNOR2_X1 port map( A => n16467, B => n3386, ZN => n15761);
   U20208 : INV_X1 port map( A => n15760, ZN => n16000);
   U20210 : XNOR2_X1 port map( A => n16418, B => n15762, ZN => n15766);
   U20211 : XNOR2_X1 port map( A => n15764, B => n15763, ZN => n15765);
   U20212 : XNOR2_X1 port map( A => n15766, B => n15765, ZN => n17312);
   U20213 : INV_X1 port map( A => n17312, ZN => n17560);
   U20214 : INV_X1 port map( A => n15769, ZN => n15771);
   U20215 : XNOR2_X1 port map( A => n16408, B => n15772, ZN => n15774);
   U20216 : XNOR2_X1 port map( A => n16444, B => n3491, ZN => n15773);
   U20217 : XNOR2_X1 port map( A => n15774, B => n15773, ZN => n15775);
   U20218 : XNOR2_X1 port map( A => n15928, B => n16052, ZN => n15778);
   U20219 : XNOR2_X1 port map( A => n16309, B => n15780, ZN => n16617);
   U20220 : XNOR2_X1 port map( A => n15781, B => n16319, ZN => n16629);
   U20221 : INV_X1 port map( A => n16629, ZN => n16011);
   U20222 : XNOR2_X1 port map( A => n16011, B => n15782, ZN => n15786);
   U20223 : XNOR2_X1 port map( A => n16416, B => n16252, ZN => n15784);
   U20224 : XNOR2_X1 port map( A => n16323, B => n2973, ZN => n15783);
   U20225 : XNOR2_X1 port map( A => n15784, B => n15783, ZN => n15785);
   U20227 : INV_X1 port map( A => n17541, ZN => n15787);
   U20228 : XNOR2_X1 port map( A => n16296, B => n15788, ZN => n16462);
   U20229 : XNOR2_X1 port map( A => n15789, B => n16462, ZN => n15794);
   U20230 : XNOR2_X1 port map( A => n16421, B => n15790, ZN => n15792);
   U20231 : XNOR2_X1 port map( A => n321, B => n1133, ZN => n15791);
   U20232 : XNOR2_X1 port map( A => n15792, B => n15791, ZN => n15793);
   U20233 : INV_X1 port map( A => n15994, ZN => n15795);
   U20234 : XNOR2_X1 port map( A => n15795, B => n15796, ZN => n15800);
   U20235 : XNOR2_X1 port map( A => n16400, B => n16283, ZN => n15798);
   U20236 : XNOR2_X1 port map( A => n15989, B => n3035, ZN => n15797);
   U20237 : XNOR2_X1 port map( A => n15798, B => n15797, ZN => n15799);
   U20238 : OAI22_X1 port map( A1 => n17542, A2 => n17545, B1 => n17543, B2 => 
                           n17540, ZN => n15807);
   U20239 : XNOR2_X1 port map( A => n15801, B => n16328, ZN => n16472);
   U20240 : XNOR2_X1 port map( A => n16472, B => n15997, ZN => n15806);
   U20241 : INV_X1 port map( A => n28585, ZN => n16386);
   U20242 : XNOR2_X1 port map( A => n15802, B => n16386, ZN => n15804);
   U20243 : XNOR2_X1 port map( A => n15999, B => n28294, ZN => n15803);
   U20244 : XNOR2_X1 port map( A => n15804, B => n15803, ZN => n15805);
   U20245 : XNOR2_X1 port map( A => n15806, B => n15805, ZN => n17539);
   U20246 : INV_X1 port map( A => n17539, ZN => n17213);
   U20247 : NAND2_X1 port map( A1 => n15807, A2 => n17213, ZN => n15809);
   U20248 : NAND2_X1 port map( A1 => n17217, A2 => n17545, ZN => n15808);
   U20250 : INV_X1 port map( A => n17413, ZN => n17297);
   U20251 : INV_X1 port map( A => n17414, ZN => n17300);
   U20252 : NAND2_X1 port map( A1 => n15812, A2 => n17300, ZN => n15816);
   U20253 : NAND3_X1 port map( A1 => n17298, A2 => n17297, A3 => n17414, ZN => 
                           n15814);
   U20254 : NAND2_X1 port map( A1 => n17298, A2 => n17411, ZN => n15813);
   U20255 : AND2_X1 port map( A1 => n15814, A2 => n15813, ZN => n15815);
   U20256 : NAND2_X1 port map( A1 => n15816, A2 => n15815, ZN => n17926);
   U20257 : INV_X1 port map( A => n17926, ZN => n18059);
   U20258 : XNOR2_X1 port map( A => n16360, B => n15817, ZN => n15819);
   U20259 : XNOR2_X1 port map( A => n16059, B => n3276, ZN => n15818);
   U20260 : XNOR2_X1 port map( A => n15819, B => n15818, ZN => n15821);
   U20262 : XNOR2_X1 port map( A => n15822, B => n29630, ZN => n15827);
   U20263 : XNOR2_X1 port map( A => n29151, B => n3654, ZN => n15824);
   U20264 : XNOR2_X1 port map( A => n15825, B => n15824, ZN => n15826);
   U20265 : XNOR2_X1 port map( A => n16203, B => n16134, ZN => n15832);
   U20266 : XNOR2_X1 port map( A => n15828, B => n15850, ZN => n15830);
   U20267 : XNOR2_X1 port map( A => n16443, B => n3695, ZN => n15829);
   U20268 : XNOR2_X1 port map( A => n15830, B => n15829, ZN => n15831);
   U20269 : INV_X1 port map( A => n16119, ZN => n15833);
   U20270 : XNOR2_X1 port map( A => n15833, B => n15834, ZN => n15838);
   U20271 : XNOR2_X1 port map( A => n16641, B => n3114, ZN => n15835);
   U20272 : XNOR2_X1 port map( A => n15836, B => n15835, ZN => n15837);
   U20273 : XNOR2_X1 port map( A => n16191, B => n16116, ZN => n15842);
   U20274 : XNOR2_X1 port map( A => n16483, B => n16232, ZN => n15840);
   U20275 : XNOR2_X1 port map( A => n15865, B => n3087, ZN => n15839);
   U20276 : XNOR2_X1 port map( A => n15840, B => n15839, ZN => n15841);
   U20277 : INV_X1 port map( A => n17554, ZN => n16911);
   U20278 : XNOR2_X1 port map( A => n16196, B => n16138, ZN => n15846);
   U20279 : XNOR2_X1 port map( A => n16618, B => n3661, ZN => n15844);
   U20280 : XNOR2_X1 port map( A => n16476, B => n900, ZN => n15843);
   U20281 : XNOR2_X1 port map( A => n15844, B => n15843, ZN => n15845);
   U20282 : INV_X1 port map( A => n16908, ZN => n17221);
   U20283 : OAI21_X1 port map( B1 => n18298, B2 => n18059, A => n29561, ZN => 
                           n15938);
   U20285 : XNOR2_X1 port map( A => n15851, B => n15850, ZN => n15853);
   U20286 : XNOR2_X1 port map( A => n16519, B => n16070, ZN => n15854);
   U20287 : XNOR2_X1 port map( A => n15855, B => n15977, ZN => n15857);
   U20288 : XNOR2_X1 port map( A => n29151, B => n2350, ZN => n15856);
   U20289 : XNOR2_X1 port map( A => n15857, B => n15856, ZN => n15861);
   U20290 : XNOR2_X1 port map( A => n15859, B => n15858, ZN => n15860);
   U20291 : XNOR2_X1 port map( A => n15863, B => n15862, ZN => n16237);
   U20292 : XNOR2_X1 port map( A => n15966, B => n28327, ZN => n15864);
   U20293 : XNOR2_X1 port map( A => n15864, B => n16090, ZN => n15867);
   U20294 : XNOR2_X1 port map( A => n15865, B => n16400, ZN => n15866);
   U20295 : XNOR2_X1 port map( A => n15867, B => n15866, ZN => n15868);
   U20296 : INV_X1 port map( A => n15949, ZN => n15870);
   U20298 : XNOR2_X1 port map( A => n15872, B => n15871, ZN => n15876);
   U20299 : XNOR2_X1 port map( A => n16241, B => n2602, ZN => n15873);
   U20300 : XNOR2_X1 port map( A => n15874, B => n15873, ZN => n15875);
   U20301 : NAND2_X1 port map( A1 => n1166, A2 => n4118, ZN => n15884);
   U20302 : INV_X1 port map( A => n15877, ZN => n15879);
   U20303 : XNOR2_X1 port map( A => n15878, B => n15879, ZN => n15883);
   U20304 : XNOR2_X1 port map( A => n16295, B => n16421, ZN => n15881);
   U20305 : XNOR2_X1 port map( A => n16534, B => n3372, ZN => n15880);
   U20306 : XNOR2_X1 port map( A => n15881, B => n15880, ZN => n15882);
   U20307 : INV_X1 port map( A => n29098, ZN => n17037);
   U20308 : XNOR2_X1 port map( A => n1967, B => n3661, ZN => n15886);
   U20309 : XNOR2_X1 port map( A => n16619, B => n16165, ZN => n15885);
   U20310 : XNOR2_X1 port map( A => n15886, B => n15885, ZN => n15891);
   U20311 : XNOR2_X1 port map( A => n15887, B => n16312, ZN => n15889);
   U20312 : XNOR2_X1 port map( A => n16313, B => n2505, ZN => n15888);
   U20313 : XNOR2_X1 port map( A => n15889, B => n15888, ZN => n15890);
   U20314 : XNOR2_X1 port map( A => n15891, B => n15890, ZN => n17566);
   U20315 : INV_X1 port map( A => n17566, ZN => n17038);
   U20317 : XNOR2_X1 port map( A => n16154, B => n15893, ZN => n15902);
   U20318 : XNOR2_X1 port map( A => n15894, B => n27956, ZN => n15897);
   U20319 : XNOR2_X1 port map( A => n15895, B => n27956, ZN => n15896);
   U20320 : XNOR2_X1 port map( A => n15898, B => n16407, ZN => n15899);
   U20321 : XNOR2_X1 port map( A => n15899, B => n15900, ZN => n15901);
   U20322 : XNOR2_X1 port map( A => n15902, B => n15901, ZN => n17571);
   U20323 : XNOR2_X1 port map( A => n16162, B => n15903, ZN => n15907);
   U20324 : XNOR2_X1 port map( A => n16575, B => n16252, ZN => n15905);
   U20325 : XNOR2_X1 port map( A => n15905, B => n15904, ZN => n15906);
   U20326 : XNOR2_X1 port map( A => n15906, B => n15907, ZN => n16904);
   U20327 : NAND2_X1 port map( A1 => n17571, A2 => n16904, ZN => n17404);
   U20328 : INV_X1 port map( A => n16179, ZN => n15908);
   U20329 : XNOR2_X1 port map( A => n15908, B => n16375, ZN => n15913);
   U20330 : XNOR2_X1 port map( A => n16387, B => n16081, ZN => n15911);
   U20331 : XNOR2_X1 port map( A => n15909, B => n3598, ZN => n15910);
   U20332 : XNOR2_X1 port map( A => n15911, B => n15910, ZN => n15912);
   U20333 : XNOR2_X1 port map( A => n15914, B => n16294, ZN => n15915);
   U20334 : XNOR2_X1 port map( A => n16183, B => n15915, ZN => n15918);
   U20335 : XNOR2_X1 port map( A => n16427, B => n3643, ZN => n15916);
   U20336 : XNOR2_X1 port map( A => n16362, B => n15916, ZN => n15917);
   U20337 : XNOR2_X1 port map( A => n15917, B => n15918, ZN => n17405);
   U20338 : NAND2_X1 port map( A1 => n17572, A2 => n17405, ZN => n17403);
   U20343 : XNOR2_X1 port map( A => n16395, B => n15668, ZN => n15920);
   U20345 : XNOR2_X1 port map( A => n16230, B => n3336, ZN => n15922);
   U20346 : XNOR2_X1 port map( A => n16367, B => n15922, ZN => n15923);
   U20347 : XNOR2_X1 port map( A => n15924, B => n15923, ZN => n16822);
   U20348 : XNOR2_X1 port map( A => n16310, B => n2523, ZN => n15926);
   U20349 : INV_X1 port map( A => n15971, ZN => n15925);
   U20350 : XNOR2_X1 port map( A => n15928, B => n15927, ZN => n15929);
   U20351 : XNOR2_X1 port map( A => n15929, B => n15777, ZN => n15930);
   U20352 : INV_X1 port map( A => n17572, ZN => n17320);
   U20353 : NAND3_X1 port map( A1 => n17707, A2 => n17570, A3 => n17320, ZN => 
                           n15933);
   U20354 : NAND3_X1 port map( A1 => n17707, A2 => n16904, A3 => n17320, ZN => 
                           n15932);
   U20355 : NOR2_X1 port map( A1 => n18298, A2 => n1861, ZN => n15935);
   U20356 : INV_X1 port map( A => n18060, ZN => n17928);
   U20357 : NAND2_X1 port map( A1 => n15935, A2 => n17928, ZN => n15936);
   U20359 : XNOR2_X1 port map( A => n15940, B => n21865, ZN => n15941);
   U20360 : XNOR2_X1 port map( A => n16654, B => n16407, ZN => n15942);
   U20361 : XNOR2_X1 port map( A => n16105, B => n16211, ZN => n16648);
   U20362 : INV_X1 port map( A => n16648, ZN => n15943);
   U20363 : XNOR2_X1 port map( A => n15943, B => n15944, ZN => n15946);
   U20364 : INV_X1 port map( A => n16514, ZN => n15947);
   U20365 : XNOR2_X1 port map( A => n15947, B => n15948, ZN => n15963);
   U20366 : XNOR2_X1 port map( A => n15949, B => n16084, ZN => n15961);
   U20367 : INV_X1 port map( A => n15955, ZN => n15950);
   U20368 : NAND2_X1 port map( A1 => n15950, A2 => n3635, ZN => n15952);
   U20369 : INV_X1 port map( A => n15954, ZN => n15951);
   U20370 : MUX2_X1 port map( A => n15952, B => n3635, S => n15951, Z => n15959
                           );
   U20371 : INV_X1 port map( A => n15956, ZN => n15953);
   U20372 : NAND3_X1 port map( A1 => n15954, A2 => n15953, A3 => n3635, ZN => 
                           n15958);
   U20373 : INV_X1 port map( A => n3635, ZN => n27384);
   U20374 : NAND3_X1 port map( A1 => n15956, A2 => n27384, A3 => n15955, ZN => 
                           n15957);
   U20375 : NAND3_X1 port map( A1 => n15959, A2 => n15958, A3 => n15957, ZN => 
                           n15960);
   U20376 : XNOR2_X1 port map( A => n15961, B => n15960, ZN => n15962);
   U20377 : XNOR2_X1 port map( A => n15963, B => n15962, ZN => n16764);
   U20378 : INV_X1 port map( A => n16764, ZN => n17278);
   U20379 : XNOR2_X1 port map( A => n15965, B => n16636, ZN => n15970);
   U20380 : XNOR2_X1 port map( A => n29084, B => n3196, ZN => n15967);
   U20381 : XNOR2_X1 port map( A => n16395, B => n15967, ZN => n15968);
   U20382 : XNOR2_X1 port map( A => n15968, B => n16506, ZN => n15969);
   U20383 : XNOR2_X1 port map( A => n15971, B => n1184, ZN => n15972);
   U20384 : INV_X1 port map( A => n16017, ZN => n15974);
   U20385 : XNOR2_X1 port map( A => n15974, B => n16619, ZN => n16198);
   U20386 : XNOR2_X1 port map( A => n16575, B => n16498, ZN => n15976);
   U20387 : XNOR2_X1 port map( A => n16497, B => n15976, ZN => n15979);
   U20388 : XNOR2_X1 port map( A => n15977, B => n3660, ZN => n15978);
   U20389 : XNOR2_X1 port map( A => n16071, B => n15982, ZN => n15984);
   U20390 : INV_X1 port map( A => n16557, ZN => n15983);
   U20391 : XNOR2_X1 port map( A => n15983, B => n16070, ZN => n16156);
   U20392 : XNOR2_X1 port map( A => n16156, B => n15984, ZN => n15988);
   U20393 : XNOR2_X1 port map( A => n16303, B => n3180, ZN => n15985);
   U20394 : XNOR2_X1 port map( A => n15986, B => n15985, ZN => n15987);
   U20395 : XNOR2_X1 port map( A => n15987, B => n15988, ZN => n17255);
   U20396 : XNOR2_X1 port map( A => n15989, B => n26531, ZN => n15990);
   U20397 : XNOR2_X1 port map( A => n15991, B => n15990, ZN => n15996);
   U20398 : XNOR2_X1 port map( A => n16170, B => n15992, ZN => n15993);
   U20399 : XNOR2_X1 port map( A => n15994, B => n15993, ZN => n15995);
   U20401 : INV_X1 port map( A => n17248, ZN => n17016);
   U20402 : XNOR2_X1 port map( A => n15998, B => n15997, ZN => n16004);
   U20403 : XNOR2_X1 port map( A => n16641, B => n1923, ZN => n16002);
   U20404 : XNOR2_X1 port map( A => n15999, B => n16000, ZN => n16001);
   U20405 : XNOR2_X1 port map( A => n16002, B => n16001, ZN => n16003);
   U20406 : XNOR2_X1 port map( A => n16004, B => n16003, ZN => n17250);
   U20407 : INV_X1 port map( A => n17250, ZN => n17017);
   U20408 : XNOR2_X1 port map( A => n16569, B => n16216, ZN => n16006);
   U20409 : XNOR2_X1 port map( A => n15914, B => n16006, ZN => n16007);
   U20410 : OAI21_X1 port map( B1 => n17016, B2 => n17017, A => n16977, ZN => 
                           n16008);
   U20411 : XNOR2_X1 port map( A => n16009, B => n16077, ZN => n16159);
   U20412 : INV_X1 port map( A => n16159, ZN => n16010);
   U20413 : XNOR2_X1 port map( A => n16010, B => n16011, ZN => n16016);
   U20414 : XNOR2_X1 port map( A => n16252, B => n16012, ZN => n16014);
   U20415 : XNOR2_X1 port map( A => n16256, B => n5490, ZN => n16013);
   U20416 : XNOR2_X1 port map( A => n16014, B => n16013, ZN => n16015);
   U20417 : AOI22_X1 port map( A1 => n17251, A2 => n17249, B1 => n16977, B2 => 
                           n29503, ZN => n17015);
   U20418 : XNOR2_X1 port map( A => n16246, B => n16617, ZN => n16021);
   U20419 : XNOR2_X1 port map( A => n16017, B => n16165, ZN => n16019);
   U20420 : XNOR2_X1 port map( A => n16607, B => n2441, ZN => n16018);
   U20421 : XNOR2_X1 port map( A => n16019, B => n16018, ZN => n16020);
   U20422 : OR2_X1 port map( A1 => n17015, A2 => n6539, ZN => n16022);
   U20424 : XNOR2_X1 port map( A => n16264, B => n16023, ZN => n16026);
   U20427 : XNOR2_X1 port map( A => n16404, B => n27298, ZN => n16027);
   U20428 : XNOR2_X1 port map( A => n16028, B => n16027, ZN => n16029);
   U20430 : INV_X1 port map( A => n16031, ZN => n16033);
   U20431 : XNOR2_X1 port map( A => n16033, B => n16032, ZN => n16037);
   U20432 : XNOR2_X1 port map( A => n16377, B => n16242, ZN => n16035);
   U20433 : XNOR2_X1 port map( A => n16035, B => n16034, ZN => n16036);
   U20434 : XNOR2_X1 port map( A => n16037, B => n16036, ZN => n17098);
   U20435 : INV_X1 port map( A => n17098, ZN => n16814);
   U20436 : XNOR2_X1 port map( A => n16038, B => n16414, ZN => n16040);
   U20437 : XNOR2_X1 port map( A => n16351, B => n16040, ZN => n16042);
   U20438 : XNOR2_X1 port map( A => n16255, B => n3751, ZN => n16041);
   U20439 : XNOR2_X1 port map( A => n16043, B => n16365, ZN => n16594);
   U20440 : INV_X1 port map( A => n16044, ZN => n16045);
   U20441 : XNOR2_X1 port map( A => n16594, B => n16045, ZN => n16049);
   U20442 : XNOR2_X1 port map( A => n16229, B => n16398, ZN => n16047);
   U20443 : XNOR2_X1 port map( A => n16047, B => n16046, ZN => n16048);
   U20445 : XNOR2_X1 port map( A => n16051, B => n16052, ZN => n16054);
   U20446 : XNOR2_X1 port map( A => n16346, B => n1248, ZN => n16053);
   U20447 : XNOR2_X1 port map( A => n16054, B => n16053, ZN => n16055);
   U20448 : XNOR2_X1 port map( A => n320, B => n3606, ZN => n16056);
   U20449 : XNOR2_X1 port map( A => n16056, B => n16567, ZN => n16057);
   U20450 : XNOR2_X1 port map( A => n16058, B => n16057, ZN => n16064);
   U20451 : INV_X1 port map( A => n16059, ZN => n16060);
   U20452 : XNOR2_X1 port map( A => n16271, B => n16060, ZN => n16061);
   U20453 : XNOR2_X1 port map( A => n16062, B => n16061, ZN => n16063);
   U20454 : NAND2_X1 port map( A1 => n16860, A2 => n17097, ZN => n16065);
   U20455 : MUX2_X1 port map( A => n16066, B => n16065, S => n17282, Z => 
                           n16067);
   U20456 : XNOR2_X1 port map( A => n16262, B => n3116, ZN => n16068);
   U20457 : XNOR2_X1 port map( A => n16068, B => n16405, ZN => n16069);
   U20458 : XNOR2_X1 port map( A => n16300, B => n16069, ZN => n16074);
   U20459 : XNOR2_X1 port map( A => n16071, B => n16070, ZN => n16072);
   U20460 : XNOR2_X1 port map( A => n16654, B => n16072, ZN => n16073);
   U20461 : XNOR2_X1 port map( A => n16252, B => n16625, ZN => n16076);
   U20462 : XNOR2_X1 port map( A => n16323, B => n16077, ZN => n16079);
   U20463 : INV_X1 port map( A => n3625, ZN => n28097);
   U20464 : XNOR2_X1 port map( A => n16257, B => n28097, ZN => n16078);
   U20465 : XNOR2_X1 port map( A => n16078, B => n16079, ZN => n16080);
   U20466 : XNOR2_X1 port map( A => n16081, B => n16470, ZN => n16083);
   U20467 : XNOR2_X1 port map( A => n16082, B => n16083, ZN => n16089);
   U20468 : XNOR2_X1 port map( A => n16328, B => n16084, ZN => n16087);
   U20469 : XNOR2_X1 port map( A => n16085, B => n2598, ZN => n16086);
   U20470 : XNOR2_X1 port map( A => n16087, B => n16086, ZN => n16088);
   U20471 : XNOR2_X1 port map( A => n16486, B => n3015, ZN => n16091);
   U20472 : XNOR2_X1 port map( A => n29571, B => n16399, ZN => n16092);
   U20473 : XNOR2_X1 port map( A => n16092, B => n16636, ZN => n16093);
   U20474 : AND2_X1 port map( A1 => n17120, A2 => n16811, ZN => n16100);
   U20475 : XNOR2_X1 port map( A => n29525, B => n3154, ZN => n16094);
   U20476 : XNOR2_X1 port map( A => n16094, B => n16480, ZN => n16097);
   U20477 : XNOR2_X1 port map( A => n16165, B => n16095, ZN => n16096);
   U20478 : XNOR2_X1 port map( A => n16097, B => n16096, ZN => n16099);
   U20479 : XNOR2_X1 port map( A => n16099, B => n16098, ZN => n17459);
   U20480 : INV_X1 port map( A => n17459, ZN => n16676);
   U20481 : OAI21_X1 port map( B1 => n16101, B2 => n16100, A => n16676, ZN => 
                           n16111);
   U20482 : AND2_X1 port map( A1 => n17459, A2 => n16812, ZN => n17113);
   U20483 : XNOR2_X1 port map( A => n16103, B => n16102, ZN => n16109);
   U20484 : INV_X1 port map( A => n3385, ZN => n16104);
   U20485 : XNOR2_X1 port map( A => n16105, B => n16104, ZN => n16106);
   U20486 : XNOR2_X1 port map( A => n16107, B => n16106, ZN => n16108);
   U20487 : XNOR2_X1 port map( A => n16108, B => n16109, ZN => n16810);
   U20488 : INV_X1 port map( A => n29083, ZN => n17457);
   U20489 : OAI21_X1 port map( B1 => n17113, B2 => n16810, A => n17457, ZN => 
                           n16110);
   U20490 : NAND2_X1 port map( A1 => n16111, A2 => n16110, ZN => n17601);
   U20491 : INV_X1 port map( A => n16598, ZN => n16113);
   U20492 : XNOR2_X1 port map( A => n16280, B => n1196, ZN => n16112);
   U20493 : XNOR2_X1 port map( A => n16113, B => n16112, ZN => n16118);
   U20494 : INV_X1 port map( A => n16366, ZN => n16114);
   U20495 : XNOR2_X1 port map( A => n16634, B => n16114, ZN => n16115);
   U20496 : XNOR2_X1 port map( A => n16116, B => n16115, ZN => n16117);
   U20497 : XNOR2_X1 port map( A => n16510, B => n3244, ZN => n16120);
   U20498 : XNOR2_X1 port map( A => n16121, B => n16120, ZN => n16122);
   U20499 : INV_X1 port map( A => n16123, ZN => n16125);
   U20500 : XNOR2_X1 port map( A => n16124, B => n16125, ZN => n16129);
   U20501 : XNOR2_X1 port map( A => n28557, B => n28693, ZN => n16127);
   U20502 : XNOR2_X1 port map( A => n16321, B => n16126, ZN => n16628);
   U20503 : XNOR2_X1 port map( A => n16127, B => n16628, ZN => n16128);
   U20504 : XNOR2_X1 port map( A => n16129, B => n16128, ZN => n16137);
   U20505 : XNOR2_X1 port map( A => n16130, B => n16131, ZN => n16132);
   U20506 : XNOR2_X1 port map( A => n16554, B => n16132, ZN => n16136);
   U20507 : XNOR2_X1 port map( A => n16653, B => n1246, ZN => n16133);
   U20508 : XNOR2_X1 port map( A => n16134, B => n16133, ZN => n16135);
   U20509 : XNOR2_X1 port map( A => n16136, B => n16135, ZN => n16668);
   U20510 : INV_X1 port map( A => n16137, ZN => n16806);
   U20511 : XNOR2_X1 port map( A => n16527, B => n16313, ZN => n16616);
   U20512 : XNOR2_X1 port map( A => n16346, B => n3062, ZN => n16141);
   U20513 : XNOR2_X1 port map( A => n16143, B => n21537, ZN => n16144);
   U20514 : XNOR2_X1 port map( A => n16145, B => n16144, ZN => n16149);
   U20515 : XNOR2_X1 port map( A => n16291, B => n16146, ZN => n16647);
   U20516 : XNOR2_X1 port map( A => n16147, B => n16647, ZN => n16148);
   U20517 : XNOR2_X1 port map( A => n16148, B => n16149, ZN => n17260);
   U20518 : NAND2_X1 port map( A1 => n17762, A2 => n17941, ZN => n16152);
   U20519 : XNOR2_X1 port map( A => n16154, B => n16302, ZN => n16158);
   U20520 : XNOR2_X1 port map( A => n16558, B => n24897, ZN => n16155);
   U20521 : XNOR2_X1 port map( A => n16156, B => n16155, ZN => n16157);
   U20522 : XNOR2_X1 port map( A => n16320, B => n16159, ZN => n16164);
   U20523 : XNOR2_X1 port map( A => n16160, B => n3697, ZN => n16161);
   U20524 : XNOR2_X1 port map( A => n16162, B => n16161, ZN => n16163);
   U20525 : XNOR2_X1 port map( A => n16477, B => n16165, ZN => n16167);
   U20526 : XNOR2_X1 port map( A => n16607, B => n3134, ZN => n16168);
   U20527 : XNOR2_X1 port map( A => n16311, B => n16168, ZN => n16169);
   U20528 : XNOR2_X1 port map( A => n16192, B => n16170, ZN => n16595);
   U20529 : XNOR2_X1 port map( A => n16171, B => n16595, ZN => n16175);
   U20530 : XNOR2_X1 port map( A => n29571, B => n2522, ZN => n16173);
   U20531 : XNOR2_X1 port map( A => n16278, B => n16173, ZN => n16174);
   U20532 : INV_X1 port map( A => n16176, ZN => n16204);
   U20533 : XNOR2_X1 port map( A => n16204, B => n2446, ZN => n16178);
   U20534 : XNOR2_X1 port map( A => n16178, B => n16177, ZN => n16181);
   U20535 : XNOR2_X1 port map( A => n16179, B => n16331, ZN => n16180);
   U20536 : XNOR2_X1 port map( A => n321, B => n3334, ZN => n16182);
   U20537 : XNOR2_X1 port map( A => n16182, B => n16294, ZN => n16184);
   U20538 : XNOR2_X1 port map( A => n16183, B => n16184, ZN => n16188);
   U20539 : XNOR2_X1 port map( A => n16569, B => n16185, ZN => n16186);
   U20540 : XNOR2_X1 port map( A => n16564, B => n16186, ZN => n16187);
   U20541 : XNOR2_X1 port map( A => n19650, B => n19607, ZN => n16698);
   U20542 : XNOR2_X1 port map( A => n16191, B => n16190, ZN => n16195);
   U20543 : XNOR2_X1 port map( A => n16192, B => n2987, ZN => n16193);
   U20545 : INV_X1 port map( A => n16888, ZN => n17140);
   U20546 : XNOR2_X1 port map( A => n16199, B => n16556, ZN => n16202);
   U20547 : XNOR2_X1 port map( A => n16558, B => n3483, ZN => n16200);
   U20548 : XNOR2_X1 port map( A => n16206, B => n16205, ZN => n16210);
   U20549 : XNOR2_X1 port map( A => n16207, B => n16208, ZN => n16209);
   U20550 : NAND2_X1 port map( A1 => n17140, A2 => n16887, ZN => n16702);
   U20551 : INV_X1 port map( A => n16211, ZN => n16212);
   U20552 : XNOR2_X1 port map( A => n16213, B => n16212, ZN => n16215);
   U20553 : XNOR2_X1 port map( A => n16215, B => n16214, ZN => n16220);
   U20554 : XNOR2_X1 port map( A => n16216, B => n26909, ZN => n16217);
   U20555 : XNOR2_X1 port map( A => n16218, B => n16217, ZN => n16219);
   U20556 : NAND2_X1 port map( A1 => n16888, A2 => n17139, ZN => n17136);
   U20557 : NAND2_X1 port map( A1 => n16702, A2 => n17136, ZN => n16227);
   U20558 : XNOR2_X1 port map( A => n16160, B => n3666, ZN => n16222);
   U20559 : XNOR2_X1 port map( A => n16221, B => n16222, ZN => n16226);
   U20560 : XNOR2_X1 port map( A => n16223, B => n16224, ZN => n16225);
   U20561 : XNOR2_X1 port map( A => n16231, B => n16230, ZN => n16235);
   U20562 : XNOR2_X1 port map( A => n16233, B => n16232, ZN => n16234);
   U20563 : XNOR2_X1 port map( A => n16235, B => n16234, ZN => n16236);
   U20564 : XNOR2_X1 port map( A => n16236, B => n16237, ZN => n16736);
   U20565 : XNOR2_X1 port map( A => n16238, B => n730, ZN => n16239);
   U20566 : XNOR2_X1 port map( A => n16240, B => n16239, ZN => n16245);
   U20567 : XNOR2_X1 port map( A => n16242, B => n16241, ZN => n16513);
   U20568 : XNOR2_X1 port map( A => n16513, B => n16243, ZN => n16244);
   U20569 : XNOR2_X1 port map( A => n16244, B => n16245, ZN => n17147);
   U20570 : NAND2_X1 port map( A1 => n16736, A2 => n17147, ZN => n17485);
   U20571 : XNOR2_X1 port map( A => n16525, B => n16246, ZN => n16251);
   U20572 : XNOR2_X1 port map( A => n16247, B => n3067, ZN => n16248);
   U20573 : XNOR2_X1 port map( A => n16249, B => n16248, ZN => n16250);
   U20574 : XNOR2_X1 port map( A => n16251, B => n16250, ZN => n17076);
   U20575 : XNOR2_X1 port map( A => n16252, B => n16498, ZN => n16254);
   U20576 : XNOR2_X1 port map( A => n16254, B => n16253, ZN => n16261);
   U20577 : XNOR2_X1 port map( A => n16256, B => n16255, ZN => n16259);
   U20578 : XNOR2_X1 port map( A => n16257, B => n27894, ZN => n16258);
   U20579 : XNOR2_X1 port map( A => n16258, B => n16259, ZN => n16260);
   U20580 : XNOR2_X2 port map( A => n16261, B => n16260, ZN => n17489);
   U20581 : OR2_X1 port map( A1 => n17076, A2 => n17489, ZN => n16735);
   U20582 : XNOR2_X1 port map( A => n16262, B => n27225, ZN => n16263);
   U20583 : XNOR2_X1 port map( A => n16263, B => n28406, ZN => n16265);
   U20584 : XNOR2_X1 port map( A => n16266, B => n16265, ZN => n16268);
   U20585 : MUX2_X1 port map( A => n17485, B => n16735, S => n17487, Z => 
                           n16277);
   U20586 : INV_X1 port map( A => n16736, ZN => n17078);
   U20587 : XNOR2_X1 port map( A => n16269, B => n16270, ZN => n16276);
   U20588 : XNOR2_X1 port map( A => n16271, B => n16272, ZN => n16274);
   U20589 : XNOR2_X1 port map( A => n16534, B => n3686, ZN => n16273);
   U20590 : XNOR2_X1 port map( A => n16274, B => n16273, ZN => n16275);
   U20592 : INV_X1 port map( A => n17487, ZN => n17153);
   U20593 : INV_X1 port map( A => n17147, ZN => n17146);
   U20594 : XNOR2_X1 port map( A => n16280, B => n16279, ZN => n16632);
   U20595 : XNOR2_X1 port map( A => n16281, B => n16632, ZN => n16288);
   U20596 : XNOR2_X1 port map( A => n16282, B => n16283, ZN => n16286);
   U20597 : XNOR2_X1 port map( A => n16284, B => n3212, ZN => n16285);
   U20598 : XNOR2_X1 port map( A => n16286, B => n16285, ZN => n16287);
   U20599 : XNOR2_X1 port map( A => n16288, B => n16287, ZN => n16612);
   U20600 : XNOR2_X1 port map( A => n320, B => n1187, ZN => n16290);
   U20601 : XNOR2_X1 port map( A => n16290, B => n16291, ZN => n16293);
   U20602 : XNOR2_X1 port map( A => n28579, B => n16649, ZN => n16358);
   U20603 : XNOR2_X1 port map( A => n16358, B => n16293, ZN => n16299);
   U20604 : XNOR2_X1 port map( A => n16295, B => n16294, ZN => n16297);
   U20605 : XNOR2_X1 port map( A => n16296, B => n16297, ZN => n16298);
   U20606 : XNOR2_X1 port map( A => n16299, B => n16298, ZN => n16730);
   U20607 : NOR2_X1 port map( A1 => n16612, A2 => n17497, ZN => n16337);
   U20608 : INV_X1 port map( A => n16300, ZN => n16301);
   U20609 : XNOR2_X1 port map( A => n16301, B => n16302, ZN => n16308);
   U20610 : XNOR2_X1 port map( A => n16304, B => n16303, ZN => n16656);
   U20611 : XNOR2_X1 port map( A => n16305, B => n3451, ZN => n16306);
   U20612 : XNOR2_X1 port map( A => n16656, B => n16306, ZN => n16307);
   U20613 : XNOR2_X1 port map( A => n16310, B => n16309, ZN => n16344);
   U20614 : XNOR2_X1 port map( A => n16344, B => n16311, ZN => n16317);
   U20615 : XNOR2_X1 port map( A => n16480, B => n16312, ZN => n16315);
   U20616 : XNOR2_X1 port map( A => n16313, B => n3414, ZN => n16314);
   U20617 : XNOR2_X1 port map( A => n16315, B => n16314, ZN => n16316);
   U20618 : XNOR2_X1 port map( A => n16319, B => n16318, ZN => n16352);
   U20619 : XNOR2_X1 port map( A => n16320, B => n16352, ZN => n16327);
   U20620 : XNOR2_X1 port map( A => n16321, B => n16322, ZN => n16325);
   U20621 : XNOR2_X1 port map( A => n16323, B => n3710, ZN => n16324);
   U20622 : XNOR2_X1 port map( A => n16325, B => n16324, ZN => n16326);
   U20623 : XNOR2_X1 port map( A => n16327, B => n16326, ZN => n17498);
   U20624 : XNOR2_X1 port map( A => n16328, B => n16329, ZN => n16330);
   U20625 : XNOR2_X1 port map( A => n16331, B => n16330, ZN => n16336);
   U20626 : INV_X1 port map( A => n16640, ZN => n16334);
   U20627 : XNOR2_X1 port map( A => n29516, B => n2510, ZN => n16333);
   U20628 : XNOR2_X1 port map( A => n16334, B => n16333, ZN => n16335);
   U20629 : NOR2_X1 port map( A1 => n6079, A2 => n18465, ZN => n16338);
   U20630 : XNOR2_X1 port map( A => n16303, B => n3742, ZN => n16341);
   U20631 : XNOR2_X1 port map( A => n16555, B => n16341, ZN => n16342);
   U20632 : INV_X1 port map( A => n16343, ZN => n16345);
   U20633 : XNOR2_X1 port map( A => n16345, B => n16344, ZN => n16350);
   U20634 : XNOR2_X1 port map( A => n16346, B => n2982, ZN => n16348);
   U20635 : XNOR2_X1 port map( A => n16348, B => n16347, ZN => n16349);
   U20636 : INV_X1 port map( A => n16712, ZN => n16381);
   U20637 : INV_X1 port map( A => n16351, ZN => n16353);
   U20638 : XNOR2_X1 port map( A => n16353, B => n16352, ZN => n16357);
   U20639 : XNOR2_X1 port map( A => n6449, B => n16579, ZN => n16355);
   U20640 : INV_X1 port map( A => n2894, ZN => n26877);
   U20641 : XNOR2_X1 port map( A => n29151, B => n26877, ZN => n16354);
   U20642 : XNOR2_X1 port map( A => n16355, B => n16354, ZN => n16356);
   U20644 : NAND2_X1 port map( A1 => n16381, A2 => n28776, ZN => n16383);
   U20646 : XNOR2_X1 port map( A => n16359, B => n16358, ZN => n16364);
   U20647 : XNOR2_X1 port map( A => n16360, B => n3493, ZN => n16361);
   U20648 : XNOR2_X1 port map( A => n16362, B => n16361, ZN => n16363);
   U20649 : INV_X1 port map( A => n17374, ZN => n17173);
   U20650 : XNOR2_X1 port map( A => n16366, B => n16365, ZN => n16368);
   U20651 : XNOR2_X1 port map( A => n16367, B => n16368, ZN => n16372);
   U20652 : XNOR2_X1 port map( A => n16369, B => n16370, ZN => n16371);
   U20653 : XNOR2_X1 port map( A => n16373, B => n16586, ZN => n16374);
   U20654 : XNOR2_X1 port map( A => n16375, B => n16374, ZN => n16380);
   U20655 : INV_X1 port map( A => n16376, ZN => n16379);
   U20656 : XNOR2_X1 port map( A => n16377, B => n3463, ZN => n16378);
   U20657 : NAND3_X1 port map( A1 => n29635, A2 => n16381, A3 => n17375, ZN => 
                           n16382);
   U20658 : XNOR2_X1 port map( A => n16509, B => n28597, ZN => n16385);
   U20659 : XNOR2_X1 port map( A => n16384, B => n16385, ZN => n16392);
   U20660 : XNOR2_X1 port map( A => n16387, B => n16386, ZN => n16390);
   U20661 : XNOR2_X1 port map( A => n16388, B => n2960, ZN => n16389);
   U20662 : XNOR2_X1 port map( A => n16390, B => n16389, ZN => n16391);
   U20663 : XNOR2_X1 port map( A => n16392, B => n16391, ZN => n16884);
   U20664 : INV_X1 port map( A => n16393, ZN => n16394);
   U20665 : XNOR2_X1 port map( A => n16395, B => n16394, ZN => n16396);
   U20666 : XNOR2_X1 port map( A => n16397, B => n16396, ZN => n16403);
   U20667 : XNOR2_X1 port map( A => n16400, B => n2306, ZN => n16401);
   U20668 : XNOR2_X1 port map( A => n16488, B => n16401, ZN => n16402);
   U20669 : XNOR2_X1 port map( A => n16404, B => n16405, ZN => n16447);
   U20670 : XNOR2_X1 port map( A => n16406, B => n16447, ZN => n16413);
   U20671 : XNOR2_X1 port map( A => n16408, B => n16407, ZN => n16411);
   U20672 : XNOR2_X1 port map( A => n16409, B => n27452, ZN => n16410);
   U20673 : XNOR2_X1 port map( A => n16411, B => n16410, ZN => n16412);
   U20674 : XNOR2_X1 port map( A => n16415, B => n16454, ZN => n16420);
   U20675 : XNOR2_X1 port map( A => n16416, B => n3527, ZN => n16417);
   U20676 : XNOR2_X1 port map( A => n16418, B => n16417, ZN => n16419);
   U20677 : NOR2_X1 port map( A1 => n17181, A2 => n17528, ZN => n17531);
   U20678 : INV_X1 port map( A => n17531, ZN => n16431);
   U20679 : XNOR2_X1 port map( A => n16422, B => n16421, ZN => n16423);
   U20680 : XNOR2_X1 port map( A => n16424, B => n16423, ZN => n16429);
   U20681 : XNOR2_X1 port map( A => n16425, B => n16426, ZN => n16464);
   U20682 : XNOR2_X1 port map( A => n16429, B => n16428, ZN => n16706);
   U20683 : INV_X1 port map( A => n16884, ZN => n17157);
   U20684 : OAI22_X1 port map( A1 => n6928, A2 => n16431, B1 => n16430, B2 => 
                           n17158, ZN => n16441);
   U20685 : XNOR2_X1 port map( A => n16433, B => n16432, ZN => n16439);
   U20686 : XNOR2_X1 port map( A => n16434, B => n16435, ZN => n16478);
   U20687 : XNOR2_X1 port map( A => n16436, B => n27462, ZN => n16437);
   U20688 : XNOR2_X1 port map( A => n16437, B => n16478, ZN => n16438);
   U20689 : XNOR2_X1 port map( A => n16438, B => n16439, ZN => n17524);
   U20690 : NAND2_X1 port map( A1 => n6928, A2 => n4979, ZN => n16440);
   U20691 : XNOR2_X1 port map( A => n16443, B => n3223, ZN => n16446);
   U20692 : INV_X1 port map( A => n16444, ZN => n16445);
   U20693 : XNOR2_X1 port map( A => n16446, B => n16445, ZN => n16448);
   U20694 : XNOR2_X1 port map( A => n16448, B => n16447, ZN => n16452);
   U20695 : XNOR2_X1 port map( A => n29511, B => n16450, ZN => n16451);
   U20696 : XNOR2_X1 port map( A => n16453, B => n16454, ZN => n16460);
   U20697 : XNOR2_X1 port map( A => n16456, B => n3211, ZN => n16457);
   U20698 : XNOR2_X1 port map( A => n16458, B => n16457, ZN => n16459);
   U20699 : XNOR2_X1 port map( A => n16460, B => n16459, ZN => n16549);
   U20700 : INV_X1 port map( A => n16549, ZN => n17508);
   U20701 : XNOR2_X1 port map( A => n16461, B => n16462, ZN => n16466);
   U20702 : XNOR2_X1 port map( A => n16059, B => n3752, ZN => n16463);
   U20703 : XNOR2_X1 port map( A => n16464, B => n16463, ZN => n16465);
   U20704 : XNOR2_X1 port map( A => n16467, B => n29247, ZN => n16469);
   U20705 : XNOR2_X1 port map( A => n16468, B => n16469, ZN => n16475);
   U20706 : XNOR2_X1 port map( A => n28597, B => n16471, ZN => n16473);
   U20707 : XNOR2_X1 port map( A => n16472, B => n16473, ZN => n16474);
   U20708 : XNOR2_X1 port map( A => n16477, B => n16476, ZN => n16479);
   U20709 : XNOR2_X1 port map( A => n16480, B => n3369, ZN => n16482);
   U20710 : XNOR2_X1 port map( A => n15070, B => n16483, ZN => n16485);
   U20711 : XNOR2_X1 port map( A => n16484, B => n16485, ZN => n16490);
   U20712 : XNOR2_X1 port map( A => n16486, B => n2381, ZN => n16487);
   U20713 : XNOR2_X1 port map( A => n16487, B => n16488, ZN => n16489);
   U20714 : OAI21_X1 port map( B1 => n4271, B2 => n17505, A => n17506, ZN => 
                           n16491);
   U20715 : INV_X1 port map( A => n18471, ZN => n18464);
   U20716 : XNOR2_X1 port map( A => n16494, B => n16495, ZN => n16496);
   U20717 : XNOR2_X1 port map( A => n16497, B => n16496, ZN => n16502);
   U20718 : XNOR2_X1 port map( A => n16498, B => n3770, ZN => n16500);
   U20719 : XNOR2_X1 port map( A => n16499, B => n16500, ZN => n16501);
   U20720 : XNOR2_X1 port map( A => n16503, B => n16504, ZN => n16508);
   U20721 : INV_X1 port map( A => n17452, ZN => n17067);
   U20722 : XNOR2_X1 port map( A => n16510, B => n16509, ZN => n16512);
   U20723 : XNOR2_X1 port map( A => n16512, B => n16511, ZN => n16516);
   U20724 : XNOR2_X1 port map( A => n16513, B => n16514, ZN => n16515);
   U20725 : INV_X1 port map( A => n17450, ZN => n17066);
   U20726 : MUX2_X1 port map( A => n6772, B => n17067, S => n17066, Z => n16539
                           );
   U20727 : XNOR2_X1 port map( A => n16517, B => n16518, ZN => n16523);
   U20728 : XNOR2_X1 port map( A => n16519, B => n3049, ZN => n16520);
   U20729 : XNOR2_X1 port map( A => n16521, B => n16520, ZN => n16522);
   U20730 : XNOR2_X1 port map( A => n16523, B => n16522, ZN => n17455);
   U20731 : XNOR2_X1 port map( A => n16524, B => n16525, ZN => n16531);
   U20732 : XNOR2_X1 port map( A => n16526, B => n16603, ZN => n16529);
   U20733 : XNOR2_X1 port map( A => n16527, B => n1062, ZN => n16528);
   U20734 : XNOR2_X1 port map( A => n16529, B => n16528, ZN => n16530);
   U20735 : XNOR2_X1 port map( A => n16531, B => n16530, ZN => n17129);
   U20736 : INV_X1 port map( A => n17129, ZN => n17068);
   U20737 : NOR2_X1 port map( A1 => n28193, A2 => n16797, ZN => n16538);
   U20738 : XNOR2_X1 port map( A => n16534, B => n3633, ZN => n16535);
   U20739 : XNOR2_X1 port map( A => n16536, B => n16535, ZN => n16537);
   U20740 : INV_X1 port map( A => n17456, ZN => n17120);
   U20741 : NAND2_X1 port map( A1 => n17120, A2 => n16810, ZN => n16540);
   U20742 : AOI21_X1 port map( B1 => n17117, B2 => n16540, A => n16676, ZN => 
                           n16545);
   U20746 : NAND2_X1 port map( A1 => n18353, A2 => n16611, ZN => n17918);
   U20747 : INV_X1 port map( A => n16728, ZN => n16546);
   U20748 : NAND2_X1 port map( A1 => n16546, A2 => n4271, ZN => n16553);
   U20749 : NAND3_X1 port map( A1 => n4271, A2 => n4270, A3 => n17505, ZN => 
                           n16548);
   U20750 : BUF_X2 port map( A => n16549, Z => n17830);
   U20751 : XNOR2_X1 port map( A => n16555, B => n16554, ZN => n16562);
   U20752 : XNOR2_X1 port map( A => n16557, B => n16556, ZN => n16560);
   U20753 : XNOR2_X1 port map( A => n16558, B => n3219, ZN => n16559);
   U20754 : XNOR2_X1 port map( A => n16560, B => n16559, ZN => n16561);
   U20755 : XNOR2_X1 port map( A => n16563, B => n16564, ZN => n16565);
   U20756 : XNOR2_X1 port map( A => n16566, B => n16565, ZN => n16573);
   U20757 : XNOR2_X1 port map( A => n16568, B => n16567, ZN => n16571);
   U20758 : XNOR2_X1 port map( A => n16569, B => n3482, ZN => n16570);
   U20759 : XNOR2_X1 port map( A => n16570, B => n16571, ZN => n16572);
   U20760 : INV_X1 port map( A => n17516, ZN => n17083);
   U20761 : XNOR2_X1 port map( A => n16574, B => n16575, ZN => n16576);
   U20762 : XNOR2_X1 port map( A => n16577, B => n16576, ZN => n16584);
   U20763 : XNOR2_X1 port map( A => n16578, B => n16579, ZN => n16582);
   U20764 : XNOR2_X1 port map( A => n16580, B => n22489, ZN => n16581);
   U20765 : XNOR2_X1 port map( A => n16582, B => n16581, ZN => n16583);
   U20767 : XNOR2_X1 port map( A => n16585, B => n16586, ZN => n16587);
   U20768 : XNOR2_X1 port map( A => n16588, B => n16587, ZN => n16593);
   U20769 : XNOR2_X1 port map( A => n16589, B => n2325, ZN => n16590);
   U20770 : XNOR2_X1 port map( A => n16591, B => n16590, ZN => n16592);
   U20771 : XNOR2_X1 port map( A => n16593, B => n16592, ZN => n17469);
   U20772 : NOR2_X1 port map( A1 => n29406, A2 => n17469, ZN => n16601);
   U20773 : XNOR2_X1 port map( A => n16596, B => n2353, ZN => n16597);
   U20774 : XNOR2_X1 port map( A => n16598, B => n16597, ZN => n16599);
   U20775 : INV_X1 port map( A => n17518, ZN => n17109);
   U20776 : INV_X1 port map( A => n16603, ZN => n16604);
   U20777 : XNOR2_X1 port map( A => n16607, B => n2912, ZN => n16608);
   U20778 : XNOR2_X1 port map( A => n16609, B => n16608, ZN => n16610);
   U20779 : NAND2_X1 port map( A1 => n536, A2 => n538, ZN => n16614);
   U20780 : NOR2_X1 port map( A1 => n29373, A2 => n17062, ZN => n16613);
   U20781 : AOI21_X1 port map( B1 => n16611, B2 => n18312, A => n18353, ZN => 
                           n16615);
   U20782 : XNOR2_X1 port map( A => n16616, B => n16617, ZN => n16624);
   U20783 : XNOR2_X1 port map( A => n16619, B => n16618, ZN => n16622);
   U20784 : XNOR2_X1 port map( A => n16620, B => n1079, ZN => n16621);
   U20785 : XNOR2_X1 port map( A => n16622, B => n16621, ZN => n16623);
   U20786 : XNOR2_X1 port map( A => n16625, B => n3644, ZN => n16626);
   U20787 : XNOR2_X1 port map( A => n16627, B => n16626, ZN => n16631);
   U20788 : XNOR2_X1 port map( A => n16629, B => n16628, ZN => n16630);
   U20789 : XNOR2_X1 port map( A => n16630, B => n16631, ZN => n17478);
   U20790 : NOR2_X1 port map( A1 => n534, A2 => n3883, ZN => n16660);
   U20791 : XNOR2_X1 port map( A => n16633, B => n16632, ZN => n16638);
   U20792 : XNOR2_X1 port map( A => n16634, B => n3650, ZN => n16635);
   U20793 : XNOR2_X1 port map( A => n16636, B => n16635, ZN => n16637);
   U20794 : INV_X1 port map( A => n16724, ZN => n17481);
   U20795 : XNOR2_X1 port map( A => n16639, B => n16640, ZN => n16646);
   U20796 : XNOR2_X1 port map( A => n16642, B => n16641, ZN => n16644);
   U20797 : XNOR2_X1 port map( A => n16644, B => n16643, ZN => n16645);
   U20798 : XNOR2_X1 port map( A => n16648, B => n16647, ZN => n16652);
   U20799 : XNOR2_X1 port map( A => n16649, B => n2986, ZN => n16650);
   U20800 : XNOR2_X1 port map( A => n16652, B => n16651, ZN => n16691);
   U20801 : INV_X1 port map( A => n16691, ZN => n16723);
   U20802 : XNOR2_X1 port map( A => n16653, B => n2477, ZN => n16655);
   U20803 : XNOR2_X1 port map( A => n16655, B => n16654, ZN => n16657);
   U20804 : XNOR2_X1 port map( A => n16657, B => n16656, ZN => n16659);
   U20805 : XNOR2_X1 port map( A => n16659, B => n16658, ZN => n17474);
   U20806 : NOR2_X1 port map( A1 => n16661, A2 => n17667, ZN => n16662);
   U20807 : NAND4_X1 port map( A1 => n2055, A2 => n16663, A3 => n518, A4 => 
                           n16662, ZN => n16664);
   U20808 : NOR2_X1 port map( A1 => n17276, A2 => n17278, ZN => n16665);
   U20811 : INV_X1 port map( A => n16685, ZN => n17663);
   U20812 : INV_X1 port map( A => n16668, ZN => n16805);
   U20813 : OAI211_X1 port map( C1 => n17259, C2 => n16805, A => n17260, B => 
                           n16669, ZN => n16671);
   U20814 : INV_X1 port map( A => n17466, ZN => n16673);
   U20815 : AOI22_X1 port map( A1 => n17090, A2 => n16675, B1 => n6830, B2 => 
                           n16674, ZN => n16693);
   U20816 : NAND2_X1 port map( A1 => n16810, A2 => n421, ZN => n16678);
   U20817 : NAND2_X1 port map( A1 => n16813, A2 => n29083, ZN => n16677);
   U20818 : NAND2_X1 port map( A1 => n29559, A2 => n16679, ZN => n17284);
   U20819 : INV_X1 port map( A => n17283, ZN => n16857);
   U20820 : OAI21_X1 port map( B1 => n17284, B2 => n16857, A => n16680, ZN => 
                           n16688);
   U20821 : NAND2_X1 port map( A1 => n16688, A2 => n17117, ZN => n16683);
   U20823 : MUX2_X1 port map( A => n29086, B => n17282, S => n17101, Z => 
                           n16681);
   U20824 : INV_X1 port map( A => n17102, ZN => n16815);
   U20825 : NAND3_X1 port map( A1 => n16681, A2 => n16815, A3 => n17117, ZN => 
                           n16682);
   U20826 : NAND2_X1 port map( A1 => n16683, A2 => n16682, ZN => n16684);
   U20827 : NAND3_X1 port map( A1 => n514, A2 => n16932, A3 => n16684, ZN => 
                           n16694);
   U20828 : OAI21_X1 port map( B1 => n16814, B2 => n17282, A => n16815, ZN => 
                           n16686);
   U20829 : NOR2_X1 port map( A1 => n16687, A2 => n16686, ZN => n16689);
   U20830 : AOI22_X1 port map( A1 => n17475, A2 => n3883, B1 => n17476, B2 => 
                           n17477, ZN => n16692);
   U20832 : XNOR2_X1 port map( A => n29505, B => n3244, ZN => n16695);
   U20833 : XNOR2_X1 port map( A => n16696, B => n16695, ZN => n16697);
   U20834 : XNOR2_X1 port map( A => n16698, B => n16697, ZN => n20551);
   U20835 : INV_X1 port map( A => n17385, ZN => n17188);
   U20836 : MUX2_X1 port map( A => n17188, B => n28497, S => n16879, Z => 
                           n16701);
   U20837 : INV_X1 port map( A => n16700, ZN => n18069);
   U20838 : AND2_X1 port map( A1 => n16702, A2 => n17139, ZN => n16705);
   U20840 : NAND2_X1 port map( A1 => n17139, A2 => n16887, ZN => n17500);
   U20841 : NOR2_X1 port map( A1 => n17500, A2 => n17502, ZN => n16703);
   U20842 : NOR2_X1 port map( A1 => n17087, A2 => n16703, ZN => n16704);
   U20844 : NOR2_X1 port map( A1 => n16706, A2 => n16883, ZN => n18221);
   U20845 : INV_X1 port map( A => n18221, ZN => n17532);
   U20846 : MUX2_X1 port map( A => n16707, B => n17532, S => n17158, Z => 
                           n16708);
   U20847 : AOI21_X1 port map( B1 => n17200, B2 => n17339, A => n28564, ZN => 
                           n16710);
   U20848 : NOR2_X1 port map( A1 => n17338, A2 => n17204, ZN => n16709);
   U20849 : NAND2_X1 port map( A1 => n17336, A2 => n17204, ZN => n16711);
   U20850 : INV_X1 port map( A => n16711, ZN => n16936);
   U20852 : INV_X1 port map( A => n17357, ZN => n17195);
   U20854 : OAI21_X1 port map( B1 => n17198, B2 => n16713, A => n17356, ZN => 
                           n16716);
   U20858 : OAI21_X1 port map( B1 => n16717, B2 => n29502, A => n18195, ZN => 
                           n16720);
   U20859 : OAI211_X1 port map( C1 => n18195, C2 => n17746, A => n16720, B => 
                           n16719, ZN => n18737);
   U20860 : NOR2_X1 port map( A1 => n17129, A2 => n16797, ZN => n16721);
   U20861 : NOR2_X1 port map( A1 => n16723, A2 => n17124, ZN => n16722);
   U20862 : INV_X1 port map( A => n17804, ZN => n16747);
   U20863 : NAND3_X1 port map( A1 => n4271, A2 => n17506, A3 => n17508, ZN => 
                           n16729);
   U20864 : NOR2_X1 port map( A1 => n17492, A2 => n17498, ZN => n17495);
   U20865 : INV_X1 port map( A => n16730, ZN => n16882);
   U20866 : NAND2_X1 port map( A1 => n16882, A2 => n17491, ZN => n16880);
   U20868 : OAI21_X1 port map( B1 => n538, B2 => n16880, A => n17493, ZN => 
                           n16733);
   U20869 : NAND3_X1 port map( A1 => n16880, A2 => n4314, A3 => n536, ZN => 
                           n16732);
   U20870 : MUX2_X1 port map( A => n16735, B => n16734, S => n17078, Z => 
                           n16739);
   U20871 : INV_X1 port map( A => n17486, ZN => n16737);
   U20872 : AOI22_X1 port map( A1 => n16737, A2 => n4655, B1 => n17488, B2 => 
                           n5737, ZN => n16738);
   U20873 : NAND3_X1 port map( A1 => n3995, A2 => n18276, A3 => n18204, ZN => 
                           n16746);
   U20874 : INV_X1 port map( A => n17110, ZN => n17520);
   U20875 : INV_X1 port map( A => n17469, ZN => n17517);
   U20876 : NAND3_X1 port map( A1 => n17109, A2 => n17106, A3 => n17517, ZN => 
                           n16742);
   U20877 : NAND3_X1 port map( A1 => n17518, A2 => n29406, A3 => n17083, ZN => 
                           n16741);
   U20878 : NAND3_X1 port map( A1 => n17106, A2 => n17470, A3 => n17469, ZN => 
                           n16740);
   U20880 : NOR2_X1 port map( A1 => n18203, A2 => n18277, ZN => n16744);
   U20881 : OAI21_X1 port map( B1 => n16744, B2 => n3994, A => n16898, ZN => 
                           n16745);
   U20882 : OAI211_X1 port map( C1 => n16747, C2 => n16898, A => n16746, B => 
                           n16745, ZN => n18899);
   U20883 : XNOR2_X1 port map( A => n18899, B => n18737, ZN => n19646);
   U20884 : NOR2_X1 port map( A1 => n17025, A2 => n17344, ZN => n17350);
   U20885 : NOR2_X1 port map( A1 => n17029, A2 => n17347, ZN => n16748);
   U20887 : NOR2_X1 port map( A1 => n17348, A2 => n17347, ZN => n16749);
   U20888 : OAI21_X1 port map( B1 => n16749, B2 => n17029, A => n17025, ZN => 
                           n18093);
   U20889 : NOR2_X1 port map( A1 => n17546, A2 => n17539, ZN => n18091);
   U20890 : AOI21_X1 port map( B1 => n18090, B2 => n18093, A => n18091, ZN => 
                           n16758);
   U20891 : OR2_X1 port map( A1 => n17542, A2 => n17543, ZN => n17215);
   U20892 : NOR2_X1 port map( A1 => n16939, A2 => n17545, ZN => n16750);
   U20893 : INV_X1 port map( A => n18096, ZN => n16757);
   U20894 : MUX2_X1 port map( A => n17555, B => n17556, S => n17554, Z => 
                           n16754);
   U20895 : OAI21_X1 port map( B1 => n16913, B2 => n17221, A => n29142, ZN => 
                           n16753);
   U20896 : NOR2_X1 port map( A1 => n16911, A2 => n16908, ZN => n16752);
   U20897 : AOI22_X1 port map( A1 => n16758, A2 => n16757, B1 => n18179, B2 => 
                           n18178, ZN => n18442);
   U20898 : INV_X1 port map( A => n17234, ZN => n17043);
   U20899 : NAND2_X1 port map( A1 => n17046, A2 => n17365, ZN => n16759);
   U20900 : INV_X1 port map( A => n17364, ZN => n16761);
   U20901 : NAND2_X1 port map( A1 => n16761, A2 => n6180, ZN => n17788);
   U20902 : NAND3_X1 port map( A1 => n16844, A2 => n17002, A3 => n17275, ZN => 
                           n16765);
   U20903 : OAI21_X1 port map( B1 => n17001, B2 => n16766, A => n16765, ZN => 
                           n16769);
   U20904 : NOR2_X1 port map( A1 => n16767, A2 => n17271, ZN => n16768);
   U20905 : INV_X1 port map( A => n18109, ZN => n17799);
   U20906 : NOR2_X1 port map( A1 => n17265, A2 => n16995, ZN => n16772);
   U20907 : INV_X1 port map( A => n29600, ZN => n16970);
   U20909 : NAND2_X1 port map( A1 => n16772, A2 => n29600, ZN => n16770);
   U20910 : OAI211_X2 port map( C1 => n16772, C2 => n16773, A => n16771, B => 
                           n16770, ZN => n18111);
   U20911 : NAND2_X1 port map( A1 => n17248, A2 => n17017, ZN => n16775);
   U20912 : NAND3_X1 port map( A1 => n16865, A2 => n16775, A3 => n17249, ZN => 
                           n16778);
   U20913 : NOR2_X1 port map( A1 => n17016, A2 => n17249, ZN => n16776);
   U20914 : NAND2_X1 port map( A1 => n16776, A2 => n17251, ZN => n16777);
   U20915 : NAND3_X1 port map( A1 => n17799, A2 => n18111, A3 => n17903, ZN => 
                           n16796);
   U20916 : NOR2_X1 port map( A1 => n17259, A2 => n16779, ZN => n16780);
   U20917 : NAND2_X1 port map( A1 => n17425, A2 => n29088, ZN => n16787);
   U20918 : NAND2_X1 port map( A1 => n17428, A2 => n28194, ZN => n16783);
   U20919 : NAND2_X1 port map( A1 => n16974, A2 => n16783, ZN => n16784);
   U20920 : NAND2_X1 port map( A1 => n16784, A2 => n2826, ZN => n16786);
   U20921 : NAND3_X1 port map( A1 => n28792, A2 => n17005, A3 => n17720, ZN => 
                           n16785);
   U20922 : NAND3_X1 port map( A1 => n17799, A2 => n17902, A3 => n18107, ZN => 
                           n16795);
   U20923 : INV_X1 port map( A => n17902, ZN => n18459);
   U20924 : NAND2_X1 port map( A1 => n17903, A2 => n18459, ZN => n16794);
   U20925 : NAND2_X1 port map( A1 => n17012, A2 => n29152, ZN => n16789);
   U20926 : XNOR2_X1 port map( A => n19252, B => n19549, ZN => n19582);
   U20927 : XNOR2_X1 port map( A => n19646, B => n19582, ZN => n16871);
   U20928 : NAND2_X1 port map( A1 => n28193, A2 => n16797, ZN => n16798);
   U20929 : NAND2_X1 port map( A1 => n16798, A2 => n17068, ZN => n16799);
   U20930 : OAI211_X1 port map( C1 => n16803, C2 => n3883, A => n17124, B => 
                           n17481, ZN => n16804);
   U20931 : NAND2_X1 port map( A1 => n16805, A2 => n29574, ZN => n16809);
   U20932 : NAND2_X1 port map( A1 => n17283, A2 => n1466, ZN => n16816);
   U20933 : MUX2_X1 port map( A => n16817, B => n16816, S => n16815, Z => 
                           n16818);
   U20934 : NOR2_X1 port map( A1 => n18174, A2 => n18168, ZN => n17689);
   U20935 : NOR2_X1 port map( A1 => n29605, A2 => n17405, ZN => n16823);
   U20937 : INV_X1 port map( A => n17401, ZN => n17394);
   U20938 : INV_X1 port map( A => n16999, ZN => n17293);
   U20939 : NOR2_X1 port map( A1 => n17394, A2 => n17293, ZN => n16824);
   U20941 : OAI211_X1 port map( C1 => n17435, C2 => n29566, A => n17437, B => 
                           n336, ZN => n16828);
   U20942 : NAND2_X1 port map( A1 => n17298, A2 => n17413, ZN => n17412);
   U20943 : NAND2_X1 port map( A1 => n15811, A2 => n17413, ZN => n16830);
   U20945 : NAND3_X1 port map( A1 => n5430, A2 => n17297, A3 => n17411, ZN => 
                           n16829);
   U20946 : NAND2_X1 port map( A1 => n16922, A2 => n15811, ZN => n16832);
   U20947 : AOI21_X1 port map( B1 => n16985, B2 => n18188, A => n29044, ZN => 
                           n16842);
   U20948 : NOR2_X1 port map( A1 => n17553, A2 => n17554, ZN => n16834);
   U20949 : NOR2_X1 port map( A1 => n17555, A2 => n16908, ZN => n16833);
   U20951 : NAND2_X1 port map( A1 => n17312, A2 => n16918, ZN => n17563);
   U20952 : INV_X1 port map( A => n17563, ZN => n16839);
   U20953 : XNOR2_X1 port map( A => n19474, B => n18395, ZN => n16869);
   U20954 : NOR2_X1 port map( A1 => n17277, A2 => n17002, ZN => n17273);
   U20955 : NOR2_X1 port map( A1 => n17428, A2 => n28194, ZN => n16845);
   U20956 : OAI21_X1 port map( B1 => n16846, B2 => n16845, A => n17425, ZN => 
                           n16849);
   U20957 : OAI21_X1 port map( B1 => n16973, B2 => n17428, A => n2826, ZN => 
                           n16848);
   U20960 : NAND2_X1 port map( A1 => n17101, A2 => n16860, ZN => n16856);
   U20961 : NAND2_X1 port map( A1 => n16856, A2 => n17284, ZN => n16858);
   U20962 : NAND2_X1 port map( A1 => n16858, A2 => n16857, ZN => n16859);
   U20963 : NOR2_X1 port map( A1 => n16863, A2 => n29298, ZN => n16864);
   U20965 : NOR2_X1 port map( A1 => n18172, A2 => n18170, ZN => n17688);
   U20966 : NOR2_X1 port map( A1 => n17688, A2 => n17780, ZN => n16872);
   U20967 : NAND2_X1 port map( A1 => n28649, A2 => n16872, ZN => n16873);
   U20969 : NAND3_X1 port map( A1 => n17375, A2 => n17374, A3 => n16874, ZN => 
                           n16875);
   U20970 : NAND3_X1 port map( A1 => n17382, A2 => n17386, A3 => n17388, ZN => 
                           n18071);
   U20971 : NAND2_X1 port map( A1 => n16879, A2 => n17385, ZN => n18070);
   U20972 : INV_X1 port map( A => n16880, ZN => n16881);
   U20973 : MUX2_X1 port map( A => n17524, B => n17527, S => n17181, Z => 
                           n16886);
   U20974 : INV_X1 port map( A => n18516, ZN => n18078);
   U20975 : OAI211_X1 port map( C1 => n29127, C2 => n17138, A => n28574, B => 
                           n17501, ZN => n18073);
   U20976 : NOR2_X1 port map( A1 => n17139, A2 => n17138, ZN => n16889);
   U20977 : NOR2_X1 port map( A1 => n18508, A2 => n18507, ZN => n16896);
   U20978 : NOR2_X1 port map( A1 => n17153, A2 => n17148, ZN => n16890);
   U20979 : NOR2_X1 port map( A1 => n17148, A2 => n17489, ZN => n16891);
   U20980 : NAND2_X1 port map( A1 => n17488, A2 => n16891, ZN => n16894);
   U20981 : INV_X1 port map( A => n17076, ZN => n17149);
   U20982 : NAND3_X1 port map( A1 => n17153, A2 => n17489, A3 => n17149, ZN => 
                           n16893);
   U20983 : NAND3_X1 port map( A1 => n17487, A2 => n17147, A3 => n17148, ZN => 
                           n16892);
   U20985 : NAND2_X1 port map( A1 => n18509, A2 => n29057, ZN => n16895);
   U20986 : XNOR2_X1 port map( A => n18906, B => n19686, ZN => n16903);
   U20987 : AND2_X1 port map( A1 => n18203, A2 => n18277, ZN => n16899);
   U20988 : OAI21_X1 port map( B1 => n3994, B2 => n18203, A => n17803, ZN => 
                           n16897);
   U20989 : OAI21_X1 port map( B1 => n17803, B2 => n16899, A => n16897, ZN => 
                           n16901);
   U20990 : AOI22_X1 port map( A1 => n16899, A2 => n18276, B1 => n18279, B2 => 
                           n17696, ZN => n16900);
   U20991 : XNOR2_X1 port map( A => n19111, B => n25044, ZN => n16902);
   U20992 : XNOR2_X1 port map( A => n16903, B => n16902, ZN => n16983);
   U20993 : MUX2_X1 port map( A => n17707, B => n17573, S => n423, Z => n16905)
                           ;
   U20994 : NAND2_X1 port map( A1 => n29605, A2 => n17572, ZN => n17406);
   U20995 : NAND2_X1 port map( A1 => n17707, A2 => n17405, ZN => n17322);
   U20996 : AND2_X1 port map( A1 => n17322, A2 => n17406, ZN => n17706);
   U20997 : NAND2_X1 port map( A1 => n17038, A2 => n17568, ZN => n16907);
   U20998 : INV_X1 port map( A => n17557, ZN => n17219);
   U20999 : NOR2_X1 port map( A1 => n17555, A2 => n17219, ZN => n16910);
   U21000 : NOR2_X1 port map( A1 => n29142, A2 => n16908, ZN => n16909);
   U21001 : AOI22_X1 port map( A1 => n16910, A2 => n16911, B1 => n16909, B2 => 
                           n17553, ZN => n16915);
   U21002 : NOR2_X1 port map( A1 => n16911, A2 => n17555, ZN => n16912);
   U21003 : NAND2_X1 port map( A1 => n16913, A2 => n16912, ZN => n16914);
   U21004 : NOR2_X1 port map( A1 => n17562, A2 => n17315, ZN => n16920);
   U21005 : NOR2_X1 port map( A1 => n17316, A2 => n17560, ZN => n16919);
   U21006 : NAND2_X1 port map( A1 => n16921, A2 => n17301, ZN => n16923);
   U21007 : NAND2_X1 port map( A1 => n18263, A2 => n18324, ZN => n17985);
   U21008 : MUX2_X1 port map( A => n17434, B => n17309, S => n17435, Z => 
                           n16928);
   U21009 : INV_X1 port map( A => n17435, ZN => n16924);
   U21010 : NAND3_X1 port map( A1 => n16924, A2 => n529, A3 => n337, ZN => 
                           n16925);
   U21011 : INV_X1 port map( A => n18324, ZN => n17895);
   U21012 : OAI22_X1 port map( A1 => n17713, A2 => n17985, B1 => n29603, B2 => 
                           n17986, ZN => n16929);
   U21013 : NAND2_X1 port map( A1 => n16932, A2 => n17117, ZN => n18341);
   U21014 : NOR2_X1 port map( A1 => n18341, A2 => n18342, ZN => n17665);
   U21015 : OAI21_X1 port map( B1 => n17043, B2 => n17368, A => n17233, ZN => 
                           n16934);
   U21016 : MUX2_X1 port map( A => n17368, B => n17365, S => n17362, Z => 
                           n16933);
   U21017 : INV_X1 port map( A => n17335, ZN => n17342);
   U21018 : NOR2_X1 port map( A1 => n17338, A2 => n17342, ZN => n16935);
   U21019 : INV_X1 port map( A => n17542, ZN => n16941);
   U21020 : OAI21_X1 port map( B1 => n16941, B2 => n17539, A => n17540, ZN => 
                           n16942);
   U21021 : INV_X1 port map( A => n16943, ZN => n17242);
   U21022 : NAND2_X1 port map( A1 => n17552, A2 => n5398, ZN => n16945);
   U21023 : AOI22_X1 port map( A1 => n1121, A2 => n16949, B1 => n16948, B2 => 
                           n17029, ZN => n16950);
   U21024 : NOR2_X1 port map( A1 => n18538, A2 => n18527, ZN => n16956);
   U21025 : NOR2_X1 port map( A1 => n17356, A2 => n2449, ZN => n16952);
   U21026 : NOR2_X1 port map( A1 => n16953, A2 => n17359, ZN => n16954);
   U21027 : AND2_X1 port map( A1 => n17358, A2 => n16954, ZN => n18530);
   U21028 : MUX2_X1 port map( A => n17402, B => n17400, S => n17394, Z => 
                           n16961);
   U21029 : NOR2_X1 port map( A1 => n17400, A2 => n17396, ZN => n16959);
   U21030 : MUX2_X1 port map( A => n16959, B => n16958, S => n17402, Z => 
                           n16960);
   U21032 : NOR2_X1 port map( A1 => n17305, A2 => n16964, ZN => n16965);
   U21034 : INV_X1 port map( A => n16995, ZN => n16969);
   U21036 : NAND2_X1 port map( A1 => n6539, A2 => n29503, ZN => n16976);
   U21037 : NAND2_X1 port map( A1 => n17018, A2 => n17249, ZN => n16975);
   U21038 : MUX2_X1 port map( A => n16976, B => n16975, S => n17248, Z => 
                           n16979);
   U21039 : NAND2_X1 port map( A1 => n17248, A2 => n16977, ZN => n16978);
   U21040 : XNOR2_X1 port map( A => n19634, B => n19598, ZN => n16982);
   U21041 : INV_X1 port map( A => n18088, ZN => n16987);
   U21042 : INV_X1 port map( A => n16985, ZN => n16986);
   U21043 : OAI21_X1 port map( B1 => n527, B2 => n16987, A => n18186, ZN => 
                           n16988);
   U21044 : NOR2_X1 port map( A1 => n29600, A2 => n16991, ZN => n16994);
   U21045 : NAND2_X1 port map( A1 => n16994, A2 => n29298, ZN => n16997);
   U21046 : NAND2_X1 port map( A1 => n16992, A2 => n16995, ZN => n17264);
   U21047 : NAND3_X1 port map( A1 => n17277, A2 => n17002, A3 => n17271, ZN => 
                           n17003);
   U21049 : NOR2_X1 port map( A1 => n2825, A2 => n17426, ZN => n17006);
   U21050 : OAI211_X1 port map( C1 => n6927, C2 => n18600, A => n17014, B => 
                           n17990, ZN => n17024);
   U21052 : NAND2_X1 port map( A1 => n2656, A2 => n28142, ZN => n17023);
   U21053 : OAI211_X1 port map( C1 => n17018, C2 => n17249, A => n17017, B => 
                           n17016, ZN => n17019);
   U21054 : INV_X1 port map( A => n17019, ZN => n17020);
   U21055 : INV_X1 port map( A => n17854, ZN => n18599);
   U21056 : AND3_X1 port map( A1 => n29065, A2 => n28142, A3 => n18599, ZN => 
                           n17022);
   U21057 : AOI21_X2 port map( B1 => n17024, B2 => n17023, A => n17022, ZN => 
                           n19507);
   U21058 : NAND2_X1 port map( A1 => n17349, A2 => n17344, ZN => n17027);
   U21059 : NAND2_X1 port map( A1 => n17029, A2 => n17347, ZN => n17026);
   U21060 : INV_X1 port map( A => n18338, ZN => n18370);
   U21061 : OR2_X1 port map( A1 => n17199, A2 => n17356, ZN => n17036);
   U21062 : NAND2_X1 port map( A1 => n29546, A2 => n17195, ZN => n17033);
   U21063 : NAND3_X1 port map( A1 => n17358, A2 => n28793, A3 => n17033, ZN => 
                           n17035);
   U21064 : NOR2_X1 port map( A1 => n18370, A2 => n18332, ZN => n18001);
   U21065 : NAND2_X1 port map( A1 => n17569, A2 => n17568, ZN => n17039);
   U21066 : AOI21_X1 port map( B1 => n17040, B2 => n17039, A => n17038, ZN => 
                           n17041);
   U21067 : MUX2_X1 port map( A => n17045, B => n17044, S => n17366, Z => 
                           n17049);
   U21068 : NOR2_X1 port map( A1 => n18338, A2 => n18332, ZN => n17060);
   U21069 : INV_X1 port map( A => n17241, ZN => n17052);
   U21070 : NOR2_X1 port map( A1 => n17052, A2 => n17051, ZN => n17053);
   U21071 : MUX2_X2 port map( A => n17054, B => n17053, S => n5398, Z => n18337
                           );
   U21072 : NAND2_X1 port map( A1 => n17540, A2 => n17539, ZN => n17057);
   U21073 : INV_X1 port map( A => n17545, ZN => n17055);
   U21074 : AOI21_X1 port map( B1 => n17057, B2 => n5695, A => n15787, ZN => 
                           n17058);
   U21075 : XNOR2_X1 port map( A => n19507, B => n19096, ZN => n19628);
   U21076 : OAI21_X1 port map( B1 => n17497, B2 => n29373, A => n17063, ZN => 
                           n17064);
   U21077 : INV_X1 port map( A => n17206, ZN => n18591);
   U21078 : NOR2_X1 port map( A1 => n18591, A2 => n18588, ZN => n18596);
   U21080 : INV_X1 port map( A => n17506, ZN => n17071);
   U21081 : AND2_X1 port map( A1 => n17074, A2 => n17071, ZN => n17831);
   U21082 : MUX2_X1 port map( A => n17072, B => n17831, S => n17830, Z => 
                           n17075);
   U21083 : OR2_X2 port map( A1 => n17075, A2 => n17828, ZN => n18124);
   U21084 : NAND2_X1 port map( A1 => n5737, A2 => n17489, ZN => n17080);
   U21085 : NAND2_X1 port map( A1 => n17076, A2 => n17489, ZN => n17077);
   U21086 : NAND2_X1 port map( A1 => n17078, A2 => n17077, ZN => n17079);
   U21087 : MUX2_X1 port map( A => n17080, B => n17079, S => n17147, Z => 
                           n17081);
   U21088 : NOR2_X1 port map( A1 => n18124, A2 => n18128, ZN => n17082);
   U21089 : INV_X1 port map( A => n17515, ZN => n17085);
   U21090 : AOI22_X1 port map( A1 => n17840, A2 => n18595, B1 => n17835, B2 => 
                           n18124, ZN => n17089);
   U21091 : NAND2_X1 port map( A1 => n17090, A2 => n28800, ZN => n17096);
   U21092 : NOR2_X1 port map( A1 => n17093, A2 => n387, ZN => n17092);
   U21093 : AOI21_X1 port map( B1 => n17094, B2 => n17093, A => n17092, ZN => 
                           n17095);
   U21094 : INV_X1 port map( A => n18144, ZN => n17627);
   U21095 : OAI21_X1 port map( B1 => n17102, B2 => n1466, A => n17099, ZN => 
                           n17285);
   U21096 : NAND2_X1 port map( A1 => n17285, A2 => n17283, ZN => n17105);
   U21097 : NAND2_X1 port map( A1 => n17110, A2 => n17106, ZN => n17107);
   U21098 : NOR2_X1 port map( A1 => n17110, A2 => n17109, ZN => n17111);
   U21100 : INV_X1 port map( A => n17117, ZN => n17121);
   U21101 : INV_X1 port map( A => n17118, ZN => n17119);
   U21102 : NAND3_X1 port map( A1 => n17481, A2 => n3883, A3 => n17476, ZN => 
                           n17123);
   U21103 : NOR2_X1 port map( A1 => n28193, A2 => n17450, ZN => n17130);
   U21104 : AND2_X1 port map( A1 => n17130, A2 => n17454, ZN => n17131);
   U21105 : XNOR2_X1 port map( A => n18695, B => n19697, ZN => n17170);
   U21106 : AOI21_X1 port map( B1 => n17136, B2 => n17135, A => n28574, ZN => 
                           n17145);
   U21107 : NAND3_X1 port map( A1 => n17140, A2 => n17139, A3 => n17138, ZN => 
                           n17141);
   U21108 : OAI21_X1 port map( B1 => n17143, B2 => n17142, A => n17141, ZN => 
                           n17144);
   U21109 : AOI21_X1 port map( B1 => n17488, B2 => n17146, A => n17148, ZN => 
                           n17154);
   U21110 : NOR2_X1 port map( A1 => n17148, A2 => n17147, ZN => n17150);
   U21111 : OAI21_X1 port map( B1 => n17151, B2 => n17150, A => n17149, ZN => 
                           n17152);
   U21112 : AOI21_X1 port map( B1 => n17156, B2 => n17338, A => n17340, ZN => 
                           n17994);
   U21113 : INV_X1 port map( A => n17181, ZN => n17183);
   U21114 : NAND2_X1 port map( A1 => n17159, A2 => n17382, ZN => n17161);
   U21115 : NAND2_X1 port map( A1 => n18069, A2 => n17385, ZN => n17160);
   U21118 : INV_X1 port map( A => n18376, ZN => n18000);
   U21120 : AOI22_X1 port map( A1 => n18383, A2 => n17166, B1 => n17165, B2 => 
                           n18382, ZN => n17167);
   U21121 : XNOR2_X1 port map( A => n19412, B => n28097, ZN => n17169);
   U21122 : XNOR2_X1 port map( A => n17170, B => n17169, ZN => n17171);
   U21123 : INV_X1 port map( A => n20551, ZN => n17172);
   U21124 : MUX2_X1 port map( A => n29294, B => n17375, S => n17173, Z => 
                           n17180);
   U21126 : NAND2_X1 port map( A1 => n29294, A2 => n17374, ZN => n17176);
   U21127 : MUX2_X1 port map( A => n17177, B => n17176, S => n28776, Z => 
                           n17178);
   U21128 : NAND2_X1 port map( A1 => n17182, A2 => n17181, ZN => n17187);
   U21129 : OAI21_X1 port map( B1 => n17527, B2 => n16884, A => n531, ZN => 
                           n17184);
   U21130 : NAND2_X1 port map( A1 => n17184, A2 => n17183, ZN => n17186);
   U21131 : INV_X1 port map( A => n18122, ZN => n18418);
   U21132 : NOR2_X1 port map( A1 => n417, A2 => n18418, ZN => n17205);
   U21133 : NAND2_X1 port map( A1 => n17386, A2 => n29045, ZN => n17190);
   U21134 : NAND3_X1 port map( A1 => n17382, A2 => n17188, A3 => n18069, ZN => 
                           n17189);
   U21135 : AOI21_X1 port map( B1 => n1121, B2 => n5420, A => n17344, ZN => 
                           n17194);
   U21136 : NAND2_X1 port map( A1 => n17348, A2 => n17349, ZN => n17193);
   U21137 : INV_X1 port map( A => n18121, ZN => n18028);
   U21138 : OAI211_X1 port map( C1 => n2449, C2 => n17196, A => n17355, B => 
                           n17195, ZN => n17197);
   U21139 : NAND2_X1 port map( A1 => n17340, A2 => n17201, ZN => n17202);
   U21140 : AOI21_X1 port map( B1 => n18128, B2 => n18126, A => n18591, ZN => 
                           n17209);
   U21141 : NOR2_X1 port map( A1 => n18126, A2 => n18124, ZN => n17208);
   U21142 : XNOR2_X1 port map( A => n19243, B => n18690, ZN => n19665);
   U21143 : INV_X1 port map( A => n18426, ZN => n17212);
   U21144 : OAI21_X1 port map( B1 => n18042, B2 => n17802, A => n17824, ZN => 
                           n17211);
   U21145 : NAND2_X1 port map( A1 => n18423, A2 => n18421, ZN => n17210);
   U21146 : MUX2_X1 port map( A => n17540, B => n15787, S => n17213, Z => 
                           n17218);
   U21147 : NAND2_X1 port map( A1 => n17540, A2 => n17545, ZN => n17214);
   U21148 : MUX2_X1 port map( A => n17215, B => n17214, S => n15787, Z => 
                           n17216);
   U21149 : OAI21_X1 port map( B1 => n29142, B2 => n17221, A => n17554, ZN => 
                           n17222);
   U21150 : MUX2_X1 port map( A => n17223, B => n17222, S => n17556, Z => 
                           n17225);
   U21151 : OAI21_X1 port map( B1 => n29550, B2 => n17314, A => n17560, ZN => 
                           n17226);
   U21152 : NAND2_X1 port map( A1 => n17228, A2 => n17229, ZN => n17231);
   U21153 : AOI21_X1 port map( B1 => n17233, B2 => n17234, A => n17232, ZN => 
                           n17238);
   U21154 : AOI21_X1 port map( B1 => n17236, B2 => n17235, A => n17369, ZN => 
                           n17237);
   U21155 : NAND2_X1 port map( A1 => n17549, A2 => n16762, ZN => n17551);
   U21156 : NAND2_X1 port map( A1 => n17241, A2 => n17240, ZN => n17244);
   U21157 : NAND3_X1 port map( A1 => n17242, A2 => n4624, A3 => n5398, ZN => 
                           n17243);
   U21160 : XNOR2_X1 port map( A => n19246, B => n19617, ZN => n18722);
   U21161 : XNOR2_X1 port map( A => n18722, B => n19665, ZN => n17334);
   U21162 : MUX2_X1 port map( A => n1880, B => n17249, S => n17248, Z => n17253
                           );
   U21163 : NOR2_X1 port map( A1 => n17251, A2 => n29503, ZN => n17252);
   U21164 : INV_X1 port map( A => n18241, ZN => n17843);
   U21165 : NAND2_X1 port map( A1 => n17264, A2 => n17263, ZN => n17270);
   U21166 : NAND2_X1 port map( A1 => n17843, A2 => n17842, ZN => n17290);
   U21167 : NOR2_X1 port map( A1 => n17271, A2 => n17275, ZN => n17274);
   U21168 : NOR2_X1 port map( A1 => n18242, A2 => n17842, ZN => n17970);
   U21169 : NOR2_X1 port map( A1 => n28800, A2 => n17280, ZN => n17281);
   U21170 : NAND2_X1 port map( A1 => n17970, A2 => n17969, ZN => n17289);
   U21171 : NAND2_X1 port map( A1 => n17285, A2 => n17284, ZN => n17286);
   U21172 : NOR2_X1 port map( A1 => n17969, A2 => n18236, ZN => n17287);
   U21173 : OAI21_X1 port map( B1 => n17607, B2 => n17287, A => n18241, ZN => 
                           n17288);
   U21175 : OAI211_X1 port map( C1 => n17400, C2 => n17294, A => n29572, B => 
                           n17293, ZN => n17295);
   U21176 : INV_X1 port map( A => n17411, ZN => n17416);
   U21178 : INV_X1 port map( A => n17423, ZN => n17615);
   U21181 : OAI21_X1 port map( B1 => n17309, B2 => n17439, A => n17308, ZN => 
                           n17311);
   U21182 : MUX2_X1 port map( A => n17435, B => n17309, S => n17438, Z => 
                           n17310);
   U21183 : INV_X1 port map( A => n18156, ZN => n18153);
   U21184 : INV_X1 port map( A => n17826, ZN => n18154);
   U21185 : INV_X1 port map( A => n17405, ZN => n17575);
   U21186 : NOR2_X1 port map( A1 => n17707, A2 => n17575, ZN => n17319);
   U21187 : MUX2_X1 port map( A => n17319, B => n17318, S => n17710, Z => 
                           n17324);
   U21188 : NAND2_X1 port map( A1 => n17320, A2 => n17575, ZN => n17321);
   U21189 : AOI21_X1 port map( B1 => n17322, B2 => n17321, A => n29513, ZN => 
                           n17323);
   U21190 : NOR2_X2 port map( A1 => n17324, A2 => n17323, ZN => n18032);
   U21191 : INV_X1 port map( A => n18032, ZN => n17745);
   U21192 : NAND3_X1 port map( A1 => n17745, A2 => n18160, A3 => n18153, ZN => 
                           n17325);
   U21193 : XNOR2_X1 port map( A => n29554, B => n29038, ZN => n17332);
   U21195 : XNOR2_X1 port map( A => n19136, B => n26531, ZN => n17331);
   U21196 : XNOR2_X1 port map( A => n17332, B => n17331, ZN => n17333);
   U21197 : NOR2_X1 port map( A1 => n17340, A2 => n17335, ZN => n17337);
   U21199 : NAND3_X1 port map( A1 => n17346, A2 => n17345, A3 => n29632, ZN => 
                           n17352);
   U21200 : OAI21_X1 port map( B1 => n17365, B2 => n17362, A => n17361, ZN => 
                           n17363);
   U21201 : NAND2_X1 port map( A1 => n17364, A2 => n17363, ZN => n17372);
   U21202 : NAND2_X1 port map( A1 => n17366, A2 => n17365, ZN => n17371);
   U21203 : NOR2_X1 port map( A1 => n17368, A2 => n15731, ZN => n17370);
   U21204 : OAI21_X1 port map( B1 => n29636, B2 => n530, A => n17374, ZN => 
                           n17380);
   U21205 : NAND2_X1 port map( A1 => n17375, A2 => n17374, ZN => n17376);
   U21206 : NAND2_X1 port map( A1 => n17377, A2 => n17376, ZN => n17378);
   U21207 : AND2_X1 port map( A1 => n28558, A2 => n18404, ZN => n17381);
   U21208 : NAND2_X1 port map( A1 => n18707, A2 => n17381, ZN => n18712);
   U21209 : OAI21_X1 port map( B1 => n17382, B2 => n29045, A => n17385, ZN => 
                           n17383);
   U21210 : NOR2_X1 port map( A1 => n17388, A2 => n29045, ZN => n17390);
   U21211 : OAI211_X1 port map( C1 => n18707, C2 => n17392, A => n18712, B => 
                           n17391, ZN => n17446);
   U21212 : OAI21_X1 port map( B1 => n17397, B2 => n17396, A => n17395, ZN => 
                           n17398);
   U21213 : NAND2_X1 port map( A1 => n17406, A2 => n17405, ZN => n17407);
   U21214 : NAND2_X1 port map( A1 => n5430, A2 => n17415, ZN => n17410);
   U21215 : NAND3_X1 port map( A1 => n17412, A2 => n17411, A3 => n17410, ZN => 
                           n17419);
   U21216 : NAND3_X1 port map( A1 => n17415, A2 => n17414, A3 => n17413, ZN => 
                           n17418);
   U21217 : NAND3_X1 port map( A1 => n18232, A2 => n17977, A3 => n18231, ZN => 
                           n17445);
   U21218 : INV_X1 port map( A => n17425, ZN => n17427);
   U21219 : NAND2_X1 port map( A1 => n17427, A2 => n17426, ZN => n17429);
   U21220 : MUX2_X1 port map( A => n17429, B => n17428, S => n28792, Z => 
                           n17430);
   U21221 : INV_X1 port map( A => n18398, ZN => n17442);
   U21222 : NAND2_X1 port map( A1 => n17438, A2 => n17437, ZN => n17441);
   U21223 : NAND3_X1 port map( A1 => n17442, A2 => n18399, A3 => n18234, ZN => 
                           n17444);
   U21224 : NAND3_X1 port map( A1 => n18232, A2 => n18400, A3 => n18233, ZN => 
                           n17443);
   U21225 : XNOR2_X1 port map( A => n19468, B => n17446, ZN => n19639);
   U21226 : NAND3_X1 port map( A1 => n17762, A2 => n519, A3 => n517, ZN => 
                           n17448);
   U21227 : AOI21_X1 port map( B1 => n17762, B2 => n17872, A => n17941, ZN => 
                           n17447);
   U21228 : XNOR2_X1 port map( A => n18942, B => n27737, ZN => n17449);
   U21229 : XNOR2_X1 port map( A => n19639, B => n17449, ZN => n17581);
   U21230 : NOR2_X1 port map( A1 => n17451, A2 => n17450, ZN => n17453);
   U21231 : NAND2_X1 port map( A1 => n17466, A2 => n17463, ZN => n17465);
   U21232 : MUX2_X1 port map( A => n17467, B => n17465, S => n17464, Z => 
                           n17468);
   U21233 : NAND2_X1 port map( A1 => n17516, A2 => n17469, ZN => n17514);
   U21234 : OR2_X1 port map( A1 => n17514, A2 => n17470, ZN => n17471);
   U21235 : NOR2_X1 port map( A1 => n17477, A2 => n17476, ZN => n17479);
   U21236 : NOR2_X1 port map( A1 => n17505, A2 => n4270, ZN => n17482);
   U21238 : NAND2_X1 port map( A1 => n17484, A2 => n17506, ZN => n17507);
   U21239 : OAI21_X1 port map( B1 => n16736, B2 => n17487, A => n17486, ZN => 
                           n17490);
   U21240 : NOR2_X1 port map( A1 => n17492, A2 => n17491, ZN => n17494);
   U21241 : OAI21_X1 port map( B1 => n17495, B2 => n17494, A => n17493, ZN => 
                           n18226);
   U21243 : NAND2_X1 port map( A1 => n18388, A2 => n18393, ZN => n18229);
   U21244 : OAI211_X1 port map( C1 => n17506, C2 => n17505, A => n17507, B => 
                           n17829, ZN => n17511);
   U21245 : INV_X1 port map( A => n17507, ZN => n17509);
   U21246 : NAND2_X1 port map( A1 => n17509, A2 => n17508, ZN => n17510);
   U21247 : NAND2_X1 port map( A1 => n17515, A2 => n17514, ZN => n17521);
   U21248 : OAI21_X1 port map( B1 => n17518, B2 => n17517, A => n17516, ZN => 
                           n17519);
   U21249 : AOI21_X1 port map( B1 => n5234, B2 => n18393, A => n18227, ZN => 
                           n17522);
   U21250 : INV_X1 port map( A => n17522, ZN => n17523);
   U21252 : OAI21_X1 port map( B1 => n17526, B2 => n16884, A => n17524, ZN => 
                           n17530);
   U21253 : OAI21_X1 port map( B1 => n17528, B2 => n17527, A => n4979, ZN => 
                           n17529);
   U21254 : INV_X1 port map( A => n18387, ZN => n18391);
   U21255 : NAND3_X1 port map( A1 => n5233, A2 => n18227, A3 => n18391, ZN => 
                           n17533);
   U21256 : XNOR2_X1 port map( A => n19122, B => n19377, ZN => n17579);
   U21258 : NOR2_X1 port map( A1 => n17969, A2 => n18243, ZN => n17536);
   U21259 : NOR2_X1 port map( A1 => n18241, A2 => n18236, ZN => n17535);
   U21260 : NAND2_X1 port map( A1 => n18243, A2 => n18241, ZN => n17966);
   U21261 : NOR2_X1 port map( A1 => n17542, A2 => n28454, ZN => n17544);
   U21262 : MUX2_X1 port map( A => n16908, B => n17554, S => n17553, Z => 
                           n17559);
   U21263 : MUX2_X1 port map( A => n17556, B => n17555, S => n17554, Z => 
                           n17558);
   U21264 : INV_X1 port map( A => n17564, ZN => n18253);
   U21265 : NAND2_X1 port map( A1 => n17573, A2 => n17572, ZN => n17574);
   U21266 : XNOR2_X1 port map( A => n19373, B => n19555, ZN => n19574);
   U21267 : XNOR2_X1 port map( A => n19574, B => n17579, ZN => n17580);
   U21268 : XNOR2_X1 port map( A => n17581, B => n17580, ZN => n19855);
   U21269 : NAND2_X1 port map( A1 => n18251, A2 => n18253, ZN => n17582);
   U21270 : INV_X1 port map( A => n6912, ZN => n17962);
   U21271 : AOI21_X1 port map( B1 => n17583, B2 => n17772, A => n18251, ZN => 
                           n17584);
   U21273 : NAND2_X1 port map( A1 => n18214, A2 => n18506, ZN => n17588);
   U21274 : NOR2_X1 port map( A1 => n18500, A2 => n520, ZN => n17586);
   U21275 : NAND2_X1 port map( A1 => n18215, A2 => n17586, ZN => n17587);
   U21276 : NAND2_X1 port map( A1 => n17588, A2 => n17587, ZN => n17591);
   U21277 : NAND2_X1 port map( A1 => n520, A2 => n2363, ZN => n17589);
   U21278 : NAND2_X1 port map( A1 => n18388, A2 => n18387, ZN => n17596);
   U21279 : INV_X1 port map( A => n18389, ZN => n17593);
   U21280 : NAND2_X1 port map( A1 => n17593, A2 => n17592, ZN => n17595);
   U21281 : MUX2_X1 port map( A => n18707, B => n18706, S => n18404, Z => 
                           n17600);
   U21282 : NOR2_X1 port map( A1 => n18707, A2 => n18404, ZN => n17599);
   U21283 : XNOR2_X1 port map( A => n19615, B => n29038, ZN => n17604);
   U21284 : XNOR2_X1 port map( A => n19490, B => n26665, ZN => n17603);
   U21285 : XNOR2_X1 port map( A => n17604, B => n17603, ZN => n17605);
   U21286 : AOI21_X1 port map( B1 => n17757, B2 => n17756, A => n18240, ZN => 
                           n17608);
   U21287 : XNOR2_X1 port map( A => n18799, B => n19256, ZN => n17623);
   U21289 : AOI21_X1 port map( B1 => n17610, B2 => n18431, A => n18148, ZN => 
                           n17611);
   U21291 : NAND3_X1 port map( A1 => n17615, A2 => n17614, A3 => n17613, ZN => 
                           n17618);
   U21292 : INV_X1 port map( A => n17616, ZN => n17617);
   U21293 : NAND2_X1 port map( A1 => n17825, A2 => n18033, ZN => n17619);
   U21294 : OAI21_X1 port map( B1 => n18160, B2 => n18156, A => n17619, ZN => 
                           n18036);
   U21295 : AOI21_X1 port map( B1 => n17621, B2 => n17620, A => n18153, ZN => 
                           n17622);
   U21296 : XNOR2_X1 port map( A => n18408, B => n18738, ZN => n19362);
   U21297 : XNOR2_X1 port map( A => n17623, B => n19362, ZN => n17631);
   U21298 : NAND2_X1 port map( A1 => n18028, A2 => n18414, ZN => n17624);
   U21299 : OAI21_X1 port map( B1 => n18413, B2 => n18122, A => n17624, ZN => 
                           n17625);
   U21300 : NAND2_X1 port map( A1 => n18137, A2 => n17847, ZN => n17626);
   U21301 : XNOR2_X1 port map( A => n18735, B => n19584, ZN => n17629);
   U21302 : XNOR2_X1 port map( A => n18949, B => n1079, ZN => n17628);
   U21303 : XNOR2_X1 port map( A => n17628, B => n17629, ZN => n17630);
   U21304 : NAND2_X1 port map( A1 => n20414, A2 => n20941, ZN => n17686);
   U21305 : INV_X1 port map( A => n20414, ZN => n20192);
   U21306 : NOR2_X1 port map( A1 => n18124, A2 => n18589, ZN => n18592);
   U21309 : NOR2_X1 port map( A1 => n17846, A2 => n18137, ZN => n17635);
   U21310 : NAND2_X1 port map( A1 => n17635, A2 => n17845, ZN => n17638);
   U21311 : NAND3_X1 port map( A1 => n18137, A2 => n526, A3 => n17847, ZN => 
                           n17637);
   U21312 : XNOR2_X1 port map( A => n19215, B => n19305, ZN => n17644);
   U21313 : NAND2_X1 port map( A1 => n18087, A2 => n18188, ZN => n17642);
   U21314 : NOR2_X1 port map( A1 => n18190, A2 => n29125, ZN => n17641);
   U21315 : OAI211_X1 port map( C1 => n17642, C2 => n17641, A => n17640, B => 
                           n17797, ZN => n19339);
   U21316 : XNOR2_X1 port map( A => n19339, B => n1187, ZN => n17643);
   U21317 : XNOR2_X1 port map( A => n17644, B => n17643, ZN => n17656);
   U21319 : INV_X1 port map( A => n18382, ZN => n17645);
   U21320 : NAND2_X1 port map( A1 => n17645, A2 => n18379, ZN => n18349);
   U21321 : NAND3_X1 port map( A1 => n17883, A2 => n17647, A3 => n18376, ZN => 
                           n17646);
   U21323 : NAND2_X1 port map( A1 => n17883, A2 => n18376, ZN => n18348);
   U21324 : NAND3_X1 port map( A1 => n18348, A2 => n17647, A3 => n18380, ZN => 
                           n17648);
   U21325 : XNOR2_X1 port map( A => n19686, B => n19108, ZN => n17654);
   U21326 : INV_X1 port map( A => n6927, ZN => n17890);
   U21327 : NOR2_X1 port map( A1 => n18338, A2 => n18372, ZN => n17653);
   U21328 : XNOR2_X1 port map( A => n18773, B => n19632, ZN => n19597);
   U21329 : XNOR2_X1 port map( A => n19597, B => n17654, ZN => n17655);
   U21331 : NOR2_X1 port map( A1 => n18465, A2 => n18471, ZN => n18008);
   U21332 : NAND2_X1 port map( A1 => n18008, A2 => n18469, ZN => n17658);
   U21333 : NAND2_X1 port map( A1 => n18314, A2 => n6079, ZN => n17657);
   U21335 : XNOR2_X1 port map( A => n18942, B => n3219, ZN => n17662);
   U21336 : XNOR2_X1 port map( A => n19123, B => n17662, ZN => n17670);
   U21337 : INV_X1 port map( A => n18341, ZN => n17908);
   U21338 : OAI21_X1 port map( B1 => n17908, B2 => n514, A => n18343, ZN => 
                           n17664);
   U21339 : INV_X1 port map( A => n17947, ZN => n18346);
   U21340 : NOR2_X1 port map( A1 => n16611, A2 => n18312, ZN => n17666);
   U21341 : INV_X1 port map( A => n18311, ZN => n18357);
   U21342 : XNOR2_X1 port map( A => n19465, B => n19232, ZN => n17669);
   U21343 : XNOR2_X1 port map( A => n17670, B => n17669, ZN => n17684);
   U21344 : NAND3_X1 port map( A1 => n29561, A2 => n18298, A3 => n18059, ZN => 
                           n17673);
   U21345 : INV_X1 port map( A => n18057, ZN => n17671);
   U21346 : NAND2_X1 port map( A1 => n18298, A2 => n1861, ZN => n17672);
   U21347 : NOR2_X1 port map( A1 => n18493, A2 => n28632, ZN => n18297);
   U21349 : MUX2_X1 port map( A => n17674, B => n28633, S => n18488, Z => 
                           n17676);
   U21350 : XNOR2_X1 port map( A => n29318, B => n18520, ZN => n17683);
   U21351 : NOR2_X1 port map( A1 => n18476, A2 => n18305, ZN => n17677);
   U21352 : NAND2_X1 port map( A1 => n17677, A2 => n18478, ZN => n17678);
   U21353 : OAI21_X1 port map( B1 => n18477, B2 => n18012, A => n17678, ZN => 
                           n17682);
   U21354 : NOR2_X1 port map( A1 => n18476, A2 => n18306, ZN => n18310);
   U21355 : INV_X1 port map( A => n18306, ZN => n18474);
   U21356 : INV_X1 port map( A => n17679, ZN => n17934);
   U21357 : NOR3_X1 port map( A1 => n18310, A2 => n18011, A3 => n17680, ZN => 
                           n17681);
   U21358 : XNOR2_X1 port map( A => n17683, B => n19637, ZN => n19336);
   U21359 : INV_X1 port map( A => n17687, ZN => n20193);
   U21360 : NOR2_X1 port map( A1 => n20414, A2 => n20193, ZN => n17753);
   U21361 : XNOR2_X1 port map( A => n19707, B => n29247, ZN => n17690);
   U21362 : NOR2_X1 port map( A1 => n510, A2 => n18078, ZN => n17692);
   U21363 : NOR2_X1 port map( A1 => n18510, A2 => n18508, ZN => n17691);
   U21365 : INV_X1 port map( A => n18277, ZN => n18275);
   U21366 : XNOR2_X1 port map( A => n19194, B => n18913, ZN => n17697);
   U21368 : NAND2_X1 port map( A1 => n17700, A2 => n17699, ZN => n17705);
   U21369 : AND2_X1 port map( A1 => n18529, A2 => n18537, ZN => n17701);
   U21370 : NOR3_X1 port map( A1 => n18260, A2 => n17864, A3 => n18529, ZN => 
                           n17702);
   U21371 : INV_X1 port map( A => n17706, ZN => n17711);
   U21372 : OAI21_X1 port map( B1 => n423, B2 => n17707, A => n17710, ZN => 
                           n17708);
   U21373 : OAI22_X1 port map( A1 => n17711, A2 => n17710, B1 => n17709, B2 => 
                           n17708, ZN => n17712);
   U21374 : INV_X1 port map( A => n18325, ZN => n18322);
   U21375 : OR2_X1 port map( A1 => n17717, A2 => n17431, ZN => n17718);
   U21377 : XNOR2_X1 port map( A => n18369, B => n28623, ZN => n17725);
   U21378 : XNOR2_X1 port map( A => n17725, B => n19603, ZN => n19357);
   U21379 : XNOR2_X1 port map( A => n17726, B => n19357, ZN => n19747);
   U21380 : BUF_X2 port map( A => n19747, Z => n20577);
   U21381 : AOI21_X2 port map( B1 => n17728, B2 => n18217, A => n17727, ZN => 
                           n19321);
   U21382 : INV_X1 port map( A => n18107, ZN => n18455);
   U21383 : XNOR2_X1 port map( A => n19321, B => n19626, ZN => n17742);
   U21385 : INV_X1 port map( A => n17592, ZN => n17732);
   U21387 : INV_X1 port map( A => n18227, ZN => n17766);
   U21388 : AND2_X1 port map( A1 => n18390, A2 => n17766, ZN => n17735);
   U21389 : NAND2_X1 port map( A1 => n5233, A2 => n17592, ZN => n17734);
   U21391 : INV_X1 port map( A => n17965, ZN => n18960);
   U21392 : NOR2_X1 port map( A1 => n18441, A2 => n18179, ZN => n17737);
   U21393 : OAI21_X1 port map( B1 => n18444, B2 => n18181, A => n17737, ZN => 
                           n17740);
   U21396 : XNOR2_X1 port map( A => n19331, B => n18960, ZN => n17741);
   U21397 : XNOR2_X1 port map( A => n17741, B => n17742, ZN => n17752);
   U21398 : NAND2_X1 port map( A1 => n18156, A2 => n18154, ZN => n18035);
   U21399 : NOR2_X1 port map( A1 => n18160, A2 => n18032, ZN => n18157);
   U21400 : NAND2_X1 port map( A1 => n18159, A2 => n18034, ZN => n17744);
   U21401 : AND2_X1 port map( A1 => n18032, A2 => n18033, ZN => n17743);
   U21402 : NAND3_X1 port map( A1 => n17746, A2 => n29502, A3 => n18193, ZN => 
                           n17748);
   U21403 : INV_X1 port map( A => n18449, ZN => n18450);
   U21404 : NOR2_X1 port map( A1 => n18450, A2 => n18198, ZN => n17747);
   U21405 : XNOR2_X1 port map( A => n19332, B => n18856, ZN => n17750);
   U21406 : XNOR2_X1 port map( A => n19697, B => n3666, ZN => n17749);
   U21407 : XNOR2_X1 port map( A => n17750, B => n17749, ZN => n17751);
   U21408 : AOI22_X1 port map( A1 => n17753, A2 => n20577, B1 => n503, B2 => 
                           n20412, ZN => n17754);
   U21409 : NOR2_X1 port map( A1 => n18506, A2 => n18500, ZN => n17755);
   U21410 : NOR2_X1 port map( A1 => n4725, A2 => n18236, ZN => n17759);
   U21411 : NAND2_X1 port map( A1 => n18240, A2 => n17842, ZN => n17758);
   U21412 : OAI211_X1 port map( C1 => n17977, C2 => n18402, A => n18399, B => 
                           n18400, ZN => n17760);
   U21413 : OAI211_X1 port map( C1 => n18397, C2 => n17977, A => n18396, B => 
                           n17760, ZN => n19535);
   U21414 : XNOR2_X1 port map( A => n19084, B => n19045, ZN => n17779);
   U21415 : INV_X1 port map( A => n17761, ZN => n17765);
   U21416 : OAI22_X1 port map( A1 => n17937, A2 => n517, B1 => n17941, B2 => 
                           n17762, ZN => n17873);
   U21417 : NAND2_X1 port map( A1 => n18393, A2 => n17592, ZN => n17769);
   U21418 : NAND3_X1 port map( A1 => n17767, A2 => n18387, A3 => n18227, ZN => 
                           n17768);
   U21420 : OAI21_X1 port map( B1 => n18019, B2 => n1888, A => n17773, ZN => 
                           n17775);
   U21421 : XNOR2_X1 port map( A => n19481, B => n19685, ZN => n18670);
   U21425 : XNOR2_X1 port map( A => n18675, B => n19378, ZN => n17801);
   U21426 : NOR2_X1 port map( A1 => n16985, A2 => n29125, ZN => n17794);
   U21427 : NAND2_X1 port map( A1 => n18087, A2 => n17794, ZN => n19564);
   U21428 : OAI21_X1 port map( B1 => n18087, B2 => n19560, A => n29044, ZN => 
                           n17795);
   U21429 : OAI21_X1 port map( B1 => n17796, B2 => n29044, A => n17795, ZN => 
                           n19559);
   U21430 : OAI211_X1 port map( C1 => n18188, C2 => n17797, A => n19564, B => 
                           n19559, ZN => n19299);
   U21432 : XNOR2_X1 port map( A => n19077, B => n17801, ZN => n17813);
   U21433 : XNOR2_X1 port map( A => n28530, B => n3622, ZN => n17811);
   U21434 : NAND3_X1 port map( A1 => n18450, A2 => n29502, A3 => n6663, ZN => 
                           n17808);
   U21436 : XNOR2_X1 port map( A => n29492, B => n19679, ZN => n19156);
   U21437 : XNOR2_X1 port map( A => n19156, B => n17811, ZN => n17812);
   U21438 : XNOR2_X1 port map( A => n17813, B => n17812, ZN => n20310);
   U21439 : INV_X1 port map( A => n20310, ZN => n20584);
   U21442 : XNOR2_X1 port map( A => n19283, B => n19278, ZN => n19105);
   U21443 : XNOR2_X1 port map( A => n19105, B => n19285, ZN => n17853);
   U21444 : INV_X1 port map( A => n17828, ZN => n17833);
   U21445 : OAI21_X1 port map( B1 => n17835, B2 => n17838, A => n17834, ZN => 
                           n17836);
   U21446 : NAND2_X1 port map( A1 => n17840, A2 => n18128, ZN => n17841);
   U21448 : NAND2_X1 port map( A1 => n18241, A2 => n17842, ZN => n18239);
   U21449 : XNOR2_X1 port map( A => n19704, B => n19354, ZN => n17851);
   U21450 : XNOR2_X1 port map( A => n17851, B => n17850, ZN => n17852);
   U21451 : XNOR2_X2 port map( A => n17853, B => n17852, ZN => n20585);
   U21452 : AOI22_X1 port map( A1 => n17890, A2 => n18366, B1 => n18367, B2 => 
                           n2656, ZN => n17855);
   U21453 : OR2_X1 port map( A1 => n17855, A2 => n17854, ZN => n17857);
   U21454 : AND2_X2 port map( A1 => n17857, A2 => n17856, ZN => n19359);
   U21455 : OAI22_X1 port map( A1 => n17858, A2 => n374, B1 => n18286, B2 => 
                           n18081, ZN => n17860);
   U21456 : XNOR2_X1 port map( A => n19359, B => n19251, ZN => n17865);
   U21457 : AOI21_X1 port map( B1 => n18508, B2 => n18507, A => n18510, ZN => 
                           n17862);
   U21458 : XNOR2_X1 port map( A => n19725, B => n19475, ZN => n18681);
   U21459 : XNOR2_X1 port map( A => n17865, B => n18681, ZN => n17879);
   U21460 : NOR2_X1 port map( A1 => n18500, A2 => n18213, ZN => n18503);
   U21461 : NOR2_X1 port map( A1 => n515, A2 => n17868, ZN => n17869);
   U21464 : AOI22_X1 port map( A1 => n18063, A2 => n18064, B1 => n18057, B2 => 
                           n17926, ZN => n18303);
   U21465 : AOI21_X1 port map( B1 => n17928, B2 => n1861, A => n18059, ZN => 
                           n17871);
   U21466 : XNOR2_X1 port map( A => n18760, B => n19727, ZN => n17877);
   U21467 : AOI21_X1 port map( B1 => n17939, B2 => n28656, A => n517, ZN => 
                           n17875);
   U21468 : INV_X1 port map( A => n17942, ZN => n17938);
   U21469 : XNOR2_X1 port map( A => n19643, B => n1175, ZN => n17876);
   U21470 : XNOR2_X1 port map( A => n17877, B => n17876, ZN => n17878);
   U21471 : XNOR2_X1 port map( A => n17879, B => n17878, ZN => n17954);
   U21472 : INV_X1 port map( A => n18350, ZN => n17882);
   U21473 : NOR2_X1 port map( A1 => n18382, A2 => n18379, ZN => n18378);
   U21474 : AOI22_X1 port map( A1 => n17882, A2 => n18000, B1 => n18378, B2 => 
                           n5383, ZN => n17886);
   U21475 : NAND3_X1 port map( A1 => n18383, A2 => n18382, A3 => n17883, ZN => 
                           n17885);
   U21476 : MUX2_X1 port map( A => n18337, B => n18372, S => n18333, Z => 
                           n17887);
   U21477 : INV_X1 port map( A => n18334, ZN => n18371);
   U21479 : NOR2_X1 port map( A1 => n17890, A2 => n29065, ZN => n17891);
   U21480 : NOR2_X1 port map( A1 => n17892, A2 => n6927, ZN => n17893);
   U21481 : MUX2_X1 port map( A => n18262, B => n17895, S => n18325, Z => 
                           n17897);
   U21482 : XNOR2_X1 port map( A => n19315, B => n19066, ZN => n17913);
   U21483 : NOR2_X1 port map( A1 => n18311, A2 => n16611, ZN => n17899);
   U21484 : INV_X1 port map( A => n18354, ZN => n17898);
   U21485 : INV_X1 port map( A => n18312, ZN => n18355);
   U21486 : NOR2_X1 port map( A1 => n17918, A2 => n18355, ZN => n17900);
   U21488 : XNOR2_X1 port map( A => n18778, B => n19346, ZN => n17911);
   U21489 : NOR2_X1 port map( A1 => n18343, A2 => n18344, ZN => n17909);
   U21490 : NOR2_X1 port map( A1 => n514, A2 => n17947, ZN => n17907);
   U21491 : XNOR2_X1 port map( A => n18646, B => n2274, ZN => n17910);
   U21492 : XNOR2_X1 port map( A => n17911, B => n17910, ZN => n17912);
   U21493 : XNOR2_X1 port map( A => n17913, B => n17912, ZN => n19827);
   U21494 : NOR2_X1 port map( A1 => n20585, A2 => n19827, ZN => n17956);
   U21496 : OAI21_X1 port map( B1 => n145, B2 => n17917, A => n18472, ZN => 
                           n19173);
   U21499 : XNOR2_X1 port map( A => n18628, B => n19692, ZN => n17932);
   U21500 : AOI21_X1 port map( B1 => n18493, B2 => n18292, A => n28633, ZN => 
                           n17925);
   U21501 : NOR2_X1 port map( A1 => n18489, A2 => n18488, ZN => n18293);
   U21502 : AOI21_X1 port map( B1 => n18015, B2 => n18489, A => n18293, ZN => 
                           n17924);
   U21503 : OR2_X1 port map( A1 => n18292, A2 => n18489, ZN => n17923);
   U21504 : OAI21_X1 port map( B1 => n17925, B2 => n17924, A => n17923, ZN => 
                           n18806);
   U21505 : NAND2_X1 port map( A1 => n17928, A2 => n18064, ZN => n17931);
   U21506 : NOR2_X1 port map( A1 => n29561, A2 => n17926, ZN => n17927);
   U21507 : XNOR2_X1 port map( A => n19508, B => n18806, ZN => n19322);
   U21508 : XNOR2_X1 port map( A => n19322, B => n17932, ZN => n17953);
   U21509 : NAND2_X1 port map( A1 => n18304, A2 => n17934, ZN => n17935);
   U21510 : INV_X1 port map( A => n18305, ZN => n18479);
   U21511 : OAI22_X1 port map( A1 => n18477, A2 => n17935, B1 => n18480, B2 => 
                           n18479, ZN => n17936);
   U21512 : NAND2_X1 port map( A1 => n17944, A2 => n17943, ZN => n17945);
   U21513 : XNOR2_X1 port map( A => n19267, B => n19323, ZN => n19095);
   U21515 : NAND3_X1 port map( A1 => n17948, A2 => n17947, A3 => n514, ZN => 
                           n17949);
   U21516 : XNOR2_X1 port map( A => n19622, B => n3654, ZN => n17951);
   U21517 : XNOR2_X1 port map( A => n19095, B => n17951, ZN => n17952);
   U21518 : XNOR2_X1 port map( A => n17953, B => n17952, ZN => n20196);
   U21519 : NOR2_X1 port map( A1 => n20196, A2 => n29144, ZN => n17955);
   U21520 : MUX2_X1 port map( A => n17956, B => n17955, S => n20311, Z => 
                           n17957);
   U21521 : NOR2_X1 port map( A1 => n17960, A2 => n17959, ZN => n17964);
   U21522 : OAI22_X1 port map( A1 => n17961, A2 => n18253, B1 => n18018, B2 => 
                           n524, ZN => n17963);
   U21523 : AOI21_X2 port map( B1 => n17964, B2 => n17963, A => n17962, ZN => 
                           n19691);
   U21524 : XNOR2_X1 port map( A => n17965, B => n19691, ZN => n19210);
   U21525 : INV_X1 port map( A => n17966, ZN => n17968);
   U21526 : OAI21_X1 port map( B1 => n17968, B2 => n17967, A => n18240, ZN => 
                           n17973);
   U21527 : AOI22_X1 port map( A1 => n29034, A2 => n17970, B1 => n17969, B2 => 
                           n4725, ZN => n17972);
   U21528 : XNOR2_X1 port map( A => n17974, B => n19409, ZN => n17975);
   U21529 : XNOR2_X1 port map( A => n17975, B => n19210, ZN => n17984);
   U21530 : NAND3_X1 port map( A1 => n17977, A2 => n18233, A3 => n18402, ZN => 
                           n17978);
   U21531 : XNOR2_X1 port map( A => n19321, B => n17982, ZN => n17983);
   U21532 : XNOR2_X1 port map( A => n17984, B => n17983, ZN => n20199);
   U21533 : NOR2_X1 port map( A1 => n18262, A2 => n18261, ZN => n17987);
   U21534 : XNOR2_X1 port map( A => n18812, B => n19462, ZN => n17991);
   U21535 : XNOR2_X1 port map( A => n18815, B => n17991, ZN => n18005);
   U21536 : OR3_X1 port map( A1 => n18383, A2 => n18382, A3 => n18376, ZN => 
                           n17999);
   U21537 : INV_X1 port map( A => n17992, ZN => n17993);
   U21538 : NAND2_X1 port map( A1 => n17993, A2 => n2048, ZN => n17995);
   U21539 : NOR3_X1 port map( A1 => n18379, A2 => n17995, A3 => n17994, ZN => 
                           n17996);
   U21540 : XNOR2_X1 port map( A => n19428, B => n19232, ZN => n19557);
   U21541 : XNOR2_X1 port map( A => n19427, B => n3483, ZN => n18003);
   U21542 : XNOR2_X1 port map( A => n19557, B => n18003, ZN => n18004);
   U21543 : NAND2_X1 port map( A1 => n20199, A2 => n20200, ZN => n20121);
   U21544 : INV_X1 port map( A => n18466, ZN => n18006);
   U21545 : NOR3_X1 port map( A1 => n18465, A2 => n18467, A3 => n18006, ZN => 
                           n18007);
   U21546 : AOI21_X1 port map( B1 => n6079, B2 => n18008, A => n18007, ZN => 
                           n18009);
   U21547 : XNOR2_X1 port map( A => n18735, B => n18762, ZN => n19548);
   U21548 : NAND2_X1 port map( A1 => n18011, A2 => n18306, ZN => n18013);
   U21551 : XNOR2_X1 port map( A => n18802, B => n19198, ZN => n19723);
   U21552 : XNOR2_X1 port map( A => n19723, B => n19548, ZN => n18025);
   U21553 : OAI21_X1 port map( B1 => n18018, B2 => n18017, A => n17771, ZN => 
                           n18022);
   U21555 : XNOR2_X1 port map( A => n19440, B => n3414, ZN => n18023);
   U21556 : XNOR2_X1 port map( A => n19473, B => n18023, ZN => n18024);
   U21557 : XNOR2_X2 port map( A => n18024, B => n18025, ZN => n20302);
   U21558 : INV_X1 port map( A => n20199, ZN => n20202);
   U21559 : XNOR2_X1 port map( A => n19273, B => n3493, ZN => n18031);
   U21560 : AOI21_X1 port map( B1 => n18413, B2 => n18027, A => n18122, ZN => 
                           n18030);
   U21561 : NAND2_X1 port map( A1 => n18028, A2 => n18122, ZN => n18029);
   U21562 : XNOR2_X1 port map( A => n19215, B => n18981, ZN => n18966);
   U21563 : XNOR2_X1 port map( A => n18966, B => n18031, ZN => n18051);
   U21564 : AND2_X1 port map( A1 => n18032, A2 => n18160, ZN => n18039);
   U21566 : INV_X1 port map( A => n18164, ZN => n18038);
   U21567 : NAND2_X1 port map( A1 => n18036, A2 => n18035, ZN => n18037);
   U21568 : OAI21_X1 port map( B1 => n18039, B2 => n18038, A => n18037, ZN => 
                           n18633);
   U21569 : XNOR2_X1 port map( A => n18633, B => n19305, ZN => n18824);
   U21570 : NOR2_X1 port map( A1 => n4805, A2 => n29507, ZN => n18043);
   U21571 : INV_X1 port map( A => n18430, ZN => n18432);
   U21572 : INV_X1 port map( A => n18146, ZN => n18046);
   U21573 : NAND2_X1 port map( A1 => n18046, A2 => n18431, ZN => n18048);
   U21574 : NAND2_X1 port map( A1 => n1758, A2 => n3467, ZN => n18047);
   U21576 : XNOR2_X1 port map( A => n19421, B => n19389, ZN => n18622);
   U21577 : XNOR2_X1 port map( A => n18622, B => n18824, ZN => n18050);
   U21578 : XNOR2_X1 port map( A => n18050, B => n18051, ZN => n20201);
   U21579 : NOR2_X1 port map( A1 => n18260, A2 => n18536, ZN => n18052);
   U21580 : MUX2_X1 port map( A => n18054, B => n18052, S => n18539, Z => 
                           n18056);
   U21581 : OAI21_X1 port map( B1 => n18535, B2 => n18537, A => n18536, ZN => 
                           n18053);
   U21582 : NOR2_X2 port map( A1 => n18056, A2 => n18055, ZN => n19229);
   U21583 : AOI21_X1 port map( B1 => n18059, B2 => n1861, A => n18063, ZN => 
                           n18058);
   U21584 : INV_X1 port map( A => n18058, ZN => n18068);
   U21585 : NOR2_X1 port map( A1 => n29561, A2 => n18059, ZN => n18067);
   U21586 : INV_X1 port map( A => n18061, ZN => n18062);
   U21587 : NAND3_X1 port map( A1 => n18063, A2 => n18298, A3 => n18062, ZN => 
                           n18066);
   U21588 : NAND2_X1 port map( A1 => n18067, A2 => n18064, ZN => n18065);
   U21589 : NAND3_X1 port map( A1 => n18071, A2 => n18070, A3 => n18069, ZN => 
                           n18072);
   U21590 : XNOR2_X1 port map( A => n19448, B => n18725, ZN => n19519);
   U21592 : XNOR2_X1 port map( A => n19717, B => n18085, ZN => n18791);
   U21593 : XNOR2_X1 port map( A => n18791, B => n19519, ZN => n18086);
   U21594 : XNOR2_X1 port map( A => n19452, B => n19278, ZN => n18099);
   U21595 : INV_X1 port map( A => n18090, ZN => n18095);
   U21596 : INV_X1 port map( A => n18091, ZN => n18092);
   U21597 : NAND2_X1 port map( A1 => n18093, A2 => n18092, ZN => n18094);
   U21598 : NOR3_X1 port map( A1 => n18096, A2 => n18095, A3 => n18094, ZN => 
                           n18097);
   U21599 : XNOR2_X1 port map( A => n18099, B => n19702, ZN => n18105);
   U21600 : NAND2_X1 port map( A1 => n18100, A2 => n18452, ZN => n18104);
   U21601 : XNOR2_X1 port map( A => n19194, B => n19004, ZN => n19541);
   U21602 : XNOR2_X1 port map( A => n18105, B => n19541, ZN => n18116);
   U21603 : MUX2_X1 port map( A => n18107, B => n18111, S => n18106, Z => 
                           n18108);
   U21604 : NAND2_X1 port map( A1 => n18108, A2 => n18456, ZN => n18112);
   U21605 : NAND2_X1 port map( A1 => n18111, A2 => n18109, ZN => n18110);
   U21606 : XNOR2_X1 port map( A => n19700, B => n2960, ZN => n18113);
   U21607 : XNOR2_X1 port map( A => n18114, B => n18113, ZN => n18115);
   U21608 : MUX2_X1 port map( A => n18118, B => n18117, S => n19947, Z => 
                           n18119);
   U21609 : AND3_X1 port map( A1 => n18410, A2 => n18122, A3 => n18121, ZN => 
                           n18123);
   U21611 : NOR3_X1 port map( A1 => n18129, A2 => n18588, A3 => n18128, ZN => 
                           n18132);
   U21612 : NOR2_X1 port map( A1 => n18591, A2 => n18130, ZN => n18131);
   U21613 : NOR3_X1 port map( A1 => n18133, A2 => n18132, A3 => n18131, ZN => 
                           n18134);
   U21614 : NAND3_X1 port map( A1 => n18137, A2 => n18136, A3 => n3264, ZN => 
                           n18139);
   U21615 : XNOR2_X1 port map( A => n18852, B => n3317, ZN => n18145);
   U21616 : AND3_X1 port map( A1 => n18147, A2 => n18148, A3 => n18146, ZN => 
                           n18152);
   U21617 : NOR2_X1 port map( A1 => n18431, A2 => n18430, ZN => n18150);
   U21618 : XNOR2_X1 port map( A => n19555, B => n19376, ZN => n18165);
   U21619 : OAI21_X1 port map( B1 => n18155, B2 => n18154, A => n18153, ZN => 
                           n18163);
   U21620 : NAND2_X1 port map( A1 => n18157, A2 => n18156, ZN => n18162);
   U21622 : XNOR2_X1 port map( A => n28530, B => n19678, ZN => n19125);
   U21623 : XNOR2_X1 port map( A => n19125, B => n18165, ZN => n18166);
   U21624 : NAND2_X1 port map( A1 => n4884, A2 => n18168, ZN => n18169);
   U21625 : NAND2_X1 port map( A1 => n18171, A2 => n18170, ZN => n18175);
   U21626 : NAND3_X1 port map( A1 => n513, A2 => n18179, A3 => n18180, ZN => 
                           n18184);
   U21627 : NOR2_X1 port map( A1 => n18181, A2 => n18180, ZN => n18182);
   U21628 : NAND2_X1 port map( A1 => n18182, A2 => n17793, ZN => n18183);
   U21629 : XNOR2_X1 port map( A => n18880, B => n19397, ZN => n19065);
   U21631 : NAND2_X1 port map( A1 => n18190, A2 => n18189, ZN => n18191);
   U21633 : XNOR2_X1 port map( A => n19141, B => n19065, ZN => n18212);
   U21635 : MUX2_X1 port map( A => n18449, B => n18195, S => n18194, Z => 
                           n18196);
   U21636 : INV_X1 port map( A => n18196, ZN => n18202);
   U21637 : NOR2_X1 port map( A1 => n18451, A2 => n18197, ZN => n18201);
   U21638 : NAND2_X1 port map( A1 => n18199, A2 => n18198, ZN => n18200);
   U21639 : MUX2_X1 port map( A => n18203, B => n18277, S => n18204, Z => 
                           n18205);
   U21640 : AND2_X1 port map( A1 => n18275, A2 => n18204, ZN => n18278);
   U21641 : AOI22_X1 port map( A1 => n18205, A2 => n16898, B1 => n18278, B2 => 
                           n18279, ZN => n18208);
   U21642 : NAND2_X1 port map( A1 => n18206, A2 => n18276, ZN => n18207);
   U21644 : XNOR2_X1 port map( A => n19617, B => n3336, ZN => n18209);
   U21645 : XNOR2_X1 port map( A => n18210, B => n18209, ZN => n18211);
   U21646 : XNOR2_X1 port map( A => n18212, B => n18211, ZN => n20544);
   U21647 : NOR3_X1 port map( A1 => n18223, A2 => n18222, A3 => n18221, ZN => 
                           n18225);
   U21648 : NAND3_X1 port map( A1 => n18226, A2 => n18225, A3 => n18224, ZN => 
                           n18228);
   U21649 : AOI21_X1 port map( B1 => n18229, B2 => n18228, A => n18227, ZN => 
                           n18230);
   U21650 : XNOR2_X1 port map( A => n19024, B => n18877, ZN => n18583);
   U21652 : OAI21_X1 port map( B1 => n18242, B2 => n18236, A => n18243, ZN => 
                           n18237);
   U21653 : AOI21_X1 port map( B1 => n18238, B2 => n18242, A => n18237, ZN => 
                           n18246);
   U21654 : NOR2_X1 port map( A1 => n18240, A2 => n18239, ZN => n18245);
   U21655 : NOR3_X1 port map( A1 => n18243, A2 => n18242, A3 => n18241, ZN => 
                           n18244);
   U21656 : NOR3_X1 port map( A1 => n18246, A2 => n18245, A3 => n18244, ZN => 
                           n18247);
   U21657 : XNOR2_X1 port map( A => n18667, B => n18247, ZN => n19130);
   U21658 : XNOR2_X1 port map( A => n19130, B => n18583, ZN => n18258);
   U21659 : XNOR2_X1 port map( A => n19402, B => n18256, ZN => n18257);
   U21660 : MUX2_X1 port map( A => n19820, B => n20544, S => n20547, Z => 
                           n18365);
   U21661 : XNOR2_X1 port map( A => n19525, B => n1193, ZN => n18269);
   U21662 : INV_X1 port map( A => n18326, ZN => n18330);
   U21663 : NAND2_X1 port map( A1 => n18330, A2 => n18261, ZN => n18267);
   U21664 : OAI21_X1 port map( B1 => n18326, B2 => n18324, A => n18263, ZN => 
                           n18264);
   U21665 : NAND2_X1 port map( A1 => n18265, A2 => n18264, ZN => n18266);
   U21666 : OAI21_X1 port map( B1 => n18268, B2 => n18267, A => n18266, ZN => 
                           n18975);
   U21667 : XNOR2_X1 port map( A => n18975, B => n19511, ZN => n19410);
   U21668 : XNOR2_X1 port map( A => n19410, B => n18269, ZN => n18290);
   U21669 : INV_X1 port map( A => n18510, ZN => n18271);
   U21670 : NAND3_X1 port map( A1 => n18276, A2 => n18279, A3 => n18275, ZN => 
                           n18284);
   U21671 : INV_X1 port map( A => n18276, ZN => n18280);
   U21672 : NAND3_X1 port map( A1 => n3995, A2 => n18280, A3 => n18277, ZN => 
                           n18283);
   U21673 : INV_X1 port map( A => n18278, ZN => n18282);
   U21674 : NAND3_X1 port map( A1 => n18280, A2 => n16898, A3 => n18279, ZN => 
                           n18281);
   U21675 : NAND4_X1 port map( A1 => n18284, A2 => n18283, A3 => n18282, A4 => 
                           n18281, ZN => n18857);
   U21676 : XNOR2_X1 port map( A => n18857, B => n19320, ZN => n18578);
   U21677 : XNOR2_X1 port map( A => n19695, B => n19622, ZN => n19116);
   U21678 : XNOR2_X1 port map( A => n19116, B => n18578, ZN => n18289);
   U21679 : XNOR2_X1 port map( A => n18290, B => n18289, ZN => n20388);
   U21680 : AND2_X1 port map( A1 => n18291, A2 => n28633, ZN => n18296);
   U21681 : NAND2_X1 port map( A1 => n18292, A2 => n28633, ZN => n18294);
   U21682 : NAND2_X1 port map( A1 => n18294, A2 => n18293, ZN => n18295);
   U21683 : NAND2_X1 port map( A1 => n18301, A2 => n18300, ZN => n18302);
   U21684 : XNOR2_X1 port map( A => n19631, B => n19482, ZN => n19391);
   U21685 : NAND3_X1 port map( A1 => n18306, A2 => n17679, A3 => n18305, ZN => 
                           n18307);
   U21686 : OAI21_X1 port map( B1 => n18011, B2 => n17679, A => n18307, ZN => 
                           n18308);
   U21687 : XNOR2_X1 port map( A => n18868, B => n19391, ZN => n18321);
   U21688 : AOI21_X1 port map( B1 => n18471, B2 => n18466, A => n18467, ZN => 
                           n18313);
   U21690 : NAND2_X1 port map( A1 => n18465, A2 => n18315, ZN => n18316);
   U21691 : OAI21_X2 port map( B1 => n18318, B2 => n18317, A => n18316, ZN => 
                           n19306);
   U21692 : XNOR2_X1 port map( A => n19087, B => n19306, ZN => n18620);
   U21693 : XNOR2_X1 port map( A => n19534, B => n1911, ZN => n18319);
   U21694 : XNOR2_X1 port map( A => n18620, B => n18319, ZN => n18320);
   U21695 : MUX2_X1 port map( A => n20388, B => n20539, S => n19820, Z => 
                           n18364);
   U21696 : NAND2_X1 port map( A1 => n18323, A2 => n18322, ZN => n18328);
   U21697 : NOR2_X1 port map( A1 => n29603, A2 => n18324, ZN => n18327);
   U21698 : XNOR2_X1 port map( A => n19359, B => n19726, ZN => n18862);
   U21699 : OAI21_X1 port map( B1 => n18337, B2 => n18332, A => n18331, ZN => 
                           n18339);
   U21701 : XNOR2_X1 port map( A => n19384, B => n18680, ZN => n19071);
   U21702 : XNOR2_X1 port map( A => n18862, B => n19071, ZN => n18363);
   U21703 : AOI21_X1 port map( B1 => n18349, B2 => n18348, A => n18380, ZN => 
                           n18352);
   U21704 : NAND2_X1 port map( A1 => n18382, A2 => n18376, ZN => n18351);
   U21705 : NOR2_X1 port map( A1 => n18355, A2 => n18353, ZN => n18360);
   U21706 : OAI21_X1 port map( B1 => n18355, B2 => n18354, A => n18356, ZN => 
                           n18359);
   U21707 : XNOR2_X1 port map( A => n18798, B => n18900, ZN => n19472);
   U21708 : XNOR2_X1 port map( A => n19549, B => n25992, ZN => n18361);
   U21709 : XNOR2_X1 port map( A => n19472, B => n18361, ZN => n18362);
   U21710 : MUX2_X1 port map( A => n18365, B => n18364, S => n20546, Z => 
                           n21346);
   U21711 : MUX2_X1 port map( A => n6314, B => n21692, S => n21346, Z => n18548
                           );
   U21712 : XNOR2_X1 port map( A => n19277, B => n18638, ZN => n18766);
   U21713 : MUX2_X2 port map( A => n18374, B => n18373, S => n18372, Z => 
                           n19191);
   U21714 : XNOR2_X1 port map( A => n19700, B => n19191, ZN => n18375);
   U21715 : XNOR2_X1 port map( A => n18766, B => n18375, ZN => n18386);
   U21716 : AND2_X1 port map( A1 => n18376, A2 => n18379, ZN => n18377);
   U21717 : NOR2_X1 port map( A1 => n18380, A2 => n18379, ZN => n18381);
   U21718 : XNOR2_X1 port map( A => n29505, B => n26032, ZN => n18384);
   U21719 : XNOR2_X1 port map( A => n19356, B => n18384, ZN => n18385);
   U21721 : AOI22_X1 port map( A1 => n29024, A2 => n18388, B1 => n17592, B2 => 
                           n18387, ZN => n18394);
   U21724 : XNOR2_X1 port map( A => n18863, B => n18395, ZN => n18987);
   U21725 : OAI21_X1 port map( B1 => n18707, B2 => n18706, A => n4757, ZN => 
                           n18407);
   U21726 : XNOR2_X1 port map( A => n28798, B => n18948, ZN => n18409);
   U21727 : NAND2_X1 port map( A1 => n20290, A2 => n20295, ZN => n20128);
   U21728 : INV_X1 port map( A => n18410, ZN => n18412);
   U21729 : MUX2_X1 port map( A => n18413, B => n18412, S => n18411, Z => 
                           n18419);
   U21730 : NAND3_X1 port map( A1 => n18410, A2 => n417, A3 => n18414, ZN => 
                           n18415);
   U21731 : XNOR2_X1 port map( A => n19409, B => n19332, ZN => n18420);
   U21732 : XNOR2_X1 port map( A => n19330, B => n18420, ZN => n18440);
   U21733 : NAND2_X1 port map( A1 => n29507, A2 => n18421, ZN => n18424);
   U21734 : AOI21_X1 port map( B1 => n1942, B2 => n18424, A => n18423, ZN => 
                           n18428);
   U21735 : XNOR2_X1 port map( A => n19697, B => n19592, ZN => n18438);
   U21736 : XNOR2_X1 port map( A => n19207, B => n3211, ZN => n18437);
   U21737 : XNOR2_X1 port map( A => n18438, B => n18437, ZN => n18439);
   U21738 : XNOR2_X1 port map( A => n18440, B => n18439, ZN => n20125);
   U21739 : NAND2_X1 port map( A1 => n18441, A2 => n523, ZN => n18447);
   U21740 : INV_X1 port map( A => n18442, ZN => n18443);
   U21741 : OAI21_X1 port map( B1 => n18445, B2 => n18444, A => n18443, ZN => 
                           n18446);
   U21742 : XNOR2_X1 port map( A => n19686, B => n19219, ZN => n18967);
   U21743 : NAND3_X1 port map( A1 => n18452, A2 => n6663, A3 => n18451, ZN => 
                           n18453);
   U21744 : XNOR2_X1 port map( A => n19338, B => n18967, ZN => n18462);
   U21745 : XNOR2_X1 port map( A => n19595, B => n19339, ZN => n18774);
   U21746 : XNOR2_X1 port map( A => n19389, B => n3633, ZN => n18460);
   U21747 : XNOR2_X1 port map( A => n18774, B => n18460, ZN => n18461);
   U21748 : XNOR2_X1 port map( A => n18462, B => n18461, ZN => n19815);
   U21749 : NAND2_X1 port map( A1 => n20125, A2 => n19815, ZN => n18463);
   U21750 : NAND2_X1 port map( A1 => n20128, A2 => n18463, ZN => n18547);
   U21751 : NOR2_X1 port map( A1 => n18465, A2 => n18464, ZN => n18470);
   U21752 : NOR2_X1 port map( A1 => n18467, A2 => n18466, ZN => n18468);
   U21753 : NOR2_X1 port map( A1 => n18472, A2 => n18471, ZN => n18473);
   U21754 : XNOR2_X1 port map( A => n19225, B => n19136, ZN => n18991);
   U21755 : AOI21_X1 port map( B1 => n18474, B2 => n18479, A => n18477, ZN => 
                           n18485);
   U21756 : AOI21_X1 port map( B1 => n18478, B2 => n18475, A => n18011, ZN => 
                           n18484);
   U21757 : NOR3_X1 port map( A1 => n18477, A2 => n18479, A3 => n18476, ZN => 
                           n18482);
   U21758 : NOR3_X1 port map( A1 => n18480, A2 => n18479, A3 => n18478, ZN => 
                           n18481);
   U21759 : NOR2_X1 port map( A1 => n18482, A2 => n18481, ZN => n18483);
   U21760 : OAI21_X1 port map( B1 => n18485, B2 => n18484, A => n18483, ZN => 
                           n19611);
   U21761 : XNOR2_X1 port map( A => n19611, B => n19245, ZN => n18779);
   U21762 : INV_X1 port map( A => n18488, ZN => n18491);
   U21763 : XNOR2_X1 port map( A => n19228, B => n2522, ZN => n18497);
   U21764 : XNOR2_X1 port map( A => n19717, B => n18935, ZN => n18496);
   U21765 : XNOR2_X1 port map( A => n18497, B => n18496, ZN => n18498);
   U21766 : XNOR2_X1 port map( A => n18499, B => n18498, ZN => n20123);
   U21767 : NOR2_X1 port map( A1 => n18500, A2 => n2363, ZN => n18501);
   U21768 : AND2_X1 port map( A1 => n18503, A2 => n18506, ZN => n18504);
   U21771 : XNOR2_X1 port map( A => n18517, B => n18652, ZN => n19333);
   U21772 : XNOR2_X1 port map( A => n18942, B => n3116, ZN => n18518);
   U21773 : XNOR2_X1 port map( A => n18518, B => n18812, ZN => n18519);
   U21774 : XNOR2_X1 port map( A => n19333, B => n18519, ZN => n18545);
   U21775 : XNOR2_X1 port map( A => n19262, B => n19577, ZN => n18755);
   U21776 : NOR2_X1 port map( A1 => n18528, A2 => n18527, ZN => n18534);
   U21779 : MUX2_X1 port map( A => n18534, B => n29327, S => n509, Z => n18543)
                           ;
   U21780 : NOR2_X1 port map( A1 => n18538, A2 => n18537, ZN => n18540);
   U21781 : XNOR2_X1 port map( A => n28144, B => n18755, ZN => n18544);
   U21782 : XNOR2_X1 port map( A => n18544, B => n18545, ZN => n20293);
   U21783 : INV_X1 port map( A => n20290, ZN => n19967);
   U21785 : INV_X1 port map( A => n19370, ZN => n18550);
   U21786 : XNOR2_X1 port map( A => n19123, B => n18550, ZN => n18894);
   U21787 : XNOR2_X1 port map( A => n19122, B => n19376, ZN => n18551);
   U21788 : XNOR2_X1 port map( A => n18894, B => n18551, ZN => n18555);
   U21789 : XNOR2_X1 port map( A => n19636, B => n19232, ZN => n18553);
   U21790 : XNOR2_X1 port map( A => n19468, B => n24897, ZN => n18552);
   U21791 : XNOR2_X1 port map( A => n18552, B => n18553, ZN => n18554);
   U21792 : XNOR2_X1 port map( A => n19346, B => n19397, ZN => n19666);
   U21793 : XNOR2_X1 port map( A => n18556, B => n19666, ZN => n18560);
   U21794 : XNOR2_X1 port map( A => n19487, B => n29554, ZN => n18558);
   U21795 : XNOR2_X1 port map( A => n19136, B => n857, ZN => n18557);
   U21796 : XNOR2_X1 port map( A => n18558, B => n18557, ZN => n18559);
   U21798 : INV_X1 port map( A => n19194, ZN => n18744);
   U21799 : XNOR2_X1 port map( A => n18744, B => n2598, ZN => n18561);
   U21800 : XNOR2_X1 port map( A => n19402, B => n18561, ZN => n18564);
   U21801 : XNOR2_X1 port map( A => n19495, B => n19655, ZN => n18562);
   U21802 : XNOR2_X1 port map( A => n18562, B => n19133, ZN => n18563);
   U21804 : XNOR2_X1 port map( A => n18695, B => n18856, ZN => n19117);
   U21805 : XNOR2_X1 port map( A => n19410, B => n19117, ZN => n18568);
   U21806 : XNOR2_X1 port map( A => n19507, B => n18960, ZN => n18566);
   U21807 : XNOR2_X1 port map( A => n19622, B => n22489, ZN => n18565);
   U21808 : XNOR2_X1 port map( A => n18566, B => n18565, ZN => n18567);
   U21809 : NOR2_X1 port map( A1 => n29315, A2 => n20077, ZN => n18573);
   U21810 : INV_X1 port map( A => n19384, ZN => n19291);
   U21811 : XNOR2_X1 port map( A => n19291, B => n19474, ZN => n18989);
   U21812 : XNOR2_X1 port map( A => n18989, B => n19359, ZN => n19649);
   U21813 : XNOR2_X1 port map( A => n18569, B => n18395, ZN => n18571);
   U21814 : XNOR2_X1 port map( A => n19162, B => n19256, ZN => n18570);
   U21815 : XNOR2_X1 port map( A => n18571, B => n18570, ZN => n18572);
   U21816 : XNOR2_X1 port map( A => n19691, B => n18628, ZN => n18576);
   U21818 : XNOR2_X1 port map( A => n18578, B => n18577, ZN => n18579);
   U21820 : BUF_X2 port map( A => n18834, Z => n20381);
   U21821 : XNOR2_X1 port map( A => n18581, B => n19702, ZN => n18582);
   U21822 : XNOR2_X1 port map( A => n18582, B => n18583, ZN => n18586);
   U21823 : XNOR2_X1 port map( A => n19700, B => n3114, ZN => n18584);
   U21824 : INV_X1 port map( A => n19004, ZN => n18769);
   U21825 : XNOR2_X1 port map( A => n18769, B => n18584, ZN => n18585);
   U21827 : XNOR2_X1 port map( A => n18852, B => n2465, ZN => n18587);
   U21828 : XNOR2_X1 port map( A => n18587, B => n19378, ZN => n18597);
   U21829 : XNOR2_X1 port map( A => n19428, B => n19300, ZN => n18754);
   U21830 : XNOR2_X1 port map( A => n18597, B => n18754, ZN => n18609);
   U21831 : OR2_X1 port map( A1 => n6927, A2 => n18598, ZN => n18606);
   U21832 : MUX2_X1 port map( A => n28142, B => n18600, S => n18599, Z => 
                           n18602);
   U21833 : NAND2_X1 port map( A1 => n18602, A2 => n6927, ZN => n18605);
   U21834 : AOI21_X1 port map( B1 => n18606, B2 => n18605, A => n18604, ZN => 
                           n18607);
   U21835 : XNOR2_X1 port map( A => n18607, B => n19427, ZN => n18608);
   U21836 : INV_X1 port map( A => n20573, ZN => n19837);
   U21837 : XNOR2_X1 port map( A => n19198, B => n18762, ZN => n19439);
   U21838 : XNOR2_X1 port map( A => n19039, B => n19439, ZN => n18612);
   U21839 : XNOR2_X1 port map( A => n18680, B => n26825, ZN => n18610);
   U21840 : XNOR2_X1 port map( A => n19727, B => n18798, ZN => n19289);
   U21841 : XNOR2_X1 port map( A => n18610, B => n19289, ZN => n18611);
   U21842 : XNOR2_X1 port map( A => n18612, B => n18611, ZN => n18613);
   U21843 : INV_X1 port map( A => n18613, ZN => n19838);
   U21844 : AOI21_X1 port map( B1 => n28637, B2 => n19837, A => n19833, ZN => 
                           n18627);
   U21846 : XNOR2_X1 port map( A => n18928, B => n19229, ZN => n19715);
   U21847 : XNOR2_X1 port map( A => n19399, B => n19715, ZN => n18617);
   U21848 : INV_X1 port map( A => n19491, ZN => n19313);
   U21849 : XNOR2_X1 port map( A => n6489, B => n18880, ZN => n18615);
   U21850 : XNOR2_X1 port map( A => n19448, B => n3035, ZN => n18614);
   U21851 : XNOR2_X1 port map( A => n18615, B => n18614, ZN => n18616);
   U21852 : NAND2_X1 port map( A1 => n29143, A2 => n20568, ZN => n18625);
   U21853 : XNOR2_X1 port map( A => n18981, B => n3722, ZN => n18619);
   U21854 : INV_X1 port map( A => n19045, ZN => n18618);
   U21855 : XNOR2_X1 port map( A => n18619, B => n18618, ZN => n18621);
   U21856 : XNOR2_X1 port map( A => n18621, B => n18620, ZN => n18623);
   U21857 : XNOR2_X1 port map( A => n18622, B => n19535, ZN => n19690);
   U21858 : MUX2_X1 port map( A => n18625, B => n18624, S => n28637, Z => 
                           n18626);
   U21859 : XNOR2_X1 port map( A => n19321, B => n18628, ZN => n18629);
   U21860 : XNOR2_X1 port map( A => n19206, B => n19692, ZN => n18730);
   U21861 : XNOR2_X1 port map( A => n18629, B => n18730, ZN => n18632);
   U21862 : XNOR2_X1 port map( A => n19592, B => n3164, ZN => n18630);
   U21863 : XNOR2_X1 port map( A => n19528, B => n18630, ZN => n18631);
   U21864 : XNOR2_X1 port map( A => n19045, B => n19595, ZN => n18634);
   U21865 : INV_X1 port map( A => n18633, ZN => n19423);
   U21866 : XNOR2_X1 port map( A => n19423, B => n19219, ZN => n19532);
   U21867 : XNOR2_X1 port map( A => n19532, B => n18634, ZN => n18637);
   U21868 : XNOR2_X1 port map( A => n19220, B => n19687, ZN => n18720);
   U21869 : XNOR2_X1 port map( A => n19305, B => n3554, ZN => n18635);
   U21870 : XNOR2_X1 port map( A => n18720, B => n18635, ZN => n18636);
   U21871 : XNOR2_X1 port map( A => n18637, B => n18636, ZN => n19849);
   U21872 : NOR2_X1 port map( A1 => n20401, A2 => n29041, ZN => n18650);
   U21873 : INV_X1 port map( A => n18114, ZN => n19166);
   U21874 : XNOR2_X1 port map( A => n19166, B => n18638, ZN => n18639);
   U21875 : XNOR2_X1 port map( A => n19192, B => n19704, ZN => n18743);
   U21876 : XNOR2_X1 port map( A => n18743, B => n18640, ZN => n18641);
   U21877 : XNOR2_X1 port map( A => n18760, B => n18863, ZN => n18643);
   U21878 : XNOR2_X1 port map( A => n19643, B => n27462, ZN => n18642);
   U21879 : XNOR2_X1 port map( A => n18643, B => n18642, ZN => n18645);
   U21880 : XNOR2_X1 port map( A => n18948, B => n19440, ZN => n19546);
   U21881 : XNOR2_X1 port map( A => n19290, B => n19546, ZN => n18644);
   U21882 : XNOR2_X1 port map( A => n18644, B => n18645, ZN => n19851);
   U21883 : NOR2_X1 port map( A1 => n20209, A2 => n19851, ZN => n20559);
   U21884 : XNOR2_X1 port map( A => n18646, B => n3374, ZN => n18647);
   U21885 : XNOR2_X1 port map( A => n19225, B => n18647, ZN => n18648);
   U21886 : XNOR2_X1 port map( A => n19518, B => n18648, ZN => n18649);
   U21887 : XNOR2_X1 port map( A => n19611, B => n19490, ZN => n19317);
   U21888 : XNOR2_X1 port map( A => n18778, B => n19317, ZN => n19183);
   U21890 : XNOR2_X1 port map( A => n19577, B => n19465, ZN => n19296);
   U21891 : XNOR2_X1 port map( A => n28144, B => n19378, ZN => n18651);
   U21892 : XNOR2_X1 port map( A => n19296, B => n18651, ZN => n18657);
   U21893 : INV_X1 port map( A => n18652, ZN => n19235);
   U21894 : XNOR2_X1 port map( A => n19568, B => n19235, ZN => n18655);
   U21895 : XNOR2_X1 port map( A => n29492, B => n3607, ZN => n18654);
   U21896 : XNOR2_X1 port map( A => n18655, B => n18654, ZN => n18656);
   U21897 : XNOR2_X1 port map( A => n18656, B => n18657, ZN => n20208);
   U21898 : NOR2_X1 port map( A1 => n20208, A2 => n29041, ZN => n20398);
   U21899 : OAI21_X1 port map( B1 => n20398, B2 => n20401, A => n20209, ZN => 
                           n18658);
   U21901 : NAND2_X1 port map( A1 => n29315, A2 => n29551, ZN => n20075);
   U21902 : INV_X1 port map( A => n19391, ZN => n18661);
   U21903 : XNOR2_X1 port map( A => n19215, B => n19108, ZN => n18660);
   U21904 : XNOR2_X1 port map( A => n18661, B => n18660, ZN => n18665);
   U21905 : XNOR2_X1 port map( A => n19111, B => n19483, ZN => n18663);
   U21906 : XNOR2_X1 port map( A => n18663, B => n18662, ZN => n18664);
   U21907 : XNOR2_X1 port map( A => n18665, B => n18664, ZN => n18838);
   U21908 : NOR2_X1 port map( A1 => n20075, A2 => n18838, ZN => n18753);
   U21909 : INV_X1 port map( A => n18753, ZN => n19914);
   U21911 : XNOR2_X1 port map( A => n19285, B => n18666, ZN => n18669);
   U21912 : XNOR2_X1 port map( A => n18912, B => n18877, ZN => n19102);
   U21913 : INV_X1 port map( A => n18667, ZN => n19709);
   U21914 : XNOR2_X1 port map( A => n19709, B => n19278, ZN => n19502);
   U21915 : XNOR2_X1 port map( A => n19102, B => n19502, ZN => n18668);
   U21916 : XNOR2_X1 port map( A => n18668, B => n18669, ZN => n18843);
   U21917 : INV_X1 port map( A => n18843, ZN => n20372);
   U21918 : XNOR2_X1 port map( A => n19688, B => n19273, ZN => n19480);
   U21919 : XNOR2_X1 port map( A => n19480, B => n18670, ZN => n18674);
   U21920 : XNOR2_X1 port map( A => n18906, B => n19087, ZN => n18672);
   U21922 : XNOR2_X1 port map( A => n18672, B => n18671, ZN => n18673);
   U21924 : INV_X1 port map( A => n20374, ZN => n19739);
   U21925 : XNOR2_X1 port map( A => n29580, B => n19679, ZN => n19298);
   U21926 : XNOR2_X1 port map( A => n18852, B => n19377, ZN => n19078);
   U21927 : XNOR2_X1 port map( A => n19298, B => n19078, ZN => n18679);
   U21928 : XNOR2_X1 port map( A => n19122, B => n19462, ZN => n18677);
   U21929 : INV_X1 port map( A => n1247, ZN => n26701);
   U21930 : XNOR2_X1 port map( A => n19464, B => n26701, ZN => n18676);
   U21931 : XNOR2_X1 port map( A => n18677, B => n18676, ZN => n18678);
   U21932 : NOR3_X1 port map( A1 => n20372, A2 => n19739, A3 => n20375, ZN => 
                           n18688);
   U21933 : INV_X1 port map( A => n18680, ZN => n19250);
   U21934 : XNOR2_X1 port map( A => n19250, B => n18395, ZN => n18682);
   U21935 : XNOR2_X1 port map( A => n18681, B => n18682, ZN => n18686);
   U21936 : XNOR2_X1 port map( A => n19251, B => n19726, ZN => n18684);
   U21937 : XNOR2_X1 port map( A => n18899, B => n2385, ZN => n18683);
   U21938 : XNOR2_X1 port map( A => n18684, B => n18683, ZN => n18685);
   U21939 : NOR2_X1 port map( A1 => n20071, A2 => n20374, ZN => n18687);
   U21940 : XNOR2_X1 port map( A => n19136, B => n1225, ZN => n18689);
   U21941 : INV_X1 port map( A => n19486, ZN => n19716);
   U21942 : XNOR2_X1 port map( A => n19716, B => n18927, ZN => n18692);
   U21943 : XNOR2_X1 port map( A => n18692, B => n18691, ZN => n18693);
   U21944 : NAND2_X1 port map( A1 => n20373, A2 => n18699, ZN => n18701);
   U21945 : XNOR2_X1 port map( A => n19267, B => n19695, ZN => n19513);
   U21946 : XNOR2_X1 port map( A => n19322, B => n19513, ZN => n18698);
   U21947 : XNOR2_X1 port map( A => n18695, B => n3660, ZN => n18696);
   U21948 : XNOR2_X1 port map( A => n18696, B => n19097, ZN => n18697);
   U21949 : XNOR2_X1 port map( A => n18698, B => n18697, ZN => n19841);
   U21950 : INV_X1 port map( A => n18699, ZN => n19740);
   U21951 : NAND3_X1 port map( A1 => n19841, A2 => n351, A3 => n19740, ZN => 
                           n18700);
   U21952 : OAI21_X1 port map( B1 => n18843, B2 => n18701, A => n18700, ZN => 
                           n18702);
   U21953 : NOR2_X2 port map( A1 => n18703, A2 => n18702, ZN => n20972);
   U21954 : INV_X1 port map( A => n20972, ZN => n21216);
   U21955 : XNOR2_X1 port map( A => n18704, B => n19637, ZN => n18705);
   U21956 : XNOR2_X1 port map( A => n18705, B => n19574, ZN => n18717);
   U21957 : MUX2_X1 port map( A => n28558, B => n18707, S => n18706, Z => 
                           n18711);
   U21958 : INV_X1 port map( A => n18712, ZN => n18713);
   U21959 : XNOR2_X1 port map( A => n19235, B => n19232, ZN => n18715);
   U21960 : XNOR2_X1 port map( A => n19075, B => n18715, ZN => n18716);
   U21961 : XNOR2_X1 port map( A => n19215, B => n3565, ZN => n18719);
   U21962 : XNOR2_X1 port map( A => n19632, B => n19085, ZN => n18718);
   U21963 : XNOR2_X1 port map( A => n18719, B => n18718, ZN => n18721);
   U21964 : INV_X1 port map( A => n18749, ZN => n18751);
   U21965 : XNOR2_X1 port map( A => n19243, B => n3212, ZN => n18724);
   U21966 : INV_X1 port map( A => n18722, ZN => n18723);
   U21967 : XNOR2_X1 port map( A => n18724, B => n18723, ZN => n18728);
   U21968 : INV_X1 port map( A => n18725, ZN => n19226);
   U21969 : XNOR2_X1 port map( A => n18726, B => n19226, ZN => n18727);
   U21970 : XNOR2_X1 port map( A => n19525, B => n19626, ZN => n18729);
   U21971 : XNOR2_X1 port map( A => n18729, B => n18730, ZN => n18734);
   U21972 : XNOR2_X1 port map( A => n18960, B => n19408, ZN => n18732);
   U21973 : XNOR2_X1 port map( A => n19096, B => n26680, ZN => n18731);
   U21974 : XNOR2_X1 port map( A => n18732, B => n18731, ZN => n18733);
   U21975 : INV_X1 port map( A => n19582, ZN => n18736);
   U21976 : XNOR2_X1 port map( A => n18735, B => n18863, ZN => n19203);
   U21977 : XNOR2_X1 port map( A => n18736, B => n19203, ZN => n18742);
   U21978 : XNOR2_X1 port map( A => n18760, B => n3369, ZN => n18740);
   U21979 : INV_X1 port map( A => n18738, ZN => n19644);
   U21980 : XNOR2_X1 port map( A => n18737, B => n19644, ZN => n18739);
   U21981 : XNOR2_X1 port map( A => n18740, B => n18739, ZN => n18741);
   U21982 : XNOR2_X1 port map( A => n19607, B => n18743, ZN => n18748);
   U21983 : XNOR2_X1 port map( A => n18744, B => n3036, ZN => n18745);
   U21984 : XNOR2_X1 port map( A => n18745, B => n18746, ZN => n18747);
   U21985 : XNOR2_X1 port map( A => n18755, B => n18754, ZN => n18759);
   U21986 : XNOR2_X1 port map( A => n29318, B => n3787, ZN => n18757);
   U21987 : XNOR2_X1 port map( A => n29492, B => n18942, ZN => n19681);
   U21988 : XNOR2_X1 port map( A => n18757, B => n19681, ZN => n18758);
   U21989 : XNOR2_X1 port map( A => n18759, B => n18758, ZN => n20064);
   U21990 : XNOR2_X1 port map( A => n18761, B => n18760, ZN => n19438);
   U21991 : XNOR2_X1 port map( A => n19585, B => n18798, ZN => n18764);
   U21992 : XNOR2_X1 port map( A => n28798, B => n3191, ZN => n18763);
   U21993 : INV_X1 port map( A => n18766, ZN => n19165);
   U21995 : XNOR2_X1 port map( A => n19165, B => n18768, ZN => n18771);
   U21996 : XNOR2_X1 port map( A => n29506, B => n19704, ZN => n18770);
   U21997 : XNOR2_X1 port map( A => n18770, B => n18769, ZN => n19455);
   U21998 : NOR2_X1 port map( A1 => n20063, A2 => n20049, ZN => n18846);
   U21999 : XNOR2_X1 port map( A => n19306, B => n19686, ZN => n18772);
   U22000 : XNOR2_X1 port map( A => n18981, B => n19687, ZN => n19420);
   U22001 : XNOR2_X1 port map( A => n18772, B => n19420, ZN => n18775);
   U22002 : INV_X1 port map( A => n18773, ZN => n19110);
   U22003 : NOR2_X1 port map( A1 => n20064, A2 => n19761, ZN => n18776);
   U22004 : XNOR2_X1 port map( A => n19448, B => n19615, ZN => n18995);
   U22005 : XNOR2_X1 port map( A => n19313, B => n5633, ZN => n18777);
   U22006 : XNOR2_X1 port map( A => n18777, B => n18995, ZN => n18781);
   U22007 : XNOR2_X1 port map( A => n18778, B => n18935, ZN => n19447);
   U22008 : XNOR2_X1 port map( A => n19447, B => n18779, ZN => n18780);
   U22009 : XNOR2_X1 port map( A => n18781, B => n18780, ZN => n18845);
   U22010 : XNOR2_X1 port map( A => n19320, B => n2350, ZN => n18783);
   U22011 : XNOR2_X1 port map( A => n19697, B => n18959, ZN => n18784);
   U22012 : XNOR2_X1 port map( A => n18784, B => n19692, ZN => n19436);
   U22013 : XNOR2_X1 port map( A => n18785, B => n19436, ZN => n20066);
   U22014 : NAND3_X1 port map( A1 => n21221, A2 => n20972, A3 => n20966, ZN => 
                           n18786);
   U22016 : INV_X1 port map( A => n20089, ZN => n19778);
   U22017 : NOR2_X1 port map( A1 => n18790, A2 => n20039, ZN => n20877);
   U22018 : INV_X1 port map( A => n18791, ZN => n18793);
   U22019 : XNOR2_X1 port map( A => n19349, B => n18937, ZN => n18792);
   U22020 : XNOR2_X1 port map( A => n18793, B => n18792, ZN => n18797);
   U22021 : XNOR2_X1 port map( A => n19491, B => n19228, ZN => n18795);
   U22022 : XNOR2_X1 port map( A => n18927, B => n2541, ZN => n18794);
   U22023 : XNOR2_X1 port map( A => n18795, B => n18794, ZN => n18796);
   U22024 : XNOR2_X1 port map( A => n18798, B => n18799, ZN => n18801);
   U22025 : XNOR2_X1 port map( A => n18899, B => n900, ZN => n18800);
   U22026 : XNOR2_X1 port map( A => n18801, B => n18800, ZN => n18805);
   U22027 : XNOR2_X1 port map( A => n18802, B => n19725, ZN => n18803);
   U22028 : XNOR2_X1 port map( A => n19546, B => n18803, ZN => n18804);
   U22029 : INV_X1 port map( A => n20098, ZN => n20096);
   U22030 : INV_X1 port map( A => n18806, ZN => n19696);
   U22031 : XNOR2_X1 port map( A => n19321, B => n19696, ZN => n18807);
   U22032 : XNOR2_X1 port map( A => n19528, B => n18807, ZN => n18811);
   U22033 : XNOR2_X1 port map( A => n19409, B => n3029, ZN => n18809);
   U22034 : XNOR2_X1 port map( A => n19320, B => n19412, ZN => n18808);
   U22035 : XNOR2_X1 port map( A => n18809, B => n18808, ZN => n18810);
   U22036 : XNOR2_X1 port map( A => n18811, B => n18810, ZN => n20150);
   U22037 : INV_X1 port map( A => n18812, ZN => n19371);
   U22038 : XNOR2_X1 port map( A => n19371, B => n19300, ZN => n18814);
   U22039 : XNOR2_X1 port map( A => n19377, B => n27956, ZN => n18813);
   U22040 : XNOR2_X1 port map( A => n18814, B => n18813, ZN => n18819);
   U22041 : XNOR2_X1 port map( A => n28144, B => n19679, ZN => n18817);
   U22042 : INV_X1 port map( A => n18815, ZN => n18816);
   U22043 : XNOR2_X1 port map( A => n18816, B => n18817, ZN => n18818);
   U22044 : XNOR2_X1 port map( A => n18912, B => n19706, ZN => n18821);
   U22045 : XNOR2_X1 port map( A => n19700, B => n2544, ZN => n18820);
   U22046 : XNOR2_X1 port map( A => n18821, B => n18820, ZN => n18823);
   U22047 : XNOR2_X1 port map( A => n18114, B => n19024, ZN => n19498);
   U22048 : XNOR2_X1 port map( A => n19498, B => n19540, ZN => n18822);
   U22049 : XNOR2_X1 port map( A => n18906, B => n19219, ZN => n18826);
   U22050 : INV_X1 port map( A => n18824, ZN => n18825);
   U22051 : XNOR2_X1 port map( A => n18826, B => n18825, ZN => n18830);
   U22052 : XNOR2_X1 port map( A => n19389, B => n19306, ZN => n18828);
   U22053 : INV_X1 port map( A => n3537, ZN => n27324);
   U22054 : XNOR2_X1 port map( A => n19685, B => n27324, ZN => n18827);
   U22055 : XNOR2_X1 port map( A => n18828, B => n18827, ZN => n18829);
   U22056 : XNOR2_X1 port map( A => n18830, B => n18829, ZN => n18887);
   U22059 : INV_X1 port map( A => n18834, ZN => n20574);
   U22061 : NOR2_X1 port map( A1 => n29145, A2 => n18838, ZN => n18836);
   U22062 : NOR2_X1 port map( A1 => n20077, A2 => n28526, ZN => n18835);
   U22063 : INV_X1 port map( A => n18838, ZN => n20083);
   U22064 : INV_X1 port map( A => n20375, ZN => n20371);
   U22065 : INV_X1 port map( A => n19841, ZN => n20377);
   U22066 : MUX2_X1 port map( A => n19739, B => n20371, S => n20377, Z => 
                           n18844);
   U22067 : INV_X1 port map( A => n20373, ZN => n20074);
   U22068 : NOR2_X1 port map( A1 => n20379, A2 => n20074, ZN => n18841);
   U22069 : NOR2_X1 port map( A1 => n19740, A2 => n19841, ZN => n18840);
   U22070 : AOI22_X1 port map( A1 => n18843, A2 => n18841, B1 => n18840, B2 => 
                           n20371, ZN => n18842);
   U22071 : NOR2_X1 port map( A1 => n21266, A2 => n20816, ZN => n18849);
   U22072 : INV_X1 port map( A => n18845, ZN => n20065);
   U22073 : INV_X1 port map( A => n20066, ZN => n20048);
   U22074 : INV_X1 port map( A => n20063, ZN => n18892);
   U22075 : INV_X1 port map( A => n18846, ZN => n19764);
   U22076 : NOR2_X1 port map( A1 => n21268, A2 => n20875, ZN => n21271);
   U22077 : AOI22_X1 port map( A1 => n21269, A2 => n18849, B1 => n21271, B2 => 
                           n21266, ZN => n18850);
   U22079 : XNOR2_X1 port map( A => n19123, B => n18852, ZN => n19575);
   U22081 : XNOR2_X1 port map( A => n19235, B => n3049, ZN => n18853);
   U22082 : XNOR2_X1 port map( A => n19125, B => n18853, ZN => n18854);
   U22083 : XNOR2_X1 port map( A => n18855, B => n18854, ZN => n20158);
   U22084 : XNOR2_X1 port map( A => n19206, B => n27894, ZN => n18858);
   U22086 : INV_X1 port map( A => n19096, ZN => n18859);
   U22087 : XNOR2_X1 port map( A => n19508, B => n18859, ZN => n19033);
   U22088 : XNOR2_X1 port map( A => n19116, B => n19033, ZN => n18860);
   U22089 : XNOR2_X1 port map( A => n18861, B => n18860, ZN => n20159);
   U22090 : NAND2_X1 port map( A1 => n20158, A2 => n20159, ZN => n19874);
   U22091 : XNOR2_X1 port map( A => n19250, B => n19256, ZN => n19583);
   U22092 : XNOR2_X1 port map( A => n19583, B => n18862, ZN => n18866);
   U22094 : XNOR2_X1 port map( A => n18863, B => n3154, ZN => n18864);
   U22095 : XNOR2_X1 port map( A => n19040, B => n18864, ZN => n18865);
   U22096 : INV_X1 port map( A => n20161, ZN => n19984);
   U22097 : NAND2_X1 port map( A1 => n19874, A2 => n19984, ZN => n18886);
   U22098 : INV_X1 port map( A => n18868, ZN => n18869);
   U22099 : XNOR2_X1 port map( A => n18869, B => n19599, ZN => n18873);
   U22100 : XNOR2_X1 port map( A => n19085, B => n19220, ZN => n18871);
   U22101 : XNOR2_X1 port map( A => n19481, B => n3752, ZN => n18870);
   U22102 : XNOR2_X1 port map( A => n18871, B => n18870, ZN => n18872);
   U22104 : INV_X1 port map( A => n20157, ZN => n20044);
   U22106 : XNOR2_X1 port map( A => n19192, B => n19103, ZN => n18876);
   U22107 : XNOR2_X1 port map( A => n19500, B => n2325, ZN => n18875);
   U22108 : INV_X1 port map( A => n19604, ZN => n19281);
   U22109 : NAND3_X1 port map( A1 => n19985, A2 => n20158, A3 => n29066, ZN => 
                           n18885);
   U22110 : XNOR2_X1 port map( A => n19243, B => n3650, ZN => n18879);
   U22111 : XNOR2_X1 port map( A => n19484, B => n19225, ZN => n18878);
   U22112 : XNOR2_X1 port map( A => n18879, B => n18878, ZN => n18882);
   U22113 : XNOR2_X1 port map( A => n18880, B => n19139, ZN => n19613);
   U22114 : XNOR2_X1 port map( A => n19141, B => n19613, ZN => n18881);
   U22115 : XNOR2_X1 port map( A => n18881, B => n18882, ZN => n20162);
   U22117 : NAND2_X1 port map( A1 => n28187, A2 => n20161, ZN => n20045);
   U22118 : INV_X1 port map( A => n21288, ZN => n20916);
   U22119 : INV_X1 port map( A => n18887, ZN => n20151);
   U22121 : NOR2_X1 port map( A1 => n18888, A2 => n28188, ZN => n18889);
   U22122 : NAND2_X1 port map( A1 => n20916, A2 => n20988, ZN => n21286);
   U22123 : OAI21_X1 port map( B1 => n18765, B2 => n19761, A => n20066, ZN => 
                           n18891);
   U22124 : XNOR2_X1 port map( A => n19462, B => n19378, ZN => n18893);
   U22125 : XNOR2_X1 port map( A => n18894, B => n18893, ZN => n18898);
   U22126 : XNOR2_X1 port map( A => n19299, B => n19377, ZN => n18896);
   U22127 : XNOR2_X1 port map( A => n19427, B => n3180, ZN => n18895);
   U22128 : XNOR2_X1 port map( A => n18896, B => n18895, ZN => n18897);
   U22129 : XNOR2_X2 port map( A => n18898, B => n18897, ZN => n18919);
   U22130 : XNOR2_X1 port map( A => n19251, B => n19256, ZN => n18901);
   U22131 : XNOR2_X1 port map( A => n18899, B => n18900, ZN => n19381);
   U22132 : XNOR2_X1 port map( A => n18901, B => n19381, ZN => n18905);
   U22133 : XNOR2_X1 port map( A => n19198, B => n19727, ZN => n18903);
   U22134 : XNOR2_X1 port map( A => n19643, B => n27105, ZN => n18902);
   U22135 : XNOR2_X1 port map( A => n18903, B => n18902, ZN => n18904);
   U22136 : XNOR2_X1 port map( A => n19086, B => n19045, ZN => n19635);
   U22137 : INV_X1 port map( A => n19635, ZN => n18907);
   U22138 : XNOR2_X1 port map( A => n19421, B => n19482, ZN => n19153);
   U22139 : XNOR2_X1 port map( A => n18907, B => n19153, ZN => n18911);
   U22140 : INV_X1 port map( A => n19084, ZN => n18909);
   U22141 : XNOR2_X1 port map( A => n19108, B => n21537, ZN => n18908);
   U22142 : XNOR2_X1 port map( A => n18909, B => n18908, ZN => n18910);
   U22143 : MUX2_X1 port map( A => n18919, B => n21091, S => n20144, Z => 
                           n18918);
   U22144 : XNOR2_X1 port map( A => n18912, B => n19025, ZN => n19651);
   U22145 : XNOR2_X1 port map( A => n19496, B => n19702, ZN => n19164);
   U22146 : XNOR2_X1 port map( A => n19651, B => n19164, ZN => n18917);
   U22147 : INV_X1 port map( A => n19105, ZN => n18915);
   U22148 : XNOR2_X1 port map( A => n18913, B => n3635, ZN => n18914);
   U22149 : XNOR2_X1 port map( A => n18915, B => n18914, ZN => n18916);
   U22150 : NOR2_X1 port map( A1 => n18918, A2 => n20145, ZN => n19011);
   U22151 : INV_X1 port map( A => n19011, ZN => n18932);
   U22152 : XNOR2_X1 port map( A => n19691, B => n19511, ZN => n18921);
   U22153 : INV_X1 port map( A => n19095, ZN => n18920);
   U22154 : XNOR2_X1 port map( A => n18920, B => n18921, ZN => n18926);
   U22155 : XNOR2_X1 port map( A => n19413, B => n18922, ZN => n18924);
   U22156 : XNOR2_X1 port map( A => n19412, B => n3697, ZN => n18923);
   U22157 : XNOR2_X1 port map( A => n18924, B => n18923, ZN => n18925);
   U22158 : INV_X1 port map( A => n18928, ZN => n19520);
   U22159 : XNOR2_X1 port map( A => n19487, B => n19229, ZN => n19181);
   U22160 : NOR2_X1 port map( A1 => n20102, A2 => n21091, ZN => n18930);
   U22161 : AOI22_X1 port map( A1 => n19010, A2 => n21091, B1 => n18930, B2 => 
                           n20145, ZN => n18931);
   U22162 : NAND2_X1 port map( A1 => n18932, A2 => n18931, ZN => n18934);
   U22163 : INV_X1 port map( A => n18934, ZN => n19014);
   U22164 : INV_X1 port map( A => n21291, ZN => n21289);
   U22165 : XNOR2_X1 port map( A => n19669, B => n29038, ZN => n18936);
   U22166 : XNOR2_X1 port map( A => n19519, B => n18936, ZN => n18941);
   U22167 : XNOR2_X1 port map( A => n19228, B => n18937, ZN => n18939);
   U22168 : XNOR2_X1 port map( A => n19246, B => n3256, ZN => n18938);
   U22169 : XNOR2_X1 port map( A => n18939, B => n18938, ZN => n18940);
   U22170 : XNOR2_X1 port map( A => n18941, B => n18940, ZN => n20165);
   U22171 : XNOR2_X1 port map( A => n28143, B => n19637, ZN => n18945);
   U22172 : XNOR2_X1 port map( A => n18942, B => n3491, ZN => n18943);
   U22173 : XNOR2_X1 port map( A => n18943, B => n19679, ZN => n18944);
   U22174 : XNOR2_X1 port map( A => n18944, B => n18945, ZN => n18947);
   U22176 : XNOR2_X1 port map( A => n19557, B => n29484, ZN => n18946);
   U22177 : XNOR2_X1 port map( A => n18946, B => n18947, ZN => n18972);
   U22178 : XNOR2_X1 port map( A => n19144, B => n19548, ZN => n18953);
   U22179 : XNOR2_X1 port map( A => n19725, B => n19644, ZN => n18951);
   U22180 : XNOR2_X1 port map( A => n18949, B => n2389, ZN => n18950);
   U22181 : XNOR2_X1 port map( A => n18951, B => n18950, ZN => n18952);
   U22182 : AOI21_X1 port map( B1 => n18972, B2 => n20165, A => n20166, ZN => 
                           n18974);
   U22183 : XNOR2_X1 port map( A => n29506, B => n2602, ZN => n18954);
   U22184 : XNOR2_X1 port map( A => n18955, B => n18954, ZN => n18957);
   U22185 : XNOR2_X1 port map( A => n19191, B => n19403, ZN => n19132);
   U22186 : XNOR2_X1 port map( A => n19132, B => n19541, ZN => n18956);
   U22187 : XNOR2_X1 port map( A => n18956, B => n18957, ZN => n19993);
   U22189 : INV_X1 port map( A => n19626, ZN => n18958);
   U22190 : XNOR2_X1 port map( A => n18958, B => n19408, ZN => n18961);
   U22191 : XNOR2_X1 port map( A => n18960, B => n18959, ZN => n19526);
   U22192 : XNOR2_X1 port map( A => n19526, B => n18961, ZN => n18965);
   U22193 : XNOR2_X1 port map( A => n19696, B => n19697, ZN => n18963);
   U22194 : XNOR2_X1 port map( A => n19207, B => n3003, ZN => n18962);
   U22195 : XNOR2_X1 port map( A => n18963, B => n18962, ZN => n18964);
   U22196 : MUX2_X1 port map( A => n29587, B => n297, S => n19989, Z => n18973)
                           ;
   U22197 : INV_X1 port map( A => n18966, ZN => n19533);
   U22198 : XNOR2_X1 port map( A => n19533, B => n18967, ZN => n18971);
   U22199 : XNOR2_X1 port map( A => n19272, B => n19632, ZN => n18969);
   U22200 : XNOR2_X1 port map( A => n19685, B => n3276, ZN => n18968);
   U22201 : XNOR2_X1 port map( A => n18969, B => n18968, ZN => n18970);
   U22202 : INV_X1 port map( A => n21290, ZN => n20986);
   U22203 : INV_X1 port map( A => n19331, ZN => n18976);
   U22204 : INV_X1 port map( A => n18975, ZN => n19625);
   U22205 : XNOR2_X1 port map( A => n18976, B => n19625, ZN => n19094);
   U22206 : XNOR2_X1 port map( A => n19094, B => n19330, ZN => n18979);
   U22207 : XNOR2_X1 port map( A => n19525, B => n19507, ZN => n19212);
   U22208 : XNOR2_X1 port map( A => n19212, B => n18977, ZN => n18978);
   U22209 : XNOR2_X1 port map( A => n18979, B => n18978, ZN => n19054);
   U22210 : XNOR2_X1 port map( A => n18981, B => n18980, ZN => n18983);
   U22211 : XNOR2_X1 port map( A => n19483, B => n3457, ZN => n18982);
   U22212 : XNOR2_X1 port map( A => n18983, B => n18982, ZN => n18986);
   U22213 : XNOR2_X1 port map( A => n19631, B => n19110, ZN => n19082);
   U22214 : XNOR2_X1 port map( A => n19082, B => n18984, ZN => n18985);
   U22215 : XNOR2_X1 port map( A => n19549, B => n3501, ZN => n18990);
   U22217 : XNOR2_X1 port map( A => n29554, B => n19397, ZN => n18992);
   U22219 : XNOR2_X1 port map( A => n19617, B => n2306, ZN => n18994);
   U22220 : XNOR2_X1 port map( A => n18995, B => n18994, ZN => n18996);
   U22221 : XNOR2_X1 port map( A => n18997, B => n18996, ZN => n20053);
   U22222 : INV_X1 port map( A => n19333, ZN => n18998);
   U22223 : XNOR2_X1 port map( A => n29318, B => n19376, ZN => n19079);
   U22224 : XNOR2_X1 port map( A => n19428, B => n3742, ZN => n18999);
   U22225 : XNOR2_X1 port map( A => n19079, B => n18999, ZN => n19000);
   U22226 : XNOR2_X1 port map( A => n19000, B => n19001, ZN => n20178);
   U22229 : OAI21_X1 port map( B1 => n20174, B2 => n4886, A => n19002, ZN => 
                           n19008);
   U22230 : XNOR2_X1 port map( A => n28516, B => n19603, ZN => n19101);
   U22231 : XNOR2_X1 port map( A => n19495, B => n19356, ZN => n19005);
   U22232 : XNOR2_X1 port map( A => n19006, B => n19005, ZN => n20176);
   U22233 : INV_X1 port map( A => n19052, ZN => n19007);
   U22234 : NOR2_X1 port map( A1 => n21291, A2 => n21287, ZN => n19013);
   U22235 : XNOR2_X1 port map( A => n22582, B => n21884, ZN => n19738);
   U22236 : XNOR2_X1 port map( A => n19371, B => n19378, ZN => n19015);
   U22237 : XNOR2_X1 port map( A => n19313, B => n24906, ZN => n19019);
   U22238 : XNOR2_X1 port map( A => n19020, B => n19019, ZN => n19023);
   U22239 : XNOR2_X1 port map( A => n19484, B => n19487, ZN => n19021);
   U22240 : XNOR2_X1 port map( A => n19399, B => n19021, ZN => n19022);
   U22241 : XNOR2_X1 port map( A => n19023, B => n19022, ZN => n20479);
   U22242 : XNOR2_X1 port map( A => n19496, B => n19024, ZN => n19027);
   U22243 : XNOR2_X1 port map( A => n19027, B => n19026, ZN => n19031);
   U22244 : XNOR2_X1 port map( A => n19700, B => n2446, ZN => n19029);
   U22245 : XNOR2_X1 port map( A => n19500, B => n19452, ZN => n19028);
   U22246 : XNOR2_X1 port map( A => n19029, B => n19028, ZN => n19030);
   U22247 : XNOR2_X1 port map( A => n19409, B => n19511, ZN => n19034);
   U22248 : XNOR2_X1 port map( A => n19033, B => n19034, ZN => n19038);
   U22249 : XNOR2_X1 port map( A => n19413, B => n3770, ZN => n19035);
   U22250 : XNOR2_X1 port map( A => n19036, B => n19035, ZN => n19037);
   U22251 : INV_X1 port map( A => n19039, ZN => n19382);
   U22252 : XNOR2_X1 port map( A => n19382, B => n19040, ZN => n19044);
   U22253 : INV_X1 port map( A => n1184, ZN => n19041);
   U22254 : XNOR2_X1 port map( A => n19440, B => n19041, ZN => n19042);
   U22255 : XNOR2_X1 port map( A => n19472, B => n19042, ZN => n19043);
   U22256 : XNOR2_X1 port map( A => n19044, B => n19043, ZN => n19995);
   U22257 : XNOR2_X1 port map( A => n19423, B => n19085, ZN => n19047);
   U22258 : XNOR2_X1 port map( A => n19045, B => n19481, ZN => n19046);
   U22259 : XNOR2_X1 port map( A => n19047, B => n19046, ZN => n19051);
   U22260 : XNOR2_X1 port map( A => n19482, B => n19306, ZN => n19049);
   U22261 : XNOR2_X1 port map( A => n19049, B => n19048, ZN => n19050);
   U22262 : INV_X1 port map( A => n19054, ZN => n19976);
   U22263 : OAI21_X1 port map( B1 => n19055, B2 => n19976, A => n20171, ZN => 
                           n19056);
   U22264 : INV_X1 port map( A => n21277, ZN => n21278);
   U22265 : NOR2_X1 port map( A1 => n297, A2 => n20219, ZN => n19059);
   U22266 : NOR3_X1 port map( A1 => n19860, A2 => n19059, A3 => n20222, ZN => 
                           n19063);
   U22267 : NAND3_X1 port map( A1 => n19989, A2 => n385, A3 => n296, ZN => 
                           n19061);
   U22268 : NAND2_X1 port map( A1 => n21278, A2 => n21703, ZN => n21378);
   U22269 : XNOR2_X1 port map( A => n19615, B => n2381, ZN => n19064);
   U22270 : XNOR2_X1 port map( A => n19665, B => n19064, ZN => n19068);
   U22271 : XNOR2_X1 port map( A => n19066, B => n19065, ZN => n19067);
   U22272 : XNOR2_X1 port map( A => n19251, B => n19727, ZN => n19070);
   U22273 : XNOR2_X1 port map( A => n19584, B => n2912, ZN => n19069);
   U22274 : XNOR2_X1 port map( A => n19070, B => n19069, ZN => n19074);
   U22275 : INV_X1 port map( A => n19071, ZN => n19072);
   U22276 : XNOR2_X1 port map( A => n19646, B => n19072, ZN => n19073);
   U22277 : INV_X1 port map( A => n19093, ZN => n20486);
   U22278 : NOR2_X1 port map( A1 => n20481, A2 => n20486, ZN => n20238);
   U22279 : XNOR2_X1 port map( A => n19075, B => n3451, ZN => n19076);
   U22280 : XNOR2_X1 port map( A => n19077, B => n19076, ZN => n19081);
   U22281 : XNOR2_X1 port map( A => n19079, B => n19078, ZN => n19080);
   U22282 : INV_X1 port map( A => n19082, ZN => n19083);
   U22283 : XNOR2_X1 port map( A => n19083, B => n19084, ZN => n19091);
   U22284 : XNOR2_X1 port map( A => n19086, B => n19085, ZN => n19089);
   U22285 : XNOR2_X1 port map( A => n19087, B => n26909, ZN => n19088);
   U22286 : XNOR2_X1 port map( A => n19089, B => n19088, ZN => n19090);
   U22287 : INV_X1 port map( A => n20483, ZN => n20000);
   U22288 : XNOR2_X1 port map( A => n19094, B => n19095, ZN => n19100);
   U22289 : XNOR2_X1 port map( A => n19096, B => n2894, ZN => n19098);
   U22290 : XNOR2_X1 port map( A => n19098, B => n19097, ZN => n19099);
   U22291 : XNOR2_X1 port map( A => n19101, B => n19102, ZN => n19107);
   U22292 : XNOR2_X1 port map( A => n19103, B => n730, ZN => n19104);
   U22293 : XNOR2_X1 port map( A => n19105, B => n19104, ZN => n19106);
   U22294 : NOR2_X1 port map( A1 => n20488, A2 => n20239, ZN => n20482);
   U22295 : XNOR2_X1 port map( A => n19272, B => n19688, ZN => n19388);
   U22296 : XNOR2_X1 port map( A => n19219, B => n19108, ZN => n19109);
   U22297 : XNOR2_X1 port map( A => n19109, B => n19388, ZN => n19115);
   U22298 : XNOR2_X1 port map( A => n19110, B => n3081, ZN => n19113);
   U22299 : XNOR2_X1 port map( A => n19113, B => n19112, ZN => n19114);
   U22300 : XNOR2_X1 port map( A => n19115, B => n19114, ZN => n20499);
   U22301 : INV_X1 port map( A => n20499, ZN => n20227);
   U22302 : XNOR2_X1 port map( A => n19116, B => n19117, ZN => n19121);
   U22303 : XNOR2_X1 port map( A => n19207, B => n24959, ZN => n19118);
   U22304 : XNOR2_X1 port map( A => n19119, B => n19118, ZN => n19120);
   U22306 : XNOR2_X1 port map( A => n28144, B => n19373, ZN => n19124);
   U22307 : XNOR2_X1 port map( A => n29318, B => n3662, ZN => n19126);
   U22308 : XNOR2_X1 port map( A => n19125, B => n19126, ZN => n19127);
   U22310 : MUX2_X1 port map( A => n20227, B => n28621, S => n20500, Z => 
                           n19151);
   U22311 : INV_X1 port map( A => n19130, ZN => n19131);
   U22312 : XNOR2_X1 port map( A => n19603, B => n2402, ZN => n19134);
   U22313 : XNOR2_X1 port map( A => n19133, B => n19134, ZN => n19135);
   U22314 : XNOR2_X1 port map( A => n19616, B => n19228, ZN => n19138);
   U22315 : XNOR2_X1 port map( A => n19136, B => n2411, ZN => n19137);
   U22316 : XNOR2_X1 port map( A => n19138, B => n19137, ZN => n19143);
   U22317 : XNOR2_X1 port map( A => n19139, B => n19615, ZN => n19140);
   U22318 : XNOR2_X1 port map( A => n19141, B => n19140, ZN => n19142);
   U22319 : XNOR2_X1 port map( A => n18395, B => n19359, ZN => n19145);
   U22320 : XNOR2_X1 port map( A => n19256, B => n19726, ZN => n19147);
   U22321 : XNOR2_X1 port map( A => n19584, B => n2404, ZN => n19146);
   U22322 : XNOR2_X1 port map( A => n19147, B => n19146, ZN => n19148);
   U22323 : NOR2_X1 port map( A1 => n20500, A2 => n20339, ZN => n19149);
   U22324 : AOI21_X2 port map( B1 => n19151, B2 => n19150, A => n19149, ZN => 
                           n21704);
   U22325 : XNOR2_X1 port map( A => n19687, B => n19305, ZN => n19152);
   U22326 : INV_X1 port map( A => n3380, ZN => n27811);
   U22327 : XNOR2_X1 port map( A => n19370, B => n2946, ZN => n19155);
   U22328 : XNOR2_X1 port map( A => n19155, B => n19234, ZN => n19158);
   U22329 : XNOR2_X1 port map( A => n19156, B => n19296, ZN => n19157);
   U22330 : INV_X1 port map( A => n20493, ZN => n20179);
   U22331 : XNOR2_X1 port map( A => n18760, B => n28798, ZN => n19161);
   U22332 : XNOR2_X1 port map( A => n19198, B => n2981, ZN => n19160);
   U22333 : XNOR2_X1 port map( A => n19161, B => n19160, ZN => n19163);
   U22334 : XNOR2_X1 port map( A => n19164, B => n19165, ZN => n19169);
   U22335 : XNOR2_X1 port map( A => n19166, B => n19706, ZN => n19167);
   U22336 : XNOR2_X1 port map( A => n19691, B => n19321, ZN => n19171);
   U22337 : XNOR2_X1 port map( A => n19696, B => n19511, ZN => n19170);
   U22338 : XNOR2_X1 port map( A => n19171, B => n19170, ZN => n19178);
   U22339 : INV_X1 port map( A => n19173, ZN => n19172);
   U22340 : NAND2_X1 port map( A1 => n19172, A2 => n5490, ZN => n19174);
   U22341 : INV_X1 port map( A => Key(26), ZN => n24166);
   U22342 : XNOR2_X1 port map( A => n19176, B => n19175, ZN => n19177);
   U22343 : INV_X1 port map( A => n20496, ZN => n19863);
   U22344 : XNOR2_X1 port map( A => n19180, B => n19348, ZN => n19182);
   U22345 : XNOR2_X1 port map( A => n19182, B => n19181, ZN => n19184);
   U22346 : XNOR2_X1 port map( A => n19184, B => n19183, ZN => n20182);
   U22348 : MUX2_X1 port map( A => n19187, B => n21374, S => n21372, Z => 
                           n19188);
   U22351 : XNOR2_X1 port map( A => n19191, B => n19702, ZN => n19193);
   U22352 : XNOR2_X1 port map( A => n19194, B => n19277, ZN => n19195);
   U22353 : XNOR2_X1 port map( A => n19495, B => n19195, ZN => n19196);
   U22354 : XNOR2_X1 port map( A => n19197, B => n19196, ZN => n20017);
   U22355 : XNOR2_X1 port map( A => n19199, B => n19198, ZN => n19201);
   U22356 : XNOR2_X1 port map( A => n19549, B => n2505, ZN => n19200);
   U22357 : XNOR2_X1 port map( A => n19201, B => n19200, ZN => n19205);
   U22358 : XNOR2_X1 port map( A => n28798, B => n19474, ZN => n19202);
   U22359 : XNOR2_X1 port map( A => n19202, B => n19203, ZN => n19204);
   U22360 : XNOR2_X1 port map( A => n19206, B => n19332, ZN => n19209);
   U22361 : XNOR2_X1 port map( A => n19207, B => n3586, ZN => n19208);
   U22362 : XNOR2_X1 port map( A => n19209, B => n19208, ZN => n19214);
   U22365 : INV_X1 port map( A => n19215, ZN => n19216);
   U22366 : XNOR2_X1 port map( A => n19216, B => n19483, ZN => n19218);
   U22367 : XNOR2_X1 port map( A => n19339, B => n2527, ZN => n19217);
   U22368 : XNOR2_X1 port map( A => n19218, B => n19217, ZN => n19224);
   U22369 : XNOR2_X1 port map( A => n19534, B => n19219, ZN => n19222);
   U22370 : XNOR2_X1 port map( A => n19421, B => n19220, ZN => n19221);
   U22371 : XNOR2_X1 port map( A => n19222, B => n19221, ZN => n19223);
   U22373 : XNOR2_X1 port map( A => n19348, B => n19226, ZN => n19227);
   U22374 : XNOR2_X1 port map( A => n19670, B => n19228, ZN => n19230);
   U22375 : XNOR2_X1 port map( A => n19230, B => n19229, ZN => n19231);
   U22376 : INV_X1 port map( A => n20342, ZN => n20509);
   U22377 : XNOR2_X1 port map( A => n19232, B => n1919, ZN => n19233);
   U22378 : XNOR2_X1 port map( A => n19234, B => n19233, ZN => n19239);
   U22379 : XNOR2_X1 port map( A => n28143, B => n19235, ZN => n19237);
   U22380 : XNOR2_X1 port map( A => n19236, B => n19237, ZN => n19238);
   U22381 : OAI21_X1 port map( B1 => n20509, B2 => n20510, A => n20343, ZN => 
                           n19240);
   U22383 : XNOR2_X1 port map( A => n19670, B => n3462, ZN => n19242);
   U22384 : XNOR2_X1 port map( A => n19242, B => n19243, ZN => n19244);
   U22385 : XNOR2_X1 port map( A => n19244, B => n19613, ZN => n19249);
   U22386 : XNOR2_X1 port map( A => n19245, B => n19246, ZN => n19247);
   U22387 : XNOR2_X1 port map( A => n19249, B => n19248, ZN => n20458);
   U22388 : INV_X1 port map( A => n20458, ZN => n20028);
   U22389 : XNOR2_X1 port map( A => n19250, B => n19251, ZN => n19254);
   U22391 : XNOR2_X1 port map( A => n19256, B => n28798, ZN => n19258);
   U22392 : XNOR2_X1 port map( A => n19474, B => n26214, ZN => n19257);
   U22393 : XNOR2_X1 port map( A => n19258, B => n19257, ZN => n19259);
   U22394 : XNOR2_X1 port map( A => n19462, B => n29484, ZN => n19261);
   U22395 : XNOR2_X1 port map( A => n19575, B => n19261, ZN => n19264);
   U22396 : XNOR2_X1 port map( A => n19262, B => n2961, ZN => n19263);
   U22397 : INV_X1 port map( A => n19628, ZN => n19266);
   U22398 : XNOR2_X1 port map( A => n19408, B => n19332, ZN => n19265);
   U22400 : XNOR2_X1 port map( A => n19267, B => n1123, ZN => n19268);
   U22401 : XNOR2_X1 port map( A => n19269, B => n19268, ZN => n19270);
   U22402 : XNOR2_X1 port map( A => n19272, B => n19273, ZN => n19275);
   U22403 : XNOR2_X1 port map( A => n19339, B => n3372, ZN => n19274);
   U22404 : XNOR2_X1 port map( A => n19275, B => n19274, ZN => n19276);
   U22405 : XNOR2_X1 port map( A => n19277, B => n28294, ZN => n19280);
   U22406 : XNOR2_X1 port map( A => n19278, B => n19403, ZN => n19279);
   U22407 : INV_X1 port map( A => n19283, ZN => n19701);
   U22408 : XNOR2_X1 port map( A => n19701, B => n3323, ZN => n19284);
   U22409 : XNOR2_X1 port map( A => n19284, B => n19285, ZN => n19288);
   U22410 : XNOR2_X1 port map( A => n28516, B => n18638, ZN => n19286);
   U22411 : XNOR2_X1 port map( A => n19498, B => n19286, ZN => n19287);
   U22414 : XNOR2_X1 port map( A => n19291, B => n28571, ZN => n19293);
   U22415 : XNOR2_X1 port map( A => n19475, B => n3134, ZN => n19292);
   U22416 : XNOR2_X1 port map( A => n19293, B => n19292, ZN => n19294);
   U22417 : XNOR2_X2 port map( A => n19295, B => n19294, ZN => n20334);
   U22418 : INV_X1 port map( A => n19296, ZN => n19297);
   U22419 : XNOR2_X1 port map( A => n19297, B => n19298, ZN => n19304);
   U22420 : XNOR2_X1 port map( A => n19299, B => n19300, ZN => n19302);
   U22421 : XNOR2_X1 port map( A => n19376, B => n2477, ZN => n19301);
   U22422 : XNOR2_X1 port map( A => n19302, B => n19301, ZN => n19303);
   U22423 : XNOR2_X2 port map( A => n19304, B => n19303, ZN => n20623);
   U22424 : XNOR2_X1 port map( A => n19631, B => n19481, ZN => n19307);
   U22425 : XNOR2_X1 port map( A => n19308, B => n19307, ZN => n19312);
   U22426 : XNOR2_X1 port map( A => n19595, B => n19535, ZN => n19310);
   U22427 : XNOR2_X1 port map( A => n19685, B => n3482, ZN => n19309);
   U22428 : XNOR2_X1 port map( A => n19310, B => n19309, ZN => n19311);
   U22430 : XNOR2_X1 port map( A => n6489, B => n19397, ZN => n19314);
   U22431 : XNOR2_X1 port map( A => n19520, B => n3015, ZN => n19316);
   U22432 : XNOR2_X1 port map( A => n19317, B => n19316, ZN => n19318);
   U22433 : INV_X1 port map( A => n20630, ZN => n20335);
   U22434 : XNOR2_X1 port map( A => n19592, B => n19323, ZN => n19529);
   U22435 : XNOR2_X1 port map( A => n19625, B => n3710, ZN => n19324);
   U22436 : XNOR2_X1 port map( A => n19529, B => n19324, ZN => n19325);
   U22438 : NAND2_X1 port map( A1 => n20625, A2 => n20623, ZN => n19327);
   U22439 : MUX2_X1 port map( A => n19328, B => n19327, S => n20005, Z => 
                           n19329);
   U22440 : OAI21_X1 port map( B1 => n21364, B2 => n21713, A => n21714, ZN => 
                           n19461);
   U22441 : INV_X1 port map( A => n21364, ZN => n21258);
   U22442 : XNOR2_X1 port map( A => n19331, B => n19626, ZN => n19591);
   U22443 : XNOR2_X1 port map( A => n19333, B => n28530, ZN => n19335);
   U22444 : XNOR2_X1 port map( A => n19568, B => n3422, ZN => n19334);
   U22445 : XNOR2_X1 port map( A => n19335, B => n19334, ZN => n19337);
   U22446 : XNOR2_X2 port map( A => n19337, B => n19336, ZN => n20617);
   U22447 : INV_X1 port map( A => n19339, ZN => n19340);
   U22448 : XNOR2_X1 port map( A => n19423, B => n19340, ZN => n19342);
   U22449 : XNOR2_X1 port map( A => n19342, B => n19341, ZN => n19343);
   U22450 : XNOR2_X1 port map( A => n19343, B => n19344, ZN => n20431);
   U22451 : NOR2_X1 port map( A1 => n20617, A2 => n29040, ZN => n19345);
   U22452 : XNOR2_X1 port map( A => n19346, B => n19669, ZN => n19347);
   U22453 : XNOR2_X1 port map( A => n19348, B => n19615, ZN => n19351);
   U22454 : XNOR2_X1 port map( A => n19349, B => n3508, ZN => n19350);
   U22455 : XNOR2_X1 port map( A => n19350, B => n19351, ZN => n19352);
   U22456 : XNOR2_X1 port map( A => n19452, B => n135, ZN => n19355);
   U22458 : INV_X1 port map( A => n20616, ZN => n20433);
   U22459 : XNOR2_X1 port map( A => n19359, B => n19440, ZN => n19361);
   U22460 : XNOR2_X1 port map( A => n29124, B => n19361, ZN => n19366);
   U22461 : XNOR2_X1 port map( A => n19584, B => n2523, ZN => n19364);
   U22462 : INV_X1 port map( A => n19362, ZN => n19363);
   U22463 : XNOR2_X1 port map( A => n19364, B => n19363, ZN => n19365);
   U22464 : OAI21_X1 port map( B1 => n20255, B2 => n20433, A => n28894, ZN => 
                           n19368);
   U22465 : NOR2_X1 port map( A1 => n19920, A2 => n20617, ZN => n19367);
   U22466 : AOI21_X2 port map( B1 => n19369, B2 => n19368, A => n19367, ZN => 
                           n21366);
   U22467 : INV_X1 port map( A => n21366, ZN => n21712);
   U22468 : AOI21_X1 port map( B1 => n21712, B2 => n5772, A => n21714, ZN => 
                           n19419);
   U22469 : XNOR2_X1 port map( A => n19370, B => n27452, ZN => n19372);
   U22470 : XNOR2_X1 port map( A => n19372, B => n19371, ZN => n19375);
   U22471 : XNOR2_X1 port map( A => n19464, B => n19373, ZN => n19374);
   U22472 : XNOR2_X1 port map( A => n19375, B => n19374, ZN => n19380);
   U22473 : XNOR2_X1 port map( A => n19377, B => n19376, ZN => n19379);
   U22475 : XNOR2_X1 port map( A => n19380, B => n19641, ZN => n20033);
   U22476 : INV_X1 port map( A => n20033, ZN => n20247);
   U22477 : XNOR2_X1 port map( A => n19726, B => n19383, ZN => n19386);
   U22478 : XNOR2_X1 port map( A => n19384, B => n3067, ZN => n19385);
   U22479 : XNOR2_X1 port map( A => n19386, B => n19385, ZN => n19387);
   U22480 : XNOR2_X1 port map( A => n19388, B => n19635, ZN => n19393);
   U22481 : XNOR2_X1 port map( A => n19389, B => n2476, ZN => n19390);
   U22482 : XNOR2_X1 port map( A => n19391, B => n19390, ZN => n19392);
   U22483 : XNOR2_X1 port map( A => n19393, B => n19392, ZN => n20453);
   U22484 : NOR2_X1 port map( A1 => n20641, A2 => n20453, ZN => n20689);
   U22485 : INV_X1 port map( A => n20689, ZN => n19394);
   U22486 : NAND2_X1 port map( A1 => n21364, A2 => n19394, ZN => n19417);
   U22487 : XNOR2_X1 port map( A => n18927, B => n2987, ZN => n19396);
   U22488 : XNOR2_X1 port map( A => n19486, B => n19616, ZN => n19395);
   U22489 : XNOR2_X1 port map( A => n19396, B => n19395, ZN => n19401);
   U22490 : XNOR2_X1 port map( A => n19487, B => n19397, ZN => n19398);
   U22491 : XNOR2_X1 port map( A => n19399, B => n19398, ZN => n19400);
   U22492 : XNOR2_X1 port map( A => n19402, B => n19651, ZN => n19407);
   U22493 : XNOR2_X1 port map( A => n19403, B => n19709, ZN => n19405);
   U22494 : XNOR2_X1 port map( A => n19700, B => n3463, ZN => n19404);
   U22495 : XNOR2_X1 port map( A => n19405, B => n19404, ZN => n19406);
   U22496 : XNOR2_X1 port map( A => n19407, B => n19406, ZN => n19787);
   U22497 : XNOR2_X1 port map( A => n19409, B => n19408, ZN => n19411);
   U22498 : XNOR2_X1 port map( A => n19410, B => n19411, ZN => n19416);
   U22499 : XNOR2_X1 port map( A => n19695, B => n27231, ZN => n19414);
   U22500 : XNOR2_X1 port map( A => n19624, B => n19414, ZN => n19415);
   U22501 : INV_X1 port map( A => n20455, ZN => n20639);
   U22502 : NOR2_X1 port map( A1 => n21716, A2 => n21258, ZN => n19460);
   U22503 : XNOR2_X1 port map( A => n19421, B => n19686, ZN => n19422);
   U22504 : XNOR2_X1 port map( A => n19632, B => n1172, ZN => n19425);
   U22505 : XNOR2_X1 port map( A => n19423, B => n19481, ZN => n19424);
   U22507 : XNOR2_X1 port map( A => n19428, B => n19427, ZN => n19429);
   U22508 : XNOR2_X1 port map( A => n19430, B => n19429, ZN => n19431);
   U22510 : XNOR2_X1 port map( A => n19433, B => n19691, ZN => n19435);
   U22511 : XNOR2_X1 port map( A => n19508, B => n19626, ZN => n19434);
   U22512 : XNOR2_X1 port map( A => n19435, B => n19434, ZN => n19437);
   U22515 : INV_X1 port map( A => n19438, ZN => n19724);
   U22516 : XNOR2_X1 port map( A => n19724, B => n19439, ZN => n19444);
   U22517 : XNOR2_X1 port map( A => n19440, B => n19644, ZN => n19442);
   U22518 : XNOR2_X1 port map( A => n19475, B => n2509, ZN => n19441);
   U22519 : XNOR2_X1 port map( A => n19442, B => n19441, ZN => n19443);
   U22520 : XNOR2_X1 port map( A => n19484, B => n19669, ZN => n19446);
   U22521 : XNOR2_X1 port map( A => n19445, B => n19446, ZN => n19451);
   U22522 : INV_X1 port map( A => n19447, ZN => n19714);
   U22523 : XNOR2_X1 port map( A => n19448, B => n1215, ZN => n19449);
   U22524 : XNOR2_X1 port map( A => n19714, B => n19449, ZN => n19450);
   U22525 : XNOR2_X1 port map( A => n19450, B => n19451, ZN => n20020);
   U22526 : INV_X1 port map( A => n20020, ZN => n20520);
   U22527 : NOR2_X1 port map( A1 => n20261, A2 => n20520, ZN => n21360);
   U22528 : XNOR2_X1 port map( A => n19452, B => n28623, ZN => n19453);
   U22529 : XNOR2_X1 port map( A => n19454, B => n19453, ZN => n19456);
   U22531 : MUX2_X1 port map( A => n19457, B => n21360, S => n28586, Z => 
                           n19459);
   U22533 : XNOR2_X1 port map( A => n22671, B => n22698, ZN => n22031);
   U22534 : INV_X1 port map( A => n22031, ZN => n21756);
   U22535 : XNOR2_X1 port map( A => n29580, B => n19462, ZN => n19467);
   U22536 : XNOR2_X1 port map( A => n19464, B => n19465, ZN => n19466);
   U22537 : XNOR2_X1 port map( A => n19466, B => n19467, ZN => n19471);
   U22538 : INV_X1 port map( A => n27422, ZN => n25250);
   U22539 : XNOR2_X1 port map( A => n19468, B => n25250, ZN => n19469);
   U22540 : XNOR2_X1 port map( A => n19474, B => n19726, ZN => n19477);
   U22541 : XNOR2_X1 port map( A => n19475, B => n2982, ZN => n19476);
   U22542 : XNOR2_X1 port map( A => n19477, B => n19476, ZN => n19478);
   U22543 : INV_X1 port map( A => n20130, ZN => n19901);
   U22544 : MUX2_X1 port map( A => n20443, B => n415, S => n19901, Z => n19506)
                           ;
   U22545 : XNOR2_X1 port map( A => n19670, B => n3673, ZN => n19485);
   U22546 : XNOR2_X1 port map( A => n19484, B => n19485, ZN => n19489);
   U22547 : XNOR2_X1 port map( A => n19486, B => n19487, ZN => n19488);
   U22548 : XNOR2_X1 port map( A => n19489, B => n19488, ZN => n19494);
   U22549 : XNOR2_X1 port map( A => n19491, B => n19490, ZN => n19492);
   U22550 : INV_X1 port map( A => n19495, ZN => n19497);
   U22551 : XNOR2_X1 port map( A => n19496, B => n19497, ZN => n19499);
   U22552 : XNOR2_X1 port map( A => n19498, B => n19499, ZN => n19504);
   U22553 : XNOR2_X1 port map( A => n19500, B => n1161, ZN => n19501);
   U22554 : XNOR2_X1 port map( A => n19502, B => n19501, ZN => n19503);
   U22555 : XNOR2_X1 port map( A => n19507, B => n19508, ZN => n19509);
   U22556 : XNOR2_X1 port map( A => n19510, B => n19509, ZN => n19515);
   U22557 : XNOR2_X1 port map( A => n19511, B => n2577, ZN => n19512);
   U22558 : XNOR2_X1 port map( A => n19513, B => n19512, ZN => n19514);
   U22559 : INV_X1 port map( A => n20125, ZN => n20294);
   U22560 : INV_X1 port map( A => n20293, ZN => n19814);
   U22561 : INV_X1 port map( A => n20123, ZN => n19969);
   U22562 : INV_X1 port map( A => n20295, ZN => n19818);
   U22563 : AOI21_X1 port map( B1 => n20290, B2 => n19969, A => n19818, ZN => 
                           n19517);
   U22564 : NAND2_X1 port map( A1 => n20123, A2 => n19814, ZN => n19516);
   U22565 : XNOR2_X1 port map( A => n19519, B => n19518, ZN => n19524);
   U22566 : XNOR2_X1 port map( A => n19520, B => n19611, ZN => n19522);
   U22567 : XNOR2_X1 port map( A => n19617, B => n3196, ZN => n19521);
   U22568 : XNOR2_X1 port map( A => n19522, B => n19521, ZN => n19523);
   U22569 : XNOR2_X1 port map( A => n19524, B => n19523, ZN => n20647);
   U22570 : XNOR2_X1 port map( A => n19525, B => n3644, ZN => n19527);
   U22571 : XNOR2_X1 port map( A => n19526, B => n19527, ZN => n19531);
   U22572 : XNOR2_X1 port map( A => n19528, B => n19529, ZN => n19530);
   U22574 : XNOR2_X1 port map( A => n19533, B => n19532, ZN => n19539);
   U22575 : XNOR2_X1 port map( A => n19595, B => n19534, ZN => n19537);
   U22576 : XNOR2_X1 port map( A => n19535, B => n3334, ZN => n19536);
   U22577 : XNOR2_X1 port map( A => n19537, B => n19536, ZN => n19538);
   U22578 : INV_X1 port map( A => n19540, ZN => n19542);
   U22579 : XNOR2_X1 port map( A => n19542, B => n19541, ZN => n19545);
   U22580 : INV_X1 port map( A => n19546, ZN => n19547);
   U22581 : XNOR2_X1 port map( A => n19547, B => n19548, ZN => n19553);
   U22582 : XNOR2_X1 port map( A => n19727, B => n19585, ZN => n19551);
   U22583 : XNOR2_X1 port map( A => n19549, B => n2441, ZN => n19550);
   U22584 : XNOR2_X1 port map( A => n19551, B => n19550, ZN => n19552);
   U22585 : XNOR2_X1 port map( A => n19555, B => n28143, ZN => n19558);
   U22586 : XNOR2_X1 port map( A => n19557, B => n19558, ZN => n19572);
   U22587 : INV_X1 port map( A => n19559, ZN => n19566);
   U22588 : NAND3_X1 port map( A1 => n29125, A2 => n29044, A3 => n123, ZN => 
                           n19563);
   U22589 : NAND2_X1 port map( A1 => n19564, A2 => n19563, ZN => n19565);
   U22590 : NOR2_X1 port map( A1 => n19566, A2 => n19565, ZN => n19567);
   U22591 : XNOR2_X1 port map( A => n19577, B => n19567, ZN => n19570);
   U22592 : XNOR2_X1 port map( A => n19570, B => n19569, ZN => n19571);
   U22593 : XNOR2_X1 port map( A => n19571, B => n19572, ZN => n19928);
   U22594 : OAI21_X1 port map( B1 => n21807, B2 => n21806, A => n21253, ZN => 
                           n19735);
   U22595 : XNOR2_X1 port map( A => n19574, B => n19575, ZN => n19581);
   U22596 : XNOR2_X1 port map( A => n19637, B => n29318, ZN => n19579);
   U22597 : XNOR2_X1 port map( A => n19577, B => n3528, ZN => n19578);
   U22598 : XNOR2_X1 port map( A => n19579, B => n19578, ZN => n19580);
   U22599 : XNOR2_X1 port map( A => n19583, B => n19582, ZN => n19589);
   U22600 : XNOR2_X1 port map( A => n19584, B => n3378, ZN => n19587);
   U22601 : XNOR2_X1 port map( A => n19644, B => n19585, ZN => n19586);
   U22602 : XNOR2_X1 port map( A => n19586, B => n19587, ZN => n19588);
   U22603 : XNOR2_X1 port map( A => n19592, B => n28693, ZN => n19593);
   U22604 : NOR2_X1 port map( A1 => n20109, A2 => n20319, ZN => n19602);
   U22605 : XNOR2_X1 port map( A => n19595, B => n3083, ZN => n19596);
   U22606 : XNOR2_X1 port map( A => n19597, B => n19596, ZN => n19601);
   U22607 : XNOR2_X1 port map( A => n19599, B => n19598, ZN => n19600);
   U22608 : MUX2_X1 port map( A => n20323, B => n19602, S => n20322, Z => 
                           n20694);
   U22609 : XNOR2_X1 port map( A => n18638, B => n19603, ZN => n19605);
   U22610 : XNOR2_X1 port map( A => n19605, B => n19604, ZN => n19610);
   U22611 : XNOR2_X1 port map( A => n19606, B => n2996, ZN => n19608);
   U22612 : XNOR2_X1 port map( A => n19607, B => n19608, ZN => n19609);
   U22613 : XNOR2_X2 port map( A => n19609, B => n19610, ZN => n20324);
   U22614 : INV_X1 port map( A => n19611, ZN => n19612);
   U22615 : XNOR2_X1 port map( A => n19612, B => n19669, ZN => n19614);
   U22616 : XNOR2_X1 port map( A => n19614, B => n19613, ZN => n19621);
   U22617 : XNOR2_X1 port map( A => n19616, B => n19615, ZN => n19619);
   U22618 : XNOR2_X1 port map( A => n19617, B => n2403, ZN => n19618);
   U22619 : XNOR2_X1 port map( A => n19619, B => n19618, ZN => n19620);
   U22620 : XNOR2_X1 port map( A => n19620, B => n19621, ZN => n19955);
   U22621 : INV_X1 port map( A => n19955, ZN => n19956);
   U22622 : NAND3_X1 port map( A1 => n19956, A2 => n20320, A3 => n2180, ZN => 
                           n20693);
   U22623 : NOR2_X1 port map( A1 => n21809, A2 => n21810, ZN => n21007);
   U22624 : XNOR2_X1 port map( A => n19622, B => n3109, ZN => n19623);
   U22625 : XNOR2_X1 port map( A => n19624, B => n19623, ZN => n19630);
   U22626 : XNOR2_X1 port map( A => n19625, B => n19626, ZN => n19627);
   U22627 : XOR2_X1 port map( A => n19628, B => n19627, Z => n19629);
   U22628 : XNOR2_X1 port map( A => n19630, B => n19629, ZN => n19810);
   U22629 : XNOR2_X1 port map( A => n19636, B => n3695, ZN => n19638);
   U22630 : XNOR2_X1 port map( A => n19638, B => n19637, ZN => n19640);
   U22631 : XNOR2_X1 port map( A => n19640, B => n19639, ZN => n19642);
   U22632 : XNOR2_X1 port map( A => n19642, B => n19641, ZN => n19938);
   U22634 : MUX2_X1 port map( A => n29166, B => n29707, S => n20281, Z => 
                           n19677);
   U22635 : XNOR2_X1 port map( A => n19643, B => n1928, ZN => n19645);
   U22636 : XNOR2_X1 port map( A => n19645, B => n19644, ZN => n19647);
   U22637 : XNOR2_X1 port map( A => n19647, B => n19646, ZN => n19648);
   U22638 : INV_X1 port map( A => n19650, ZN => n19652);
   U22639 : INV_X1 port map( A => n28516, ZN => n19654);
   U22640 : XNOR2_X1 port map( A => n19655, B => n19654, ZN => n19663);
   U22641 : INV_X1 port map( A => n19659, ZN => n19657);
   U22642 : NAND2_X1 port map( A1 => n19657, A2 => n3386, ZN => n19661);
   U22643 : OAI21_X1 port map( B1 => n19656, B2 => n19659, A => n19658, ZN => 
                           n19660);
   U22644 : OAI21_X1 port map( B1 => n19656, B2 => n19661, A => n19660, ZN => 
                           n19662);
   U22645 : XNOR2_X1 port map( A => n19663, B => n19662, ZN => n19664);
   U22646 : INV_X1 port map( A => n19665, ZN => n19667);
   U22647 : XNOR2_X1 port map( A => n19667, B => n19666, ZN => n19674);
   U22648 : XNOR2_X1 port map( A => n19668, B => n19669, ZN => n19672);
   U22649 : XNOR2_X1 port map( A => n29554, B => n28327, ZN => n19671);
   U22650 : XNOR2_X1 port map( A => n19672, B => n19671, ZN => n19673);
   U22651 : INV_X1 port map( A => n20283, ZN => n20285);
   U22652 : NAND2_X1 port map( A1 => n20285, A2 => n20281, ZN => n19675);
   U22653 : NAND2_X1 port map( A1 => n20289, A2 => n19675, ZN => n19676);
   U22654 : XNOR2_X1 port map( A => n19678, B => n3223, ZN => n19680);
   U22655 : XNOR2_X1 port map( A => n19680, B => n19679, ZN => n19682);
   U22656 : XNOR2_X1 port map( A => n19682, B => n19681, ZN => n19684);
   U22658 : INV_X1 port map( A => n20440, ZN => n20608);
   U22659 : XNOR2_X1 port map( A => n19691, B => n19692, ZN => n19694);
   U22660 : XNOR2_X1 port map( A => n19695, B => n19696, ZN => n19699);
   U22661 : XNOR2_X1 port map( A => n19697, B => n3527, ZN => n19698);
   U22662 : MUX2_X1 port map( A => n29625, B => n20608, S => n20441, Z => 
                           n19731);
   U22663 : XNOR2_X1 port map( A => n19701, B => n19700, ZN => n19703);
   U22664 : XNOR2_X1 port map( A => n19703, B => n19702, ZN => n19713);
   U22665 : INV_X1 port map( A => n19704, ZN => n19705);
   U22666 : XNOR2_X1 port map( A => n19706, B => n19705, ZN => n19711);
   U22667 : XNOR2_X1 port map( A => n19707, B => n2510, ZN => n19708);
   U22668 : XNOR2_X1 port map( A => n19708, B => n19709, ZN => n19710);
   U22669 : XNOR2_X1 port map( A => n19710, B => n19711, ZN => n19712);
   U22670 : XNOR2_X1 port map( A => n19712, B => n19713, ZN => n20609);
   U22672 : XNOR2_X1 port map( A => n19714, B => n19715, ZN => n19722);
   U22673 : XNOR2_X1 port map( A => n19716, B => n19717, ZN => n19720);
   U22674 : XNOR2_X1 port map( A => n19718, B => n2353, ZN => n19719);
   U22675 : XNOR2_X1 port map( A => n19720, B => n19719, ZN => n19721);
   U22676 : XNOR2_X1 port map( A => n19726, B => n28571, ZN => n19729);
   U22677 : XNOR2_X1 port map( A => n19727, B => n1062, ZN => n19728);
   U22678 : XNOR2_X1 port map( A => n19729, B => n19728, ZN => n19730);
   U22679 : NOR2_X1 port map( A1 => n21811, A2 => n21253, ZN => n20698);
   U22680 : OAI211_X2 port map( C1 => n21007, C2 => n19735, A => n19734, B => 
                           n19733, ZN => n22295);
   U22681 : XNOR2_X1 port map( A => n22295, B => n1133, ZN => n19736);
   U22682 : XNOR2_X1 port map( A => n21756, B => n19736, ZN => n19737);
   U22683 : MUX2_X1 port map( A => n19739, B => n20377, S => n351, Z => n19742)
                           ;
   U22684 : MUX2_X1 port map( A => n20371, B => n20373, S => n20372, Z => 
                           n19741);
   U22685 : INV_X1 port map( A => n20401, ZN => n20558);
   U22686 : INV_X1 port map( A => n20208, ZN => n20400);
   U22687 : OAI21_X1 port map( B1 => n20558, B2 => n29041, A => n20209, ZN => 
                           n19746);
   U22688 : NAND2_X1 port map( A1 => n20394, A2 => n20563, ZN => n19744);
   U22689 : INV_X1 port map( A => n19851, ZN => n20562);
   U22690 : MUX2_X1 port map( A => n19744, B => n19743, S => n20562, Z => 
                           n19745);
   U22691 : INV_X1 port map( A => n19747, ZN => n20417);
   U22693 : NAND2_X1 port map( A1 => n20412, A2 => n20414, ZN => n19749);
   U22694 : NAND2_X1 port map( A1 => n503, A2 => n20577, ZN => n19748);
   U22695 : INV_X1 port map( A => n22140, ZN => n22142);
   U22696 : MUX2_X1 port map( A => n20383, B => n19837, S => n20567, Z => 
                           n19751);
   U22697 : INV_X1 port map( A => n19836, ZN => n19750);
   U22698 : INV_X1 port map( A => n28526, ZN => n19844);
   U22699 : NOR2_X1 port map( A1 => n18837, A2 => n19844, ZN => n19754);
   U22700 : OAI211_X1 port map( C1 => n6495, C2 => n29551, A => n29582, B => 
                           n20083, ZN => n19753);
   U22701 : INV_X1 port map( A => n20041, ZN => n20092);
   U22702 : NAND2_X1 port map( A1 => n20092, A2 => n414, ZN => n19756);
   U22703 : AOI21_X1 port map( B1 => n19756, B2 => n19755, A => n20039, ZN => 
                           n19759);
   U22704 : NAND2_X1 port map( A1 => n20041, A2 => n29114, ZN => n19757);
   U22705 : MUX2_X1 port map( A => n29540, B => n22145, S => n22143, Z => 
                           n19760);
   U22706 : NAND2_X1 port map( A1 => n29540, A2 => n6532, ZN => n21626);
   U22707 : NAND2_X1 port map( A1 => n20069, A2 => n20049, ZN => n19762);
   U22708 : NAND3_X1 port map( A1 => n20048, A2 => n18765, A3 => n20049, ZN => 
                           n19763);
   U22709 : INV_X1 port map( A => n19766, ZN => n20146);
   U22710 : NOR2_X1 port map( A1 => n20146, A2 => n28479, ZN => n19767);
   U22711 : AOI22_X1 port map( A1 => n20146, A2 => n29134, B1 => n19767, B2 => 
                           n20144, ZN => n19768);
   U22713 : INV_X1 port map( A => n20158, ZN => n20160);
   U22716 : OAI21_X1 port map( B1 => n20163, B2 => n19769, A => n28187, ZN => 
                           n19772);
   U22717 : AOI21_X1 port map( B1 => n19984, B2 => n20162, A => n20159, ZN => 
                           n19770);
   U22718 : OR2_X1 port map( A1 => n19770, A2 => n20158, ZN => n19771);
   U22719 : OAI21_X1 port map( B1 => n28188, B2 => n19773, A => n20043, ZN => 
                           n19774);
   U22720 : OAI21_X1 port map( B1 => n20092, B2 => n29114, A => n20093, ZN => 
                           n19777);
   U22722 : NOR2_X1 port map( A1 => n20851, A2 => n21143, ZN => n19783);
   U22723 : AND2_X1 port map( A1 => n21118, A2 => n21143, ZN => n19782);
   U22724 : XNOR2_X1 port map( A => n22194, B => n22784, ZN => n19805);
   U22725 : INV_X1 port map( A => n20349, ZN => n19785);
   U22726 : NOR2_X1 port map( A1 => n20013, A2 => n20342, ZN => n19786);
   U22727 : INV_X1 port map( A => n20017, ZN => n20345);
   U22728 : INV_X1 port map( A => n20343, ZN => n20014);
   U22729 : NOR2_X1 port map( A1 => n20247, A2 => n20453, ZN => n19788);
   U22731 : OAI21_X1 port map( B1 => n19788, B2 => n20032, A => n20637, ZN => 
                           n19790);
   U22732 : NAND2_X1 port map( A1 => n20247, A2 => n28538, ZN => n19789);
   U22734 : INV_X1 port map( A => n20481, ZN => n20001);
   U22735 : NAND2_X1 port map( A1 => n19793, A2 => n28155, ZN => n19803);
   U22736 : INV_X1 port map( A => n21356, ZN => n20023);
   U22738 : AND2_X1 port map( A1 => n28610, A2 => n21355, ZN => n20024);
   U22739 : INV_X1 port map( A => n21359, ZN => n21354);
   U22740 : NAND2_X1 port map( A1 => n21354, A2 => n19796, ZN => n19797);
   U22741 : OAI21_X1 port map( B1 => n20024, B2 => n21354, A => n19797, ZN => 
                           n19798);
   U22742 : NOR2_X1 port map( A1 => n20498, A2 => n20499, ZN => n19800);
   U22744 : NAND2_X1 port map( A1 => n20333, A2 => n20334, ZN => n20631);
   U22745 : INV_X1 port map( A => n20625, ZN => n20628);
   U22746 : INV_X1 port map( A => n20626, ZN => n20330);
   U22747 : NAND3_X1 port map( A1 => n20628, A2 => n20005, A3 => n20330, ZN => 
                           n19802);
   U22748 : XNOR2_X1 port map( A => n28449, B => n27605, ZN => n19804);
   U22749 : XNOR2_X1 port map( A => n19805, B => n19804, ZN => n19909);
   U22750 : INV_X1 port map( A => n20201, ZN => n20305);
   U22751 : MUX2_X1 port map( A => n20202, B => n20305, S => n20200, Z => 
                           n19807);
   U22752 : NOR2_X1 port map( A1 => n416, A2 => n20200, ZN => n19806);
   U22753 : NAND2_X1 port map( A1 => n20205, A2 => n20302, ZN => n20306);
   U22754 : NAND2_X1 port map( A1 => n19810, A2 => n20284, ZN => n19939);
   U22755 : INV_X1 port map( A => n19939, ZN => n19809);
   U22756 : OAI21_X1 port map( B1 => n2081, B2 => n19809, A => n2152, ZN => 
                           n19813);
   U22757 : INV_X1 port map( A => n19810, ZN => n20286);
   U22758 : AOI21_X1 port map( B1 => n20281, B2 => n20284, A => n20286, ZN => 
                           n19811);
   U22759 : NAND2_X1 port map( A1 => n19967, A2 => n20123, ZN => n20292);
   U22760 : INV_X1 port map( A => n19815, ZN => n19968);
   U22761 : OAI22_X1 port map( A1 => n20292, A2 => n19818, B1 => n19967, B2 => 
                           n20122, ZN => n19817);
   U22762 : AND2_X1 port map( A1 => n19818, A2 => n19815, ZN => n20124);
   U22763 : INV_X1 port map( A => n20124, ZN => n19816);
   U22765 : INV_X1 port map( A => n20546, ZN => n20191);
   U22766 : NOR2_X1 port map( A1 => n19820, A2 => n20389, ZN => n19819);
   U22767 : AND2_X1 port map( A1 => n20544, A2 => n20546, ZN => n20190);
   U22768 : OAI21_X1 port map( B1 => n20190, B2 => n20388, A => n19820, ZN => 
                           n19821);
   U22769 : INV_X1 port map( A => n20319, ZN => n19940);
   U22770 : NAND2_X1 port map( A1 => n19940, A2 => n20323, ZN => n19822);
   U22771 : MUX2_X1 port map( A => n19822, B => n20112, S => n20324, Z => 
                           n19826);
   U22772 : NOR2_X1 port map( A1 => n20323, A2 => n20320, ZN => n19824);
   U22773 : NOR2_X1 port map( A1 => n19940, A2 => n20322, ZN => n19823);
   U22774 : AOI22_X1 port map( A1 => n19824, A2 => n19940, B1 => n19823, B2 => 
                           n502, ZN => n19825);
   U22775 : NAND2_X1 port map( A1 => n20311, A2 => n19949, ZN => n19829);
   U22776 : INV_X1 port map( A => n20196, ZN => n20588);
   U22777 : OR2_X1 port map( A1 => n21495, A2 => n21496, ZN => n19830);
   U22778 : NAND2_X1 port map( A1 => n19834, A2 => n19838, ZN => n19839);
   U22779 : OAI211_X1 port map( C1 => n20379, C2 => n20373, A => n351, B => 
                           n20374, ZN => n19842);
   U22780 : OAI21_X1 port map( B1 => n6495, B2 => n20083, A => n29582, ZN => 
                           n19848);
   U22781 : NOR2_X1 port map( A1 => n6495, A2 => n19844, ZN => n19846);
   U22782 : AND2_X1 port map( A1 => n19851, A2 => n20208, ZN => n20396);
   U22783 : NAND2_X1 port map( A1 => n20401, A2 => n20396, ZN => n19854);
   U22784 : INV_X1 port map( A => n19849, ZN => n19850);
   U22785 : NAND3_X1 port map( A1 => n20209, A2 => n20562, A3 => n20563, ZN => 
                           n19852);
   U22786 : NAND2_X1 port map( A1 => n20749, A2 => n21574, ZN => n21487);
   U22787 : MUX2_X1 port map( A => n20941, B => n20577, S => n28140, Z => 
                           n19858);
   U22789 : XNOR2_X1 port map( A => n22661, B => n21758, ZN => n22575);
   U22790 : INV_X1 port map( A => n22575, ZN => n19907);
   U22793 : OAI21_X1 port map( B1 => n5303, B2 => n29616, A => n20218, ZN => 
                           n19864);
   U22794 : OAI21_X1 port map( B1 => n19865, B2 => n20218, A => n19864, ZN => 
                           n19866);
   U22795 : INV_X1 port map( A => n21155, ZN => n21158);
   U22796 : NAND2_X1 port map( A1 => n19032, A2 => n382, ZN => n20737);
   U22797 : INV_X1 port map( A => n20176, ZN => n20054);
   U22798 : NOR2_X1 port map( A1 => n19868, A2 => n20171, ZN => n19869);
   U22800 : INV_X1 port map( A => n20144, ZN => n20106);
   U22801 : NAND2_X1 port map( A1 => n20527, A2 => n20858, ZN => n19871);
   U22802 : INV_X1 port map( A => n20159, ZN => n19981);
   U22803 : MUX2_X1 port map( A => n20160, B => n20157, S => n19981, Z => 
                           n19876);
   U22804 : NOR2_X1 port map( A1 => n19981, A2 => n29066, ZN => n19873);
   U22805 : AOI22_X1 port map( A1 => n19874, A2 => n19873, B1 => n19985, B2 => 
                           n19872, ZN => n19875);
   U22806 : NAND2_X1 port map( A1 => n494, A2 => n21159, ZN => n21111);
   U22808 : OAI21_X1 port map( B1 => n21111, B2 => n20858, A => n19877, ZN => 
                           n19878);
   U22809 : NOR2_X2 port map( A1 => n19879, A2 => n19878, ZN => n22218);
   U22810 : NAND2_X1 port map( A1 => n20603, A2 => n1915, ZN => n19880);
   U22811 : NOR2_X1 port map( A1 => n20601, A2 => n20272, ZN => n19883);
   U22812 : NOR2_X1 port map( A1 => n20603, A2 => n20272, ZN => n19882);
   U22813 : NOR3_X1 port map( A1 => n19882, A2 => n28408, A3 => n19883, ZN => 
                           n19884);
   U22814 : NOR2_X1 port map( A1 => n19886, A2 => n20607, ZN => n19888);
   U22815 : INV_X1 port map( A => n20618, ZN => n19889);
   U22816 : AOI21_X1 port map( B1 => n19889, B2 => n6567, A => n20616, ZN => 
                           n19891);
   U22820 : NOR2_X1 port map( A1 => n20622, A2 => n19920, ZN => n19893);
   U22821 : NOR2_X1 port map( A1 => n20137, A2 => n19808, ZN => n19895);
   U22823 : NOR2_X1 port map( A1 => n20281, A2 => n20137, ZN => n19897);
   U22824 : NOR2_X1 port map( A1 => n20449, A2 => n20265, ZN => n20450);
   U22825 : NAND2_X1 port map( A1 => n20450, A2 => n5377, ZN => n19900);
   U22826 : AOI211_X1 port map( C1 => n415, C2 => n20444, A => n3247, B => 
                           n19901, ZN => n19902);
   U22827 : INV_X1 port map( A => n21459, ZN => n20842);
   U22828 : NAND2_X1 port map( A1 => n1814, A2 => n20842, ZN => n19904);
   U22830 : XNOR2_X1 port map( A => n22218, B => n22279, ZN => n19906);
   U22831 : XNOR2_X1 port map( A => n19907, B => n19906, ZN => n19908);
   U22832 : NOR2_X1 port map( A1 => n23535, A2 => n23529, ZN => n20473);
   U22833 : NAND2_X1 port map( A1 => n22139, A2 => n22145, ZN => n21029);
   U22834 : INV_X1 port map( A => n29540, ZN => n22146);
   U22835 : NAND3_X1 port map( A1 => n22146, A2 => n22139, A3 => n22143, ZN => 
                           n19911);
   U22836 : NOR2_X1 port map( A1 => n5939, A2 => n22139, ZN => n21623);
   U22838 : MUX2_X1 port map( A => n20972, B => n21217, S => n21000, Z => 
                           n19912);
   U22839 : NOR2_X1 port map( A1 => n19912, A2 => n21220, ZN => n19918);
   U22841 : NAND2_X1 port map( A1 => n28980, A2 => n21218, ZN => n19916);
   U22842 : NAND2_X1 port map( A1 => n20966, A2 => n19914, ZN => n20701);
   U22843 : OAI21_X1 port map( B1 => n19916, B2 => n20701, A => n19915, ZN => 
                           n19917);
   U22844 : XNOR2_X1 port map( A => n21875, B => n22330, ZN => n19945);
   U22845 : NAND3_X1 port map( A1 => n20255, A2 => n28894, A3 => n20616, ZN => 
                           n19919);
   U22846 : OAI21_X1 port map( B1 => n19901, B2 => n20443, A => n19924, ZN => 
                           n19925);
   U22847 : INV_X1 port map( A => n21748, ZN => n21401);
   U22849 : NAND2_X1 port map( A1 => n28555, A2 => n20440, ZN => n19935);
   U22850 : NAND3_X1 port map( A1 => n20441, A2 => n29508, A3 => n20607, ZN => 
                           n19937);
   U22851 : NAND2_X1 port map( A1 => n21642, A2 => n20658, ZN => n21040);
   U22852 : AOI22_X1 port map( A1 => n502, A2 => n20109, B1 => n20323, B2 => 
                           n20322, ZN => n19942);
   U22853 : AND2_X1 port map( A1 => n20109, A2 => n19955, ZN => n20325);
   U22854 : OAI21_X1 port map( B1 => n20325, B2 => n19940, A => n2181, ZN => 
                           n19941);
   U22856 : NAND2_X1 port map( A1 => n20659, A2 => n497, ZN => n19943);
   U22857 : XNOR2_X1 port map( A => n22265, B => n2960, ZN => n19944);
   U22858 : XNOR2_X1 port map( A => n19945, B => n19944, ZN => n20062);
   U22859 : NOR2_X1 port map( A1 => n20205, A2 => n20302, ZN => n19946);
   U22860 : INV_X1 port map( A => n20302, ZN => n20119);
   U22861 : NOR2_X1 port map( A1 => n19949, A2 => n20584, ZN => n19950);
   U22862 : INV_X1 port map( A => n20585, ZN => n20315);
   U22863 : MUX2_X1 port map( A => n20315, B => n20196, S => n20314, Z => 
                           n19952);
   U22864 : NOR2_X1 port map( A1 => n19952, A2 => n3973, ZN => n19953);
   U22865 : NOR2_X1 port map( A1 => n21472, A2 => n1930, ZN => n21733);
   U22866 : NAND2_X1 port map( A1 => n502, A2 => n20319, ZN => n19957);
   U22867 : OAI21_X1 port map( B1 => n20546, B2 => n20544, A => n20188, ZN => 
                           n19961);
   U22868 : AOI22_X2 port map( A1 => n20392, A2 => n19961, B1 => n19960, B2 => 
                           n19959, ZN => n21473);
   U22869 : MUX2_X1 port map( A => n21733, B => n21388, S => n21473, Z => 
                           n19975);
   U22870 : INV_X1 port map( A => n19962, ZN => n19966);
   U22871 : INV_X1 port map( A => n20405, ZN => n20553);
   U22872 : NOR2_X1 port map( A1 => n20556, A2 => n20553, ZN => n19964);
   U22873 : OAI21_X1 port map( B1 => n19964, B2 => n20404, A => n505, ZN => 
                           n21032);
   U22874 : OAI21_X1 port map( B1 => n19968, B2 => n20125, A => n19967, ZN => 
                           n19972);
   U22875 : NOR2_X1 port map( A1 => n19969, A2 => n20295, ZN => n19970);
   U22877 : OAI21_X1 port map( B1 => n21471, B2 => n21731, A => n21477, ZN => 
                           n19974);
   U22878 : INV_X1 port map( A => n20055, ZN => n19980);
   U22879 : MUX2_X1 port map( A => n20178, B => n20173, S => n19976, Z => 
                           n19978);
   U22880 : MUX2_X1 port map( A => n19978, B => n19977, S => n20054, Z => 
                           n19979);
   U22881 : OAI21_X1 port map( B1 => n19982, B2 => n19981, A => n20164, ZN => 
                           n19988);
   U22882 : AOI21_X1 port map( B1 => n19985, B2 => n19984, A => n19983, ZN => 
                           n20047);
   U22884 : NOR2_X1 port map( A1 => n297, A2 => n19989, ZN => n19990);
   U22885 : NOR2_X1 port map( A1 => n385, A2 => n19992, ZN => n19994);
   U22886 : OAI211_X1 port map( C1 => n20479, C2 => n19997, A => n20475, B => 
                           n383, ZN => n19999);
   U22887 : NAND2_X1 port map( A1 => n5408, A2 => n20478, ZN => n19996);
   U22888 : NOR2_X1 port map( A1 => n19996, A2 => n20477, ZN => n19998);
   U22889 : NOR2_X1 port map( A1 => n28620, A2 => n20000, ZN => n20002);
   U22890 : AOI22_X1 port map( A1 => n20002, A2 => n20001, B1 => n29527, B2 => 
                           n20485, ZN => n20004);
   U22891 : XNOR2_X1 port map( A => n21956, B => n22633, ZN => n20060);
   U22893 : INV_X1 port map( A => n20623, ZN => n20258);
   U22895 : NOR2_X1 port map( A1 => n28515, A2 => n20012, ZN => n20670);
   U22896 : NOR3_X1 port map( A1 => n20675, A2 => n21638, A3 => n20670, ZN => 
                           n20031);
   U22897 : INV_X1 port map( A => n20013, ZN => n20344);
   U22898 : MUX2_X1 port map( A => n28489, B => n19785, S => n20344, Z => 
                           n20016);
   U22899 : NOR2_X1 port map( A1 => n20345, A2 => n20342, ZN => n20015);
   U22900 : INV_X1 port map( A => n20347, ZN => n20019);
   U22901 : NAND2_X1 port map( A1 => n20511, A2 => n20349, ZN => n20018);
   U22902 : NOR2_X1 port map( A1 => n20019, A2 => n20018, ZN => n20671);
   U22903 : NOR2_X2 port map( A1 => n20669, A2 => n20671, ZN => n21639);
   U22905 : MUX2_X1 port map( A => n20518, B => n20021, S => n21359, Z => 
                           n20026);
   U22906 : NOR2_X1 port map( A1 => n28610, A2 => n28491, ZN => n20022);
   U22907 : AOI22_X1 port map( A1 => n20024, A2 => n20023, B1 => n20022, B2 => 
                           n28586, ZN => n20025);
   U22908 : NAND3_X1 port map( A1 => n386, A2 => n20603, A3 => n20028, ZN => 
                           n20029);
   U22909 : AND2_X1 port map( A1 => n20033, A2 => n20453, ZN => n20252);
   U22912 : NOR2_X1 port map( A1 => n21092, A2 => n20146, ZN => n20038);
   U22913 : NOR2_X1 port map( A1 => n21091, A2 => n21095, ZN => n20036);
   U22914 : AOI22_X1 port map( A1 => n20038, A2 => n20148, B1 => n20036, B2 => 
                           n18919, ZN => n20037);
   U22916 : NAND3_X1 port map( A1 => n20045, A2 => n20158, A3 => n20044, ZN => 
                           n20046);
   U22917 : OAI21_X1 port map( B1 => n20047, B2 => n20163, A => n20046, ZN => 
                           n21211);
   U22919 : NAND2_X1 port map( A1 => n20052, A2 => n28448, ZN => n21209);
   U22920 : INV_X1 port map( A => n20053, ZN => n20056);
   U22921 : NAND3_X1 port map( A1 => n20056, A2 => n504, A3 => n20173, ZN => 
                           n20057);
   U22922 : XNOR2_X1 port map( A => n22643, B => n22690, ZN => n20059);
   U22923 : XNOR2_X1 port map( A => n20060, B => n20059, ZN => n20061);
   U22924 : MUX2_X1 port map( A => n20065, B => n20064, S => n20063, Z => 
                           n20067);
   U22925 : OAI21_X1 port map( B1 => n351, B2 => n20374, A => n20377, ZN => 
                           n20072);
   U22926 : NAND2_X1 port map( A1 => n20372, A2 => n20072, ZN => n20073);
   U22927 : INV_X1 port map( A => n20075, ZN => n20079);
   U22928 : NOR2_X1 port map( A1 => n18837, A2 => n29315, ZN => n20078);
   U22930 : NOR2_X1 port map( A1 => n20081, A2 => n29551, ZN => n20082);
   U22931 : AOI22_X1 port map( A1 => n20084, A2 => n20083, B1 => n20082, B2 => 
                           n18837, ZN => n20085);
   U22932 : NOR2_X1 port map( A1 => n22013, A2 => n20532, ZN => n21818);
   U22933 : NOR2_X1 port map( A1 => n20155, A2 => n20096, ZN => n20101);
   U22934 : NAND2_X1 port map( A1 => n20097, A2 => n18887, ZN => n20100);
   U22935 : NAND2_X1 port map( A1 => n21078, A2 => n495, ZN => n20108);
   U22936 : NAND2_X1 port map( A1 => n18919, A2 => n20102, ZN => n20107);
   U22937 : AOI21_X1 port map( B1 => n29134, B2 => n20102, A => n21091, ZN => 
                           n20104);
   U22938 : NOR2_X1 port map( A1 => n18919, A2 => n28479, ZN => n20103);
   U22939 : OAI22_X1 port map( A1 => n20104, A2 => n20103, B1 => n20102, B2 => 
                           n4877, ZN => n20105);
   U22940 : NOR2_X1 port map( A1 => n20320, A2 => n20319, ZN => n20110);
   U22941 : NOR2_X1 port map( A1 => n20112, A2 => n20324, ZN => n20897);
   U22942 : NOR2_X1 port map( A1 => n20607, A2 => n20440, ZN => n20113);
   U22943 : NOR2_X1 port map( A1 => n20113, A2 => n20441, ZN => n20116);
   U22944 : NOR2_X1 port map( A1 => n20441, A2 => n20440, ZN => n20114);
   U22945 : NOR2_X1 port map( A1 => n20609, A2 => n29508, ZN => n20435);
   U22946 : OAI21_X1 port map( B1 => n20114, B2 => n20435, A => n20614, ZN => 
                           n20115);
   U22947 : INV_X1 port map( A => n20898, ZN => n20129);
   U22948 : INV_X1 port map( A => n20897, ZN => n20118);
   U22949 : OAI21_X1 port map( B1 => n20295, B2 => n20123, A => n20122, ZN => 
                           n20127);
   U22950 : NAND2_X1 port map( A1 => n20125, A2 => n20124, ZN => n20126);
   U22951 : INV_X1 port map( A => n20299, ZN => n20131);
   U22952 : NOR2_X1 port map( A1 => n20131, A2 => n20130, ZN => n20132);
   U22953 : NOR2_X1 port map( A1 => n20446, A2 => n20132, ZN => n20134);
   U22954 : NAND3_X1 port map( A1 => n19938, A2 => n19808, A3 => n20286, ZN => 
                           n20136);
   U22955 : NAND2_X1 port map( A1 => n20141, A2 => n20140, ZN => n20142);
   U22956 : XNOR2_X1 port map( A => n22098, B => n22270, ZN => n20215);
   U22957 : NOR2_X1 port map( A1 => n29134, A2 => n20144, ZN => n21096);
   U22958 : NAND2_X1 port map( A1 => n20149, A2 => n20148, ZN => n21097);
   U22959 : INV_X1 port map( A => n21097, ZN => n20953);
   U22960 : AOI21_X1 port map( B1 => n20152, B2 => n20151, A => n20150, ZN => 
                           n20153);
   U22961 : NOR3_X1 port map( A1 => n20954, A2 => n20953, A3 => n21932, ZN => 
                           n20187);
   U22962 : NOR2_X1 port map( A1 => n20165, A2 => n385, ZN => n20170);
   U22963 : AND3_X1 port map( A1 => n20166, A2 => n297, A3 => n20219, ZN => 
                           n20167);
   U22964 : NOR2_X1 port map( A1 => n20168, A2 => n20167, ZN => n20169);
   U22965 : INV_X1 port map( A => n21089, ZN => n20802);
   U22966 : NOR2_X1 port map( A1 => n504, A2 => n20173, ZN => n20175);
   U22967 : NAND2_X1 port map( A1 => n20786, A2 => n21932, ZN => n20951);
   U22968 : NAND2_X1 port map( A1 => n20494, A2 => n20179, ZN => n20181);
   U22969 : NAND2_X1 port map( A1 => n21090, A2 => n21089, ZN => n20466);
   U22970 : NAND2_X1 port map( A1 => n20191, A2 => n20539, ZN => n20189);
   U22971 : INV_X1 port map( A => n20388, ZN => n20541);
   U22973 : NAND2_X1 port map( A1 => n28779, A2 => n20416, ZN => n20823);
   U22974 : NAND2_X1 port map( A1 => n20823, A2 => n20418, ZN => n20195);
   U22975 : NAND2_X1 port map( A1 => n20192, A2 => n20193, ZN => n20821);
   U22976 : NAND2_X1 port map( A1 => n20193, A2 => n20580, ZN => n20194);
   U22977 : NOR2_X1 port map( A1 => n20413, A2 => n20194, ZN => n20824);
   U22978 : NAND2_X1 port map( A1 => n21675, A2 => n21677, ZN => n21447);
   U22979 : MUX2_X1 port map( A => n20585, B => n20311, S => n29144, Z => 
                           n20198);
   U22980 : NOR2_X1 port map( A1 => n20585, A2 => n20196, ZN => n20586);
   U22981 : NOR2_X1 port map( A1 => n20315, A2 => n20314, ZN => n20197);
   U22982 : AND2_X1 port map( A1 => n20199, A2 => n20201, ZN => n20303);
   U22983 : OAI21_X1 port map( B1 => n6935, B2 => n20202, A => n416, ZN => 
                           n20203);
   U22985 : OAI21_X1 port map( B1 => n20558, B2 => n20208, A => n20560, ZN => 
                           n20211);
   U22986 : OAI21_X1 port map( B1 => n20209, B2 => n20563, A => n20562, ZN => 
                           n20210);
   U22989 : OAI22_X1 port map( A1 => n21448, A2 => n21678, B1 => n21677, B2 => 
                           n21676, ZN => n21004);
   U22990 : XNOR2_X1 port map( A => n20215, B => n20214, ZN => n20280);
   U22991 : NAND3_X1 port map( A1 => n29488, A2 => n20878, A3 => n20875, ZN => 
                           n20216);
   U22992 : XNOR2_X1 port map( A => n28483, B => n1193, ZN => n20278);
   U22993 : INV_X1 port map( A => n21655, ZN => n21074);
   U22994 : NAND2_X1 port map( A1 => n20498, A2 => n20504, ZN => n20229);
   U22995 : NAND2_X1 port map( A1 => n20226, A2 => n20503, ZN => n20228);
   U22997 : NAND2_X1 port map( A1 => n20480, A2 => n20475, ZN => n20231);
   U22998 : OAI211_X1 port map( C1 => n21074, C2 => n6275, A => n21442, B => 
                           n21654, ZN => n20246);
   U22999 : INV_X1 port map( A => n20511, ZN => n20235);
   U23000 : AOI21_X1 port map( B1 => n20345, B2 => n20235, A => n20349, ZN => 
                           n20234);
   U23001 : NOR2_X1 port map( A1 => n20014, A2 => n20510, ZN => n20233);
   U23002 : OAI22_X1 port map( A1 => n20234, A2 => n20233, B1 => n20344, B2 => 
                           n20235, ZN => n20237);
   U23003 : NAND3_X1 port map( A1 => n20235, A2 => n20342, A3 => n20510, ZN => 
                           n20236);
   U23004 : AND2_X2 port map( A1 => n20237, A2 => n20236, ZN => n21653);
   U23005 : INV_X1 port map( A => n21442, ZN => n21661);
   U23007 : NAND2_X1 port map( A1 => n20488, A2 => n28620, ZN => n20243);
   U23008 : AOI21_X1 port map( B1 => n20240, B2 => n29527, A => n20239, ZN => 
                           n20242);
   U23011 : NOR2_X1 port map( A1 => n20635, A2 => n20637, ZN => n20250);
   U23012 : NOR2_X1 port map( A1 => n20247, A2 => n28538, ZN => n20249);
   U23013 : MUX2_X1 port map( A => n20250, B => n20249, S => n20248, Z => 
                           n20254);
   U23014 : OAI21_X1 port map( B1 => n20636, B2 => n20453, A => n20635, ZN => 
                           n20251);
   U23017 : NOR2_X1 port map( A1 => n22402, A2 => n21429, ZN => n20271);
   U23018 : NOR2_X1 port map( A1 => n20630, A2 => n20334, ZN => n20259);
   U23019 : NAND2_X1 port map( A1 => n28515, A2 => n20259, ZN => n20260);
   U23020 : NAND2_X1 port map( A1 => n19795, A2 => n21359, ZN => n20329);
   U23021 : AOI21_X1 port map( B1 => n20329, B2 => n20262, A => n20520, ZN => 
                           n20264);
   U23022 : INV_X1 port map( A => n21067, ZN => n20270);
   U23023 : NOR2_X1 port map( A1 => n22397, A2 => n22401, ZN => n20269);
   U23025 : NAND2_X1 port map( A1 => n28552, A2 => n6203, ZN => n21062);
   U23026 : OAI21_X1 port map( B1 => n21061, B2 => n21063, A => n21062, ZN => 
                           n20268);
   U23027 : NAND2_X1 port map( A1 => n20268, A2 => n21065, ZN => n21665);
   U23028 : NOR2_X1 port map( A1 => n28408, A2 => n20275, ZN => n21431);
   U23029 : NOR2_X2 port map( A1 => n21432, A2 => n21431, ZN => n22404);
   U23030 : XNOR2_X1 port map( A => n20277, B => n20278, ZN => n20279);
   U23031 : MUX2_X1 port map( A => n20283, B => n28657, S => n20281, Z => 
                           n20288);
   U23032 : NOR2_X1 port map( A1 => n20285, A2 => n20284, ZN => n20287);
   U23033 : AND2_X1 port map( A1 => n20289, A2 => n2152, ZN => n20766);
   U23034 : NOR2_X2 port map( A1 => n20767, A2 => n20766, ZN => n21304);
   U23035 : NAND2_X1 port map( A1 => n20290, A2 => n20293, ZN => n20291);
   U23036 : NAND2_X1 port map( A1 => n20292, A2 => n20291, ZN => n20297);
   U23037 : AOI21_X1 port map( B1 => n3247, B2 => n19901, A => n20299, ZN => 
                           n20300);
   U23038 : NAND2_X1 port map( A1 => n20303, A2 => n20302, ZN => n20309);
   U23039 : NAND3_X1 port map( A1 => n20306, A2 => n20305, A3 => n20304, ZN => 
                           n20308);
   U23040 : NOR2_X1 port map( A1 => n20587, A2 => n29144, ZN => n20313);
   U23041 : NOR2_X1 port map( A1 => n20311, A2 => n20584, ZN => n20312);
   U23042 : MUX2_X1 port map( A => n20313, B => n20312, S => n20589, Z => 
                           n20318);
   U23043 : NAND2_X1 port map( A1 => n20315, A2 => n20314, ZN => n20316);
   U23044 : OAI22_X1 port map( A1 => n20316, A2 => n20589, B1 => n20588, B2 => 
                           n20584, ZN => n20317);
   U23045 : OAI21_X1 port map( B1 => n21311, B2 => n21309, A => n21307, ZN => 
                           n20326);
   U23046 : NAND2_X1 port map( A1 => n20326, A2 => n20771, ZN => n20327);
   U23048 : NAND2_X1 port map( A1 => n1881, A2 => n20334, ZN => n20332);
   U23050 : OAI21_X1 port map( B1 => n28515, B2 => n20332, A => n20331, ZN => 
                           n20337);
   U23051 : NAND2_X1 port map( A1 => n20335, A2 => n20334, ZN => n20336);
   U23052 : NOR2_X1 port map( A1 => n21550, A2 => n21177, ZN => n20365);
   U23053 : MUX2_X1 port map( A => n20503, B => n20504, S => n20499, Z => 
                           n20338);
   U23055 : NOR2_X1 port map( A1 => n20500, A2 => n20498, ZN => n20340);
   U23056 : MUX2_X1 port map( A => n20343, B => n20342, S => n20344, Z => 
                           n20350);
   U23057 : AOI21_X1 port map( B1 => n20345, B2 => n20344, A => n19785, ZN => 
                           n20346);
   U23058 : OAI21_X1 port map( B1 => n20350, B2 => n20349, A => n20348, ZN => 
                           n20351);
   U23059 : OAI21_X1 port map( B1 => n21549, B2 => n21177, A => n21553, ZN => 
                           n20364);
   U23060 : NOR2_X1 port map( A1 => n20783, A2 => n21177, ZN => n21520);
   U23061 : AOI21_X1 port map( B1 => n20353, B2 => n20352, A => n4557, ZN => 
                           n20357);
   U23062 : OAI22_X1 port map( A1 => n20355, A2 => n20354, B1 => n20480, B2 => 
                           n382, ZN => n20356);
   U23063 : INV_X1 port map( A => n20782, ZN => n21547);
   U23064 : INV_X1 port map( A => n20484, ZN => n20358);
   U23065 : OAI21_X1 port map( B1 => n20488, B2 => n20483, A => n20358, ZN => 
                           n20360);
   U23066 : AOI22_X1 port map( A1 => n20361, A2 => n20360, B1 => n20481, B2 => 
                           n20359, ZN => n21519);
   U23068 : XNOR2_X1 port map( A => n22301, B => n22472, ZN => n20424);
   U23069 : INV_X1 port map( A => n20848, ZN => n20366);
   U23070 : NOR2_X1 port map( A1 => n20366, A2 => n21576, ZN => n20370);
   U23071 : AND2_X1 port map( A1 => n20749, A2 => n21483, ZN => n20367);
   U23072 : AOI22_X1 port map( A1 => n5142, A2 => n20368, B1 => n20367, B2 => 
                           n21575, ZN => n20369);
   U23073 : OAI21_X1 port map( B1 => n5142, B2 => n20370, A => n20369, ZN => 
                           n22116);
   U23074 : MUX2_X1 port map( A => n20372, B => n20371, S => n20373, Z => 
                           n20380);
   U23075 : NOR2_X1 port map( A1 => n20374, A2 => n20373, ZN => n20376);
   U23078 : INV_X1 port map( A => n20571, ZN => n20387);
   U23079 : OAI21_X1 port map( B1 => n20567, B2 => n20381, A => n20383, ZN => 
                           n20386);
   U23080 : INV_X1 port map( A => n20567, ZN => n20382);
   U23082 : NAND2_X1 port map( A1 => n20383, A2 => n97, ZN => n20384);
   U23084 : OAI21_X1 port map( B1 => n29644, B2 => n20389, A => n20388, ZN => 
                           n20390);
   U23085 : NAND2_X1 port map( A1 => n20390, A2 => n20547, ZN => n20391);
   U23088 : NOR2_X1 port map( A1 => n6086, A2 => n505, ZN => n20411);
   U23089 : OAI21_X1 port map( B1 => n20552, B2 => n28501, A => n20404, ZN => 
                           n20410);
   U23090 : MUX2_X1 port map( A => n20408, B => n20407, S => n20551, Z => 
                           n20409);
   U23092 : OAI21_X1 port map( B1 => n21504, B2 => n21499, A => n21503, ZN => 
                           n20422);
   U23093 : INV_X1 port map( A => n20412, ZN => n20413);
   U23094 : INV_X1 port map( A => n20583, ZN => n20415);
   U23095 : NAND2_X1 port map( A1 => n20577, A2 => n20414, ZN => n20939);
   U23096 : MUX2_X1 port map( A => n20415, B => n20939, S => n20941, Z => 
                           n20776);
   U23097 : NAND2_X1 port map( A1 => n20419, A2 => n20823, ZN => n20777);
   U23098 : AOI21_X1 port map( B1 => n20776, B2 => n20777, A => n28619, ZN => 
                           n20420);
   U23099 : OAI21_X1 port map( B1 => n21192, B2 => n20420, A => n21539, ZN => 
                           n20421);
   U23100 : AND2_X1 port map( A1 => n20422, A2 => n20421, ZN => n21949);
   U23101 : INV_X1 port map( A => n21949, ZN => n22327);
   U23102 : XNOR2_X1 port map( A => n22327, B => n22116, ZN => n20423);
   U23103 : XNOR2_X1 port map( A => n20423, B => n20424, ZN => n20472);
   U23104 : NOR2_X1 port map( A1 => n22012, A2 => n20934, ZN => n20427);
   U23107 : NOR2_X1 port map( A1 => n20618, A2 => n20617, ZN => n20429);
   U23108 : INV_X1 port map( A => n20435, ZN => n20439);
   U23109 : NAND2_X1 port map( A1 => n20607, A2 => n20440, ZN => n20438);
   U23110 : INV_X1 port map( A => n20614, ZN => n20436);
   U23111 : NOR2_X1 port map( A1 => n21514, A2 => n21513, ZN => n21531);
   U23112 : AND3_X1 port map( A1 => n20444, A2 => n19901, A3 => n20443, ZN => 
                           n20445);
   U23113 : NOR2_X1 port map( A1 => n20446, A2 => n20445, ZN => n20447);
   U23114 : OAI21_X1 port map( B1 => n20448, B2 => n415, A => n20447, ZN => 
                           n21199);
   U23115 : INV_X1 port map( A => n21199, ZN => n21516);
   U23116 : NOR2_X1 port map( A1 => n21531, A2 => n21516, ZN => n20465);
   U23117 : NAND2_X1 port map( A1 => n20634, A2 => n20453, ZN => n20454);
   U23118 : NOR2_X1 port map( A1 => n21516, A2 => n21513, ZN => n20462);
   U23119 : OR2_X1 port map( A1 => n20597, A2 => n1916, ZN => n20457);
   U23121 : OAI21_X1 port map( B1 => n20463, B2 => n20462, A => n21509, ZN => 
                           n20464);
   U23123 : XNOR2_X1 port map( A => n22302, B => n28162, ZN => n22157);
   U23124 : AND2_X1 port map( A1 => n20951, A2 => n20466, ZN => n20469);
   U23125 : OAI21_X1 port map( B1 => n20955, B2 => n20802, A => n21090, ZN => 
                           n20467);
   U23126 : NAND2_X1 port map( A1 => n20467, A2 => n29586, ZN => n20468);
   U23127 : OAI21_X2 port map( B1 => n21934, B2 => n20469, A => n20468, ZN => 
                           n22601);
   U23128 : XNOR2_X1 port map( A => n22601, B => n2403, ZN => n20470);
   U23129 : MUX2_X1 port map( A => n20473, B => n23136, S => n23531, Z => 
                           n20657);
   U23130 : NAND3_X1 port map( A1 => n20480, A2 => n20479, A3 => n20478, ZN => 
                           n21330);
   U23131 : NAND2_X1 port map( A1 => n20482, A2 => n20481, ZN => n21610);
   U23132 : MUX2_X1 port map( A => n28620, B => n20486, S => n20483, Z => 
                           n20489);
   U23133 : NOR3_X1 port map( A1 => n20486, A2 => n20485, A3 => n20484, ZN => 
                           n20487);
   U23134 : NAND2_X1 port map( A1 => n20496, A2 => n20494, ZN => n20490);
   U23135 : AOI21_X1 port map( B1 => n20491, B2 => n20490, A => n499, ZN => 
                           n20492);
   U23136 : AOI21_X1 port map( B1 => n20503, B2 => n20498, A => n20504, ZN => 
                           n20502);
   U23137 : NAND2_X1 port map( A1 => n20500, A2 => n20499, ZN => n20501);
   U23138 : NAND2_X1 port map( A1 => n20502, A2 => n20501, ZN => n20508);
   U23139 : NAND3_X1 port map( A1 => n1624, A2 => n20504, A3 => n20503, ZN => 
                           n20507);
   U23140 : OAI211_X1 port map( C1 => n20511, C2 => n19785, A => n20510, B => 
                           n20509, ZN => n20512);
   U23142 : NAND3_X1 port map( A1 => n21610, A2 => n21611, A3 => n21612, ZN => 
                           n20515);
   U23143 : NAND2_X1 port map( A1 => n21618, A2 => n20515, ZN => n20516);
   U23144 : NAND2_X1 port map( A1 => n21619, A2 => n20516, ZN => n20524);
   U23145 : NOR2_X1 port map( A1 => n28610, A2 => n28586, ZN => n20521);
   U23146 : AOI22_X1 port map( A1 => n20521, A2 => n20520, B1 => n28133, B2 => 
                           n501, ZN => n20522);
   U23147 : NAND2_X1 port map( A1 => n21326, A2 => n21334, ZN => n20523);
   U23148 : NOR2_X1 port map( A1 => n20744, A2 => n21159, ZN => n20531);
   U23149 : INV_X1 port map( A => n21159, ZN => n20526);
   U23150 : NAND3_X1 port map( A1 => n20526, A2 => n21157, A3 => n21155, ZN => 
                           n20529);
   U23151 : INV_X1 port map( A => n20527, ZN => n20528);
   U23153 : XNOR2_X1 port map( A => n22750, B => n22609, ZN => n22714);
   U23154 : INV_X1 port map( A => n20532, ZN => n22011);
   U23155 : AND2_X1 port map( A1 => n22011, A2 => n22013, ZN => n20537);
   U23156 : NOR2_X1 port map( A1 => n20933, A2 => n21078, ZN => n20535);
   U23157 : NAND2_X1 port map( A1 => n22011, A2 => n20533, ZN => n20534);
   U23160 : MUX2_X1 port map( A => n20546, B => n20547, S => n29644, Z => 
                           n20543);
   U23161 : NOR2_X1 port map( A1 => n6261, A2 => n20539, ZN => n20542);
   U23162 : INV_X1 port map( A => n20544, ZN => n20545);
   U23163 : NOR2_X1 port map( A1 => n21586, A2 => n21585, ZN => n20889);
   U23164 : NAND2_X1 port map( A1 => n20553, A2 => n20549, ZN => n20550);
   U23165 : NAND3_X1 port map( A1 => n20554, A2 => n20553, A3 => n20552, ZN => 
                           n20555);
   U23166 : INV_X1 port map( A => n20559, ZN => n20565);
   U23167 : OAI21_X1 port map( B1 => n20563, B2 => n20562, A => n20561, ZN => 
                           n20564);
   U23168 : NAND2_X1 port map( A1 => n6932, A2 => n97, ZN => n20572);
   U23169 : NAND2_X1 port map( A1 => n20574, A2 => n28508, ZN => n20713);
   U23170 : NOR2_X1 port map( A1 => n28779, A2 => n20941, ZN => n20579);
   U23171 : INV_X1 port map( A => n21585, ZN => n20591);
   U23172 : NOR2_X1 port map( A1 => n3789, A2 => n21322, ZN => n20593);
   U23173 : OAI21_X1 port map( B1 => n20591, B2 => n21322, A => n20886, ZN => 
                           n20592);
   U23174 : NOR3_X1 port map( A1 => n20594, A2 => n20593, A3 => n20592, ZN => 
                           n20595);
   U23178 : NAND2_X1 port map( A1 => n20601, A2 => n20597, ZN => n20599);
   U23179 : MUX2_X1 port map( A => n20600, B => n20599, S => n28408, Z => 
                           n20606);
   U23180 : NOR3_X1 port map( A1 => n20601, A2 => n4569, A3 => n1915, ZN => 
                           n20602);
   U23181 : AOI21_X1 port map( B1 => n20604, B2 => n20603, A => n20602, ZN => 
                           n20605);
   U23182 : INV_X1 port map( A => n21599, ZN => n21603);
   U23183 : AOI22_X1 port map( A1 => n20609, A2 => n20611, B1 => n20608, B2 => 
                           n20607, ZN => n20615);
   U23184 : NAND3_X1 port map( A1 => n20614, A2 => n20611, A3 => n29625, ZN => 
                           n20613);
   U23185 : INV_X1 port map( A => n21600, ZN => n20720);
   U23186 : AND2_X1 port map( A1 => n20617, A2 => n20616, ZN => n20621);
   U23187 : MUX2_X1 port map( A => n20618, B => n6567, S => n20617, Z => n20620
                           );
   U23188 : INV_X1 port map( A => n20722, ZN => n21316);
   U23189 : NOR2_X1 port map( A1 => n1881, A2 => n20626, ZN => n20627);
   U23190 : NAND2_X1 port map( A1 => n20628, A2 => n20627, ZN => n20629);
   U23191 : NAND2_X1 port map( A1 => n21316, A2 => n21601, ZN => n21138);
   U23192 : INV_X1 port map( A => n21138, ZN => n20643);
   U23193 : INV_X1 port map( A => n28538, ZN => n20642);
   U23194 : OAI21_X1 port map( B1 => n20637, B2 => n20636, A => n20635, ZN => 
                           n20638);
   U23195 : OAI21_X1 port map( B1 => n20642, B2 => n20641, A => n20640, ZN => 
                           n21314);
   U23196 : INV_X1 port map( A => n21314, ZN => n21605);
   U23197 : NAND2_X1 port map( A1 => n21314, A2 => n21601, ZN => n20649);
   U23198 : NAND2_X1 port map( A1 => n21308, A2 => n29531, ZN => n21150);
   U23199 : XNOR2_X1 port map( A => n22681, B => n22240, ZN => n20655);
   U23200 : OAI21_X1 port map( B1 => n21119, B2 => n21140, A => n21143, ZN => 
                           n20653);
   U23201 : NAND2_X1 port map( A1 => n21141, A2 => n20650, ZN => n20652);
   U23202 : NOR2_X1 port map( A1 => n20851, A2 => n21118, ZN => n20651);
   U23203 : AOI21_X2 port map( B1 => n20652, B2 => n20653, A => n20651, ZN => 
                           n22855);
   U23204 : XNOR2_X1 port map( A => n22855, B => n1079, ZN => n20654);
   U23206 : XNOR2_X1 port map( A => n22227, B => n3334, ZN => n20660);
   U23207 : XNOR2_X1 port map( A => n20660, B => n22773, ZN => n20665);
   U23210 : OAI21_X1 port map( B1 => n21472, B2 => n21473, A => n21731, ZN => 
                           n20661);
   U23211 : MUX2_X2 port map( A => n20662, B => n20661, S => n21471, Z => 
                           n22697);
   U23212 : XNOR2_X1 port map( A => n22697, B => n22882, ZN => n20664);
   U23213 : XNOR2_X1 port map( A => n20665, B => n20664, ZN => n20682);
   U23214 : MUX2_X1 port map( A => n22286, B => n22026, S => n22023, Z => 
                           n20667);
   U23215 : INV_X1 port map( A => n22286, ZN => n22291);
   U23218 : NAND2_X1 port map( A1 => n22286, A2 => n22290, ZN => n21208);
   U23220 : NAND2_X1 port map( A1 => n20668, A2 => n22294, ZN => n22879);
   U23221 : INV_X1 port map( A => n22879, ZN => n21848);
   U23222 : NOR2_X1 port map( A1 => n21394, A2 => n21632, ZN => n20679);
   U23223 : INV_X1 port map( A => n20669, ZN => n20673);
   U23224 : NOR2_X1 port map( A1 => n20671, A2 => n20670, ZN => n20672);
   U23225 : NAND2_X1 port map( A1 => n20673, A2 => n20672, ZN => n20674);
   U23226 : OAI21_X1 port map( B1 => n20675, B2 => n20674, A => n21638, ZN => 
                           n20678);
   U23227 : NAND2_X1 port map( A1 => n21637, A2 => n21392, ZN => n21226);
   U23228 : NAND2_X1 port map( A1 => n21632, A2 => n21227, ZN => n21393);
   U23229 : NAND2_X1 port map( A1 => n21226, A2 => n21393, ZN => n20676);
   U23230 : NAND2_X1 port map( A1 => n20676, A2 => n21631, ZN => n20677);
   U23231 : OAI21_X1 port map( B1 => n20679, B2 => n20678, A => n20677, ZN => 
                           n22226);
   U23232 : INV_X1 port map( A => n22226, ZN => n22073);
   U23233 : XNOR2_X1 port map( A => n21848, B => n20680, ZN => n20681);
   U23234 : INV_X1 port map( A => n22568, ZN => n21841);
   U23235 : OAI21_X1 port map( B1 => n29227, B2 => n6934, A => n29526, ZN => 
                           n20684);
   U23236 : AOI22_X1 port map( A1 => n21704, A2 => n21273, B1 => n6934, B2 => 
                           n21703, ZN => n20683);
   U23237 : NAND2_X1 port map( A1 => n20684, A2 => n20683, ZN => n22821);
   U23238 : XNOR2_X1 port map( A => n21841, B => n22821, ZN => n20687);
   U23239 : INV_X1 port map( A => n21287, ZN => n20726);
   U23240 : NOR2_X1 port map( A1 => n21288, A2 => n21291, ZN => n20989);
   U23241 : OAI211_X1 port map( C1 => n20914, C2 => n29313, A => n21287, B => 
                           n21292, ZN => n20685);
   U23242 : XNOR2_X1 port map( A => n22890, B => n3527, ZN => n20686);
   U23243 : XNOR2_X1 port map( A => n20687, B => n20686, ZN => n20709);
   U23244 : OAI21_X1 port map( B1 => n20688, B2 => n20689, A => n5772, ZN => 
                           n20975);
   U23245 : INV_X1 port map( A => n20975, ZN => n21261);
   U23246 : INV_X1 port map( A => n20688, ZN => n20691);
   U23247 : NOR2_X1 port map( A1 => n20689, A2 => n21364, ZN => n20690);
   U23248 : INV_X1 port map( A => n21717, ZN => n21260);
   U23249 : NOR2_X1 port map( A1 => n21714, A2 => n21713, ZN => n21263);
   U23250 : OAI21_X1 port map( B1 => n21260, B2 => n21258, A => n21263, ZN => 
                           n20692);
   U23251 : NAND2_X1 port map( A1 => n21809, A2 => n21810, ZN => n20699);
   U23252 : NAND2_X1 port map( A1 => n20694, A2 => n20693, ZN => n21250);
   U23253 : INV_X1 port map( A => n21250, ZN => n20695);
   U23254 : INV_X1 port map( A => n21254, ZN => n20696);
   U23255 : INV_X1 port map( A => n21806, ZN => n21379);
   U23256 : AOI21_X1 port map( B1 => n20696, B2 => n21379, A => n21253, ZN => 
                           n20697);
   U23257 : XNOR2_X1 port map( A => n22796, B => n1858, ZN => n22249);
   U23258 : NOR2_X1 port map( A1 => n21346, A2 => n21343, ZN => n21691);
   U23261 : NOR2_X1 port map( A1 => n21695, A2 => n21242, ZN => n20700);
   U23262 : INV_X1 port map( A => n21696, ZN => n21348);
   U23263 : NOR2_X1 port map( A1 => n20702, A2 => n20701, ZN => n20969);
   U23264 : NAND2_X1 port map( A1 => n20969, A2 => n20704, ZN => n20707);
   U23265 : OAI21_X1 port map( B1 => n20703, B2 => n381, A => n21217, ZN => 
                           n20706);
   U23266 : INV_X1 port map( A => n21218, ZN => n20967);
   U23267 : XNOR2_X1 port map( A => n22798, B => n22248, ZN => n22486);
   U23268 : XOR2_X1 port map( A => n22249, B => n22486, Z => n20708);
   U23269 : INV_X1 port map( A => n20875, ZN => n20710);
   U23270 : OAI21_X1 port map( B1 => n21268, B2 => n20710, A => n20878, ZN => 
                           n20712);
   U23271 : NAND3_X1 port map( A1 => n20816, A2 => n20878, A3 => n20875, ZN => 
                           n20711);
   U23272 : XNOR2_X1 port map( A => n22327, B => n22913, ZN => n21838);
   U23273 : INV_X1 port map( A => n21591, ZN => n20717);
   U23274 : AND2_X1 port map( A1 => n21322, A2 => n5983, ZN => n20716);
   U23275 : OAI21_X1 port map( B1 => n20717, B2 => n20716, A => n28584, ZN => 
                           n20718);
   U23276 : AND2_X1 port map( A1 => n21086, A2 => n21426, ZN => n20719);
   U23277 : XNOR2_X1 port map( A => n22232, B => n22759, ZN => n22474);
   U23278 : XNOR2_X1 port map( A => n22474, B => n21838, ZN => n20735);
   U23279 : AOI21_X1 port map( B1 => n21599, B2 => n20721, A => n20720, ZN => 
                           n20725);
   U23280 : NAND2_X1 port map( A1 => n21598, A2 => n21601, ZN => n20724);
   U23281 : NAND2_X1 port map( A1 => n20916, A2 => n20726, ZN => n20728);
   U23282 : INV_X1 port map( A => n20917, ZN => n20727);
   U23283 : XNOR2_X1 port map( A => n22845, B => n22762, ZN => n22358);
   U23287 : NAND3_X1 port map( A1 => n21326, A2 => n21327, A3 => n21612, ZN => 
                           n20730);
   U23289 : XNOR2_X1 port map( A => n22763, B => n2987, ZN => n20733);
   U23290 : XNOR2_X1 port map( A => n22358, B => n20733, ZN => n20734);
   U23291 : INV_X1 port map( A => n20736, ZN => n20738);
   U23292 : NAND2_X1 port map( A1 => n20738, A2 => n20737, ZN => n20742);
   U23293 : INV_X1 port map( A => n20739, ZN => n20740);
   U23294 : NOR3_X1 port map( A1 => n20742, A2 => n20741, A3 => n20740, ZN => 
                           n20743);
   U23295 : NAND2_X1 port map( A1 => n494, A2 => n21155, ZN => n20745);
   U23296 : AOI21_X1 port map( B1 => n20746, B2 => n20745, A => n4960, ZN => 
                           n20747);
   U23297 : NOR2_X2 port map( A1 => n20748, A2 => n20747, ZN => n22812);
   U23298 : INV_X1 port map( A => n22437, ZN => n20750);
   U23299 : XNOR2_X1 port map( A => n20750, B => n22812, ZN => n20753);
   U23300 : NOR2_X1 port map( A1 => n28789, A2 => n6752, ZN => n20751);
   U23301 : AOI21_X1 port map( B1 => n2037, B2 => n1946, A => n21496, ZN => 
                           n20752);
   U23302 : XNOR2_X1 port map( A => n22898, B => n22245, ZN => n22688);
   U23303 : XNOR2_X1 port map( A => n22688, B => n20753, ZN => n20761);
   U23304 : XNOR2_X1 port map( A => n21728, B => n22330, ZN => n20759);
   U23305 : XNOR2_X1 port map( A => n22778, B => n135, ZN => n20758);
   U23306 : XNOR2_X1 port map( A => n20759, B => n20758, ZN => n20760);
   U23307 : NOR2_X1 port map( A1 => n20762, A2 => n4828, ZN => n20764);
   U23308 : NOR3_X1 port map( A1 => n22012, A2 => n22011, A3 => n22013, ZN => 
                           n20763);
   U23309 : NOR3_X1 port map( A1 => n22014, A2 => n20764, A3 => n20763, ZN => 
                           n20765);
   U23310 : XNOR2_X1 port map( A => n20765, B => n28499, ZN => n21856);
   U23312 : INV_X1 port map( A => n21308, ZN => n20769);
   U23313 : NOR2_X1 port map( A1 => n20769, A2 => n29530, ZN => n21305);
   U23314 : NOR2_X1 port map( A1 => n21153, A2 => n21305, ZN => n20775);
   U23315 : NAND2_X1 port map( A1 => n20938, A2 => n21306, ZN => n20770);
   U23316 : NAND2_X1 port map( A1 => n21308, A2 => n20770, ZN => n20772);
   U23317 : INV_X1 port map( A => n21500, ZN => n21543);
   U23319 : AOI21_X1 port map( B1 => n21500, B2 => n21539, A => n21192, ZN => 
                           n20778);
   U23320 : INV_X1 port map( A => n21539, ZN => n20945);
   U23321 : INV_X1 port map( A => n28619, ZN => n20948);
   U23322 : OAI21_X1 port map( B1 => n20945, B2 => n20948, A => n21192, ZN => 
                           n20781);
   U23323 : INV_X1 port map( A => n21503, ZN => n21540);
   U23324 : NOR3_X1 port map( A1 => n21540, A2 => n21539, A3 => n28185, ZN => 
                           n20780);
   U23325 : XNOR2_X1 port map( A => n20885, B => n22219, ZN => n22461);
   U23327 : INV_X1 port map( A => n22792, ZN => n22086);
   U23328 : XNOR2_X1 port map( A => n22086, B => n2961, ZN => n20797);
   U23329 : NOR2_X1 port map( A1 => n21930, A2 => n21932, ZN => n20785);
   U23330 : NAND2_X1 port map( A1 => n20785, A2 => n20954, ZN => n20791);
   U23331 : INV_X1 port map( A => n20801, ZN => n20788);
   U23332 : NOR2_X1 port map( A1 => n21932, A2 => n21097, ZN => n20787);
   U23333 : AOI22_X1 port map( A1 => n20788, A2 => n21932, B1 => n20787, B2 => 
                           n20786, ZN => n20790);
   U23334 : INV_X1 port map( A => n21513, ZN => n21512);
   U23335 : NAND3_X1 port map( A1 => n21534, A2 => n21530, A3 => n21509, ZN => 
                           n20795);
   U23336 : INV_X1 port map( A => n21514, ZN => n21533);
   U23337 : NAND3_X1 port map( A1 => n21533, A2 => n21199, A3 => n21532, ZN => 
                           n20794);
   U23338 : XNOR2_X1 port map( A => n22790, B => n22835, ZN => n22383);
   U23339 : NAND2_X1 port map( A1 => n23353, A2 => n4231, ZN => n20840);
   U23340 : INV_X1 port map( A => n20798, ZN => n22340);
   U23341 : INV_X1 port map( A => n20954, ZN => n20800);
   U23342 : XNOR2_X1 port map( A => n22340, B => n22903, ZN => n20813);
   U23343 : NAND2_X1 port map( A1 => n20899, A2 => n21424, ZN => n20808);
   U23344 : NAND2_X1 port map( A1 => n21087, A2 => n21425, ZN => n20806);
   U23345 : OAI21_X1 port map( B1 => n28602, B2 => n20808, A => n20807, ZN => 
                           n22553);
   U23346 : INV_X1 port map( A => n21665, ZN => n21015);
   U23347 : NAND3_X1 port map( A1 => n22404, A2 => n21662, A3 => n22401, ZN => 
                           n20811);
   U23348 : INV_X1 port map( A => n21018, ZN => n20809);
   U23349 : NAND2_X1 port map( A1 => n22402, A2 => n20809, ZN => n20810);
   U23350 : AND3_X1 port map( A1 => n20812, A2 => n20811, A3 => n20810, ZN => 
                           n21805);
   U23351 : INV_X1 port map( A => n21805, ZN => n22066);
   U23352 : XNOR2_X1 port map( A => n22066, B => n22553, ZN => n22748);
   U23353 : XNOR2_X1 port map( A => n20813, B => n22748, ZN => n20839);
   U23354 : NOR2_X1 port map( A1 => n29488, A2 => n20816, ZN => n20815);
   U23355 : INV_X1 port map( A => n20816, ZN => n20874);
   U23356 : NAND3_X1 port map( A1 => n21268, A2 => n20874, A3 => n20875, ZN => 
                           n20817);
   U23357 : NAND2_X1 port map( A1 => n21272, A2 => n20817, ZN => n20820);
   U23358 : INV_X1 port map( A => n20878, ZN => n21267);
   U23359 : AOI21_X1 port map( B1 => n20818, B2 => n21267, A => n21268, ZN => 
                           n20819);
   U23360 : INV_X1 port map( A => n21676, ZN => n21673);
   U23361 : INV_X1 port map( A => n20821, ZN => n20822);
   U23362 : NOR2_X1 port map( A1 => n20823, A2 => n20822, ZN => n20828);
   U23363 : INV_X1 port map( A => n20824, ZN => n20825);
   U23364 : NAND2_X1 port map( A1 => n20825, A2 => n20418, ZN => n20827);
   U23365 : OAI21_X1 port map( B1 => n20828, B2 => n20827, A => n28215, ZN => 
                           n20829);
   U23366 : XNOR2_X1 port map( A => n22718, B => n22426, ZN => n22497);
   U23367 : INV_X1 port map( A => n21653, ZN => n21660);
   U23371 : XNOR2_X1 port map( A => n22497, B => n20837, ZN => n20838);
   U23372 : NAND3_X1 port map( A1 => n21125, A2 => n21458, A3 => n21567, ZN => 
                           n20845);
   U23373 : XNOR2_X1 port map( A => n22703, B => n22033, ZN => n20850);
   U23374 : XNOR2_X1 port map( A => n22773, B => n20850, ZN => n20873);
   U23375 : INV_X1 port map( A => n21118, ZN => n20854);
   U23376 : MUX2_X1 port map( A => n20854, B => n20851, S => n21119, Z => 
                           n20856);
   U23378 : OAI21_X1 port map( B1 => n494, B2 => n20858, A => n20857, ZN => 
                           n20859);
   U23379 : AOI21_X1 port map( B1 => n21158, B2 => n20858, A => n20859, ZN => 
                           n20860);
   U23380 : XNOR2_X1 port map( A => n22670, B => n22526, ZN => n21339);
   U23381 : XNOR2_X1 port map( A => n22387, B => n3081, ZN => n20870);
   U23382 : MUX2_X1 port map( A => n21497, B => n21495, S => n20864, Z => 
                           n20869);
   U23383 : NOR2_X1 port map( A1 => n28789, A2 => n21496, ZN => n20866);
   U23386 : XNOR2_X1 port map( A => n20870, B => n22523, ZN => n20871);
   U23387 : XNOR2_X1 port map( A => n20871, B => n21339, ZN => n20872);
   U23388 : OR3_X1 port map( A1 => n21269, A2 => n20874, A3 => n21266, ZN => 
                           n20884);
   U23389 : NAND3_X1 port map( A1 => n21269, A2 => n21268, A3 => n20878, ZN => 
                           n20883);
   U23390 : NOR2_X1 port map( A1 => n20876, A2 => n20875, ZN => n20881);
   U23391 : NOR2_X1 port map( A1 => n21268, A2 => n21267, ZN => n20880);
   U23392 : INV_X1 port map( A => n20890, ZN => n20893);
   U23393 : INV_X1 port map( A => n20891, ZN => n20892);
   U23394 : NOR4_X1 port map( A1 => n20898, A2 => n20897, A3 => n20893, A4 => 
                           n20892, ZN => n20894);
   U23395 : NAND2_X1 port map( A1 => n1925, A2 => n21085, ZN => n20901);
   U23396 : NOR3_X1 port map( A1 => n20898, A2 => n20897, A3 => n21424, ZN => 
                           n21084);
   U23397 : INV_X1 port map( A => n20899, ZN => n20900);
   U23398 : XNOR2_X1 port map( A => n21760, B => n22545, ZN => n20925);
   U23399 : OAI21_X1 port map( B1 => n28442, B2 => n21600, A => n21316, ZN => 
                           n20904);
   U23400 : INV_X1 port map( A => n21601, ZN => n21315);
   U23401 : NOR2_X1 port map( A1 => n21598, A2 => n21601, ZN => n21320);
   U23402 : INV_X1 port map( A => n21320, ZN => n20902);
   U23403 : OAI211_X1 port map( C1 => n20905, C2 => n21315, A => n1941, B => 
                           n20902, ZN => n20903);
   U23405 : INV_X1 port map( A => n20906, ZN => n20908);
   U23406 : NOR2_X1 port map( A1 => n20908, A2 => n20907, ZN => n20912);
   U23407 : INV_X1 port map( A => n21334, ZN => n21607);
   U23408 : INV_X1 port map( A => n21612, ZN => n21609);
   U23409 : AOI22_X1 port map( A1 => n20910, A2 => n21163, B1 => n20909, B2 => 
                           n21609, ZN => n20911);
   U23410 : NAND2_X1 port map( A1 => n20915, A2 => n20914, ZN => n20920);
   U23411 : NAND3_X1 port map( A1 => n21292, A2 => n20916, A3 => n20986, ZN => 
                           n20919);
   U23412 : NAND4_X2 port map( A1 => n20918, A2 => n20921, A3 => n20920, A4 => 
                           n20919, ZN => n22664);
   U23413 : XNOR2_X1 port map( A => n22664, B => n27298, ZN => n20922);
   U23414 : XNOR2_X1 port map( A => n20923, B => n20922, ZN => n20924);
   U23415 : XNOR2_X1 port map( A => n20925, B => n20924, ZN => n23167);
   U23416 : NOR2_X1 port map( A1 => n28457, A2 => n23167, ZN => n21027);
   U23417 : MUX2_X1 port map( A => n21530, B => n21514, S => n21513, Z => 
                           n20928);
   U23419 : NAND2_X1 port map( A1 => n21516, A2 => n21514, ZN => n20926);
   U23420 : MUX2_X1 port map( A => n21535, B => n20926, S => n21530, Z => 
                           n20927);
   U23421 : NAND2_X1 port map( A1 => n20931, A2 => n21549, ZN => n20929);
   U23422 : INV_X1 port map( A => n22689, ZN => n20937);
   U23423 : INV_X1 port map( A => n20934, ZN => n20935);
   U23424 : XNOR2_X1 port map( A => n22897, B => n22437, ZN => n20936);
   U23425 : XNOR2_X1 port map( A => n20937, B => n20936, ZN => n20960);
   U23426 : INV_X1 port map( A => n21192, ZN => n21538);
   U23427 : NAND2_X1 port map( A1 => n21500, A2 => n28611, ZN => n20950);
   U23429 : INV_X1 port map( A => n20939, ZN => n20942);
   U23430 : NOR2_X1 port map( A1 => n503, A2 => n20941, ZN => n20940);
   U23431 : AOI22_X1 port map( A1 => n20942, A2 => n20941, B1 => n20940, B2 => 
                           n20413, ZN => n20943);
   U23432 : NAND2_X1 port map( A1 => n20777, A2 => n20943, ZN => n20944);
   U23436 : NOR3_X1 port map( A1 => n20954, A2 => n28916, A3 => n20953, ZN => 
                           n20956);
   U23437 : XNOR2_X1 port map( A => n22811, B => n730, ZN => n20958);
   U23438 : XNOR2_X1 port map( A => n22502, B => n20958, ZN => n20959);
   U23441 : NAND2_X1 port map( A1 => n21347, A2 => n20961, ZN => n20965);
   U23442 : NOR3_X1 port map( A1 => n3260, A2 => n28440, A3 => n21692, ZN => 
                           n20964);
   U23443 : NOR3_X2 port map( A1 => n20965, A2 => n20964, A3 => n20963, ZN => 
                           n22338);
   U23444 : NOR2_X1 port map( A1 => n20999, A2 => n21221, ZN => n20971);
   U23445 : OAI21_X1 port map( B1 => n20969, B2 => n20968, A => n20967, ZN => 
                           n20970);
   U23446 : OAI21_X1 port map( B1 => n20972, B2 => n20971, A => n20970, ZN => 
                           n22717);
   U23447 : XNOR2_X1 port map( A => n29562, B => n3134, ZN => n20973);
   U23448 : XNOR2_X1 port map( A => n22519, B => n20973, ZN => n20997);
   U23449 : NAND2_X1 port map( A1 => n21713, A2 => n20976, ZN => n20974);
   U23450 : AOI21_X1 port map( B1 => n20975, B2 => n20974, A => n21260, ZN => 
                           n20979);
   U23451 : OAI22_X1 port map( A1 => n20977, A2 => n21717, B1 => n20976, B2 => 
                           n21712, ZN => n20978);
   U23452 : NOR2_X1 port map( A1 => n20979, A2 => n20978, ZN => n22104);
   U23454 : INV_X1 port map( A => n21811, ZN => n20982);
   U23455 : NOR2_X1 port map( A1 => n21809, A2 => n21806, ZN => n21380);
   U23456 : INV_X1 port map( A => n21380, ZN => n20984);
   U23457 : XNOR2_X1 port map( A => n22713, B => n29591, ZN => n20995);
   U23458 : NOR2_X1 port map( A1 => n20988, A2 => n21291, ZN => n20987);
   U23459 : OAI21_X1 port map( B1 => n20987, B2 => n20986, A => n20985, ZN => 
                           n20991);
   U23460 : OAI21_X1 port map( B1 => n20989, B2 => n6911, A => n20988, ZN => 
                           n20990);
   U23461 : INV_X1 port map( A => n21703, ZN => n20992);
   U23462 : NAND2_X1 port map( A1 => n20992, A2 => n29526, ZN => n21281);
   U23463 : INV_X1 port map( A => n21372, ZN => n21702);
   U23464 : NAND3_X1 port map( A1 => n21705, A2 => n20992, A3 => n21372, ZN => 
                           n20993);
   U23465 : XNOR2_X1 port map( A => n22006, B => n22856, ZN => n21470);
   U23466 : XNOR2_X1 port map( A => n21470, B => n20995, ZN => n20996);
   U23467 : XNOR2_X1 port map( A => n20996, B => n20997, ZN => n23168);
   U23468 : NOR2_X1 port map( A1 => n23683, A2 => n23168, ZN => n21026);
   U23469 : NAND2_X1 port map( A1 => n20998, A2 => n21221, ZN => n21003);
   U23470 : INV_X1 port map( A => n20999, ZN => n21002);
   U23471 : NAND3_X1 port map( A1 => n21221, A2 => n21000, A3 => n21218, ZN => 
                           n21001);
   U23472 : XNOR2_X1 port map( A => n22759, B => n22912, ZN => n21766);
   U23473 : INV_X1 port map( A => n21004, ZN => n21006);
   U23474 : NOR2_X1 port map( A1 => n21675, A2 => n21677, ZN => n21079);
   U23475 : OAI21_X1 port map( B1 => n21079, B2 => n21676, A => n21448, ZN => 
                           n21005);
   U23476 : AND2_X1 port map( A1 => n21808, A2 => n19732, ZN => n21011);
   U23477 : NOR2_X1 port map( A1 => n19732, A2 => n21806, ZN => n21010);
   U23478 : INV_X1 port map( A => n21810, ZN => n21008);
   U23479 : NAND3_X1 port map( A1 => n21811, A2 => n21008, A3 => n21379, ZN => 
                           n21009);
   U23480 : XNOR2_X1 port map( A => n22910, B => n22734, ZN => n22532);
   U23481 : XNOR2_X1 port map( A => n22532, B => n21766, ZN => n21025);
   U23482 : XNOR2_X1 port map( A => n22731, B => n22735, ZN => n21023);
   U23483 : OAI21_X1 port map( B1 => n22291, B2 => n29364, A => n21213, ZN => 
                           n21021);
   U23484 : INV_X1 port map( A => n22290, ZN => n21019);
   U23485 : INV_X1 port map( A => n21917, ZN => n22844);
   U23486 : XNOR2_X1 port map( A => n22844, B => n3423, ZN => n21022);
   U23487 : XNOR2_X1 port map( A => n21023, B => n21022, ZN => n21024);
   U23488 : XNOR2_X2 port map( A => n21025, B => n21024, ZN => n23016);
   U23490 : INV_X1 port map( A => n23168, ZN => n23682);
   U23491 : NOR2_X1 port map( A1 => n22140, A2 => n22139, ZN => n21106);
   U23492 : NOR2_X1 port map( A1 => n21030, A2 => n5339, ZN => n21031);
   U23493 : NAND2_X1 port map( A1 => n21736, A2 => n21389, ZN => n21033);
   U23494 : XNOR2_X1 port map( A => n22271, B => n22888, ZN => n22511);
   U23495 : XNOR2_X1 port map( A => n22798, B => n3586, ZN => n21035);
   U23496 : XNOR2_X1 port map( A => n22511, B => n21035, ZN => n21057);
   U23497 : NOR2_X1 port map( A1 => n21639, A2 => n21036, ZN => n21038);
   U23498 : NAND2_X1 port map( A1 => n21227, A2 => n21392, ZN => n21395);
   U23499 : NAND2_X1 port map( A1 => n21395, A2 => n21638, ZN => n21037);
   U23500 : INV_X1 port map( A => n21040, ZN => n21041);
   U23501 : NAND2_X1 port map( A1 => n21041, A2 => n21400, ZN => n21045);
   U23502 : NAND3_X1 port map( A1 => n21042, A2 => n21402, A3 => n21750, ZN => 
                           n21044);
   U23503 : NAND2_X1 port map( A1 => n21410, A2 => n21409, ZN => n21051);
   U23505 : AND2_X1 port map( A1 => n21408, A2 => n21171, ZN => n21413);
   U23507 : NAND2_X1 port map( A1 => n21053, A2 => n21187, ZN => n21054);
   U23508 : NAND2_X1 port map( A1 => n21055, A2 => n21054, ZN => n22509);
   U23509 : XNOR2_X1 port map( A => n22820, B => n22509, ZN => n21525);
   U23510 : XNOR2_X1 port map( A => n22727, B => n21525, ZN => n21056);
   U23511 : NAND2_X1 port map( A1 => n23679, A2 => n23168, ZN => n21058);
   U23513 : NOR2_X2 port map( A1 => n21060, A2 => n21059, ZN => n24617);
   U23515 : NAND2_X1 port map( A1 => n21061, A2 => n21062, ZN => n21066);
   U23516 : NAND2_X1 port map( A1 => n21063, A2 => n21062, ZN => n21064);
   U23517 : INV_X1 port map( A => n21663, ZN => n21433);
   U23518 : AND2_X1 port map( A1 => n21433, A2 => n22401, ZN => n21068);
   U23519 : NAND2_X1 port map( A1 => n22404, A2 => n21067, ZN => n22403);
   U23520 : NAND2_X1 port map( A1 => n21656, A2 => n21657, ZN => n21075);
   U23521 : NAND3_X1 port map( A1 => n21654, A2 => n6275, A3 => n21012, ZN => 
                           n21072);
   U23522 : NAND2_X1 port map( A1 => n20833, A2 => n21657, ZN => n21071);
   U23523 : AND2_X1 port map( A1 => n21077, A2 => n21076, ZN => n21819);
   U23524 : XNOR2_X1 port map( A => n21847, B => n22594, ZN => n21105);
   U23525 : INV_X1 port map( A => n21079, ZN => n21082);
   U23526 : AOI21_X1 port map( B1 => n21675, B2 => n21673, A => n21678, ZN => 
                           n21081);
   U23527 : INV_X1 port map( A => n21448, ZN => n21680);
   U23528 : XNOR2_X1 port map( A => n22199, B => n2986, ZN => n21083);
   U23529 : OAI211_X1 port map( C1 => n21087, C2 => n21425, A => n21424, B => 
                           n21086, ZN => n21088);
   U23530 : AOI21_X1 port map( B1 => n4877, B2 => n21091, A => n28479, ZN => 
                           n21094);
   U23531 : NAND2_X1 port map( A1 => n29134, A2 => n18919, ZN => n21093);
   U23532 : AOI22_X1 port map( A1 => n21096, A2 => n28479, B1 => n21094, B2 => 
                           n21093, ZN => n21098);
   U23533 : NAND2_X1 port map( A1 => n21098, A2 => n21097, ZN => n21099);
   U23534 : XNOR2_X1 port map( A => n22298, B => n22768, ZN => n21946);
   U23536 : NAND3_X1 port map( A1 => n22141, A2 => n22145, A3 => n6532, ZN => 
                           n21108);
   U23537 : NAND2_X1 port map( A1 => n21106, A2 => n22141, ZN => n21107);
   U23538 : INV_X1 port map( A => n22116, ZN => n21871);
   U23539 : XNOR2_X1 port map( A => n21871, B => n22052, ZN => n21116);
   U23540 : NAND3_X1 port map( A1 => n21156, A2 => n21155, A3 => n21159, ZN => 
                           n21110);
   U23541 : OAI21_X1 port map( B1 => n21111, B2 => n4960, A => n21110, ZN => 
                           n21112);
   U23542 : NAND2_X1 port map( A1 => n21113, A2 => n21464, ZN => n21564);
   U23544 : XNOR2_X1 port map( A => n28486, B => n22410, ZN => n22159);
   U23545 : XNOR2_X1 port map( A => n22159, B => n21116, ZN => n21133);
   U23546 : AOI21_X1 port map( B1 => n21143, B2 => n21140, A => n21119, ZN => 
                           n21123);
   U23547 : AOI22_X1 port map( A1 => n21119, A2 => n21118, B1 => n21144, B2 => 
                           n21140, ZN => n21121);
   U23548 : OAI22_X1 port map( A1 => n21123, A2 => n21122, B1 => n21121, B2 => 
                           n21120, ZN => n22760);
   U23549 : INV_X1 port map( A => n22760, ZN => n22328);
   U23550 : XNOR2_X1 port map( A => n22328, B => n3374, ZN => n21131);
   U23551 : NAND3_X1 port map( A1 => n1832, A2 => n21496, A3 => n21495, ZN => 
                           n21128);
   U23553 : XNOR2_X1 port map( A => n22409, B => n22414, ZN => n21130);
   U23554 : XNOR2_X1 port map( A => n21131, B => n21130, ZN => n21132);
   U23555 : XNOR2_X1 port map( A => n21133, B => n21132, ZN => n23678);
   U23556 : NOR2_X1 port map( A1 => n23360, A2 => n23678, ZN => n23367);
   U23557 : XNOR2_X1 port map( A => n22418, B => n22822, ZN => n21149);
   U23558 : NOR2_X1 port map( A1 => n21140, A2 => n21143, ZN => n21142);
   U23559 : NOR2_X1 port map( A1 => n21142, A2 => n21141, ZN => n21147);
   U23560 : XNOR2_X1 port map( A => n22059, B => n26680, ZN => n21148);
   U23561 : XNOR2_X1 port map( A => n21149, B => n21148, ZN => n21170);
   U23562 : NAND2_X1 port map( A1 => n21311, A2 => n21309, ZN => n21152);
   U23564 : INV_X1 port map( A => n22419, ZN => n21154);
   U23565 : XNOR2_X1 port map( A => n22098, B => n21154, ZN => n21168);
   U23566 : NAND3_X1 port map( A1 => n21156, A2 => n4960, A3 => n21155, ZN => 
                           n21161);
   U23567 : INV_X1 port map( A => n21618, ZN => n21166);
   U23568 : AND2_X1 port map( A1 => n21162, A2 => n21613, ZN => n21165);
   U23569 : INV_X1 port map( A => n21326, ZN => n21608);
   U23570 : XNOR2_X1 port map( A => n22656, B => n22506, ZN => n22801);
   U23571 : INV_X1 port map( A => n22801, ZN => n21167);
   U23572 : XNOR2_X1 port map( A => n21167, B => n21168, ZN => n21169);
   U23573 : NAND3_X1 port map( A1 => n21412, A2 => n21414, A3 => n28184, ZN => 
                           n21175);
   U23574 : AND2_X1 port map( A1 => n21410, A2 => n21171, ZN => n21173);
   U23575 : INV_X1 port map( A => n21410, ZN => n21172);
   U23576 : AOI22_X1 port map( A1 => n21414, A2 => n21173, B1 => n21172, B2 => 
                           n21408, ZN => n21174);
   U23578 : NAND2_X1 port map( A1 => n21549, A2 => n1875, ZN => n21179);
   U23579 : NAND3_X1 port map( A1 => n21180, A2 => n21549, A3 => n21547, ZN => 
                           n21178);
   U23580 : XNOR2_X1 port map( A => n21182, B => n22678, ZN => n22752);
   U23581 : INV_X1 port map( A => n22752, ZN => n21191);
   U23582 : NOR2_X1 port map( A1 => n1832, A2 => n28789, ZN => n21184);
   U23584 : NAND2_X1 port map( A1 => n22286, A2 => n21213, ZN => n21189);
   U23585 : XNOR2_X1 port map( A => n22427, B => n22068, ZN => n21190);
   U23586 : XNOR2_X1 port map( A => n21191, B => n21190, ZN => n21206);
   U23588 : NAND2_X1 port map( A1 => n21503, A2 => n21500, ZN => n21196);
   U23589 : NOR2_X1 port map( A1 => n21503, A2 => n28619, ZN => n21194);
   U23591 : XNOR2_X1 port map( A => n29489, B => n22855, ZN => n21204);
   U23592 : AOI22_X1 port map( A1 => n21198, A2 => n21532, B1 => n21514, B2 => 
                           n21512, ZN => n21202);
   U23593 : NOR2_X1 port map( A1 => n21514, A2 => n21530, ZN => n21200);
   U23594 : AOI22_X1 port map( A1 => n21200, A2 => n21509, B1 => n21533, B2 => 
                           n21199, ZN => n21201);
   U23595 : XNOR2_X1 port map( A => n22854, B => n900, ZN => n21203);
   U23596 : XNOR2_X1 port map( A => n21204, B => n21203, ZN => n21205);
   U23597 : NOR2_X1 port map( A1 => n23672, A2 => n23131, ZN => n21207);
   U23598 : NOR2_X1 port map( A1 => n23367, A2 => n21207, ZN => n23108);
   U23599 : INV_X1 port map( A => n23678, ZN => n23363);
   U23600 : OAI21_X1 port map( B1 => n28790, B2 => n22286, A => n21208, ZN => 
                           n21214);
   U23601 : AOI21_X1 port map( B1 => n21210, B2 => n21209, A => n22290, ZN => 
                           n21212);
   U23602 : AND2_X1 port map( A1 => n21215, A2 => n21221, ZN => n21225);
   U23603 : OR2_X1 port map( A1 => n21220, A2 => n21216, ZN => n21224);
   U23604 : NAND2_X1 port map( A1 => n21220, A2 => n381, ZN => n21222);
   U23605 : NAND2_X1 port map( A1 => n21218, A2 => n21217, ZN => n21219);
   U23606 : OAI22_X1 port map( A1 => n21222, A2 => n21221, B1 => n21220, B2 => 
                           n21219, ZN => n21223);
   U23607 : XNOR2_X1 port map( A => n29079, B => n28517, ZN => n21671);
   U23608 : XNOR2_X1 port map( A => n22164, B => n21671, ZN => n21241);
   U23609 : XNOR2_X1 port map( A => n22194, B => n2465, ZN => n21239);
   U23610 : INV_X1 port map( A => n21472, ZN => n21478);
   U23611 : MUX2_X1 port map( A => n1930, B => n21471, S => n21478, Z => n21234
                           );
   U23612 : NOR2_X1 port map( A1 => n21389, A2 => n21473, ZN => n21231);
   U23613 : NAND2_X1 port map( A1 => n21231, A2 => n1930, ZN => n21232);
   U23615 : NAND2_X1 port map( A1 => n21748, A2 => n20658, ZN => n21235);
   U23616 : NAND2_X1 port map( A1 => n21645, A2 => n21400, ZN => n21646);
   U23617 : OAI22_X1 port map( A1 => n21235, A2 => n21749, B1 => n20658, B2 => 
                           n21646, ZN => n21238);
   U23618 : NAND2_X1 port map( A1 => n21402, A2 => n497, ZN => n21236);
   U23619 : XNOR2_X1 port map( A => n22195, B => n22278, ZN => n22442);
   U23620 : XNOR2_X1 port map( A => n22442, B => n21239, ZN => n21240);
   U23621 : XNOR2_X1 port map( A => n21241, B => n21240, ZN => n23673);
   U23622 : NOR2_X1 port map( A1 => n21346, A2 => n29101, ZN => n21244);
   U23623 : NOR2_X1 port map( A1 => n21242, A2 => n21698, ZN => n21243);
   U23624 : NOR2_X1 port map( A1 => n21348, A2 => n28440, ZN => n21245);
   U23626 : NAND3_X1 port map( A1 => n21251, A2 => n21250, A3 => n21249, ZN => 
                           n21252);
   U23627 : OAI211_X1 port map( C1 => n21254, C2 => n21253, A => n19732, B => 
                           n21252, ZN => n21256);
   U23628 : OAI211_X1 port map( C1 => n21808, C2 => n19732, A => n21256, B => 
                           n21255, ZN => n21955);
   U23629 : XNOR2_X1 port map( A => n22204, B => n21955, ZN => n22436);
   U23630 : INV_X1 port map( A => n21713, ZN => n21257);
   U23631 : NOR3_X1 port map( A1 => n21714, A2 => n21366, A3 => n21258, ZN => 
                           n21259);
   U23632 : AOI21_X1 port map( B1 => n21261, B2 => n21260, A => n21259, ZN => 
                           n21262);
   U23633 : XNOR2_X1 port map( A => n22093, B => n22561, ZN => n22810);
   U23635 : XNOR2_X1 port map( A => n28432, B => n22436, ZN => n21300);
   U23636 : INV_X1 port map( A => n21269, ZN => n21270);
   U23637 : XNOR2_X1 port map( A => n22363, B => n3516, ZN => n21298);
   U23639 : NAND2_X1 port map( A1 => n21274, A2 => n29227, ZN => n21285);
   U23640 : INV_X1 port map( A => n21275, ZN => n21276);
   U23641 : NAND2_X1 port map( A1 => n29526, A2 => n21276, ZN => n21282);
   U23642 : NAND2_X1 port map( A1 => n21372, A2 => n496, ZN => n21279);
   U23643 : NAND2_X1 port map( A1 => n21279, A2 => n21278, ZN => n21280);
   U23644 : OAI211_X1 port map( C1 => n21283, C2 => n21282, A => n21281, B => 
                           n21280, ZN => n21284);
   U23645 : NAND2_X1 port map( A1 => n21288, A2 => n21287, ZN => n21294);
   U23646 : NAND2_X1 port map( A1 => n21294, A2 => n29313, ZN => n21296);
   U23647 : NAND2_X1 port map( A1 => n21291, A2 => n21290, ZN => n21293);
   U23648 : MUX2_X1 port map( A => n21294, B => n21293, S => n21292, Z => 
                           n21295);
   U23649 : XNOR2_X1 port map( A => n22501, B => n22644, ZN => n22776);
   U23650 : XNOR2_X1 port map( A => n22776, B => n21298, ZN => n21299);
   U23652 : OAI211_X1 port map( C1 => n23363, C2 => n23673, A => n23672, B => 
                           n28604, ZN => n21301);
   U23653 : OAI21_X1 port map( B1 => n21302, B2 => n23108, A => n21301, ZN => 
                           n24748);
   U23654 : INV_X1 port map( A => n24748, ZN => n21303);
   U23655 : INV_X1 port map( A => n22594, ZN => n22077);
   U23656 : OAI21_X1 port map( B1 => n29328, B2 => n21307, A => n21311, ZN => 
                           n21313);
   U23657 : NOR2_X1 port map( A1 => n21308, A2 => n29531, ZN => n21312);
   U23658 : NAND3_X1 port map( A1 => n21316, A2 => n21315, A3 => n21314, ZN => 
                           n21318);
   U23659 : NAND3_X1 port map( A1 => n21603, A2 => n21601, A3 => n21600, ZN => 
                           n21317);
   U23660 : AOI21_X1 port map( B1 => n21613, B2 => n21327, A => n21326, ZN => 
                           n21337);
   U23661 : NAND2_X1 port map( A1 => n21328, A2 => n21327, ZN => n21333);
   U23662 : NAND3_X1 port map( A1 => n21331, A2 => n20497, A3 => n21330, ZN => 
                           n21332);
   U23663 : XNOR2_X1 port map( A => n29514, B => n3276, ZN => n21338);
   U23664 : XNOR2_X1 port map( A => n21339, B => n21338, ZN => n21340);
   U23665 : XNOR2_X1 port map( A => n22664, B => n3049, ZN => n21342);
   U23666 : XNOR2_X1 port map( A => n21342, B => n28517, ZN => n21371);
   U23667 : NAND2_X1 port map( A1 => n21692, A2 => n28440, ZN => n21345);
   U23668 : OAI21_X1 port map( B1 => n21346, B2 => n21345, A => n21344, ZN => 
                           n21352);
   U23670 : NOR2_X1 port map( A1 => n21348, A2 => n21698, ZN => n21349);
   U23672 : NOR2_X2 port map( A1 => n21352, A2 => n21351, ZN => n22380);
   U23673 : MUX2_X1 port map( A => n21713, B => n21714, S => n21366, Z => 
                           n21369);
   U23674 : NAND2_X1 port map( A1 => n28491, A2 => n21354, ZN => n21358);
   U23675 : NAND2_X1 port map( A1 => n28126, A2 => n21354, ZN => n21357);
   U23676 : MUX2_X1 port map( A => n21358, B => n21357, S => n28133, Z => 
                           n21363);
   U23677 : NAND2_X1 port map( A1 => n21360, A2 => n28586, ZN => n21361);
   U23678 : NAND3_X1 port map( A1 => n21363, A2 => n21362, A3 => n21361, ZN => 
                           n21365);
   U23679 : AND2_X1 port map( A1 => n21364, A2 => n21365, ZN => n21368);
   U23680 : XNOR2_X1 port map( A => n22380, B => n22628, ZN => n21370);
   U23681 : XNOR2_X1 port map( A => n21371, B => n21370, ZN => n21386);
   U23682 : MUX2_X1 port map( A => n21373, B => n21372, S => n21704, Z => 
                           n21376);
   U23685 : INV_X1 port map( A => n22625, ZN => n21383);
   U23686 : XNOR2_X1 port map( A => n21384, B => n21383, ZN => n21385);
   U23687 : INV_X1 port map( A => n21389, ZN => n21476);
   U23688 : NAND2_X1 port map( A1 => n1930, A2 => n21476, ZN => n21390);
   U23689 : XNOR2_X1 port map( A => n22326, B => n22052, ZN => n21407);
   U23690 : NOR3_X1 port map( A1 => n21394, A2 => n21638, A3 => n21639, ZN => 
                           n21397);
   U23691 : NOR2_X1 port map( A1 => n21639, A2 => n21395, ZN => n21396);
   U23692 : NOR2_X1 port map( A1 => n21397, A2 => n21396, ZN => n21398);
   U23693 : NAND3_X1 port map( A1 => n21401, A2 => n21400, A3 => n21399, ZN => 
                           n21405);
   U23694 : OAI21_X1 port map( B1 => n21749, B2 => n20658, A => n21748, ZN => 
                           n21404);
   U23695 : NOR3_X1 port map( A1 => n21749, A2 => n21402, A3 => n497, ZN => 
                           n21403);
   U23696 : XNOR2_X1 port map( A => n22158, B => n22411, ZN => n22325);
   U23697 : INV_X1 port map( A => n22325, ZN => n21406);
   U23698 : XNOR2_X1 port map( A => n21407, B => n21406, ZN => n21419);
   U23699 : OAI21_X1 port map( B1 => n21410, B2 => n21409, A => n21408, ZN => 
                           n21411);
   U23700 : XNOR2_X1 port map( A => n22912, B => n22473, ZN => n21417);
   U23701 : XNOR2_X1 port map( A => n22844, B => n1179, ZN => n21416);
   U23702 : XNOR2_X1 port map( A => n21417, B => n21416, ZN => n21418);
   U23704 : OAI21_X1 port map( B1 => n23344, B2 => n23338, A => n28570, ZN => 
                           n21529);
   U23705 : NAND2_X1 port map( A1 => n21421, A2 => n21425, ZN => n21423);
   U23706 : NAND2_X1 port map( A1 => n21423, A2 => n21422, ZN => n21427);
   U23707 : XNOR2_X1 port map( A => n22897, B => n22434, ZN => n21446);
   U23708 : MUX2_X1 port map( A => n21664, B => n22398, S => n21429, Z => 
                           n21430);
   U23709 : NOR2_X1 port map( A1 => n21430, A2 => n22404, ZN => n21434);
   U23710 : NOR2_X1 port map( A1 => n21014, A2 => n21433, ZN => n22396);
   U23711 : NAND2_X1 port map( A1 => n21653, A2 => n21657, ZN => n21445);
   U23712 : INV_X1 port map( A => n21435, ZN => n21436);
   U23713 : NOR2_X1 port map( A1 => n21437, A2 => n21436, ZN => n21438);
   U23714 : NAND2_X1 port map( A1 => n21443, A2 => n21656, ZN => n21444);
   U23715 : XNOR2_X1 port map( A => n22333, B => n22479, ZN => n21876);
   U23716 : XNOR2_X1 port map( A => n21446, B => n21876, ZN => n21456);
   U23717 : INV_X1 port map( A => n21447, ZN => n21452);
   U23718 : OAI21_X1 port map( B1 => n21677, B2 => n21674, A => n21680, ZN => 
                           n21451);
   U23719 : NOR2_X1 port map( A1 => n21673, A2 => n21674, ZN => n21450);
   U23720 : INV_X1 port map( A => n891, ZN => n27788);
   U23721 : XNOR2_X1 port map( A => n22334, B => n27788, ZN => n21453);
   U23722 : XNOR2_X1 port map( A => n21454, B => n21453, ZN => n21455);
   U23725 : XNOR2_X1 port map( A => n22605, B => n22677, ZN => n21970);
   U23726 : XNOR2_X1 port map( A => n21470, B => n21970, ZN => n21492);
   U23727 : NAND2_X1 port map( A1 => n21473, A2 => n21472, ZN => n21474);
   U23728 : NAND2_X1 port map( A1 => n21475, A2 => n21474, ZN => n21480);
   U23729 : NAND2_X1 port map( A1 => n21477, A2 => n21476, ZN => n21479);
   U23730 : XNOR2_X1 port map( A => n22610, B => n22068, ZN => n21490);
   U23734 : XNOR2_X1 port map( A => n21889, B => n2912, ZN => n21489);
   U23735 : XNOR2_X1 port map( A => n21490, B => n21489, ZN => n21491);
   U23737 : AOI21_X1 port map( B1 => n21501, B2 => n21500, A => n21499, ZN => 
                           n21508);
   U23739 : NOR2_X1 port map( A1 => n21503, A2 => n28185, ZN => n21506);
   U23740 : INV_X1 port map( A => n21504, ZN => n21505);
   U23742 : XNOR2_X1 port map( A => n22374, B => n22619, ZN => n21523);
   U23743 : NAND3_X1 port map( A1 => n21509, A2 => n21513, A3 => n21514, ZN => 
                           n21510);
   U23744 : NAND2_X1 port map( A1 => n21511, A2 => n21510, ZN => n21518);
   U23745 : NAND2_X1 port map( A1 => n21520, A2 => n21551, ZN => n21521);
   U23746 : INV_X1 port map( A => n22567, ZN => n22487);
   U23747 : XNOR2_X1 port map( A => n22487, B => n22615, ZN => n21881);
   U23748 : XNOR2_X1 port map( A => n21881, B => n21523, ZN => n21527);
   U23749 : XNOR2_X1 port map( A => n22059, B => n5490, ZN => n21524);
   U23750 : XNOR2_X1 port map( A => n21525, B => n21524, ZN => n21526);
   U23751 : XNOR2_X1 port map( A => n21527, B => n21526, ZN => n23138);
   U23752 : OAI21_X1 port map( B1 => n29108, B2 => n28659, A => n23139, ZN => 
                           n21528);
   U23753 : XNOR2_X1 port map( A => n22522, B => n21537, ZN => n21546);
   U23754 : NAND2_X1 port map( A1 => n21540, A2 => n21539, ZN => n21542);
   U23755 : XNOR2_X1 port map( A => n22594, B => n21980, ZN => n21545);
   U23757 : OAI21_X1 port map( B1 => n21551, B2 => n21550, A => n21549, ZN => 
                           n21555);
   U23758 : INV_X1 port map( A => n21552, ZN => n21554);
   U23759 : XNOR2_X1 port map( A => n22768, B => n22829, ZN => n22313);
   U23760 : XNOR2_X1 port map( A => n21982, B => n22033, ZN => n21557);
   U23761 : XNOR2_X1 port map( A => n22313, B => n21557, ZN => n21558);
   U23762 : XNOR2_X2 port map( A => n21558, B => n21559, ZN => n23662);
   U23763 : AND2_X1 port map( A1 => n21561, A2 => n21560, ZN => n21562);
   U23764 : XNOR2_X1 port map( A => n22887, B => n27894, ZN => n21566);
   U23765 : INV_X1 port map( A => n21568, ZN => n21569);
   U23766 : XNOR2_X1 port map( A => n22656, B => n22891, ZN => n21573);
   U23767 : NOR2_X1 port map( A1 => n21575, A2 => n21574, ZN => n21578);
   U23768 : XNOR2_X1 port map( A => n21987, B => n22059, ZN => n21582);
   U23769 : XNOR2_X1 port map( A => n21582, B => n22619, ZN => n21583);
   U23770 : INV_X1 port map( A => n22644, ZN => n21593);
   U23771 : XNOR2_X1 port map( A => n21998, B => n21593, ZN => n21595);
   U23772 : XNOR2_X1 port map( A => n22692, B => n2544, ZN => n21594);
   U23773 : XNOR2_X1 port map( A => n21595, B => n21594, ZN => n21622);
   U23774 : NOR2_X1 port map( A1 => n21601, A2 => n21600, ZN => n21602);
   U23775 : NAND2_X1 port map( A1 => n21603, A2 => n21602, ZN => n21604);
   U23776 : NAND3_X1 port map( A1 => n21608, A2 => n21607, A3 => n21613, ZN => 
                           n21617);
   U23777 : INV_X1 port map( A => n21611, ZN => n21615);
   U23778 : NAND2_X1 port map( A1 => n21613, A2 => n21612, ZN => n21614);
   U23779 : XNOR2_X1 port map( A => n22500, B => n22813, ZN => n22899);
   U23780 : XNOR2_X1 port map( A => n22899, B => n21620, ZN => n21621);
   U23781 : XNOR2_X1 port map( A => n21621, B => n21622, ZN => n23162);
   U23782 : AOI21_X1 port map( B1 => n22146, B2 => n22145, A => n21623, ZN => 
                           n21628);
   U23783 : INV_X1 port map( A => n22717, ZN => n21800);
   U23784 : XNOR2_X1 port map( A => n21800, B => n22606, ZN => n21630);
   U23785 : XNOR2_X1 port map( A => n22068, B => n2389, ZN => n21629);
   U23786 : XNOR2_X1 port map( A => n21630, B => n21629, ZN => n21652);
   U23787 : NOR2_X1 port map( A1 => n21633, A2 => n21632, ZN => n21636);
   U23788 : AOI21_X1 port map( B1 => n21639, B2 => n21636, A => n21635, ZN => 
                           n21641);
   U23789 : OR3_X1 port map( A1 => n21639, A2 => n21638, A3 => n21637, ZN => 
                           n21640);
   U23790 : XNOR2_X1 port map( A => n22180, B => n22678, ZN => n22341);
   U23791 : NAND2_X1 port map( A1 => n21042, A2 => n21642, ZN => n21644);
   U23792 : NAND2_X1 port map( A1 => n21750, A2 => n21645, ZN => n21647);
   U23793 : XNOR2_X1 port map( A => n22067, B => n21649, ZN => n22181);
   U23794 : INV_X1 port map( A => n22181, ZN => n21650);
   U23795 : XNOR2_X1 port map( A => n22341, B => n21650, ZN => n21651);
   U23796 : XNOR2_X1 port map( A => n21651, B => n21652, ZN => n23006);
   U23797 : INV_X1 port map( A => n23006, ZN => n23665);
   U23798 : OAI21_X1 port map( B1 => n23666, B2 => n23162, A => n23665, ZN => 
                           n21690);
   U23799 : NOR2_X1 port map( A1 => n23666, A2 => n23006, ZN => n23164);
   U23800 : NOR2_X1 port map( A1 => n21654, A2 => n21653, ZN => n21659);
   U23801 : NOR2_X1 port map( A1 => n21656, A2 => n21655, ZN => n21658);
   U23802 : NOR2_X1 port map( A1 => n21662, A2 => n22401, ZN => n21668);
   U23803 : NOR2_X1 port map( A1 => n21664, A2 => n21663, ZN => n21669);
   U23804 : NOR2_X1 port map( A1 => n21665, A2 => n22397, ZN => n21666);
   U23805 : NOR2_X1 port map( A1 => n21669, A2 => n21666, ZN => n21667);
   U23807 : XNOR2_X1 port map( A => n22574, B => n22542, ZN => n22193);
   U23808 : XNOR2_X1 port map( A => n21671, B => n22193, ZN => n21689);
   U23809 : XNOR2_X1 port map( A => n22710, B => n22625, ZN => n21687);
   U23810 : INV_X1 port map( A => n21672, ZN => n21685);
   U23811 : OAI21_X1 port map( B1 => n21675, B2 => n21674, A => n21673, ZN => 
                           n21684);
   U23812 : NAND2_X1 port map( A1 => n21677, A2 => n21676, ZN => n21682);
   U23813 : NAND2_X1 port map( A1 => n21679, A2 => n21678, ZN => n21681);
   U23814 : MUX2_X1 port map( A => n21682, B => n21681, S => n21680, Z => 
                           n21683);
   U23815 : XNOR2_X1 port map( A => n22221, B => n3787, ZN => n21686);
   U23816 : XNOR2_X1 port map( A => n21687, B => n21686, ZN => n21688);
   U23817 : XNOR2_X1 port map( A => n21689, B => n21688, ZN => n23163);
   U23818 : AOI22_X1 port map( A1 => n23662, A2 => n21690, B1 => n23164, B2 => 
                           n23163, ZN => n21725);
   U23819 : INV_X1 port map( A => n21691, ZN => n21693);
   U23820 : INV_X1 port map( A => n21692, ZN => n21694);
   U23821 : NOR2_X1 port map( A1 => n21693, A2 => n21694, ZN => n21701);
   U23822 : NOR2_X1 port map( A1 => n21695, A2 => n21694, ZN => n21700);
   U23823 : AOI21_X1 port map( B1 => n21698, B2 => n21697, A => n3260, ZN => 
                           n21699);
   U23824 : XNOR2_X1 port map( A => n21872, B => n22734, ZN => n21719);
   U23825 : NAND3_X1 port map( A1 => n21705, A2 => n21704, A3 => n21703, ZN => 
                           n21706);
   U23826 : NOR2_X1 port map( A1 => n21709, A2 => n21708, ZN => n21710);
   U23827 : NOR2_X2 port map( A1 => n21711, A2 => n21710, ZN => n22589);
   U23828 : AOI21_X1 port map( B1 => n21714, B2 => n21713, A => n21712, ZN => 
                           n21715);
   U23829 : OAI22_X1 port map( A1 => n21718, A2 => n21717, B1 => n21716, B2 => 
                           n21715, ZN => n22535);
   U23830 : XNOR2_X1 port map( A => n22589, B => n22535, ZN => n22908);
   U23831 : XNOR2_X1 port map( A => n22908, B => n21719, ZN => n21723);
   U23832 : XNOR2_X1 port map( A => n22052, B => n22411, ZN => n21721);
   U23833 : INV_X1 port map( A => n3212, ZN => n27936);
   U23834 : XNOR2_X1 port map( A => n22328, B => n27936, ZN => n21720);
   U23835 : XNOR2_X1 port map( A => n21720, B => n21721, ZN => n21722);
   U23836 : XNOR2_X1 port map( A => n21723, B => n21722, ZN => n23525);
   U23837 : NAND2_X1 port map( A1 => n29123, A2 => n23163, ZN => n21898);
   U23839 : MUX2_X1 port map( A => n493, B => n29314, S => n1930, Z => n21737);
   U23840 : INV_X1 port map( A => n21731, ZN => n21732);
   U23841 : NAND2_X1 port map( A1 => n21732, A2 => n21736, ZN => n21735);
   U23842 : NAND2_X1 port map( A1 => n21733, A2 => n493, ZN => n21734);
   U23843 : OAI211_X1 port map( C1 => n21737, C2 => n21736, A => n21735, B => 
                           n21734, ZN => n21738);
   U23844 : XNOR2_X1 port map( A => n22643, B => n3323, ZN => n21740);
   U23845 : XNOR2_X1 port map( A => n21739, B => n21740, ZN => n21741);
   U23846 : XNOR2_X1 port map( A => n21741, B => n21742, ZN => n23783);
   U23847 : INV_X1 port map( A => n23783, ZN => n23785);
   U23848 : INV_X1 port map( A => n22426, ZN => n21743);
   U23849 : XNOR2_X1 port map( A => n21743, B => n21801, ZN => n22749);
   U23850 : XNOR2_X1 port map( A => n22609, B => n22553, ZN => n22037);
   U23851 : XNOR2_X1 port map( A => n22749, B => n22037, ZN => n21747);
   U23852 : XNOR2_X1 port map( A => n22681, B => n29490, ZN => n21745);
   U23853 : INV_X1 port map( A => n22006, ZN => n22515);
   U23854 : INV_X1 port map( A => n2441, ZN => n26314);
   U23855 : XNOR2_X1 port map( A => n22515, B => n26314, ZN => n21744);
   U23856 : XNOR2_X1 port map( A => n21745, B => n21744, ZN => n21746);
   U23858 : INV_X1 port map( A => n21825, ZN => n22285);
   U23859 : XNOR2_X1 port map( A => n22285, B => n22526, ZN => n21755);
   U23860 : MUX2_X1 port map( A => n21749, B => n21042, S => n21748, Z => 
                           n21752);
   U23861 : MUX2_X1 port map( A => n21752, B => n21751, S => n21750, Z => 
                           n22584);
   U23862 : XNOR2_X1 port map( A => n22199, B => n2476, ZN => n21753);
   U23863 : XNOR2_X1 port map( A => n21753, B => n22584, ZN => n21754);
   U23864 : XNOR2_X1 port map( A => n21755, B => n21754, ZN => n21757);
   U23865 : INV_X1 port map( A => n21758, ZN => n22786);
   U23866 : INV_X1 port map( A => n22195, ZN => n21759);
   U23867 : XNOR2_X1 port map( A => n22786, B => n21759, ZN => n21761);
   U23868 : XNOR2_X1 port map( A => n22218, B => n22790, ZN => n22015);
   U23869 : XNOR2_X1 port map( A => n28449, B => n72, ZN => n21762);
   U23870 : XNOR2_X1 port map( A => n22015, B => n21762, ZN => n21763);
   U23871 : XNOR2_X1 port map( A => n21764, B => n21763, ZN => n23784);
   U23872 : XNOR2_X1 port map( A => n22409, B => n3087, ZN => n21765);
   U23873 : XNOR2_X1 port map( A => n22601, B => n28589, ZN => n21767);
   U23874 : XNOR2_X1 port map( A => n22472, B => n21767, ZN => n22048);
   U23875 : XNOR2_X1 port map( A => n21768, B => n22048, ZN => n21775);
   U23876 : INV_X1 port map( A => n22798, ZN => n22422);
   U23877 : XNOR2_X1 port map( A => n22422, B => n22418, ZN => n21770);
   U23878 : XNOR2_X1 port map( A => n22796, B => n21959, ZN => n22569);
   U23879 : XNOR2_X1 port map( A => n21770, B => n22569, ZN => n21774);
   U23880 : XNOR2_X1 port map( A => n28492, B => n1123, ZN => n21772);
   U23882 : XNOR2_X1 port map( A => n22509, B => n22724, ZN => n21771);
   U23883 : XNOR2_X1 port map( A => n21772, B => n21771, ZN => n21773);
   U23884 : XNOR2_X1 port map( A => n21774, B => n21773, ZN => n23786);
   U23885 : INV_X1 port map( A => n23786, ZN => n23005);
   U23886 : INV_X1 port map( A => n21775, ZN => n23482);
   U23887 : AOI211_X1 port map( C1 => n23005, C2 => n23482, A => n23484, B => 
                           n23036, ZN => n21776);
   U23888 : XNOR2_X1 port map( A => n22710, B => n22086, ZN => n21778);
   U23889 : XNOR2_X1 port map( A => n28517, B => n22786, ZN => n21777);
   U23890 : XNOR2_X1 port map( A => n21778, B => n21777, ZN => n21782);
   U23891 : INV_X1 port map( A => n22835, ZN => n21995);
   U23892 : XNOR2_X1 port map( A => n21995, B => n22219, ZN => n21780);
   U23893 : XNOR2_X1 port map( A => n21780, B => n21779, ZN => n21781);
   U23894 : XNOR2_X1 port map( A => n22757, B => n22052, ZN => n21784);
   U23895 : XNOR2_X1 port map( A => n28461, B => n22734, ZN => n21783);
   U23896 : XNOR2_X1 port map( A => n21784, B => n21783, ZN => n21788);
   U23897 : XNOR2_X1 port map( A => n22763, B => n3650, ZN => n21785);
   U23898 : XNOR2_X1 port map( A => n21786, B => n21785, ZN => n21787);
   U23899 : XNOR2_X2 port map( A => n21788, B => n21787, ZN => n23765);
   U23900 : AND2_X1 port map( A1 => n23767, A2 => n23765, ZN => n21829);
   U23901 : XNOR2_X1 port map( A => n21789, B => n22245, ZN => n21792);
   U23902 : INV_X1 port map( A => n22363, ZN => n21790);
   U23903 : XNOR2_X1 port map( A => n21956, B => n21790, ZN => n21791);
   U23904 : XNOR2_X1 port map( A => n22812, B => n22692, ZN => n21794);
   U23905 : XNOR2_X1 port map( A => n22778, B => n2602, ZN => n21793);
   U23906 : XNOR2_X1 port map( A => n21794, B => n21793, ZN => n21795);
   U23907 : XNOR2_X1 port map( A => n22821, B => n22059, ZN => n22617);
   U23908 : XNOR2_X1 port map( A => n22728, B => n22617, ZN => n21799);
   U23909 : XNOR2_X1 port map( A => n21959, B => n1859, ZN => n21797);
   U23910 : XNOR2_X1 port map( A => n22488, B => n3770, ZN => n21796);
   U23911 : XNOR2_X1 port map( A => n21797, B => n21796, ZN => n21798);
   U23912 : XNOR2_X1 port map( A => n22068, B => n2404, ZN => n21804);
   U23913 : XNOR2_X1 port map( A => n21800, B => n21801, ZN => n22259);
   U23914 : INV_X1 port map( A => n22718, ZN => n21802);
   U23915 : XNOR2_X1 port map( A => n22259, B => n21802, ZN => n21803);
   U23916 : NAND3_X1 port map( A1 => n21808, A2 => n21807, A3 => n21806, ZN => 
                           n21815);
   U23917 : OAI21_X1 port map( B1 => n21811, B2 => n21810, A => n21809, ZN => 
                           n21814);
   U23918 : INV_X1 port map( A => n21812, ZN => n21813);
   U23919 : AOI21_X1 port map( B1 => n21815, B2 => n21814, A => n21813, ZN => 
                           n22370);
   U23920 : XNOR2_X1 port map( A => n21816, B => n22370, ZN => n22008);
   U23921 : INV_X1 port map( A => n22703, ZN => n21817);
   U23923 : INV_X1 port map( A => n21818, ZN => n21822);
   U23924 : NOR2_X1 port map( A1 => n491, A2 => n22013, ZN => n21820);
   U23925 : AOI22_X1 port map( A1 => n21823, A2 => n21820, B1 => n21819, B2 => 
                           n22013, ZN => n21821);
   U23926 : OAI21_X1 port map( B1 => n21823, B2 => n21822, A => n21821, ZN => 
                           n21824);
   U23927 : XNOR2_X1 port map( A => n21979, B => n21824, ZN => n22390);
   U23928 : INV_X1 port map( A => n22390, ZN => n21828);
   U23929 : XNOR2_X1 port map( A => n22033, B => n22226, ZN => n22524);
   U23930 : XNOR2_X1 port map( A => n22524, B => n21826, ZN => n21827);
   U23931 : NOR2_X1 port map( A1 => n23501, A2 => n23499, ZN => n21830);
   U23932 : XNOR2_X1 port map( A => n22204, B => n22265, ZN => n22642);
   U23933 : XNOR2_X1 port map( A => n28387, B => n22898, ZN => n21831);
   U23934 : XNOR2_X1 port map( A => n22642, B => n21831, ZN => n21835);
   U23935 : XNOR2_X1 port map( A => n22330, B => n22501, ZN => n21833);
   U23936 : XNOR2_X1 port map( A => n22334, B => n3386, ZN => n21832);
   U23937 : XNOR2_X1 port map( A => n21833, B => n21832, ZN => n21834);
   U23939 : XNOR2_X1 port map( A => n22326, B => n2353, ZN => n21836);
   U23941 : XNOR2_X1 port map( A => n22302, B => n22409, ZN => n22650);
   U23942 : XNOR2_X1 port map( A => n21838, B => n22650, ZN => n21839);
   U23943 : XNOR2_X1 port map( A => n22374, B => n21841, ZN => n21842);
   U23944 : XNOR2_X1 port map( A => n22100, B => n21842, ZN => n21846);
   U23945 : XNOR2_X1 port map( A => n22822, B => n22890, ZN => n21844);
   U23946 : XNOR2_X1 port map( A => n22506, B => n3211, ZN => n21843);
   U23947 : XNOR2_X1 port map( A => n21844, B => n21843, ZN => n21845);
   U23948 : NOR2_X1 port map( A1 => n339, A2 => n23772, ZN => n21853);
   U23949 : XNOR2_X1 port map( A => n22386, B => n3083, ZN => n21849);
   U23950 : XNOR2_X1 port map( A => n22199, B => n21850, ZN => n22675);
   U23951 : INV_X1 port map( A => n22675, ZN => n21851);
   U23952 : INV_X1 port map( A => n23156, ZN => n23512);
   U23953 : AOI22_X1 port map( A1 => n23488, A2 => n23513, B1 => n21853, B2 => 
                           n23512, ZN => n21864);
   U23954 : XNOR2_X1 port map( A => n22240, B => n29489, ZN => n21854);
   U23955 : XNOR2_X1 port map( A => n21854, B => n22340, ZN => n22684);
   U23956 : XNOR2_X1 port map( A => n22514, B => n22854, ZN => n21855);
   U23957 : XNOR2_X1 port map( A => n22164, B => n21856, ZN => n21860);
   U23958 : XNOR2_X1 port map( A => n22380, B => n27422, ZN => n21858);
   U23959 : INV_X1 port map( A => n22279, ZN => n21857);
   U23960 : XNOR2_X1 port map( A => n22195, B => n21857, ZN => n22663);
   U23961 : XNOR2_X1 port map( A => n22663, B => n21858, ZN => n21859);
   U23962 : XNOR2_X1 port map( A => n21859, B => n21860, ZN => n23771);
   U23963 : INV_X1 port map( A => n23771, ZN => n23487);
   U23964 : NOR2_X1 port map( A1 => n23487, A2 => n23772, ZN => n21861);
   U23967 : XNOR2_X1 port map( A => n22194, B => n22221, ZN => n21912);
   U23968 : XNOR2_X1 port map( A => n22278, B => n22380, ZN => n22839);
   U23969 : XNOR2_X1 port map( A => n22839, B => n21912, ZN => n21868);
   U23970 : XNOR2_X1 port map( A => n22464, B => n22784, ZN => n22578);
   U23971 : XNOR2_X1 port map( A => n22628, B => n21865, ZN => n21866);
   U23972 : XNOR2_X1 port map( A => n22578, B => n21866, ZN => n21867);
   U23973 : XNOR2_X1 port map( A => n21868, B => n21867, ZN => n23802);
   U23974 : INV_X1 port map( A => n23802, ZN => n23541);
   U23975 : XNOR2_X1 port map( A => n22158, B => n3336, ZN => n21870);
   U23976 : XNOR2_X1 port map( A => n22326, B => n22414, ZN => n22843);
   U23978 : XNOR2_X1 port map( A => n21870, B => n28613, ZN => n21874);
   U23979 : XNOR2_X1 port map( A => n21871, B => n21872, ZN => n21918);
   U23980 : XNOR2_X1 port map( A => n28162, B => n22473, ZN => n22588);
   U23981 : XNOR2_X1 port map( A => n22588, B => n21918, ZN => n21873);
   U23982 : XNOR2_X1 port map( A => n21998, B => n21875, ZN => n21940);
   U23983 : INV_X1 port map( A => n21940, ZN => n21877);
   U23984 : XNOR2_X1 port map( A => n22690, B => n29247, ZN => n21878);
   U23985 : XNOR2_X1 port map( A => n21987, B => n22098, ZN => n21880);
   U23986 : XNOR2_X1 port map( A => n22723, B => n2511, ZN => n21879);
   U23987 : XNOR2_X1 port map( A => n21880, B => n21879, ZN => n21883);
   U23988 : XNOR2_X1 port map( A => n22374, B => n22419, ZN => n22819);
   U23989 : INV_X1 port map( A => n22819, ZN => n22057);
   U23990 : XNOR2_X1 port map( A => n22057, B => n21881, ZN => n21882);
   U23991 : XNOR2_X1 port map( A => n22298, B => n22386, ZN => n22827);
   U23992 : XNOR2_X1 port map( A => n22827, B => n21884, ZN => n21887);
   U23993 : XNOR2_X1 port map( A => n21980, B => n3554, ZN => n21885);
   U23994 : XNOR2_X1 port map( A => n22152, B => n29514, ZN => n21947);
   U23995 : XNOR2_X1 port map( A => n21885, B => n21947, ZN => n21886);
   U23996 : XNOR2_X2 port map( A => n21887, B => n21886, ZN => n23689);
   U23997 : XNOR2_X1 port map( A => n22606, B => n22855, ZN => n21888);
   U23998 : XNOR2_X1 port map( A => n21970, B => n21888, ZN => n21892);
   U23999 : INV_X1 port map( A => n22852, ZN => n22065);
   U24000 : XNOR2_X1 port map( A => n22750, B => n3062, ZN => n21890);
   U24001 : XNOR2_X1 port map( A => n22065, B => n21890, ZN => n21891);
   U24002 : INV_X1 port map( A => n23800, ZN => n21893);
   U24003 : OAI22_X1 port map( A1 => n21895, A2 => n23690, B1 => n23803, B2 => 
                           n21894, ZN => n23932);
   U24004 : INV_X1 port map( A => n23932, ZN => n24728);
   U24005 : OR2_X1 port map( A1 => n24596, A2 => n24728, ZN => n24732);
   U24007 : INV_X1 port map( A => n23666, ZN => n21896);
   U24008 : NAND2_X1 port map( A1 => n28577, A2 => n21896, ZN => n21897);
   U24009 : MUX2_X1 port map( A => n21898, B => n21897, S => n23162, Z => 
                           n21901);
   U24010 : NOR2_X1 port map( A1 => n23163, A2 => n23663, ZN => n21899);
   U24011 : NOR2_X1 port map( A1 => n23162, A2 => n23006, ZN => n23669);
   U24012 : AOI21_X1 port map( B1 => n23662, B2 => n21899, A => n23669, ZN => 
                           n21900);
   U24013 : NAND2_X1 port map( A1 => n21901, A2 => n21900, ZN => n24595);
   U24014 : INV_X1 port map( A => n24595, ZN => n24288);
   U24015 : NAND2_X1 port map( A1 => n24732, A2 => n24724, ZN => n21943);
   U24016 : XNOR2_X1 port map( A => n22820, B => n22891, ZN => n22061);
   U24017 : XNOR2_X1 port map( A => n22061, B => n22098, ZN => n22213);
   U24018 : XNOR2_X1 port map( A => n21902, B => n22888, ZN => n21904);
   U24019 : XNOR2_X1 port map( A => n21904, B => n22620, ZN => n21905);
   U24020 : XNOR2_X1 port map( A => n29591, B => n22606, ZN => n21907);
   U24021 : XNOR2_X1 port map( A => n22338, B => n22067, ZN => n22905);
   U24022 : INV_X1 port map( A => n22905, ZN => n21906);
   U24023 : XNOR2_X1 port map( A => n21906, B => n21907, ZN => n21911);
   U24024 : XNOR2_X1 port map( A => n22718, B => n22856, ZN => n21909);
   U24025 : XNOR2_X1 port map( A => n22855, B => n27105, ZN => n21908);
   U24026 : XNOR2_X1 port map( A => n21909, B => n21908, ZN => n21910);
   U24027 : XNOR2_X1 port map( A => n22320, B => n22542, ZN => n22920);
   U24028 : XNOR2_X1 port map( A => n21912, B => n22920, ZN => n21916);
   U24029 : XNOR2_X1 port map( A => n22123, B => n22219, ZN => n21914);
   U24030 : XNOR2_X1 port map( A => n22664, B => n1247, ZN => n21913);
   U24031 : XNOR2_X1 port map( A => n21914, B => n21913, ZN => n21915);
   U24034 : XNOR2_X1 port map( A => n21917, B => n22535, ZN => n22187);
   U24035 : XNOR2_X1 port map( A => n21918, B => n22187, ZN => n21922);
   U24036 : XNOR2_X1 port map( A => n22731, B => n28461, ZN => n21920);
   U24037 : XNOR2_X1 port map( A => n28472, B => n3035, ZN => n21919);
   U24038 : XNOR2_X1 port map( A => n21920, B => n21919, ZN => n21921);
   U24039 : XNOR2_X1 port map( A => n21922, B => n21921, ZN => n23793);
   U24040 : XNOR2_X1 port map( A => n22697, B => n22523, ZN => n21924);
   U24041 : XNOR2_X1 port map( A => n22828, B => n21924, ZN => n21928);
   U24042 : XNOR2_X1 port map( A => n21980, B => n22387, ZN => n22595);
   U24043 : INV_X1 port map( A => n22595, ZN => n21926);
   U24044 : XNOR2_X1 port map( A => n22522, B => n3565, ZN => n21925);
   U24045 : XNOR2_X1 port map( A => n21926, B => n21925, ZN => n21927);
   U24046 : NAND2_X1 port map( A1 => n29586, A2 => n21932, ZN => n21933);
   U24047 : OAI22_X1 port map( A1 => n21934, A2 => n21933, B1 => n21932, B2 => 
                           n21931, ZN => n21935);
   U24048 : INV_X1 port map( A => n22205, ZN => n22080);
   U24049 : XNOR2_X1 port map( A => n22094, B => n22245, ZN => n21938);
   U24050 : XNOR2_X1 port map( A => n22080, B => n21938, ZN => n21942);
   U24051 : XNOR2_X1 port map( A => n22896, B => n2598, ZN => n21939);
   U24052 : XOR2_X1 port map( A => n21940, B => n21939, Z => n21941);
   U24055 : XNOR2_X1 port map( A => n22582, B => n21946, ZN => n21948);
   U24056 : XNOR2_X1 port map( A => n22158, B => n22760, ZN => n22117);
   U24057 : XNOR2_X1 port map( A => n21949, B => n22301, ZN => n22587);
   U24058 : XNOR2_X1 port map( A => n22117, B => n22587, ZN => n21953);
   U24059 : XNOR2_X1 port map( A => n22535, B => n22473, ZN => n21951);
   U24060 : XNOR2_X1 port map( A => n22414, B => n1215, ZN => n21950);
   U24061 : XNOR2_X1 port map( A => n21951, B => n21950, ZN => n21952);
   U24063 : NAND2_X1 port map( A1 => n23606, A2 => n23247, ZN => n23211);
   U24065 : XNOR2_X1 port map( A => n22479, B => n22330, ZN => n22641);
   U24066 : XNOR2_X1 port map( A => n22500, B => n3463, ZN => n21954);
   U24067 : XNOR2_X1 port map( A => n22641, B => n21954, ZN => n21958);
   U24068 : XNOR2_X1 port map( A => n21956, B => n21955, ZN => n22264);
   U24069 : XNOR2_X1 port map( A => n22333, B => n22644, ZN => n22092);
   U24070 : XNOR2_X1 port map( A => n22264, B => n22092, ZN => n21957);
   U24071 : XNOR2_X1 port map( A => n21957, B => n21958, ZN => n23245);
   U24072 : XNOR2_X1 port map( A => n22419, B => n21959, ZN => n22272);
   U24073 : XNOR2_X1 port map( A => n22272, B => n22350, ZN => n21963);
   U24074 : XNOR2_X1 port map( A => n22567, B => n22891, ZN => n21961);
   U24075 : XNOR2_X1 port map( A => n28483, B => n3728, ZN => n21960);
   U24076 : XNOR2_X1 port map( A => n21961, B => n21960, ZN => n21962);
   U24077 : XNOR2_X1 port map( A => n21963, B => n21962, ZN => n23246);
   U24078 : INV_X1 port map( A => n23246, ZN => n23603);
   U24081 : XNOR2_X1 port map( A => n22278, B => n22542, ZN => n21967);
   U24082 : INV_X1 port map( A => n2477, ZN => n26287);
   U24083 : XNOR2_X1 port map( A => n22464, B => n26287, ZN => n21966);
   U24084 : XNOR2_X1 port map( A => n21967, B => n21966, ZN => n21969);
   U24085 : XNOR2_X1 port map( A => n22783, B => n22628, ZN => n22318);
   U24086 : XNOR2_X1 port map( A => n22575, B => n22318, ZN => n21968);
   U24087 : INV_X1 port map( A => n23607, ZN => n22985);
   U24088 : INV_X1 port map( A => n23247, ZN => n23578);
   U24089 : XNOR2_X1 port map( A => n21970, B => n21971, ZN => n21975);
   U24090 : XNOR2_X1 port map( A => n22678, B => n22067, ZN => n21973);
   U24091 : XNOR2_X1 port map( A => n6504, B => n1062, ZN => n21972);
   U24092 : XNOR2_X1 port map( A => n21973, B => n21972, ZN => n21974);
   U24093 : XNOR2_X1 port map( A => n21974, B => n21975, ZN => n23602);
   U24094 : INV_X1 port map( A => n23602, ZN => n23583);
   U24095 : OAI21_X1 port map( B1 => n22985, B2 => n23578, A => n23583, ZN => 
                           n21976);
   U24096 : NAND2_X1 port map( A1 => n21976, A2 => n23577, ZN => n21977);
   U24099 : XNOR2_X1 port map( A => n22671, B => n25044, ZN => n21984);
   U24100 : XNOR2_X1 port map( A => n21982, B => n22226, ZN => n21983);
   U24101 : XNOR2_X1 port map( A => n21984, B => n21983, ZN => n21985);
   U24102 : XNOR2_X1 port map( A => n21987, B => n22509, ZN => n22252);
   U24103 : XNOR2_X1 port map( A => n22252, B => n22821, ZN => n22886);
   U24104 : XNOR2_X1 port map( A => n22488, B => n1858, ZN => n21988);
   U24105 : XNOR2_X1 port map( A => n22886, B => n21989, ZN => n23258);
   U24106 : XNOR2_X1 port map( A => n22411, B => n22735, ZN => n22188);
   U24107 : XNOR2_X1 port map( A => n22599, B => n22188, ZN => n21993);
   U24108 : INV_X1 port map( A => n22472, ZN => n22300);
   U24109 : XNOR2_X1 port map( A => n22300, B => n4029, ZN => n21991);
   U24110 : XNOR2_X1 port map( A => n22533, B => n21991, ZN => n21992);
   U24111 : XNOR2_X1 port map( A => n22459, B => n22625, ZN => n22192);
   U24112 : XNOR2_X1 port map( A => n21994, B => n22792, ZN => n22220);
   U24113 : XNOR2_X1 port map( A => n22192, B => n22220, ZN => n21997);
   U24114 : XNOR2_X1 port map( A => n21995, B => n22221, ZN => n22922);
   U24115 : NAND2_X1 port map( A1 => n23735, A2 => n23227, ZN => n23734);
   U24116 : INV_X1 port map( A => n21998, ZN => n21999);
   U24117 : XNOR2_X1 port map( A => n22000, B => n21789, ZN => n22001);
   U24118 : XNOR2_X1 port map( A => n29136, B => n22001, ZN => n22005);
   U24119 : XNOR2_X1 port map( A => n22643, B => n22434, ZN => n22003);
   U24120 : XNOR2_X1 port map( A => n22778, B => n2916, ZN => n22002);
   U24121 : XNOR2_X1 port map( A => n22003, B => n22002, ZN => n22004);
   U24122 : XNOR2_X1 port map( A => n22606, B => n22006, ZN => n22238);
   U24123 : XNOR2_X1 port map( A => n22681, B => n26825, ZN => n22007);
   U24124 : AOI21_X1 port map( B1 => n22010, B2 => n23734, A => n22009, ZN => 
                           n23962);
   U24125 : AND2_X1 port map( A1 => n24583, A2 => n23962, ZN => n24586);
   U24126 : XNOR2_X1 port map( A => n22923, B => n22015, ZN => n22018);
   U24127 : XNOR2_X1 port map( A => n28450, B => n24897, ZN => n22016);
   U24128 : XNOR2_X1 port map( A => n22017, B => n22018, ZN => n22976);
   U24129 : INV_X1 port map( A => n22976, ZN => n23408);
   U24130 : XNOR2_X1 port map( A => n22633, B => n28387, ZN => n22020);
   U24131 : XNOR2_X1 port map( A => n21728, B => n3036, ZN => n22019);
   U24132 : XNOR2_X1 port map( A => n22020, B => n22019, ZN => n22021);
   U24136 : OAI211_X1 port map( C1 => n489, C2 => n21019, A => n22291, B => 
                           n22025, ZN => n22030);
   U24138 : INV_X1 port map( A => n1927, ZN => n28108);
   U24139 : OAI21_X1 port map( B1 => n22027, B2 => n22028, A => n28108, ZN => 
                           n22029);
   U24140 : XNOR2_X1 port map( A => n22031, B => n22032, ZN => n22036);
   U24141 : XNOR2_X1 port map( A => n22830, B => n22033, ZN => n22034);
   U24142 : XNOR2_X1 port map( A => n22034, B => n22523, ZN => n22035);
   U24143 : XNOR2_X1 port map( A => n22036, B => n22035, ZN => n22977);
   U24144 : MUX2_X1 port map( A => n23408, B => n23406, S => n23252, Z => 
                           n22051);
   U24146 : XNOR2_X1 port map( A => n22495, B => n22037, ZN => n22040);
   U24147 : XNOR2_X1 port map( A => n22854, B => n3154, ZN => n22038);
   U24148 : XNOR2_X1 port map( A => n22519, B => n22038, ZN => n22039);
   U24149 : XNOR2_X1 port map( A => n22040, B => n22039, ZN => n22979);
   U24150 : XNOR2_X1 port map( A => n22041, B => n22511, ZN => n22045);
   U24151 : XNOR2_X1 port map( A => n22796, B => n22822, ZN => n22043);
   U24152 : XNOR2_X1 port map( A => n22890, B => n3029, ZN => n22042);
   U24153 : XNOR2_X1 port map( A => n22043, B => n22042, ZN => n22044);
   U24154 : XNOR2_X1 port map( A => n22045, B => n22044, ZN => n23213);
   U24155 : INV_X1 port map( A => n23213, ZN => n22980);
   U24156 : MUX2_X1 port map( A => n22979, B => n22980, S => n28527, Z => 
                           n22050);
   U24157 : XNOR2_X1 port map( A => n29519, B => n1225, ZN => n22046);
   U24158 : XNOR2_X1 port map( A => n22046, B => n22913, ZN => n22047);
   U24159 : XNOR2_X1 port map( A => n22532, B => n22047, ZN => n22049);
   U24160 : INV_X1 port map( A => n24584, ZN => n24581);
   U24161 : XNOR2_X1 port map( A => n29087, B => n22187, ZN => n22056);
   U24162 : XNOR2_X1 port map( A => n22763, B => n3508, ZN => n22055);
   U24163 : XNOR2_X1 port map( A => n22057, B => n22058, ZN => n22063);
   U24164 : XNOR2_X1 port map( A => n22059, B => n3109, ZN => n22060);
   U24165 : XNOR2_X1 port map( A => n22061, B => n22060, ZN => n22062);
   U24166 : XNOR2_X1 port map( A => n22063, B => n22062, ZN => n23706);
   U24167 : XNOR2_X1 port map( A => n22856, B => n1248, ZN => n22064);
   U24168 : XNOR2_X1 port map( A => n22065, B => n22064, ZN => n22071);
   U24169 : XNOR2_X1 port map( A => n22066, B => n22067, ZN => n22518);
   U24170 : INV_X1 port map( A => n22518, ZN => n22069);
   U24171 : XNOR2_X1 port map( A => n22068, B => n22104, ZN => n22607);
   U24172 : XNOR2_X1 port map( A => n22069, B => n22607, ZN => n22070);
   U24173 : XNOR2_X1 port map( A => n22387, B => n22072, ZN => n22074);
   U24174 : XNOR2_X1 port map( A => n22074, B => n22073, ZN => n22075);
   U24175 : XNOR2_X1 port map( A => n22827, B => n22075, ZN => n22079);
   U24176 : XNOR2_X1 port map( A => n22670, B => n22522, ZN => n22076);
   U24177 : XNOR2_X1 port map( A => n22077, B => n22076, ZN => n22078);
   U24178 : XNOR2_X1 port map( A => n22079, B => n22078, ZN => n22451);
   U24180 : XNOR2_X1 port map( A => n22363, B => n22094, ZN => n22634);
   U24181 : XNOR2_X1 port map( A => n22080, B => n22634, ZN => n22083);
   U24182 : XNOR2_X1 port map( A => n22778, B => n2510, ZN => n22081);
   U24183 : XNOR2_X1 port map( A => n22081, B => n22809, ZN => n22082);
   U24185 : XNOR2_X1 port map( A => n22086, B => n22542, ZN => n22088);
   U24186 : XNOR2_X1 port map( A => n22123, B => n28517, ZN => n22626);
   U24187 : XNOR2_X1 port map( A => n22626, B => n22088, ZN => n22091);
   U24188 : XNOR2_X1 port map( A => n22664, B => n1246, ZN => n22089);
   U24189 : XNOR2_X1 port map( A => n22839, B => n22089, ZN => n22090);
   U24190 : XNOR2_X1 port map( A => n22091, B => n22090, ZN => n22452);
   U24191 : INV_X1 port map( A => n22452, ZN => n23220);
   U24192 : XNOR2_X1 port map( A => n22642, B => n22092, ZN => n22097);
   U24193 : XNOR2_X1 port map( A => n22093, B => n22813, ZN => n22207);
   U24194 : XNOR2_X1 port map( A => n22094, B => n3598, ZN => n22095);
   U24195 : XNOR2_X1 port map( A => n22207, B => n22095, ZN => n22096);
   U24196 : XNOR2_X1 port map( A => n22097, B => n22096, ZN => n22953);
   U24197 : XNOR2_X1 port map( A => n28409, B => n22099, ZN => n22818);
   U24198 : XNOR2_X1 port map( A => n22100, B => n22818, ZN => n22103);
   U24199 : XNOR2_X1 port map( A => n22350, B => n22101, ZN => n22102);
   U24200 : XNOR2_X1 port map( A => n22103, B => n22102, ZN => n22455);
   U24201 : XNOR2_X1 port map( A => n22104, B => n22240, ZN => n22105);
   U24202 : XNOR2_X1 port map( A => n22341, B => n22105, ZN => n22109);
   U24203 : XNOR2_X1 port map( A => n22428, B => n22605, ZN => n22107);
   U24204 : XNOR2_X1 port map( A => n22855, B => n26214, ZN => n22106);
   U24205 : XNOR2_X1 port map( A => n22107, B => n22106, ZN => n22108);
   U24206 : XNOR2_X1 port map( A => n22109, B => n22108, ZN => n23843);
   U24208 : INV_X1 port map( A => n22199, ZN => n22110);
   U24209 : XNOR2_X1 port map( A => n22313, B => n22111, ZN => n22115);
   U24210 : XNOR2_X1 port map( A => n22387, B => n22295, ZN => n22113);
   U24211 : XNOR2_X1 port map( A => n22152, B => n1172, ZN => n22112);
   U24212 : XNOR2_X1 port map( A => n22113, B => n22112, ZN => n22114);
   U24214 : XNOR2_X1 port map( A => n22589, B => n22116, ZN => n22842);
   U24215 : INV_X1 port map( A => n22842, ZN => n22118);
   U24217 : XNOR2_X1 port map( A => n22731, B => n2381, ZN => n22119);
   U24218 : XNOR2_X1 port map( A => n22119, B => n22650, ZN => n22120);
   U24221 : INV_X1 port map( A => n22455, ZN => n23722);
   U24222 : XNOR2_X1 port map( A => n22194, B => n3662, ZN => n22122);
   U24223 : XNOR2_X1 port map( A => n22663, B => n22122, ZN => n22126);
   U24224 : XNOR2_X1 port map( A => n22574, B => n22123, ZN => n22124);
   U24225 : XNOR2_X1 port map( A => n22318, B => n22124, ZN => n22125);
   U24226 : XNOR2_X1 port map( A => n22126, B => n22125, ZN => n22954);
   U24227 : NAND2_X1 port map( A1 => n22127, A2 => n23845, ZN => n22128);
   U24229 : INV_X1 port map( A => n24577, ZN => n23963);
   U24230 : MUX2_X1 port map( A => n24586, B => n22130, S => n23963, Z => 
                           n22179);
   U24231 : XNOR2_X1 port map( A => n22615, B => n22270, ZN => n22131);
   U24232 : XNOR2_X1 port map( A => n22486, B => n22131, ZN => n22135);
   U24233 : XNOR2_X1 port map( A => n22506, B => n2894, ZN => n22133);
   U24234 : XNOR2_X1 port map( A => n22571, B => n22133, ZN => n22134);
   U24235 : XNOR2_X1 port map( A => n22134, B => n22135, ZN => n22174);
   U24236 : INV_X1 port map( A => n22174, ZN => n23710);
   U24237 : XNOR2_X1 port map( A => n22514, B => n22240, ZN => n22261);
   U24238 : XNOR2_X1 port map( A => n22497, B => n22261, ZN => n22138);
   U24239 : XNOR2_X1 port map( A => n22605, B => n2505, ZN => n22136);
   U24240 : XNOR2_X1 port map( A => n22854, B => n22750, ZN => n22558);
   U24241 : XNOR2_X1 port map( A => n22136, B => n22558, ZN => n22137);
   U24242 : INV_X1 port map( A => n23712, ZN => n22971);
   U24243 : OAI21_X1 port map( B1 => n22140, B2 => n5339, A => n22139, ZN => 
                           n22149);
   U24244 : NOR2_X1 port map( A1 => n22142, A2 => n22141, ZN => n22148);
   U24245 : NAND2_X1 port map( A1 => n22146, A2 => n22143, ZN => n22144);
   U24246 : OAI211_X1 port map( C1 => n22146, C2 => n22145, A => n22144, B => 
                           n21624, ZN => n22147);
   U24247 : XNOR2_X1 port map( A => n22295, B => n22525, ZN => n22150);
   U24248 : XNOR2_X1 port map( A => n22151, B => n22150, ZN => n22156);
   U24249 : XNOR2_X1 port map( A => n22830, B => n29548, ZN => n22154);
   U24250 : XNOR2_X1 port map( A => n22152, B => n3385, ZN => n22153);
   U24251 : XNOR2_X1 port map( A => n22154, B => n22153, ZN => n22155);
   U24252 : XNOR2_X1 port map( A => n22157, B => n22474, ZN => n22162);
   U24253 : XNOR2_X1 port map( A => n22158, B => n2306, ZN => n22160);
   U24254 : XNOR2_X1 port map( A => n22159, B => n22160, ZN => n22161);
   U24255 : XNOR2_X1 port map( A => n22162, B => n22161, ZN => n23262);
   U24257 : XNOR2_X1 port map( A => n22164, B => n22461, ZN => n22168);
   U24258 : XNOR2_X1 port map( A => n22279, B => n22628, ZN => n22166);
   U24259 : XNOR2_X1 port map( A => n22784, B => n3491, ZN => n22165);
   U24260 : XNOR2_X1 port map( A => n22166, B => n22165, ZN => n22167);
   U24261 : XNOR2_X1 port map( A => n22168, B => n22167, ZN => n23233);
   U24262 : INV_X1 port map( A => n23233, ZN => n23585);
   U24263 : XNOR2_X1 port map( A => n22333, B => n22169, ZN => n22170);
   U24264 : XNOR2_X1 port map( A => n22265, B => n2995, ZN => n22171);
   U24265 : XNOR2_X1 port map( A => n22172, B => n22245, ZN => n22483);
   U24266 : OAI211_X1 port map( C1 => n23716, C2 => n23585, A => n23715, B => 
                           n23260, ZN => n22175);
   U24267 : MUX2_X1 port map( A => n24584, B => n24054, S => n29026, Z => 
                           n22177);
   U24269 : XNOR2_X1 port map( A => n22713, B => n22180, ZN => n22182);
   U24270 : XNOR2_X1 port map( A => n22181, B => n22182, ZN => n22186);
   U24271 : XNOR2_X1 port map( A => n22428, B => n22856, ZN => n22184);
   U24272 : XNOR2_X1 port map( A => n22855, B => Key(19), ZN => n22183);
   U24273 : XNOR2_X1 port map( A => n22184, B => n22183, ZN => n22185);
   U24274 : XNOR2_X1 port map( A => n22186, B => n22185, ZN => n23266);
   U24275 : XNOR2_X1 port map( A => n22188, B => n22187, ZN => n22191);
   U24276 : XNOR2_X1 port map( A => n22409, B => n3673, ZN => n22189);
   U24277 : XNOR2_X1 port map( A => n22842, B => n22189, ZN => n22190);
   U24278 : XNOR2_X1 port map( A => n22193, B => n22192, ZN => n22198);
   U24279 : XNOR2_X1 port map( A => n22664, B => n22194, ZN => n22837);
   U24280 : XNOR2_X1 port map( A => n22195, B => n3695, ZN => n22196);
   U24281 : XNOR2_X1 port map( A => n22837, B => n22196, ZN => n22197);
   U24282 : XNOR2_X1 port map( A => n22198, B => n22197, ZN => n23267);
   U24283 : XNOR2_X1 port map( A => n22828, B => n22395, ZN => n22203);
   U24284 : XNOR2_X1 port map( A => n22522, B => n355, ZN => n22201);
   U24285 : XNOR2_X1 port map( A => n22703, B => n3633, ZN => n22200);
   U24286 : XNOR2_X1 port map( A => n22201, B => n22200, ZN => n22202);
   U24287 : MUX2_X1 port map( A => n379, B => n23217, S => n406, Z => n22217);
   U24288 : XNOR2_X1 port map( A => n28514, B => n22206, ZN => n22210);
   U24289 : XNOR2_X1 port map( A => n22434, B => n2996, ZN => n22208);
   U24290 : XNOR2_X1 port map( A => n22208, B => n22207, ZN => n22209);
   U24291 : INV_X1 port map( A => n23562, ZN => n23615);
   U24292 : OAI22_X1 port map( A1 => n23615, A2 => n406, B1 => n23267, B2 => 
                           n23266, ZN => n22215);
   U24293 : XNOR2_X1 port map( A => n22488, B => n6319, ZN => n22211);
   U24294 : XNOR2_X1 port map( A => n22211, B => n22418, ZN => n22212);
   U24295 : XNOR2_X1 port map( A => n22619, B => n28409, ZN => n22348);
   U24296 : XNOR2_X1 port map( A => n22212, B => n22348, ZN => n22214);
   U24297 : XNOR2_X1 port map( A => n22213, B => n22214, ZN => n23611);
   U24298 : INV_X1 port map( A => n23611, ZN => n23216);
   U24299 : NAND2_X1 port map( A1 => n22215, A2 => n23216, ZN => n22216);
   U24301 : INV_X1 port map( A => n24735, ZN => n24280);
   U24302 : INV_X1 port map( A => n22218, ZN => n22624);
   U24304 : INV_X1 port map( A => n22220, ZN => n22546);
   U24305 : XNOR2_X1 port map( A => n22712, B => n22546, ZN => n22225);
   U24306 : XNOR2_X1 port map( A => n22221, B => n22790, ZN => n22223);
   U24307 : XNOR2_X1 port map( A => n22279, B => n27956, ZN => n22222);
   U24308 : XNOR2_X1 port map( A => n22223, B => n22222, ZN => n22224);
   U24309 : XNOR2_X1 port map( A => n22225, B => n22224, ZN => n23563);
   U24310 : XNOR2_X1 port map( A => n22226, B => n22227, ZN => n22772);
   U24311 : XNOR2_X1 port map( A => n22880, B => n22772, ZN => n22231);
   U24312 : XNOR2_X1 port map( A => n22295, B => n22697, ZN => n22229);
   U24313 : XNOR2_X1 port map( A => n22698, B => n3752, ZN => n22228);
   U24314 : XNOR2_X1 port map( A => n22229, B => n22228, ZN => n22230);
   U24315 : XNOR2_X1 port map( A => n22232, B => n22601, ZN => n22733);
   U24316 : INV_X1 port map( A => n22733, ZN => n22233);
   U24317 : XNOR2_X1 port map( A => n22533, B => n22233, ZN => n22237);
   U24318 : XNOR2_X1 port map( A => n22762, B => Key(66), ZN => n22234);
   U24319 : XNOR2_X1 port map( A => n22235, B => n22234, ZN => n22236);
   U24320 : INV_X1 port map( A => n22609, ZN => n22239);
   U24321 : XNOR2_X1 port map( A => n22240, B => n22239, ZN => n22242);
   U24322 : XNOR2_X1 port map( A => n22718, B => n2981, ZN => n22241);
   U24323 : XNOR2_X1 port map( A => n22242, B => n22241, ZN => n22243);
   U24324 : XNOR2_X1 port map( A => n22633, B => n22778, ZN => n22247);
   U24325 : XNOR2_X1 port map( A => n22247, B => n22897, ZN => n22504);
   U24327 : XNOR2_X1 port map( A => n22248, B => n22270, ZN => n22250);
   U24328 : XNOR2_X1 port map( A => n22249, B => n22250, ZN => n22254);
   U24329 : XNOR2_X1 port map( A => n22724, B => n2984, ZN => n22251);
   U24330 : XNOR2_X1 port map( A => n22251, B => n22252, ZN => n22253);
   U24332 : INV_X1 port map( A => n23640, ZN => n23314);
   U24333 : NAND2_X1 port map( A1 => n2138, A2 => n23640, ZN => n22255);
   U24335 : OAI211_X1 port map( C1 => n28963, C2 => n23564, A => n22258, B => 
                           n22257, ZN => n22311);
   U24336 : NOR2_X1 port map( A1 => n24280, A2 => n22311, ZN => n24737);
   U24337 : XNOR2_X1 port map( A => n22495, B => n22259, ZN => n22263);
   U24338 : XNOR2_X1 port map( A => n6504, B => n3067, ZN => n22260);
   U24339 : XNOR2_X1 port map( A => n22261, B => n22260, ZN => n22262);
   U24340 : XNOR2_X1 port map( A => n22263, B => n22262, ZN => n23309);
   U24341 : INV_X1 port map( A => n23309, ZN => n23632);
   U24342 : XNOR2_X1 port map( A => n22264, B => n22481, ZN => n22269);
   U24343 : XNOR2_X1 port map( A => n22501, B => n2402, ZN => n22267);
   U24344 : XNOR2_X1 port map( A => n22265, B => n22692, ZN => n22266);
   U24345 : XNOR2_X1 port map( A => n22267, B => n22266, ZN => n22268);
   U24346 : XNOR2_X1 port map( A => n22271, B => n22270, ZN => n22274);
   U24347 : INV_X1 port map( A => n22272, ZN => n22273);
   U24348 : XNOR2_X1 port map( A => n22273, B => n22274, ZN => n22276);
   U24349 : XNOR2_X1 port map( A => n22506, B => n22890, ZN => n22485);
   U24350 : XNOR2_X1 port map( A => n28492, B => n3751, ZN => n22275);
   U24352 : XNOR2_X1 port map( A => n22786, B => n22278, ZN => n22281);
   U24353 : XNOR2_X1 port map( A => n22279, B => n22791, ZN => n22280);
   U24354 : XNOR2_X1 port map( A => n22281, B => n22280, ZN => n22282);
   U24355 : XNOR2_X1 port map( A => n22283, B => n22282, ZN => n23630);
   U24356 : XNOR2_X1 port map( A => n22285, B => n22525, ZN => n22771);
   U24357 : AOI21_X1 port map( B1 => n22286, B2 => n28790, A => n22290, ZN => 
                           n22287);
   U24358 : OAI21_X1 port map( B1 => n28790, B2 => n22288, A => n22287, ZN => 
                           n22293);
   U24359 : NAND3_X1 port map( A1 => n22291, A2 => n489, A3 => n22290, ZN => 
                           n22292);
   U24360 : NAND3_X1 port map( A1 => n22294, A2 => n22293, A3 => n22292, ZN => 
                           n22699);
   U24361 : XNOR2_X1 port map( A => n22699, B => n22295, ZN => n22297);
   U24362 : XNOR2_X1 port map( A => n22671, B => n2527, ZN => n22296);
   U24363 : XNOR2_X1 port map( A => n22033, B => n22394, ZN => n22299);
   U24364 : MUX2_X1 port map( A => n23630, B => n23558, S => n23557, Z => 
                           n22310);
   U24365 : XNOR2_X1 port map( A => n22300, B => n22734, ZN => n22304);
   U24366 : XNOR2_X1 port map( A => n22301, B => n22302, ZN => n22303);
   U24367 : XNOR2_X1 port map( A => n22304, B => n22303, ZN => n22309);
   U24368 : XNOR2_X1 port map( A => n22913, B => n22414, ZN => n22307);
   U24369 : INV_X1 port map( A => n22756, ZN => n22305);
   U24370 : XNOR2_X1 port map( A => n22305, B => n1196, ZN => n22306);
   U24371 : XNOR2_X1 port map( A => n22307, B => n22306, ZN => n22308);
   U24372 : XNOR2_X1 port map( A => n22309, B => n22308, ZN => n23631);
   U24373 : INV_X1 port map( A => n23631, ZN => n23629);
   U24374 : INV_X1 port map( A => n22311, ZN => n24736);
   U24375 : XNOR2_X1 port map( A => n22312, B => n22523, ZN => n22314);
   U24376 : XNOR2_X1 port map( A => n22314, B => n22313, ZN => n22317);
   U24377 : INV_X1 port map( A => n22315, ZN => n22316);
   U24378 : XNOR2_X1 port map( A => n22574, B => n22625, ZN => n22319);
   U24379 : XNOR2_X1 port map( A => n22319, B => n22318, ZN => n22324);
   U24380 : XNOR2_X1 port map( A => n22380, B => n3483, ZN => n22322);
   U24381 : XNOR2_X1 port map( A => n22379, B => n28499, ZN => n22321);
   U24382 : XNOR2_X1 port map( A => n22321, B => n22322, ZN => n22323);
   U24383 : XNOR2_X1 port map( A => n22326, B => n22910, ZN => n22357);
   U24384 : XNOR2_X1 port map( A => n22357, B => n22325, ZN => n22329);
   U24386 : OAI21_X1 port map( B1 => n23761, B2 => n23762, A => n23474, ZN => 
                           n22346);
   U24387 : XNOR2_X1 port map( A => n22330, B => n22644, ZN => n22332);
   U24388 : XNOR2_X1 port map( A => n22813, B => n3232, ZN => n22331);
   U24389 : XNOR2_X1 port map( A => n22332, B => n22331, ZN => n22336);
   U24390 : XNOR2_X1 port map( A => n22333, B => n22434, ZN => n22635);
   U24391 : XNOR2_X1 port map( A => n22635, B => n22362, ZN => n22335);
   U24393 : XNOR2_X1 port map( A => n22338, B => n22337, ZN => n22369);
   U24394 : XNOR2_X1 port map( A => n22610, B => n27462, ZN => n22339);
   U24395 : XNOR2_X1 port map( A => n22339, B => n22369, ZN => n22345);
   U24396 : XNOR2_X1 port map( A => n22605, B => n22340, ZN => n22343);
   U24397 : INV_X1 port map( A => n22341, ZN => n22342);
   U24398 : XNOR2_X1 port map( A => n22342, B => n22343, ZN => n22344);
   U24400 : NAND2_X1 port map( A1 => n22346, A2 => n23475, ZN => n22355);
   U24401 : NAND2_X1 port map( A1 => n23762, A2 => n23760, ZN => n22354);
   U24402 : XNOR2_X1 port map( A => n22374, B => n22888, ZN => n22347);
   U24403 : XNOR2_X1 port map( A => n22348, B => n22347, ZN => n22352);
   U24404 : XNOR2_X1 port map( A => n28483, B => n3625, ZN => n22349);
   U24405 : XNOR2_X1 port map( A => n22350, B => n22349, ZN => n22351);
   U24406 : XNOR2_X1 port map( A => n22351, B => n22352, ZN => n23326);
   U24407 : INV_X1 port map( A => n23762, ZN => n23034);
   U24409 : AOI22_X1 port map( A1 => n22356, A2 => n24735, B1 => n24736, B2 => 
                           n24602, ZN => n22450);
   U24410 : XNOR2_X1 port map( A => n22735, B => n26531, ZN => n22359);
   U24411 : XNOR2_X1 port map( A => n22358, B => n22359, ZN => n22360);
   U24412 : XNOR2_X1 port map( A => n22689, B => n22362, ZN => n22367);
   U24413 : XNOR2_X1 port map( A => n22363, B => n22812, ZN => n22365);
   U24414 : XNOR2_X1 port map( A => n21728, B => n1119, ZN => n22364);
   U24415 : XNOR2_X1 port map( A => n22365, B => n22364, ZN => n22366);
   U24416 : XNOR2_X1 port map( A => n22369, B => n22368, ZN => n22373);
   U24417 : XNOR2_X1 port map( A => n22370, B => n22553, ZN => n22371);
   U24418 : XNOR2_X1 port map( A => n22607, B => n22371, ZN => n22372);
   U24419 : XNOR2_X1 port map( A => n22372, B => n22373, ZN => n23620);
   U24420 : NAND2_X1 port map( A1 => n23621, A2 => n23620, ZN => n23273);
   U24421 : XNOR2_X1 port map( A => n22374, B => n3660, ZN => n22375);
   U24422 : XNOR2_X1 port map( A => n22617, B => n22375, ZN => n22378);
   U24423 : XNOR2_X1 port map( A => n22796, B => n22888, ZN => n22376);
   U24424 : XNOR2_X1 port map( A => n22727, B => n22376, ZN => n22377);
   U24425 : XNOR2_X1 port map( A => n22377, B => n22378, ZN => n23619);
   U24426 : INV_X1 port map( A => n23619, ZN => n22987);
   U24427 : OAI21_X1 port map( B1 => n23620, B2 => n22987, A => n23273, ZN => 
                           n22392);
   U24428 : XNOR2_X1 port map( A => n22379, B => n22380, ZN => n22381);
   U24429 : XNOR2_X1 port map( A => n22626, B => n22381, ZN => n22385);
   U24430 : XNOR2_X1 port map( A => n22383, B => n22382, ZN => n22384);
   U24432 : NAND2_X1 port map( A1 => n23622, A2 => n23566, ZN => n22391);
   U24433 : XNOR2_X1 port map( A => n22386, B => n22584, ZN => n22389);
   U24434 : XNOR2_X1 port map( A => n22387, B => n3722, ZN => n22388);
   U24435 : INV_X1 port map( A => n23618, ZN => n23567);
   U24436 : OAI21_X1 port map( B1 => n23622, B2 => n23273, A => n22393, ZN => 
                           n24739);
   U24437 : INV_X1 port map( A => n24739, ZN => n24282);
   U24438 : AND2_X1 port map( A1 => n3310, A2 => n22311, ZN => n24603);
   U24439 : INV_X1 port map( A => n22396, ZN => n22400);
   U24440 : NAND2_X1 port map( A1 => n22402, A2 => n22397, ZN => n22399);
   U24441 : AOI21_X1 port map( B1 => n22400, B2 => n22399, A => n22398, ZN => 
                           n22406);
   U24442 : OAI21_X1 port map( B1 => n6940, B2 => n22404, A => n22403, ZN => 
                           n22405);
   U24443 : NOR2_X1 port map( A1 => n22406, A2 => n22405, ZN => n22407);
   U24444 : INV_X1 port map( A => n22581, ZN => n22408);
   U24445 : INV_X1 port map( A => n23049, ZN => n23472);
   U24446 : XNOR2_X1 port map( A => n22759, B => n22409, ZN => n22413);
   U24447 : XNOR2_X1 port map( A => n22414, B => n22473, ZN => n22415);
   U24448 : XNOR2_X1 port map( A => n28162, B => n22415, ZN => n22416);
   U24449 : XNOR2_X1 port map( A => n22418, B => n2577, ZN => n22421);
   U24450 : XNOR2_X1 port map( A => n22567, B => n22419, ZN => n22420);
   U24451 : XNOR2_X1 port map( A => n22421, B => n22420, ZN => n22425);
   U24452 : XNOR2_X1 port map( A => n22422, B => n22619, ZN => n22423);
   U24453 : XNOR2_X1 port map( A => n22423, B => n22571, ZN => n22424);
   U24454 : XNOR2_X1 port map( A => n22610, B => n29562, ZN => n22430);
   U24455 : XNOR2_X1 port map( A => n29490, B => n22427, ZN => n22429);
   U24456 : INV_X1 port map( A => n3378, ZN => n26545);
   U24457 : XNOR2_X1 port map( A => n22556, B => n26545, ZN => n22431);
   U24458 : XNOR2_X1 port map( A => n22558, B => n22431, ZN => n22432);
   U24459 : OAI21_X1 port map( B1 => n23318, B2 => n23472, A => n22433, ZN => 
                           n23473);
   U24460 : INV_X1 port map( A => n23473, ZN => n22448);
   U24461 : XNOR2_X1 port map( A => n22561, B => n22434, ZN => n22435);
   U24462 : XNOR2_X1 port map( A => n22436, B => n22435, ZN => n22440);
   U24463 : XNOR2_X1 port map( A => n22690, B => n22437, ZN => n22780);
   U24464 : XNOR2_X1 port map( A => n22479, B => n1046, ZN => n22438);
   U24465 : XNOR2_X1 port map( A => n22780, B => n22438, ZN => n22439);
   U24466 : XNOR2_X1 port map( A => n22784, B => n3422, ZN => n22441);
   U24467 : XNOR2_X1 port map( A => n22443, B => n22442, ZN => n22446);
   U24468 : XNOR2_X1 port map( A => n22464, B => n22787, ZN => n22444);
   U24469 : XNOR2_X1 port map( A => n22444, B => n22625, ZN => n22445);
   U24470 : XNOR2_X1 port map( A => n22446, B => n22445, ZN => n23648);
   U24471 : AOI22_X1 port map( A1 => n24744, A2 => n24604, B1 => n24603, B2 => 
                           n24734, ZN => n22449);
   U24472 : OAI21_X1 port map( B1 => n24737, B2 => n22450, A => n22449, ZN => 
                           n25428);
   U24473 : XNOR2_X1 port map( A => n26044, B => n25428, ZN => n25803);
   U24474 : XNOR2_X1 port map( A => n24885, B => n25803, ZN => n22943);
   U24476 : OAI21_X1 port map( B1 => n29618, B2 => n23700, A => n23705, ZN => 
                           n22453);
   U24477 : NOR2_X1 port map( A1 => n22953, A2 => n22455, ZN => n23396);
   U24478 : NOR2_X1 port map( A1 => n23396, A2 => n23726, ZN => n22458);
   U24479 : NOR2_X1 port map( A1 => n28484, A2 => n23843, ZN => n22456);
   U24480 : AOI22_X1 port map( A1 => n23396, A2 => n23845, B1 => n22456, B2 => 
                           n22455, ZN => n22457);
   U24482 : XNOR2_X1 port map( A => n22791, B => n3607, ZN => n22460);
   U24483 : XNOR2_X1 port map( A => n22460, B => n22459, ZN => n22462);
   U24484 : XNOR2_X1 port map( A => n22462, B => n22461, ZN => n22466);
   U24485 : XNOR2_X1 port map( A => n22464, B => n28450, ZN => n22666);
   U24486 : XNOR2_X1 port map( A => n22923, B => n22666, ZN => n22465);
   U24487 : XNOR2_X1 port map( A => n22703, B => n2889, ZN => n22467);
   U24488 : XNOR2_X1 port map( A => n22671, B => n29514, ZN => n22469);
   U24489 : XNOR2_X1 port map( A => n22472, B => n22473, ZN => n22652);
   U24490 : XNOR2_X1 port map( A => n22652, B => n22474, ZN => n22478);
   U24491 : XNOR2_X1 port map( A => n22913, B => n22735, ZN => n22476);
   U24492 : XNOR2_X1 port map( A => n28486, B => n26665, ZN => n22475);
   U24493 : XNOR2_X1 port map( A => n22476, B => n22475, ZN => n22477);
   U24494 : INV_X1 port map( A => n22494, ZN => n23837);
   U24496 : XNOR2_X1 port map( A => n22479, B => n3114, ZN => n22480);
   U24497 : XNOR2_X1 port map( A => n22480, B => n21789, ZN => n22482);
   U24498 : XNOR2_X1 port map( A => n22481, B => n22482, ZN => n22484);
   U24499 : XNOR2_X1 port map( A => n22485, B => n22486, ZN => n22493);
   U24500 : XNOR2_X1 port map( A => n22487, B => n22488, ZN => n22491);
   U24501 : XNOR2_X1 port map( A => n22657, B => n22489, ZN => n22490);
   U24502 : XNOR2_X1 port map( A => n22491, B => n22490, ZN => n22492);
   U24503 : XNOR2_X1 port map( A => n22493, B => n22492, ZN => n23078);
   U24504 : INV_X1 port map( A => n23078, ZN => n23390);
   U24505 : XNOR2_X1 port map( A => n22514, B => n22713, ZN => n22496);
   U24506 : XNOR2_X1 port map( A => n22556, B => n3191, ZN => n22498);
   U24507 : NAND3_X1 port map( A1 => n28460, A2 => n23839, A3 => n28418, ZN => 
                           n22499);
   U24508 : MUX2_X1 port map( A => n24614, B => n24610, S => n29109, Z => 
                           n22640);
   U24509 : XNOR2_X1 port map( A => n22503, B => n22502, ZN => n22505);
   U24510 : XNOR2_X1 port map( A => n22891, B => n22724, ZN => n22508);
   U24511 : XNOR2_X1 port map( A => n22506, B => n3654, ZN => n22507);
   U24512 : XNOR2_X1 port map( A => n22508, B => n22507, ZN => n22513);
   U24513 : XNOR2_X1 port map( A => n1858, B => n22509, ZN => n22510);
   U24514 : XNOR2_X1 port map( A => n22514, B => n22609, ZN => n22517);
   U24515 : XNOR2_X1 port map( A => n22515, B => n5059, ZN => n22516);
   U24516 : XNOR2_X1 port map( A => n22517, B => n22516, ZN => n22521);
   U24517 : XNOR2_X1 port map( A => n22519, B => n22518, ZN => n22520);
   U24518 : XNOR2_X1 port map( A => n22520, B => n22521, ZN => n23295);
   U24519 : MUX2_X1 port map( A => n22531, B => n23077, S => n23295, Z => 
                           n22552);
   U24520 : XNOR2_X1 port map( A => n22523, B => n22522, ZN => n22884);
   U24521 : XNOR2_X1 port map( A => n22884, B => n22524, ZN => n22530);
   U24522 : XNOR2_X1 port map( A => n22526, B => n22525, ZN => n22528);
   U24523 : XNOR2_X1 port map( A => n22698, B => n3493, ZN => n22527);
   U24524 : XNOR2_X1 port map( A => n22528, B => n22527, ZN => n22529);
   U24525 : INV_X1 port map( A => n23297, ZN => n22962);
   U24526 : INV_X1 port map( A => n23295, ZN => n23832);
   U24527 : XNOR2_X1 port map( A => n22532, B => n22533, ZN => n22540);
   U24528 : XNOR2_X1 port map( A => n28486, B => n22534, ZN => n22538);
   U24529 : INV_X1 port map( A => n22601, ZN => n22536);
   U24530 : XNOR2_X1 port map( A => n22536, B => n22535, ZN => n22537);
   U24531 : XNOR2_X1 port map( A => n22537, B => n22538, ZN => n22539);
   U24532 : NAND2_X1 port map( A1 => n23832, A2 => n29602, ZN => n22541);
   U24533 : NOR2_X1 port map( A1 => n23833, A2 => n22541, ZN => n22550);
   U24534 : NOR2_X1 port map( A1 => n29020, A2 => n29602, ZN => n22549);
   U24535 : XNOR2_X1 port map( A => n22624, B => n22542, ZN => n22544);
   U24536 : XNOR2_X1 port map( A => n22791, B => n3528, ZN => n22543);
   U24537 : XNOR2_X1 port map( A => n22544, B => n22543, ZN => n22548);
   U24538 : XNOR2_X1 port map( A => n22546, B => n22545, ZN => n22547);
   U24539 : XNOR2_X1 port map( A => n22547, B => n22548, ZN => n22864);
   U24540 : INV_X1 port map( A => n23831, ZN => n23296);
   U24541 : OAI21_X1 port map( B1 => n22550, B2 => n22549, A => n23298, ZN => 
                           n22551);
   U24542 : OAI21_X1 port map( B1 => n22552, B2 => n22962, A => n22551, ZN => 
                           n24017);
   U24543 : XNOR2_X1 port map( A => n22180, B => n22553, ZN => n22554);
   U24544 : XNOR2_X1 port map( A => n22555, B => n22554, ZN => n22560);
   U24545 : XNOR2_X1 port map( A => n22556, B => n1184, ZN => n22557);
   U24546 : XNOR2_X1 port map( A => n22558, B => n22557, ZN => n22559);
   U24548 : XNOR2_X1 port map( A => n22813, B => n2325, ZN => n22562);
   U24550 : XNOR2_X1 port map( A => n22567, B => n22568, ZN => n22655);
   U24551 : XNOR2_X1 port map( A => n22569, B => n22655, ZN => n22573);
   U24552 : XNOR2_X1 port map( A => n28409, B => n3003, ZN => n22570);
   U24553 : XNOR2_X1 port map( A => n22571, B => n22570, ZN => n22572);
   U24554 : XNOR2_X1 port map( A => n22575, B => n22838, ZN => n22580);
   U24555 : INV_X1 port map( A => n22790, ZN => n22576);
   U24556 : XNOR2_X1 port map( A => n22576, B => n3180, ZN => n22577);
   U24557 : XNOR2_X1 port map( A => n22578, B => n22577, ZN => n22579);
   U24558 : XNOR2_X2 port map( A => n22579, B => n22580, ZN => n23382);
   U24559 : XNOR2_X1 port map( A => n22582, B => n22581, ZN => n22586);
   U24560 : INV_X1 port map( A => n22829, ZN => n22881);
   U24561 : XNOR2_X1 port map( A => n22881, B => n3457, ZN => n22583);
   U24562 : XNOR2_X1 port map( A => n22584, B => n22583, ZN => n22585);
   U24563 : XNOR2_X1 port map( A => n22586, B => n22585, ZN => n22946);
   U24564 : XNOR2_X1 port map( A => n22589, B => n28589, ZN => n22591);
   U24565 : XNOR2_X1 port map( A => n22410, B => n2541, ZN => n22590);
   U24566 : MUX2_X1 port map( A => n24017, B => n29109, S => n24612, Z => 
                           n22639);
   U24567 : XNOR2_X1 port map( A => n22596, B => n22595, ZN => n22597);
   U24568 : XNOR2_X1 port map( A => n22598, B => n22597, ZN => n22742);
   U24569 : INV_X1 port map( A => n22599, ZN => n22909);
   U24570 : XNOR2_X1 port map( A => n22909, B => n22600, ZN => n22604);
   U24571 : XNOR2_X1 port map( A => n22601, B => n3015, ZN => n22602);
   U24572 : XNOR2_X1 port map( A => n22325, B => n22602, ZN => n22603);
   U24574 : XNOR2_X1 port map( A => n22605, B => n22606, ZN => n22608);
   U24575 : XNOR2_X1 port map( A => n22607, B => n22608, ZN => n22614);
   U24576 : XNOR2_X1 port map( A => n22610, B => n2982, ZN => n22611);
   U24577 : XNOR2_X1 port map( A => n22611, B => n22612, ZN => n22613);
   U24578 : XNOR2_X1 port map( A => n22613, B => n22614, ZN => n23810);
   U24579 : XNOR2_X1 port map( A => n22615, B => n3644, ZN => n22616);
   U24580 : XNOR2_X1 port map( A => n22617, B => n22616, ZN => n22623);
   U24581 : XNOR2_X1 port map( A => n22618, B => n22619, ZN => n22621);
   U24582 : XNOR2_X1 port map( A => n22620, B => n22621, ZN => n22622);
   U24583 : XNOR2_X1 port map( A => n22624, B => n22625, ZN => n22627);
   U24584 : XNOR2_X1 port map( A => n22626, B => n22627, ZN => n22631);
   U24585 : XNOR2_X1 port map( A => n22628, B => n27452, ZN => n22629);
   U24586 : XNOR2_X1 port map( A => n22922, B => n22629, ZN => n22630);
   U24587 : XNOR2_X1 port map( A => n22630, B => n22631, ZN => n23285);
   U24588 : XNOR2_X1 port map( A => n22635, B => n22634, ZN => n22636);
   U24589 : XNOR2_X1 port map( A => n22637, B => n22636, ZN => n22877);
   U24590 : INV_X1 port map( A => n22877, ZN => n23074);
   U24591 : MUX2_X1 port map( A => n22640, B => n22639, S => n5137, Z => n25727
                           );
   U24592 : XNOR2_X1 port map( A => n22641, B => n22642, ZN => n22648);
   U24593 : XNOR2_X1 port map( A => n22811, B => n22643, ZN => n22646);
   U24594 : XNOR2_X1 port map( A => n22644, B => n1887, ZN => n22645);
   U24595 : XNOR2_X1 port map( A => n22646, B => n22645, ZN => n22647);
   U24596 : XNOR2_X1 port map( A => n22844, B => n857, ZN => n22649);
   U24597 : XNOR2_X1 port map( A => n22650, B => n22649, ZN => n22654);
   U24598 : XNOR2_X1 port map( A => n22651, B => n22652, ZN => n22653);
   U24599 : XNOR2_X1 port map( A => n22656, B => n22820, ZN => n22659);
   U24600 : XNOR2_X1 port map( A => n28492, B => n3697, ZN => n22658);
   U24601 : XNOR2_X1 port map( A => n22659, B => n22658, ZN => n22660);
   U24602 : MUX2_X1 port map( A => n1829, B => n22686, S => n408, Z => n22676);
   U24603 : XNOR2_X1 port map( A => n22661, B => n29079, ZN => n22662);
   U24604 : XNOR2_X1 port map( A => n22663, B => n22662, ZN => n22667);
   U24605 : XNOR2_X1 port map( A => n22664, B => n27225, ZN => n22665);
   U24606 : XNOR2_X1 port map( A => n22668, B => n3537, ZN => n22669);
   U24607 : XNOR2_X1 port map( A => n22670, B => n22669, ZN => n22673);
   U24608 : XNOR2_X1 port map( A => n22768, B => n22671, ZN => n22672);
   U24609 : XNOR2_X1 port map( A => n22673, B => n22672, ZN => n22674);
   U24610 : XNOR2_X1 port map( A => n22674, B => n22675, ZN => n23302);
   U24611 : INV_X1 port map( A => n22678, ZN => n22679);
   U24612 : XNOR2_X1 port map( A => n22679, B => n22680, ZN => n22683);
   U24613 : XNOR2_X1 port map( A => n22681, B => n22856, ZN => n22682);
   U24614 : XNOR2_X1 port map( A => n22683, B => n22682, ZN => n22685);
   U24615 : XNOR2_X1 port map( A => n22685, B => n22684, ZN => n23433);
   U24616 : XNOR2_X1 port map( A => n22688, B => n22689, ZN => n22696);
   U24617 : XNOR2_X1 port map( A => n22691, B => n22690, ZN => n22694);
   U24618 : XNOR2_X1 port map( A => n22692, B => n1161, ZN => n22693);
   U24619 : XNOR2_X1 port map( A => n22694, B => n22693, ZN => n22695);
   U24621 : INV_X1 port map( A => n23450, ZN => n23447);
   U24622 : XNOR2_X1 port map( A => n22697, B => n22033, ZN => n22702);
   U24625 : XNOR2_X1 port map( A => n22701, B => n22702, ZN => n22709);
   U24626 : XNOR2_X1 port map( A => n22703, B => n22387, ZN => n22707);
   U24627 : XNOR2_X1 port map( A => n22707, B => n22706, ZN => n22708);
   U24628 : XNOR2_X1 port map( A => n22784, B => n3223, ZN => n22711);
   U24629 : XNOR2_X1 port map( A => n22713, B => n22903, ZN => n22715);
   U24630 : XNOR2_X1 port map( A => n22715, B => n22714, ZN => n22722);
   U24631 : XNOR2_X1 port map( A => n22717, B => n29591, ZN => n22720);
   U24632 : XNOR2_X1 port map( A => n22718, B => n3414, ZN => n22719);
   U24633 : XNOR2_X1 port map( A => n22720, B => n22719, ZN => n22721);
   U24634 : XNOR2_X1 port map( A => n22722, B => n22721, ZN => n22935);
   U24635 : INV_X1 port map( A => n22935, ZN => n23109);
   U24636 : AOI22_X1 port map( A1 => n23447, A2 => n23442, B1 => n23370, B2 => 
                           n23109, ZN => n22741);
   U24637 : XNOR2_X1 port map( A => n22723, B => n28693, ZN => n22726);
   U24638 : XNOR2_X1 port map( A => n22724, B => n22890, ZN => n22725);
   U24639 : XNOR2_X1 port map( A => n22725, B => n22726, ZN => n22730);
   U24640 : XNOR2_X2 port map( A => n22729, B => n22730, ZN => n23445);
   U24641 : XNOR2_X1 port map( A => n22731, B => n28162, ZN => n22732);
   U24642 : XNOR2_X1 port map( A => n22732, B => n22733, ZN => n22739);
   U24643 : XNOR2_X1 port map( A => n22735, B => n22734, ZN => n22737);
   U24644 : XNOR2_X1 port map( A => n22913, B => n3196, ZN => n22736);
   U24645 : XNOR2_X1 port map( A => n22736, B => n22737, ZN => n22738);
   U24646 : INV_X1 port map( A => n24552, ZN => n23205);
   U24647 : INV_X1 port map( A => n23809, ZN => n23075);
   U24648 : INV_X1 port map( A => n24551, ZN => n22746);
   U24649 : NOR2_X1 port map( A1 => n22747, A2 => n22746, ZN => n22872);
   U24650 : XNOR2_X1 port map( A => n22748, B => n22749, ZN => n22754);
   U24651 : XNOR2_X1 port map( A => n22750, B => n2385, ZN => n22751);
   U24652 : XNOR2_X1 port map( A => n22752, B => n22751, ZN => n22753);
   U24653 : XNOR2_X1 port map( A => n22754, B => n22753, ZN => n23099);
   U24654 : XNOR2_X1 port map( A => n22756, B => n22755, ZN => n22758);
   U24655 : XNOR2_X1 port map( A => n22759, B => n22760, ZN => n22761);
   U24656 : XNOR2_X1 port map( A => n22763, B => n28589, ZN => n22764);
   U24657 : XNOR2_X1 port map( A => n28162, B => n22764, ZN => n22766);
   U24658 : XNOR2_X2 port map( A => n22767, B => n22766, ZN => n23419);
   U24659 : XNOR2_X1 port map( A => n22769, B => n22768, ZN => n22770);
   U24660 : XNOR2_X1 port map( A => n22770, B => n22771, ZN => n22775);
   U24661 : XNOR2_X1 port map( A => n22773, B => n22772, ZN => n22774);
   U24662 : XNOR2_X1 port map( A => n22777, B => n22776, ZN => n22782);
   U24663 : XNOR2_X1 port map( A => n22778, B => n3244, ZN => n22779);
   U24664 : XNOR2_X1 port map( A => n22780, B => n22779, ZN => n22781);
   U24665 : XNOR2_X1 port map( A => n22782, B => n22781, ZN => n23073);
   U24666 : INV_X1 port map( A => n23073, ZN => n23417);
   U24667 : XNOR2_X1 port map( A => n22785, B => n22784, ZN => n22789);
   U24668 : XNOR2_X1 port map( A => n22787, B => n22786, ZN => n22788);
   U24669 : XNOR2_X1 port map( A => n22789, B => n22788, ZN => n22795);
   U24670 : XNOR2_X1 port map( A => n22791, B => n22790, ZN => n22793);
   U24671 : XNOR2_X1 port map( A => n22792, B => n22793, ZN => n22794);
   U24672 : INV_X1 port map( A => n22796, ZN => n22797);
   U24673 : XNOR2_X1 port map( A => n22797, B => n22798, ZN => n22799);
   U24674 : XNOR2_X1 port map( A => n22799, B => n22800, ZN => n22804);
   U24675 : XNOR2_X1 port map( A => n1859, B => n3164, ZN => n22802);
   U24676 : XNOR2_X1 port map( A => n22801, B => n22802, ZN => n22803);
   U24677 : NAND2_X1 port map( A1 => n480, A2 => n23418, ZN => n22805);
   U24678 : MUX2_X1 port map( A => n22806, B => n22805, S => n23415, Z => 
                           n22807);
   U24680 : NOR2_X1 port map( A1 => n24556, A2 => n24552, ZN => n23207);
   U24681 : INV_X1 port map( A => n23207, ZN => n22870);
   U24682 : XNOR2_X1 port map( A => n22810, B => n22809, ZN => n22817);
   U24683 : XNOR2_X1 port map( A => n22811, B => n22812, ZN => n22815);
   U24684 : XNOR2_X1 port map( A => n22813, B => n2446, ZN => n22814);
   U24685 : XNOR2_X1 port map( A => n22815, B => n22814, ZN => n22816);
   U24686 : XNOR2_X1 port map( A => n22819, B => n22818, ZN => n22826);
   U24687 : XNOR2_X1 port map( A => n22820, B => n22821, ZN => n22824);
   U24688 : XNOR2_X1 port map( A => n22822, B => n2973, ZN => n22823);
   U24689 : XNOR2_X1 port map( A => n22824, B => n22823, ZN => n22825);
   U24690 : XNOR2_X1 port map( A => n22826, B => n22825, ZN => n22931);
   U24691 : NOR2_X1 port map( A1 => n23820, A2 => n22931, ZN => n22851);
   U24692 : XNOR2_X1 port map( A => n22828, B => n22827, ZN => n22834);
   U24693 : XNOR2_X1 port map( A => n355, B => n22882, ZN => n22832);
   U24694 : XNOR2_X1 port map( A => n22830, B => n26909, ZN => n22831);
   U24695 : XNOR2_X1 port map( A => n22832, B => n22831, ZN => n22833);
   U24696 : XNOR2_X1 port map( A => n22835, B => n2946, ZN => n22836);
   U24697 : XNOR2_X1 port map( A => n22837, B => n22836, ZN => n22841);
   U24699 : XNOR2_X1 port map( A => n22842, B => n22843, ZN => n22850);
   U24700 : XNOR2_X1 port map( A => n22844, B => n22845, ZN => n22848);
   U24701 : XNOR2_X1 port map( A => n22410, B => n3256, ZN => n22847);
   U24702 : XNOR2_X1 port map( A => n22848, B => n22847, ZN => n22849);
   U24703 : XNOR2_X1 port map( A => n22852, B => n22902, ZN => n22860);
   U24704 : INV_X1 port map( A => n2509, ZN => n22853);
   U24705 : XNOR2_X1 port map( A => n22854, B => n22853, ZN => n22858);
   U24706 : XNOR2_X1 port map( A => n22856, B => n22855, ZN => n22857);
   U24707 : XNOR2_X1 port map( A => n22858, B => n22857, ZN => n22859);
   U24708 : XNOR2_X1 port map( A => n22860, B => n22859, ZN => n23291);
   U24709 : MUX2_X1 port map( A => n23290, B => n23291, S => n28182, Z => 
                           n22861);
   U24710 : INV_X1 port map( A => n22864, ZN => n23835);
   U24711 : NAND2_X1 port map( A1 => n23835, A2 => n29602, ZN => n22865);
   U24712 : AOI21_X1 port map( B1 => n22865, B2 => n23295, A => n23833, ZN => 
                           n22866);
   U24714 : INV_X1 port map( A => n24555, ZN => n24178);
   U24715 : OAI22_X1 port map( A1 => n22870, A2 => n22869, B1 => n22868, B2 => 
                           n24178, ZN => n22871);
   U24716 : XNOR2_X1 port map( A => n28576, B => n25727, ZN => n22941);
   U24717 : NOR2_X1 port map( A1 => n1829, A2 => n23433, ZN => n22874);
   U24718 : NOR2_X1 port map( A1 => n23302, A2 => n4020, ZN => n22873);
   U24719 : MUX2_X1 port map( A => n22874, B => n22873, S => n23431, Z => 
                           n22876);
   U24720 : INV_X1 port map( A => n23430, ZN => n23301);
   U24721 : INV_X1 port map( A => n24592, ZN => n23929);
   U24722 : XNOR2_X1 port map( A => n22879, B => n22880, ZN => n22885);
   U24723 : XNOR2_X1 port map( A => n22881, B => n3482, ZN => n22883);
   U24724 : INV_X1 port map( A => n23145, ZN => n23465);
   U24725 : INV_X1 port map( A => n22886, ZN => n22895);
   U24726 : XNOR2_X1 port map( A => n22887, B => n27231, ZN => n22889);
   U24727 : XNOR2_X1 port map( A => n22889, B => n22888, ZN => n22893);
   U24728 : XNOR2_X1 port map( A => n22891, B => n22890, ZN => n22892);
   U24729 : XNOR2_X1 port map( A => n22893, B => n22892, ZN => n22894);
   U24730 : XNOR2_X1 port map( A => n22895, B => n22894, ZN => n23148);
   U24731 : XNOR2_X1 port map( A => n22898, B => n1923, ZN => n22900);
   U24732 : XNOR2_X1 port map( A => n22900, B => n22899, ZN => n22901);
   U24733 : XNOR2_X1 port map( A => n22903, B => n2523, ZN => n22904);
   U24734 : XNOR2_X1 port map( A => n22905, B => n22904, ZN => n22906);
   U24735 : XNOR2_X1 port map( A => n22907, B => n22906, ZN => n23454);
   U24736 : AOI21_X1 port map( B1 => n23455, B2 => n23456, A => n23454, ZN => 
                           n22926);
   U24737 : XNOR2_X1 port map( A => n22909, B => n22908, ZN => n22917);
   U24738 : INV_X1 port map( A => n28472, ZN => n22911);
   U24739 : XNOR2_X1 port map( A => n22912, B => n22911, ZN => n22915);
   U24740 : XNOR2_X1 port map( A => n22913, B => n2411, ZN => n22914);
   U24741 : XNOR2_X1 port map( A => n22915, B => n22914, ZN => n22916);
   U24742 : NOR2_X1 port map( A1 => n23454, A2 => n23148, ZN => n22925);
   U24743 : XNOR2_X1 port map( A => n22919, B => n22918, ZN => n22921);
   U24744 : XNOR2_X1 port map( A => n22921, B => n22920, ZN => n22924);
   U24745 : NOR2_X1 port map( A1 => n23099, A2 => n23073, ZN => n22927);
   U24746 : MUX2_X1 port map( A => n22928, B => n22927, S => n23419, Z => 
                           n22930);
   U24749 : INV_X1 port map( A => n24593, ZN => n23853);
   U24750 : NOR2_X1 port map( A1 => n23289, A2 => n28182, ZN => n22934);
   U24753 : NOR2_X1 port map( A1 => n23290, A2 => n28609, ZN => n23818);
   U24754 : AND3_X1 port map( A1 => n22931, A2 => n28609, A3 => n23291, ZN => 
                           n22932);
   U24755 : NOR2_X1 port map( A1 => n23818, A2 => n22932, ZN => n22933);
   U24756 : OAI21_X1 port map( B1 => n22934, B2 => n23090, A => n22933, ZN => 
                           n24141);
   U24757 : INV_X1 port map( A => n23442, ZN => n23446);
   U24758 : MUX2_X1 port map( A => n292, B => n23446, S => n29296, Z => n22939)
                           ;
   U24759 : NAND2_X1 port map( A1 => n23370, A2 => n292, ZN => n22937);
   U24760 : NAND2_X1 port map( A1 => n23445, A2 => n23449, ZN => n22936);
   U24761 : MUX2_X1 port map( A => n22937, B => n22936, S => n23442, Z => 
                           n22938);
   U24762 : XNOR2_X1 port map( A => n25369, B => n3527, ZN => n22940);
   U24763 : XNOR2_X1 port map( A => n22941, B => n22940, ZN => n22942);
   U24765 : NOR2_X1 port map( A1 => n885, A2 => n23382, ZN => n22945);
   U24766 : NOR2_X1 port map( A1 => n24542, A2 => n2823, ZN => n22952);
   U24767 : INV_X1 port map( A => n23733, ZN => n23257);
   U24768 : AOI21_X1 port map( B1 => n23399, B2 => n23228, A => n23257, ZN => 
                           n22951);
   U24769 : NOR2_X1 port map( A1 => n22949, A2 => n23736, ZN => n23401);
   U24770 : INV_X1 port map( A => n24001, ZN => n24541);
   U24771 : NOR2_X1 port map( A1 => n22952, A2 => n24541, ZN => n22970);
   U24772 : INV_X1 port map( A => n22953, ZN => n23721);
   U24773 : INV_X1 port map( A => n22954, ZN => n23849);
   U24774 : INV_X1 port map( A => n23843, ZN => n23720);
   U24775 : NOR2_X1 port map( A1 => n23846, A2 => n23720, ZN => n22955);
   U24776 : NAND2_X1 port map( A1 => n23846, A2 => n28484, ZN => n23724);
   U24777 : INV_X1 port map( A => n24547, ZN => n22969);
   U24778 : MUX2_X1 port map( A => n6279, B => n23839, S => n487, Z => n22961);
   U24780 : NAND2_X1 port map( A1 => n28551, A2 => n23839, ZN => n22959);
   U24781 : NAND2_X1 port map( A1 => n23280, A2 => n23078, ZN => n22958);
   U24782 : NAND2_X1 port map( A1 => n22962, A2 => n23831, ZN => n22964);
   U24783 : NAND2_X1 port map( A1 => n23832, A2 => n23077, ZN => n22963);
   U24784 : NAND2_X1 port map( A1 => n22531, A2 => n23077, ZN => n23294);
   U24785 : NAND2_X1 port map( A1 => n23294, A2 => n23832, ZN => n22965);
   U24786 : NOR2_X1 port map( A1 => n24547, A2 => n24019, ZN => n22967);
   U24787 : NAND2_X1 port map( A1 => n24538, A2 => n24001, ZN => n23127);
   U24788 : INV_X1 port map( A => n22972, ZN => n22975);
   U24789 : OAI21_X1 port map( B1 => n23260, B2 => n22971, A => n380, ZN => 
                           n22974);
   U24790 : NAND2_X1 port map( A1 => n23585, A2 => n23587, ZN => n23586);
   U24791 : MUX2_X1 port map( A => n23586, B => n22972, S => n23716, Z => 
                           n22973);
   U24792 : NOR2_X1 port map( A1 => n22977, A2 => n22976, ZN => n23251);
   U24793 : INV_X1 port map( A => n23251, ZN => n22978);
   U24794 : NAND2_X1 port map( A1 => n22980, A2 => n22979, ZN => n23747);
   U24795 : NAND2_X1 port map( A1 => n22980, A2 => n28527, ZN => n22981);
   U24796 : AOI21_X1 port map( B1 => n22979, B2 => n22981, A => n23252, ZN => 
                           n22982);
   U24798 : INV_X1 port map( A => n22984, ZN => n23208);
   U24799 : INV_X1 port map( A => n23245, ZN => n23604);
   U24800 : INV_X1 port map( A => n23621, ZN => n23270);
   U24801 : NAND2_X1 port map( A1 => n23270, A2 => n22987, ZN => n23624);
   U24802 : OR2_X1 port map( A1 => n23624, A2 => n22986, ZN => n22990);
   U24803 : INV_X1 port map( A => n23620, ZN => n23569);
   U24804 : OAI22_X1 port map( A1 => n23618, A2 => n23622, B1 => n22987, B2 => 
                           n23569, ZN => n23184);
   U24805 : INV_X1 port map( A => n23184, ZN => n22989);
   U24806 : INV_X1 port map( A => n23626, ZN => n22988);
   U24808 : NAND2_X1 port map( A1 => n22991, A2 => n1838, ZN => n23183);
   U24809 : INV_X1 port map( A => n23183, ZN => n22994);
   U24810 : INV_X1 port map( A => n23563, ZN => n23317);
   U24812 : NAND2_X1 port map( A1 => n23180, A2 => n29074, ZN => n22998);
   U24814 : NOR2_X1 port map( A1 => n23615, A2 => n23216, ZN => n23000);
   U24815 : INV_X1 port map( A => n23267, ZN => n23610);
   U24816 : NOR2_X1 port map( A1 => n23610, A2 => n406, ZN => n22999);
   U24817 : MUX2_X1 port map( A => n23000, B => n22999, S => n28581, Z => 
                           n23003);
   U24818 : NOR2_X1 port map( A1 => n23001, A2 => n760, ZN => n23002);
   U24819 : NOR2_X2 port map( A1 => n23003, A2 => n23002, ZN => n24435);
   U24820 : AND3_X1 port map( A1 => n29128, A2 => n24437, A3 => n24434, ZN => 
                           n23004);
   U24821 : XNOR2_X1 port map( A => n28645, B => n25681, ZN => n24834);
   U24822 : NOR2_X1 port map( A1 => n23787, A2 => n23786, ZN => n23480);
   U24823 : OAI21_X1 port map( B1 => n23486, B2 => n23480, A => n473, ZN => 
                           n24686);
   U24824 : INV_X1 port map( A => n23162, ZN => n23522);
   U24825 : NOR2_X1 port map( A1 => n23006, A2 => n23522, ZN => n23007);
   U24826 : INV_X1 port map( A => n23662, ZN => n23667);
   U24830 : INV_X1 port map( A => n23014, ZN => n23015);
   U24831 : INV_X1 port map( A => n23016, ZN => n23680);
   U24832 : INV_X1 port map( A => n23134, ZN => n23019);
   U24833 : NOR2_X1 port map( A1 => n23516, A2 => n23680, ZN => n23018);
   U24834 : NAND2_X1 port map( A1 => n24682, A2 => n24688, ZN => n23020);
   U24835 : NAND2_X1 port map( A1 => n23513, A2 => n29641, ZN => n23022);
   U24836 : MUX2_X1 port map( A => n23022, B => n23021, S => n23512, Z => 
                           n24684);
   U24837 : NOR2_X1 port map( A1 => n23512, A2 => n339, ZN => n23023);
   U24838 : OAI21_X1 port map( B1 => n23023, B2 => n23488, A => n6424, ZN => 
                           n24685);
   U24839 : NAND2_X1 port map( A1 => n24684, A2 => n24685, ZN => n24310);
   U24840 : NAND2_X1 port map( A1 => n24391, A2 => n24688, ZN => n23025);
   U24841 : AOI21_X1 port map( B1 => n24682, B2 => n23025, A => n24390, ZN => 
                           n23026);
   U24842 : AND2_X1 port map( A1 => n23764, A2 => n23763, ZN => n23028);
   U24843 : NAND2_X1 port map( A1 => n23028, A2 => n23767, ZN => n23031);
   U24844 : NAND2_X1 port map( A1 => n23028, A2 => n23766, ZN => n23030);
   U24845 : NAND3_X1 port map( A1 => n23769, A2 => n23765, A3 => n28554, ZN => 
                           n23029);
   U24846 : NOR2_X1 port map( A1 => n23768, A2 => n23765, ZN => n23151);
   U24847 : INV_X1 port map( A => n23190, ZN => n23035);
   U24848 : INV_X1 port map( A => n23326, ZN => n23759);
   U24849 : INV_X1 port map( A => n23474, ZN => n23033);
   U24850 : NOR2_X1 port map( A1 => n23036, A2 => n473, ZN => n23154);
   U24851 : AOI21_X1 port map( B1 => n23785, B2 => n23787, A => n23484, ZN => 
                           n23038);
   U24852 : NAND2_X1 port map( A1 => n23783, A2 => n473, ZN => n23037);
   U24853 : AOI21_X1 port map( B1 => n24706, B2 => n29043, A => n24707, ZN => 
                           n23051);
   U24854 : INV_X1 port map( A => n23793, ZN => n23493);
   U24855 : NAND2_X1 port map( A1 => n23795, A2 => n23493, ZN => n23321);
   U24856 : INV_X1 port map( A => n23799, ZN => n23497);
   U24857 : NOR2_X1 port map( A1 => n23799, A2 => n23789, ZN => n23039);
   U24858 : INV_X1 port map( A => n23555, ZN => n23045);
   U24859 : NAND2_X1 port map( A1 => n23041, A2 => n477, ZN => n23044);
   U24860 : INV_X1 port map( A => n23630, ZN => n23559);
   U24861 : NAND2_X1 port map( A1 => n23559, A2 => n29061, ZN => n23042);
   U24862 : INV_X1 port map( A => n23194, ZN => n23046);
   U24863 : AOI21_X1 port map( B1 => n23470, B2 => n23472, A => n23046, ZN => 
                           n23047);
   U24864 : MUX2_X1 port map( A => n23048, B => n23047, S => n23469, Z => 
                           n24339);
   U24865 : NOR2_X1 port map( A1 => n23648, A2 => n661, ZN => n23050);
   U24866 : NAND2_X1 port map( A1 => n23193, A2 => n23050, ZN => n24334);
   U24867 : XNOR2_X1 port map( A => n25910, B => n28593, ZN => n24890);
   U24868 : XNOR2_X1 port map( A => n24834, B => n24890, ZN => n23125);
   U24869 : NAND2_X1 port map( A1 => n29295, A2 => n23445, ZN => n23052);
   U24870 : AOI21_X1 port map( B1 => n23052, B2 => n23442, A => n292, ZN => 
                           n23056);
   U24871 : INV_X1 port map( A => n23445, ZN => n23053);
   U24872 : NAND3_X1 port map( A1 => n23109, A2 => n23053, A3 => n292, ZN => 
                           n23055);
   U24873 : NAND3_X1 port map( A1 => n23370, A2 => n29295, A3 => n23445, ZN => 
                           n23054);
   U24874 : INV_X1 port map( A => n23138, ZN => n23057);
   U24875 : NAND2_X1 port map( A1 => n28570, A2 => n23057, ZN => n23058);
   U24876 : AND2_X1 port map( A1 => n23341, A2 => n23058, ZN => n23061);
   U24877 : NOR2_X1 port map( A1 => n28570, A2 => n28659, ZN => n23059);
   U24878 : NAND2_X1 port map( A1 => n23416, A2 => n485, ZN => n23062);
   U24879 : AOI21_X1 port map( B1 => n24713, B2 => n24716, A => n4136, ZN => 
                           n23072);
   U24880 : MUX2_X1 port map( A => n23454, B => n23148, S => n23456, Z => 
                           n23066);
   U24881 : INV_X1 port map( A => n23456, ZN => n23147);
   U24882 : MUX2_X2 port map( A => n23066, B => n23065, S => n23460, Z => 
                           n24712);
   U24883 : INV_X1 port map( A => n23676, ZN => n23364);
   U24884 : INV_X1 port map( A => n23672, ZN => n23366);
   U24885 : INV_X1 port map( A => n23673, ZN => n23107);
   U24886 : NOR2_X1 port map( A1 => n23107, A2 => n23363, ZN => n23068);
   U24887 : NOR2_X1 port map( A1 => n28604, A2 => n23131, ZN => n23674);
   U24888 : AND2_X1 port map( A1 => n24409, A2 => n24711, ZN => n24351);
   U24889 : INV_X1 port map( A => n24711, ZN => n24715);
   U24891 : XNOR2_X1 port map( A => n28769, B => n27737, ZN => n23123);
   U24892 : AND2_X1 port map( A1 => n28653, A2 => n23285, ZN => n23805);
   U24893 : INV_X1 port map( A => n23810, ZN => n23807);
   U24894 : NAND2_X1 port map( A1 => n22877, A2 => n23806, ZN => n23286);
   U24895 : INV_X1 port map( A => n24374, ZN => n24372);
   U24896 : NOR2_X1 port map( A1 => n24373, A2 => n24372, ZN => n23083);
   U24897 : OAI211_X1 port map( C1 => n23392, C2 => n23839, A => n487, B => 
                           n28418, ZN => n23080);
   U24898 : OAI21_X1 port map( B1 => n28551, B2 => n23078, A => n28460, ZN => 
                           n23079);
   U24899 : NOR2_X1 port map( A1 => n23995, A2 => n23994, ZN => n23082);
   U24900 : NOR2_X1 port map( A1 => n23301, A2 => n23433, ZN => n23085);
   U24901 : NOR2_X1 port map( A1 => n4178, A2 => n4020, ZN => n23084);
   U24902 : MUX2_X1 port map( A => n23085, B => n23084, S => n201, Z => n23088)
                           ;
   U24903 : MUX2_X1 port map( A => n1829, B => n408, S => n23433, Z => n23086);
   U24904 : NOR2_X1 port map( A1 => n23086, A2 => n5699, ZN => n23087);
   U24905 : NAND2_X1 port map( A1 => n22931, A2 => n28609, ZN => n23089);
   U24906 : NAND3_X1 port map( A1 => n23441, A2 => n23090, A3 => n23089, ZN => 
                           n23091);
   U24908 : OAI211_X1 port map( C1 => n23994, C2 => n23906, A => n23093, B => 
                           n24372, ZN => n23094);
   U24910 : OAI21_X1 port map( B1 => n23415, B2 => n23419, A => n23101, ZN => 
                           n23968);
   U24911 : INV_X1 port map( A => n23968, ZN => n23972);
   U24912 : NOR2_X1 port map( A1 => n1829, A2 => n29018, ZN => n23103);
   U24913 : NOR2_X1 port map( A1 => n23302, A2 => n23102, ZN => n23434);
   U24914 : OAI21_X1 port map( B1 => n23103, B2 => n23434, A => n4020, ZN => 
                           n23104);
   U24915 : INV_X1 port map( A => n24209, ZN => n24046);
   U24916 : AOI21_X1 port map( B1 => n23364, B2 => n23366, A => n23131, ZN => 
                           n23106);
   U24917 : NAND2_X1 port map( A1 => n29296, A2 => n23109, ZN => n23110);
   U24918 : NOR2_X1 port map( A1 => n469, A2 => n24479, ZN => n23970);
   U24919 : INV_X1 port map( A => n23422, ZN => n23428);
   U24920 : INV_X1 port map( A => n23338, ZN => n23426);
   U24921 : MUX2_X1 port map( A => n23138, B => n23427, S => n28659, Z => 
                           n23114);
   U24922 : INV_X1 port map( A => n23343, ZN => n23339);
   U24924 : NOR2_X1 port map( A1 => n23339, A2 => n28122, ZN => n23113);
   U24925 : INV_X1 port map( A => n29108, ZN => n23112);
   U24926 : AOI22_X1 port map( A1 => n23344, A2 => n23114, B1 => n23113, B2 => 
                           n23112, ZN => n23115);
   U24927 : OAI21_X1 port map( B1 => n23116, B2 => n23970, A => n24483, ZN => 
                           n23121);
   U24929 : NOR2_X1 port map( A1 => n23456, A2 => n29042, ZN => n23117);
   U24930 : INV_X1 port map( A => n23460, ZN => n23458);
   U24931 : AND2_X1 port map( A1 => n23455, A2 => n23460, ZN => n23355);
   U24932 : NAND2_X1 port map( A1 => n24484, A2 => n24209, ZN => n23119);
   U24933 : XNOR2_X1 port map( A => n28628, B => n25845, ZN => n23122);
   U24934 : XNOR2_X1 port map( A => n23122, B => n23123, ZN => n23124);
   U24935 : INV_X1 port map( A => n26789, ZN => n26575);
   U24936 : NAND2_X1 port map( A1 => n24542, A2 => n2823, ZN => n24540);
   U24937 : OAI21_X1 port map( B1 => n24540, B2 => n24160, A => n23128, ZN => 
                           n23130);
   U24939 : INV_X1 port map( A => n23683, ZN => n23517);
   U24940 : NOR2_X1 port map( A1 => n4232, A2 => n4231, ZN => n23142);
   U24941 : INV_X1 port map( A => n24891, ZN => n23144);
   U24942 : NAND2_X1 port map( A1 => n24631, A2 => n24629, ZN => n24530);
   U24943 : OAI21_X1 port map( B1 => n1837, B2 => n23461, A => n23458, ZN => 
                           n23146);
   U24944 : NAND2_X1 port map( A1 => n29042, A2 => n23456, ZN => n23457);
   U24945 : INV_X1 port map( A => n23767, ZN => n23329);
   U24946 : OAI21_X1 port map( B1 => n23764, B2 => n23763, A => n23769, ZN => 
                           n23152);
   U24947 : NAND2_X1 port map( A1 => n23768, A2 => n23152, ZN => n23153);
   U24948 : INV_X1 port map( A => n24642, ZN => n24568);
   U24949 : NAND3_X1 port map( A1 => n23785, A2 => n475, A3 => n23788, ZN => 
                           n23155);
   U24950 : NAND2_X1 port map( A1 => n24568, A2 => n24237, ZN => n24641);
   U24951 : NAND2_X1 port map( A1 => n23156, A2 => n23771, ZN => n23157);
   U24952 : INV_X1 port map( A => n23157, ZN => n23489);
   U24953 : OAI21_X1 port map( B1 => n23779, B2 => n23776, A => n23772, ZN => 
                           n23161);
   U24954 : NOR2_X1 port map( A1 => n23514, A2 => n23776, ZN => n23159);
   U24955 : AND2_X1 port map( A1 => n23666, A2 => n23162, ZN => n23527);
   U24956 : OAI21_X1 port map( B1 => n29123, B2 => n23163, A => n23527, ZN => 
                           n23166);
   U24957 : NAND2_X1 port map( A1 => n23164, A2 => n23663, ZN => n23165);
   U24958 : OAI211_X1 port map( C1 => n23662, C2 => n23663, A => n23166, B => 
                           n23165, ZN => n24638);
   U24959 : NAND2_X1 port map( A1 => n23169, A2 => n23016, ZN => n23171);
   U24962 : AOI21_X1 port map( B1 => n23801, B2 => n23800, A => n1913, ZN => 
                           n23174);
   U24963 : NOR2_X1 port map( A1 => n23537, A2 => n28444, ZN => n23172);
   U24965 : NOR3_X1 port map( A1 => n29074, A2 => n23177, A3 => n23563, ZN => 
                           n23179);
   U24966 : NAND2_X1 port map( A1 => n23621, A2 => n23619, ZN => n23568);
   U24967 : NAND2_X1 port map( A1 => n23568, A2 => n23620, ZN => n23185);
   U24968 : NAND2_X1 port map( A1 => n23185, A2 => n726, ZN => n23186);
   U24969 : NOR2_X1 port map( A1 => n24241, A2 => n24240, ZN => n23990);
   U24970 : NOR2_X1 port map( A1 => n5775, A2 => n23629, ZN => n23187);
   U24971 : NOR2_X1 port map( A1 => n23309, A2 => n28644, ZN => n23188);
   U24973 : MUX2_X1 port map( A => n23193, B => n23649, S => n23651, Z => 
                           n23195);
   U24974 : NAND2_X1 port map( A1 => n23196, A2 => n23492, ZN => n23197);
   U24975 : NAND2_X1 port map( A1 => n23197, A2 => n23792, ZN => n23200);
   U24979 : NAND2_X1 port map( A1 => n24239, A2 => n25794, ZN => n23201);
   U24980 : XNOR2_X1 port map( A => n25775, B => n26004, ZN => n25216);
   U24981 : XNOR2_X1 port map( A => n25216, B => n25563, ZN => n23244);
   U24982 : AOI21_X1 port map( B1 => n23202, B2 => n1883, A => n24377, ZN => 
                           n23204);
   U24983 : NOR3_X1 port map( A1 => n24373, A2 => n24374, A3 => n1883, ZN => 
                           n23203);
   U24984 : NAND2_X1 port map( A1 => n23936, A2 => n24553, ZN => n23206);
   U24985 : XNOR2_X1 port map( A => n29534, B => n25565, ZN => n23242);
   U24986 : NOR2_X1 port map( A1 => n23607, A2 => n23247, ZN => n23209);
   U24988 : NAND2_X1 port map( A1 => n23602, A2 => n23246, ZN => n23210);
   U24989 : OAI21_X1 port map( B1 => n23606, B2 => n23578, A => n23210, ZN => 
                           n23608);
   U24990 : INV_X1 port map( A => n23406, ZN => n23214);
   U24991 : OAI21_X1 port map( B1 => n23403, B2 => n23250, A => n23252, ZN => 
                           n23215);
   U24992 : AOI22_X1 port map( A1 => n23615, A2 => n23216, B1 => n28225, B2 => 
                           n28544, ZN => n23219);
   U24996 : NAND2_X1 port map( A1 => n1862, A2 => n23398, ZN => n23230);
   U24997 : INV_X1 port map( A => n23736, ZN => n23228);
   U24999 : NAND2_X1 port map( A1 => n24524, A2 => n28481, ZN => n23238);
   U25000 : NAND2_X1 port map( A1 => n380, A2 => n23714, ZN => n23713);
   U25004 : NAND2_X1 port map( A1 => n23238, A2 => n24245, ZN => n23239);
   U25005 : NOR2_X2 port map( A1 => n23240, A2 => n23239, ZN => n25346);
   U25006 : XNOR2_X1 port map( A => n25346, B => n1079, ZN => n23241);
   U25007 : XNOR2_X1 port map( A => n23242, B => n23241, ZN => n23243);
   U25008 : MUX2_X1 port map( A => n23602, B => n23246, S => n23245, Z => 
                           n23248);
   U25009 : AND2_X1 port map( A1 => n23406, A2 => n22979, ZN => n23254);
   U25010 : NOR2_X1 port map( A1 => n23213, A2 => n22979, ZN => n23253);
   U25011 : INV_X1 port map( A => n23258, ZN => n23256);
   U25012 : NAND2_X1 port map( A1 => n23732, A2 => n23257, ZN => n23259);
   U25014 : NOR2_X1 port map( A1 => n28528, A2 => n28415, ZN => n23269);
   U25015 : AOI21_X1 port map( B1 => n23267, B2 => n28582, A => n29115, ZN => 
                           n23268);
   U25016 : NOR2_X1 port map( A1 => n24368, A2 => n24369, ZN => n24064);
   U25019 : OAI21_X1 port map( B1 => n29564, B2 => n23382, A => n23825, ZN => 
                           n23276);
   U25020 : AOI21_X1 port map( B1 => n23385, B2 => n23382, A => n23276, ZN => 
                           n23279);
   U25021 : NAND3_X1 port map( A1 => n28181, A2 => n23382, A3 => n2187, ZN => 
                           n23277);
   U25022 : OAI21_X1 port map( B1 => n23738, B2 => n28181, A => n23277, ZN => 
                           n23278);
   U25024 : INV_X1 port map( A => n24083, ZN => n24084);
   U25025 : INV_X1 port map( A => n23281, ZN => n23282);
   U25026 : INV_X1 port map( A => n23285, ZN => n23287);
   U25027 : MUX2_X1 port map( A => n24084, B => n6265, S => n24403, Z => n23307
                           );
   U25028 : INV_X1 port map( A => n23291, ZN => n23816);
   U25029 : NOR3_X1 port map( A1 => n4950, A2 => n28182, A3 => n23290, ZN => 
                           n23292);
   U25030 : OAI22_X1 port map( A1 => n23292, A2 => n23821, B1 => n23819, B2 => 
                           n5591, ZN => n23293);
   U25031 : INV_X1 port map( A => n23294, ZN => n23300);
   U25032 : OAI21_X1 port map( B1 => n22531, B2 => n23295, A => n29602, ZN => 
                           n23299);
   U25033 : OAI21_X1 port map( B1 => n23301, B2 => n29018, A => n5530, ZN => 
                           n23304);
   U25034 : XNOR2_X1 port map( A => n26011, B => n25884, ZN => n23337);
   U25035 : NOR2_X1 port map( A1 => n23637, A2 => n23630, ZN => n23308);
   U25036 : OAI21_X1 port map( B1 => n23309, B2 => n5775, A => n477, ZN => 
                           n23311);
   U25038 : NAND2_X1 port map( A1 => n22992, A2 => n23640, ZN => n23313);
   U25039 : OAI21_X1 port map( B1 => n22996, B2 => n23314, A => n1838, ZN => 
                           n23316);
   U25041 : NOR2_X1 port map( A1 => n24395, A2 => n28635, ZN => n24068);
   U25042 : NOR2_X1 port map( A1 => n23320, A2 => n23792, ZN => n23322);
   U25043 : NOR2_X1 port map( A1 => n24678, A2 => n24672, ZN => n23324);
   U25044 : NOR2_X1 port map( A1 => n24068, A2 => n23324, ZN => n23334);
   U25045 : INV_X1 port map( A => n28635, ZN => n24676);
   U25046 : MUX2_X1 port map( A => n23758, B => n23326, S => n29131, Z => 
                           n23327);
   U25048 : NAND2_X1 port map( A1 => n4759, A2 => n23769, ZN => n23332);
   U25049 : NAND2_X1 port map( A1 => n23764, A2 => n28554, ZN => n23330);
   U25050 : MUX2_X1 port map( A => n23330, B => n23501, S => n23767, Z => 
                           n23331);
   U25052 : AND2_X1 port map( A1 => n29471, A2 => n24688, ZN => n23335);
   U25053 : AOI22_X1 port map( A1 => n466, A2 => n23335, B1 => n24682, B2 => 
                           n24391, ZN => n23336);
   U25054 : XNOR2_X1 port map( A => n25761, B => n25444, ZN => n25234);
   U25055 : XNOR2_X1 port map( A => n25234, B => n23337, ZN => n23414);
   U25056 : NAND2_X1 port map( A1 => n23339, A2 => n23338, ZN => n23342);
   U25057 : NOR3_X1 port map( A1 => n23344, A2 => n29108, A3 => n28570, ZN => 
                           n23345);
   U25059 : MUX2_X1 port map( A => n23535, B => n5030, S => n28164, Z => n23350
                           );
   U25060 : NAND2_X1 port map( A1 => n23696, A2 => n23529, ZN => n23347);
   U25061 : MUX2_X1 port map( A => n23348, B => n23347, S => n23535, Z => 
                           n23349);
   U25062 : INV_X1 port map( A => n24665, ZN => n24382);
   U25063 : AOI21_X1 port map( B1 => n23657, B2 => n23351, A => n29583, ZN => 
                           n23352);
   U25064 : NAND2_X1 port map( A1 => n4605, A2 => n4195, ZN => n23375);
   U25065 : NAND2_X1 port map( A1 => n23355, A2 => n29042, ZN => n23359);
   U25066 : INV_X1 port map( A => n23356, ZN => n23358);
   U25067 : NOR2_X1 port map( A1 => n24665, A2 => n24666, ZN => n23373);
   U25069 : MUX2_X1 port map( A => n23362, B => n23361, S => n23360, Z => 
                           n23369);
   U25070 : AOI21_X1 port map( B1 => n23367, B2 => n23366, A => n23365, ZN => 
                           n23368);
   U25071 : NOR2_X1 port map( A1 => n24382, A2 => n24668, ZN => n24073);
   U25072 : INV_X1 port map( A => n23370, ZN => n23371);
   U25073 : NAND2_X1 port map( A1 => n24316, A2 => n24383, ZN => n23372);
   U25075 : AOI21_X1 port map( B1 => n24374, B2 => n1828, A => n24373, ZN => 
                           n23376);
   U25076 : NAND2_X1 port map( A1 => n23906, A2 => n24376, ZN => n23380);
   U25077 : NAND2_X1 port map( A1 => n1828, A2 => n24380, ZN => n23378);
   U25078 : XNOR2_X1 port map( A => n25933, B => n25931, ZN => n23412);
   U25079 : NAND2_X1 port map( A1 => n23738, A2 => n23827, ZN => n23384);
   U25080 : OAI21_X1 port map( B1 => n22451, B2 => n29618, A => n23702, ZN => 
                           n23388);
   U25081 : OAI21_X1 port map( B1 => n23722, B2 => n28484, A => n23726, ZN => 
                           n23395);
   U25082 : NOR2_X1 port map( A1 => n28484, A2 => n23720, ZN => n23394);
   U25083 : INV_X1 port map( A => n24388, ZN => n23911);
   U25084 : OAI211_X1 port map( C1 => n23228, C2 => n23399, A => n23398, B => 
                           n23397, ZN => n23400);
   U25085 : NOR2_X1 port map( A1 => n23403, A2 => n28527, ZN => n23404);
   U25086 : NAND3_X1 port map( A1 => n24133, A2 => n24388, A3 => n24078, ZN => 
                           n23409);
   U25087 : XNOR2_X1 port map( A => n25179, B => n622, ZN => n23411);
   U25088 : XNOR2_X1 port map( A => n23412, B => n23411, ZN => n23413);
   U25090 : NAND2_X1 port map( A1 => n23422, A2 => n28659, ZN => n23423);
   U25091 : NAND2_X1 port map( A1 => n23424, A2 => n23423, ZN => n23429);
   U25092 : NOR2_X1 port map( A1 => n1829, A2 => n408, ZN => n23437);
   U25093 : NAND2_X1 port map( A1 => n4020, A2 => n23431, ZN => n23436);
   U25094 : OAI21_X1 port map( B1 => n23433, B2 => n29018, A => n23431, ZN => 
                           n23435);
   U25095 : NAND2_X1 port map( A1 => n4950, A2 => n28182, ZN => n23440);
   U25096 : NAND3_X1 port map( A1 => n2281, A2 => n4950, A3 => n22931, ZN => 
                           n23438);
   U25097 : NOR2_X1 port map( A1 => n23445, A2 => n23442, ZN => n23443);
   U25098 : NAND3_X1 port map( A1 => n23447, A2 => n23446, A3 => n23445, ZN => 
                           n23452);
   U25099 : NAND3_X1 port map( A1 => n29296, A2 => n23449, A3 => n292, ZN => 
                           n23451);
   U25100 : MUX2_X1 port map( A => n23456, B => n23455, S => n23454, Z => 
                           n23466);
   U25101 : INV_X1 port map( A => n23457, ZN => n23459);
   U25102 : AND2_X1 port map( A1 => n23460, A2 => n23461, ZN => n23462);
   U25103 : NAND2_X1 port map( A1 => n23462, A2 => n23465, ZN => n23463);
   U25105 : OR2_X1 port map( A1 => n24012, A2 => n23597, ZN => n23468);
   U25106 : INV_X1 port map( A => n23475, ZN => n23479);
   U25107 : OAI21_X1 port map( B1 => n23758, B2 => n23759, A => n23761, ZN => 
                           n23478);
   U25108 : MUX2_X1 port map( A => n23476, B => n23475, S => n23474, Z => 
                           n23477);
   U25109 : NOR2_X1 port map( A1 => n24775, A2 => n470, ZN => n23502);
   U25110 : INV_X1 port map( A => n23480, ZN => n23481);
   U25111 : NOR2_X1 port map( A1 => n23481, A2 => n23788, ZN => n23485);
   U25112 : NAND2_X1 port map( A1 => n23482, A2 => n23784, ZN => n23483);
   U25113 : INV_X1 port map( A => n24777, ZN => n24780);
   U25114 : OAI22_X1 port map( A1 => n23157, A2 => n23778, B1 => n23514, B2 => 
                           n29641, ZN => n23490);
   U25115 : NAND3_X1 port map( A1 => n23493, A2 => n23789, A3 => n23492, ZN => 
                           n23494);
   U25116 : OAI21_X1 port map( B1 => n23495, B2 => n23795, A => n23494, ZN => 
                           n23496);
   U25117 : AOI21_X2 port map( B1 => n23498, B2 => n23497, A => n23496, ZN => 
                           n24776);
   U25118 : NOR2_X1 port map( A1 => n23946, A2 => n24776, ZN => n24454);
   U25119 : OAI21_X1 port map( B1 => n23499, B2 => n23765, A => n23764, ZN => 
                           n23500);
   U25120 : XNOR2_X1 port map( A => n25282, B => n26029, ZN => n23511);
   U25121 : NAND2_X1 port map( A1 => n24083, A2 => n24408, ZN => n23504);
   U25122 : MUX2_X1 port map( A => n23504, B => n23503, S => n24404, Z => 
                           n23505);
   U25123 : MUX2_X1 port map( A => n24077, B => n24388, S => n24387, Z => 
                           n23510);
   U25125 : XNOR2_X1 port map( A => n25324, B => n25751, ZN => n24307);
   U25126 : XNOR2_X1 port map( A => n23511, B => n24307, ZN => n23596);
   U25128 : MUX2_X2 port map( A => n23521, B => n23520, S => n23016, Z => 
                           n24772);
   U25130 : MUX2_X1 port map( A => n23524, B => n23523, S => n23663, Z => 
                           n23528);
   U25131 : NOR2_X1 port map( A1 => n23666, A2 => n23525, ZN => n23526);
   U25132 : MUX2_X1 port map( A => n24697, B => n24772, S => n24765, Z => 
                           n23550);
   U25133 : NAND2_X1 port map( A1 => n23531, A2 => n23697, ZN => n23534);
   U25135 : INV_X1 port map( A => n23689, ZN => n23539);
   U25136 : INV_X1 port map( A => n23540, ZN => n23542);
   U25138 : NOR2_X1 port map( A1 => n24769, A2 => n29624, ZN => n23547);
   U25139 : AOI21_X2 port map( B1 => n23550, B2 => n28598, A => n23549, ZN => 
                           n25037);
   U25142 : INV_X1 port map( A => n24484, ZN => n24213);
   U25143 : NAND3_X1 port map( A1 => n24213, A2 => n29597, A3 => n24209, ZN => 
                           n23552);
   U25144 : NAND3_X1 port map( A1 => n24480, A2 => n24210, A3 => n24483, ZN => 
                           n23551);
   U25145 : OAI211_X2 port map( C1 => n24482, C2 => n23553, A => n23552, B => 
                           n23551, ZN => n25209);
   U25146 : XNOR2_X1 port map( A => n25037, B => n25209, ZN => n25939);
   U25147 : NAND2_X1 port map( A1 => n23559, A2 => n23558, ZN => n23560);
   U25148 : NOR3_X1 port map( A1 => n29115, A2 => n379, A3 => n28225, ZN => 
                           n23955);
   U25149 : INV_X1 port map( A => n23955, ZN => n24218);
   U25150 : NAND2_X1 port map( A1 => n24447, A2 => n24218, ZN => n23576);
   U25151 : NAND2_X1 port map( A1 => n23641, A2 => n23563, ZN => n23646);
   U25152 : NOR2_X1 port map( A1 => n23618, A2 => n23621, ZN => n23574);
   U25153 : OAI21_X1 port map( B1 => n23567, B2 => n23566, A => n23622, ZN => 
                           n23573);
   U25154 : INV_X1 port map( A => n23568, ZN => n23571);
   U25155 : NOR2_X1 port map( A1 => n23621, A2 => n23569, ZN => n23570);
   U25156 : INV_X1 port map( A => n24760, ZN => n23588);
   U25157 : AOI21_X1 port map( B1 => n29592, B2 => n24761, A => n23588, ZN => 
                           n23575);
   U25158 : MUX2_X1 port map( A => n5347, B => n23578, S => n23577, Z => n23582
                           );
   U25159 : NAND2_X1 port map( A1 => n23583, A2 => n23603, ZN => n23580);
   U25160 : NAND2_X1 port map( A1 => n23607, A2 => n23578, ZN => n23579);
   U25161 : MUX2_X1 port map( A => n23580, B => n23579, S => n5347, Z => n23581
                           );
   U25162 : INV_X1 port map( A => n24757, ZN => n24220);
   U25163 : OAI21_X1 port map( B1 => n24220, B2 => n24756, A => n23588, ZN => 
                           n23591);
   U25164 : INV_X1 port map( A => n23956, ZN => n23589);
   U25165 : AOI21_X1 port map( B1 => n23589, B2 => n24218, A => n28509, ZN => 
                           n23590);
   U25167 : INV_X1 port map( A => n2544, ZN => n23593);
   U25168 : XNOR2_X1 port map( A => n25785, B => n23593, ZN => n23594);
   U25169 : XNOR2_X1 port map( A => n25939, B => n23594, ZN => n23595);
   U25170 : XNOR2_X1 port map( A => n23595, B => n23596, ZN => n26791);
   U25172 : NOR2_X1 port map( A1 => n24972, A2 => n24256, ZN => n23598);
   U25173 : OAI21_X1 port map( B1 => n23604, B2 => n23603, A => n23602, ZN => 
                           n23605);
   U25175 : NAND3_X1 port map( A1 => n4599, A2 => n23610, A3 => n28581, ZN => 
                           n23617);
   U25176 : MUX2_X1 port map( A => n23611, B => n23615, S => n379, Z => n23613)
                           ;
   U25177 : NOR2_X1 port map( A1 => n24790, A2 => n24791, ZN => n24507);
   U25178 : AOI21_X1 port map( B1 => n23622, B2 => n23619, A => n23618, ZN => 
                           n23625);
   U25179 : NOR2_X1 port map( A1 => n23621, A2 => n23620, ZN => n23623);
   U25180 : INV_X1 port map( A => n24790, ZN => n24792);
   U25181 : AOI21_X1 port map( B1 => n23630, B2 => n23629, A => n23628, ZN => 
                           n23635);
   U25182 : NOR2_X1 port map( A1 => n23632, A2 => n28644, ZN => n23634);
   U25183 : MUX2_X1 port map( A => n23635, B => n23634, S => n29061, Z => 
                           n23639);
   U25184 : NOR2_X1 port map( A1 => n23637, A2 => n23636, ZN => n23638);
   U25185 : OR2_X2 port map( A1 => n23639, A2 => n23638, ZN => n24269);
   U25186 : NOR2_X1 port map( A1 => n23641, A2 => n23640, ZN => n23644);
   U25187 : NAND2_X1 port map( A1 => n23648, A2 => n23647, ZN => n23650);
   U25188 : XNOR2_X1 port map( A => n25944, B => n25826, ZN => n23756);
   U25189 : NOR2_X1 port map( A1 => n23656, A2 => n23657, ZN => n23660);
   U25190 : NOR2_X1 port map( A1 => n23662, A2 => n28577, ZN => n23664);
   U25191 : NOR2_X1 port map( A1 => n23666, A2 => n23665, ZN => n23668);
   U25192 : NOR3_X1 port map( A1 => n23669, A2 => n23668, A3 => n23667, ZN => 
                           n23670);
   U25194 : NOR2_X1 port map( A1 => n23673, A2 => n23672, ZN => n23675);
   U25195 : AOI21_X1 port map( B1 => n28604, B2 => n23675, A => n23674, ZN => 
                           n23677);
   U25196 : INV_X1 port map( A => n23681, ZN => n23685);
   U25197 : NOR2_X1 port map( A1 => n23016, A2 => n23682, ZN => n23684);
   U25198 : NOR2_X1 port map( A1 => n24808, A2 => n24817, ZN => n23691);
   U25199 : OAI21_X1 port map( B1 => n23801, B2 => n23687, A => n23800, ZN => 
                           n23688);
   U25200 : MUX2_X1 port map( A => n23692, B => n23691, S => n5004, Z => n23699
                           );
   U25201 : INV_X1 port map( A => n24817, ZN => n24461);
   U25202 : NAND2_X1 port map( A1 => n484, A2 => n23067, ZN => n23695);
   U25203 : NOR2_X2 port map( A1 => n23699, A2 => n23698, ZN => n25943);
   U25204 : NOR2_X1 port map( A1 => n22084, A2 => n23700, ZN => n23703);
   U25205 : MUX2_X1 port map( A => n23704, B => n23703, S => n23387, Z => 
                           n23709);
   U25206 : NOR2_X2 port map( A1 => n23709, A2 => n23708, ZN => n24111);
   U25207 : INV_X1 port map( A => n24111, ZN => n24179);
   U25208 : NAND2_X1 port map( A1 => n23714, A2 => n23710, ZN => n23711);
   U25209 : MUX2_X1 port map( A => n23712, B => n23711, S => n23715, Z => 
                           n23719);
   U25210 : OAI21_X1 port map( B1 => n23715, B2 => n23714, A => n23713, ZN => 
                           n23717);
   U25211 : NAND2_X1 port map( A1 => n23717, A2 => n23716, ZN => n23718);
   U25212 : INV_X1 port map( A => n24517, ZN => n24113);
   U25213 : MUX2_X1 port map( A => n23722, B => n23721, S => n23720, Z => 
                           n23723);
   U25214 : NOR2_X1 port map( A1 => n23724, A2 => n23843, ZN => n23729);
   U25215 : NOR2_X1 port map( A1 => n23849, A2 => n28484, ZN => n23727);
   U25217 : INV_X1 port map( A => n23745, ZN => n24515);
   U25218 : NOR2_X1 port map( A1 => n24520, A2 => n24515, ZN => n23744);
   U25219 : INV_X1 port map( A => n23738, ZN => n23739);
   U25220 : OAI21_X1 port map( B1 => n28181, B2 => n23827, A => n23739, ZN => 
                           n23740);
   U25221 : OAI21_X2 port map( B1 => n23743, B2 => n23382, A => n23742, ZN => 
                           n24514);
   U25222 : NAND2_X1 port map( A1 => n24515, A2 => n24514, ZN => n24424);
   U25223 : NOR2_X1 port map( A1 => n24516, A2 => n24111, ZN => n23752);
   U25224 : INV_X1 port map( A => n23746, ZN => n23751);
   U25226 : XNOR2_X1 port map( A => n25943, B => n26056, ZN => n23755);
   U25227 : XNOR2_X1 port map( A => n23756, B => n23755, ZN => n23861);
   U25228 : NAND2_X1 port map( A1 => n23764, A2 => n23765, ZN => n23770);
   U25229 : NOR2_X1 port map( A1 => n339, A2 => n23771, ZN => n23775);
   U25230 : NOR2_X1 port map( A1 => n29641, A2 => n23772, ZN => n23774);
   U25231 : MUX2_X1 port map( A => n23775, B => n23774, S => n23776, Z => 
                           n23782);
   U25232 : AOI21_X1 port map( B1 => n23780, B2 => n23779, A => n23778, ZN => 
                           n23781);
   U25234 : MUX2_X1 port map( A => n24162, B => n24503, S => n24801, Z => 
                           n23804);
   U25236 : MUX2_X1 port map( A => n23790, B => n23789, S => n23791, Z => 
                           n23798);
   U25237 : NAND3_X1 port map( A1 => n6608, A2 => n23792, A3 => n23791, ZN => 
                           n23794);
   U25238 : OAI21_X1 port map( B1 => n23796, B2 => n23795, A => n23794, ZN => 
                           n23797);
   U25239 : NOR2_X1 port map( A1 => n22742, A2 => n23808, ZN => n23812);
   U25240 : OAI21_X1 port map( B1 => n23812, B2 => n23811, A => n23810, ZN => 
                           n23813);
   U25241 : NOR2_X1 port map( A1 => n23819, A2 => n23816, ZN => n23817);
   U25244 : AND2_X1 port map( A1 => n23842, A2 => n24472, ZN => n24475);
   U25245 : OAI211_X1 port map( C1 => n23829, C2 => n482, A => n28181, B => 
                           n23827, ZN => n24091);
   U25246 : NOR2_X1 port map( A1 => n23832, A2 => n29602, ZN => n23834);
   U25247 : NOR2_X1 port map( A1 => n24471, A2 => n29051, ZN => n23841);
   U25248 : NAND3_X1 port map( A1 => n6279, A2 => n28460, A3 => n23839, ZN => 
                           n23840);
   U25249 : INV_X1 port map( A => n23842, ZN => n24100);
   U25250 : XNOR2_X1 port map( A => n24949, B => n26054, ZN => n23859);
   U25251 : NOR2_X1 port map( A1 => n23853, A2 => n24141, ZN => n23857);
   U25252 : INV_X1 port map( A => n24591, ZN => n24143);
   U25253 : NOR2_X1 port map( A1 => n24143, A2 => n24592, ZN => n23854);
   U25254 : XNOR2_X1 port map( A => n25858, B => n3081, ZN => n23858);
   U25255 : XNOR2_X1 port map( A => n23858, B => n23859, ZN => n23860);
   U25256 : INV_X1 port map( A => n26793, ZN => n26572);
   U25257 : NOR2_X1 port map( A1 => n23863, A2 => n6826, ZN => n23864);
   U25258 : INV_X1 port map( A => n307, ZN => n24364);
   U25259 : INV_X1 port map( A => n24767, ZN => n24426);
   U25260 : MUX2_X1 port map( A => n1856, B => n24426, S => n24765, Z => n23866
                           );
   U25261 : MUX2_X1 port map( A => n24765, B => n24427, S => n24772, Z => 
                           n23865);
   U25262 : MUX2_X1 port map( A => n24711, B => n24716, S => n24712, Z => 
                           n23868);
   U25263 : INV_X1 port map( A => n24409, ZN => n24720);
   U25265 : INV_X1 port map( A => n24514, ZN => n24421);
   U25266 : NOR2_X1 port map( A1 => n24111, A2 => n24420, ZN => n24518);
   U25267 : INV_X1 port map( A => n24518, ZN => n23871);
   U25270 : XNOR2_X1 port map( A => n26073, B => n26040, ZN => n25687);
   U25271 : XNOR2_X1 port map( A => n25687, B => n25260, ZN => n23893);
   U25272 : INV_X1 port map( A => n23874, ZN => n24474);
   U25273 : NAND2_X1 port map( A1 => n24474, A2 => n24471, ZN => n24490);
   U25274 : INV_X1 port map( A => n24490, ZN => n23879);
   U25275 : INV_X1 port map( A => n24472, ZN => n24491);
   U25276 : NAND2_X1 port map( A1 => n24491, A2 => n24100, ZN => n23876);
   U25277 : MUX2_X1 port map( A => n24408, B => n24085, S => n24405, Z => 
                           n23883);
   U25278 : NAND2_X1 port map( A1 => n24403, A2 => n24084, ZN => n23881);
   U25279 : MUX2_X1 port map( A => n23881, B => n23880, S => n24405, Z => 
                           n23882);
   U25280 : OAI21_X2 port map( B1 => n23883, B2 => n24403, A => n23882, ZN => 
                           n26045);
   U25281 : XNOR2_X1 port map( A => n1922, B => n26045, ZN => n23891);
   U25282 : NAND2_X1 port map( A1 => n24347, A2 => n29726, ZN => n23884);
   U25284 : XNOR2_X1 port map( A => n28540, B => n624, ZN => n23890);
   U25285 : XNOR2_X1 port map( A => n23891, B => n23890, ZN => n23892);
   U25286 : INV_X1 port map( A => n26179, ZN => n26456);
   U25287 : NAND2_X1 port map( A1 => n24323, A2 => n28635, ZN => n23896);
   U25288 : NAND2_X1 port map( A1 => n24678, A2 => n24672, ZN => n24396);
   U25289 : NAND2_X1 port map( A1 => n24396, A2 => n6944, ZN => n23894);
   U25290 : NAND2_X1 port map( A1 => n24068, A2 => n24677, ZN => n23895);
   U25291 : AND3_X1 port map( A1 => n24369, A2 => n24304, A3 => n25005, ZN => 
                           n23898);
   U25292 : XNOR2_X1 port map( A => n25532, B => n25855, ZN => n25150);
   U25293 : INV_X1 port map( A => n24691, ZN => n23899);
   U25295 : NOR2_X1 port map( A1 => n24682, A2 => n24391, ZN => n23902);
   U25296 : NOR2_X1 port map( A1 => n466, A2 => n29567, ZN => n23901);
   U25297 : NOR2_X1 port map( A1 => n23905, A2 => n24372, ZN => n23907);
   U25298 : XNOR2_X1 port map( A => n25246, B => n26055, ZN => n23908);
   U25299 : XNOR2_X1 port map( A => n25150, B => n23908, ZN => n23920);
   U25300 : XNOR2_X1 port map( A => n25375, B => n27978, ZN => n23918);
   U25301 : INV_X1 port map( A => n24387, ZN => n24079);
   U25302 : NOR2_X1 port map( A1 => n28424, A2 => n24072, ZN => n23917);
   U25303 : NAND2_X1 port map( A1 => n23914, A2 => n4195, ZN => n23916);
   U25304 : NAND2_X1 port map( A1 => n24668, A2 => n24383, ZN => n23913);
   U25306 : XNOR2_X1 port map( A => n26060, B => n25372, ZN => n25698);
   U25307 : XNOR2_X1 port map( A => n23918, B => n25698, ZN => n23919);
   U25308 : NAND2_X1 port map( A1 => n26456, A2 => n26449, ZN => n25622);
   U25309 : INV_X1 port map( A => n24610, ZN => n23953);
   U25310 : OAI21_X1 port map( B1 => n23953, B2 => n24057, A => n24614, ZN => 
                           n23923);
   U25311 : XNOR2_X1 port map( A => n25848, B => n29543, ZN => n25310);
   U25313 : NOR2_X1 port map( A1 => n24617, A2 => n24747, ZN => n24022);
   U25314 : NOR2_X1 port map( A1 => n21303, A2 => n24617, ZN => n23926);
   U25315 : AOI22_X1 port map( A1 => n28223, A2 => n24022, B1 => n23926, B2 => 
                           n24751, ZN => n23927);
   U25316 : OAI21_X1 port map( B1 => n24593, B2 => n24277, A => n24590, ZN => 
                           n23930);
   U25317 : XNOR2_X1 port map( A => n25328, B => n25249, ZN => n26021);
   U25318 : XNOR2_X1 port map( A => n26021, B => n25310, ZN => n23941);
   U25319 : OAI21_X1 port map( B1 => n24596, B2 => n24597, A => n24595, ZN => 
                           n23934);
   U25320 : XNOR2_X1 port map( A => n25808, B => n2477, ZN => n23939);
   U25321 : INV_X1 port map( A => n24734, ZN => n24601);
   U25322 : OAI21_X1 port map( B1 => n24601, B2 => n24736, A => n24602, ZN => 
                           n23935);
   U25324 : OAI21_X1 port map( B1 => n24555, B2 => n24551, A => n28519, ZN => 
                           n23937);
   U25325 : XNOR2_X1 port map( A => n25133, B => n25396, ZN => n23938);
   U25326 : XNOR2_X1 port map( A => n23939, B => n23938, ZN => n23940);
   U25327 : INV_X1 port map( A => n24471, ZN => n23942);
   U25329 : NOR2_X1 port map( A1 => n23945, A2 => n29308, ZN => n24040);
   U25330 : INV_X1 port map( A => n24040, ZN => n24456);
   U25331 : OAI21_X1 port map( B1 => n23946, B2 => n24777, A => n29308, ZN => 
                           n23947);
   U25332 : NAND2_X1 port map( A1 => n24456, A2 => n23947, ZN => n23949);
   U25333 : OAI211_X1 port map( C1 => n24779, C2 => n24775, A => n24777, B => 
                           n24776, ZN => n23948);
   U25334 : XNOR2_X1 port map( A => n25708, B => n25922, ZN => n23952);
   U25335 : AOI21_X1 port map( B1 => n5004, B2 => n24808, A => n24499, ZN => 
                           n23950);
   U25337 : XNOR2_X1 port map( A => n23952, B => n29111, ZN => n25258);
   U25338 : OAI211_X1 port map( C1 => n5168, C2 => n24017, A => n24057, B => 
                           n23953, ZN => n23954);
   U25339 : AOI21_X1 port map( B1 => n24220, B2 => n28509, A => n378, ZN => 
                           n23959);
   U25340 : AND2_X1 port map( A1 => n24760, A2 => n24756, ZN => n24450);
   U25341 : INV_X1 port map( A => n24450, ZN => n23957);
   U25342 : XNOR2_X1 port map( A => n25868, B => n27515, ZN => n23960);
   U25343 : XNOR2_X1 port map( A => n23960, B => n25773, ZN => n23961);
   U25344 : INV_X1 port map( A => n23962, ZN => n24467);
   U25347 : INV_X1 port map( A => n24055, ZN => n23966);
   U25349 : MUX2_X1 port map( A => n24484, B => n469, S => n23968, Z => n24050)
                           ;
   U25350 : NAND2_X1 port map( A1 => n24050, A2 => n23969, ZN => n23975);
   U25351 : INV_X1 port map( A => n23970, ZN => n23974);
   U25352 : INV_X1 port map( A => n24483, ZN => n23971);
   U25353 : AND3_X1 port map( A1 => n23972, A2 => n24480, A3 => n23971, ZN => 
                           n23973);
   U25355 : XNOR2_X1 port map( A => n25187, B => n28485, ZN => n25713);
   U25356 : INV_X1 port map( A => n24556, ZN => n24174);
   U25357 : NOR2_X1 port map( A1 => n24174, A2 => n24552, ZN => n23977);
   U25358 : MUX2_X1 port map( A => n24555, B => n24551, S => n24173, Z => 
                           n23976);
   U25359 : NAND2_X1 port map( A1 => n23981, A2 => n23980, ZN => n25270);
   U25361 : NAND2_X1 port map( A1 => n29642, A2 => n24642, ZN => n24639);
   U25362 : NOR2_X1 port map( A1 => n24237, A2 => n24644, ZN => n24231);
   U25363 : NAND2_X1 port map( A1 => n24231, A2 => n24568, ZN => n23987);
   U25364 : INV_X1 port map( A => n24645, ZN => n24232);
   U25365 : NAND2_X1 port map( A1 => n2209, A2 => n24638, ZN => n23985);
   U25366 : OAI211_X1 port map( C1 => n24232, C2 => n2209, A => n29645, B => 
                           n23985, ZN => n23986);
   U25367 : OAI211_X1 port map( C1 => n2209, C2 => n24639, A => n23987, B => 
                           n23986, ZN => n24984);
   U25368 : XNOR2_X1 port map( A => n28534, B => n25781, ZN => n23988);
   U25369 : XNOR2_X1 port map( A => n25056, B => n23988, ZN => n24011);
   U25370 : INV_X1 port map( A => n24634, ZN => n24557);
   U25371 : NOR2_X1 port map( A1 => n24637, A2 => n23990, ZN => n23991);
   U25372 : NOR2_X2 port map( A1 => n23992, A2 => n23991, ZN => n25516);
   U25373 : NAND2_X1 port map( A1 => n24380, A2 => n24372, ZN => n23993);
   U25374 : OAI21_X1 port map( B1 => n24373, B2 => n24380, A => n23993, ZN => 
                           n23999);
   U25375 : NAND2_X1 port map( A1 => n24373, A2 => n24374, ZN => n23997);
   U25378 : XNOR2_X1 port map( A => n28654, B => n2996, ZN => n24000);
   U25379 : XNOR2_X1 port map( A => n25516, B => n24000, ZN => n24009);
   U25380 : MUX2_X1 port map( A => n24542, B => n2823, S => n24541, Z => n24004
                           );
   U25381 : OAI22_X1 port map( A1 => n24547, A2 => n24002, B1 => n24542, B2 => 
                           n24159, ZN => n24003);
   U25384 : XNOR2_X1 port map( A => n26109, B => n25577, ZN => n24008);
   U25385 : XNOR2_X1 port map( A => n24009, B => n24008, ZN => n24010);
   U25386 : XNOR2_X1 port map( A => n24011, B => n24010, ZN => n26454);
   U25387 : NAND2_X1 port map( A1 => n26452, A2 => n26454, ZN => n25415);
   U25388 : NOR2_X1 port map( A1 => n26456, A2 => n25415, ZN => n24038);
   U25389 : NOR2_X1 port map( A1 => n24972, A2 => n471, ZN => n24974);
   U25390 : INV_X1 port map( A => n24012, ZN => n24980);
   U25391 : AOI21_X1 port map( B1 => n24976, B2 => n24974, A => n24980, ZN => 
                           n24013);
   U25392 : OAI21_X1 port map( B1 => n24014, B2 => n23597, A => n24013, ZN => 
                           n24018);
   U25393 : MUX2_X1 port map( A => n24610, B => n24614, S => n24613, Z => 
                           n24015);
   U25394 : INV_X1 port map( A => n24015, ZN => n24016);
   U25395 : INV_X1 port map( A => n24017, ZN => n24609);
   U25396 : XNOR2_X1 port map( A => n24018, B => n24852, ZN => n26013);
   U25398 : XNOR2_X1 port map( A => n25381, B => n2522, ZN => n24021);
   U25399 : XNOR2_X1 port map( A => n26013, B => n24021, ZN => n24036);
   U25402 : NAND2_X1 port map( A1 => n462, A2 => n24751, ZN => n24618);
   U25403 : OAI21_X1 port map( B1 => n28223, B2 => n24024, A => n24618, ZN => 
                           n24025);
   U25404 : INV_X1 port map( A => n28785, ZN => n24029);
   U25405 : AOI21_X1 port map( B1 => n1955, B2 => n24792, A => n24507, ZN => 
                           n24034);
   U25406 : MUX2_X1 port map( A => n24789, B => n24794, S => n28455, Z => 
                           n24033);
   U25407 : NOR2_X1 port map( A1 => n28455, A2 => n24791, ZN => n24032);
   U25409 : XNOR2_X1 port map( A => n25703, B => n29073, ZN => n25408);
   U25410 : XNOR2_X1 port map( A => n25412, B => n25408, ZN => n24035);
   U25411 : XNOR2_X1 port map( A => n24035, B => n24036, ZN => n26450);
   U25412 : INV_X1 port map( A => n26450, ZN => n26162);
   U25413 : NAND3_X1 port map( A1 => n26162, A2 => n26448, A3 => n26449, ZN => 
                           n24037);
   U25414 : MUX2_X1 port map( A => n29308, B => n24776, S => n24777, Z => 
                           n24043);
   U25415 : NAND2_X1 port map( A1 => n24040, A2 => n24779, ZN => n24042);
   U25416 : NAND3_X1 port map( A1 => n23946, A2 => n24776, A3 => n29308, ZN => 
                           n24041);
   U25417 : OAI211_X1 port map( C1 => n24043, C2 => n463, A => n24042, B => 
                           n24041, ZN => n26084);
   U25418 : XNOR2_X1 port map( A => n26084, B => n25943, ZN => n25569);
   U25419 : NAND2_X1 port map( A1 => n24758, A2 => n29592, ZN => n24449);
   U25420 : INV_X1 port map( A => n24449, ZN => n24045);
   U25421 : OAI21_X1 port map( B1 => n29592, B2 => n24756, A => n23588, ZN => 
                           n24044);
   U25422 : NAND2_X1 port map( A1 => n24479, A2 => n24483, ZN => n24048);
   U25424 : OAI21_X2 port map( B1 => n24050, B2 => n24479, A => n24049, ZN => 
                           n25454);
   U25425 : XNOR2_X1 port map( A => n25454, B => n26053, ZN => n24051);
   U25426 : XNOR2_X1 port map( A => n25569, B => n24051, ZN => n24063);
   U25427 : NOR2_X1 port map( A1 => n24584, A2 => n24582, ZN => n24053);
   U25428 : NOR2_X1 port map( A1 => n24583, A2 => n29025, ZN => n24052);
   U25429 : NAND2_X1 port map( A1 => n24577, A2 => n24584, ZN => n24466);
   U25431 : MUX2_X1 port map( A => n24057, B => n23922, S => n24610, Z => 
                           n24058);
   U25433 : XNOR2_X1 port map( A => n25722, B => n24061, ZN => n24062);
   U25435 : NOR2_X1 port map( A1 => n25006, A2 => n25005, ZN => n24366);
   U25436 : NOR2_X1 port map( A1 => n24366, A2 => n24304, ZN => n24066);
   U25437 : OAI21_X1 port map( B1 => n23897, B2 => n24066, A => n24065, ZN => 
                           n26019);
   U25438 : XNOR2_X1 port map( A => n26019, B => n25190, ZN => n24070);
   U25439 : XNOR2_X1 port map( A => n25910, B => n25809, ZN => n25590);
   U25440 : XNOR2_X1 port map( A => n25590, B => n24070, ZN => n24089);
   U25441 : NOR2_X1 port map( A1 => n24666, A2 => n24072, ZN => n24071);
   U25442 : INV_X1 port map( A => n24074, ZN => n24669);
   U25443 : AOI22_X1 port map( A1 => n28424, A2 => n24075, B1 => n24383, B2 => 
                           n24669, ZN => n24076);
   U25444 : AOI21_X1 port map( B1 => n24077, B2 => n24388, A => n24079, ZN => 
                           n24082);
   U25445 : XNOR2_X1 port map( A => n25398, B => n25251, ZN => n25743);
   U25446 : OAI21_X1 port map( B1 => n24403, B2 => n24408, A => n24084, ZN => 
                           n24086);
   U25447 : INV_X1 port map( A => n2961, ZN => n27333);
   U25448 : XNOR2_X1 port map( A => n29039, B => n27333, ZN => n24087);
   U25449 : XNOR2_X1 port map( A => n24087, B => n25743, ZN => n24088);
   U25450 : INV_X1 port map( A => n24090, ZN => n24098);
   U25451 : INV_X1 port map( A => n24093, ZN => n24094);
   U25452 : XNOR2_X1 port map( A => n25037, B => n25509, ZN => n24110);
   U25453 : INV_X1 port map( A => n24712, ZN => n24104);
   U25454 : AOI21_X1 port map( B1 => n24720, B2 => n24711, A => n24104, ZN => 
                           n24108);
   U25455 : AOI21_X1 port map( B1 => n4136, B2 => n24412, A => n24712, ZN => 
                           n24107);
   U25456 : NOR2_X1 port map( A1 => n24716, A2 => n4136, ZN => n24105);
   U25457 : XNOR2_X1 port map( A => n25385, B => n2960, ZN => n24109);
   U25458 : XNOR2_X1 port map( A => n24110, B => n24109, ZN => n24131);
   U25459 : NOR2_X1 port map( A1 => n24520, A2 => n24516, ZN => n24112);
   U25460 : NOR2_X1 port map( A1 => n24111, A2 => n24517, ZN => n24180);
   U25461 : MUX2_X1 port map( A => n24112, B => n24180, S => n24514, Z => 
                           n24116);
   U25462 : OAI21_X1 port map( B1 => n24420, B2 => n24113, A => n24516, ZN => 
                           n24114);
   U25463 : NOR2_X1 port map( A1 => n24180, A2 => n24114, ZN => n24115);
   U25464 : XNOR2_X1 port map( A => n28402, B => n25751, ZN => n24129);
   U25465 : NAND2_X1 port map( A1 => n24347, A2 => n24433, ZN => n24119);
   U25466 : INV_X1 port map( A => n24434, ZN => n24117);
   U25467 : NAND2_X1 port map( A1 => n24338, A2 => n29043, ZN => n24123);
   U25468 : NAND3_X1 port map( A1 => n24707, A2 => n24417, A3 => n5571, ZN => 
                           n24126);
   U25469 : XNOR2_X1 port map( A => n25513, B => n26110, ZN => n25387);
   U25470 : XNOR2_X1 port map( A => n25387, B => n24129, ZN => n24130);
   U25471 : XNOR2_X1 port map( A => n24130, B => n24131, ZN => n25317);
   U25472 : INV_X1 port map( A => n25317, ZN => n26181);
   U25473 : NOR2_X1 port map( A1 => n811, A2 => n29470, ZN => n24136);
   U25474 : XNOR2_X1 port map( A => n25563, B => n24137, ZN => n24152);
   U25475 : NOR2_X1 port map( A1 => n24367, A2 => n24369, ZN => n25009);
   U25476 : AOI211_X1 port map( C1 => n24369, C2 => n24368, A => n28415, B => 
                           n24138, ZN => n24140);
   U25477 : NAND2_X1 port map( A1 => n24278, A2 => n24141, ZN => n24588);
   U25478 : INV_X1 port map( A => n24142, ZN => n24146);
   U25479 : NOR2_X1 port map( A1 => n22356, A2 => n24735, ZN => n24740);
   U25480 : OAI211_X1 port map( C1 => n29050, C2 => n24280, A => n24736, B => 
                           n24601, ZN => n24150);
   U25481 : XNOR2_X1 port map( A => n25735, B => n26007, ZN => n24151);
   U25482 : XNOR2_X1 port map( A => n24151, B => n24152, ZN => n25666);
   U25483 : INV_X1 port map( A => n25666, ZN => n26180);
   U25484 : NAND3_X1 port map( A1 => n26181, A2 => n26180, A3 => n28561, ZN => 
                           n24202);
   U25485 : NOR2_X1 port map( A1 => n26186, A2 => n29528, ZN => n24171);
   U25486 : INV_X1 port map( A => n24256, ZN => n24508);
   U25487 : MUX2_X1 port map( A => n24651, B => n28785, S => n24653, Z => 
                           n24156);
   U25488 : INV_X1 port map( A => n24248, ZN => n24526);
   U25489 : OAI21_X1 port map( B1 => n24526, B2 => n28785, A => n24249, ZN => 
                           n24649);
   U25490 : MUX2_X1 port map( A => n24794, B => n24789, S => n28455, Z => 
                           n24158);
   U25491 : MUX2_X1 port map( A => n24793, B => n24791, S => n1955, Z => n24157
                           );
   U25492 : XNOR2_X1 port map( A => n25901, B => n26041, ZN => n25015);
   U25493 : XNOR2_X1 port map( A => n25903, B => n25727, ZN => n24168);
   U25497 : NOR2_X1 port map( A1 => n29120, A2 => n24162, ZN => n24163);
   U25498 : NAND2_X1 port map( A1 => n24163, A2 => n6600, ZN => n24164);
   U25499 : XNOR2_X1 port map( A => n26039, B => n24166, ZN => n24167);
   U25500 : XNOR2_X1 port map( A => n24167, B => n24168, ZN => n24169);
   U25501 : NAND2_X1 port map( A1 => n24171, A2 => n28547, ZN => n24201);
   U25502 : NOR2_X1 port map( A1 => n28519, A2 => n24552, ZN => n24554);
   U25503 : AOI21_X1 port map( B1 => n24174, B2 => n24173, A => n24554, ZN => 
                           n24177);
   U25504 : OAI22_X1 port map( A1 => n24175, A2 => n24178, B1 => n24556, B2 => 
                           n24553, ZN => n24176);
   U25506 : NAND2_X1 port map( A1 => n24179, A2 => n24514, ZN => n24185);
   U25507 : NOR2_X1 port map( A1 => n24179, A2 => n24420, ZN => n24181);
   U25508 : AOI21_X1 port map( B1 => n24181, B2 => n24520, A => n24180, ZN => 
                           n24184);
   U25509 : AND2_X1 port map( A1 => n24516, A2 => n24514, ZN => n24182);
   U25510 : NAND2_X1 port map( A1 => n24520, A2 => n24182, ZN => n24183);
   U25511 : OAI211_X1 port map( C1 => n24520, C2 => n24185, A => n24184, B => 
                           n24183, ZN => n25932);
   U25512 : XNOR2_X1 port map( A => n25932, B => n28520, ZN => n24187);
   U25513 : XNOR2_X1 port map( A => n25931, B => n2274, ZN => n24186);
   U25514 : XNOR2_X1 port map( A => n24187, B => n24186, ZN => n24199);
   U25515 : MUX2_X1 port map( A => n24436, B => n24437, S => n24347, Z => 
                           n24191);
   U25516 : OAI21_X1 port map( B1 => n403, B2 => n29726, A => n24188, ZN => 
                           n24190);
   U25518 : NAND2_X1 port map( A1 => n2619, A2 => n24434, ZN => n24189);
   U25519 : XNOR2_X1 port map( A => n25179, B => n25440, ZN => n25763);
   U25520 : INV_X1 port map( A => n24241, ZN => n24242);
   U25521 : MUX2_X1 port map( A => n24557, B => n24192, S => n24633, Z => 
                           n24193);
   U25522 : OAI21_X2 port map( B1 => n24194, B2 => n25794, A => n24193, ZN => 
                           n25702);
   U25523 : XNOR2_X1 port map( A => n26102, B => n25702, ZN => n26015);
   U25524 : XNOR2_X1 port map( A => n25763, B => n26015, ZN => n24198);
   U25525 : OAI21_X1 port map( B1 => n24204, B2 => n26181, A => n24203, ZN => 
                           n27032);
   U25526 : INV_X1 port map( A => n24205, ZN => n24460);
   U25528 : NOR2_X1 port map( A1 => n24816, A2 => n24817, ZN => n24206);
   U25529 : AOI21_X2 port map( B1 => n24207, B2 => n24208, A => n24206, ZN => 
                           n26046);
   U25530 : XNOR2_X1 port map( A => n26046, B => n25107, ZN => n25429);
   U25531 : INV_X1 port map( A => n24776, ZN => n24457);
   U25532 : XNOR2_X1 port map( A => n25429, B => n25081, ZN => n24226);
   U25533 : XNOR2_X1 port map( A => n26044, B => n25727, ZN => n24224);
   U25534 : NOR2_X1 port map( A1 => n24758, A2 => n24216, ZN => n24222);
   U25535 : NOR2_X1 port map( A1 => n24222, A2 => n24221, ZN => n25498);
   U25536 : XNOR2_X1 port map( A => n25498, B => n3211, ZN => n24223);
   U25537 : XNOR2_X1 port map( A => n24224, B => n24223, ZN => n24225);
   U25538 : XNOR2_X2 port map( A => n24226, B => n24225, ZN => n27395);
   U25539 : INV_X1 port map( A => n27395, ZN => n26195);
   U25540 : OAI21_X1 port map( B1 => n24630, B2 => n24293, A => n24295, ZN => 
                           n24228);
   U25542 : XNOR2_X1 port map( A => n26023, B => n25134, ZN => n25806);
   U25543 : XNOR2_X1 port map( A => n28628, B => n25396, ZN => n24230);
   U25544 : XNOR2_X1 port map( A => n25806, B => n24230, ZN => n24255);
   U25545 : NAND2_X1 port map( A1 => n24231, A2 => n24642, ZN => n24235);
   U25546 : INV_X1 port map( A => n24638, ZN => n24564);
   U25547 : OAI21_X1 port map( B1 => n24232, B2 => n24564, A => n24643, ZN => 
                           n24233);
   U25548 : NAND2_X1 port map( A1 => n24233, A2 => n29645, ZN => n24234);
   U25550 : OAI21_X1 port map( B1 => n24633, B2 => n465, A => n24634, ZN => 
                           n24238);
   U25552 : XNOR2_X1 port map( A => n25065, B => n25745, ZN => n25449);
   U25553 : NAND2_X1 port map( A1 => n24247, A2 => n28481, ZN => n24252);
   U25554 : NAND2_X1 port map( A1 => n24249, A2 => n24248, ZN => n24250);
   U25555 : INV_X1 port map( A => n24653, ZN => n24655);
   U25556 : NAND2_X1 port map( A1 => n24250, A2 => n24655, ZN => n24251);
   U25557 : NAND2_X1 port map( A1 => n24252, A2 => n24251, ZN => n24963);
   U25558 : XNOR2_X1 port map( A => n26120, B => n26701, ZN => n24253);
   U25559 : XNOR2_X1 port map( A => n25449, B => n24253, ZN => n24254);
   U25560 : XNOR2_X1 port map( A => n25346, B => n25059, ZN => n25772);
   U25561 : XNOR2_X1 port map( A => n25773, B => n300, ZN => n24264);
   U25562 : XNOR2_X1 port map( A => n25772, B => n24264, ZN => n24276);
   U25563 : NAND3_X1 port map( A1 => n24748, A2 => n24751, A3 => n24747, ZN => 
                           n24267);
   U25564 : OAI211_X1 port map( C1 => n28550, C2 => n24747, A => n24267, B => 
                           n24266, ZN => n25736);
   U25565 : XNOR2_X1 port map( A => n25738, B => n29017, ZN => n24274);
   U25566 : INV_X1 port map( A => n24791, ZN => n24268);
   U25567 : OAI211_X1 port map( C1 => n24792, C2 => n24268, A => n24793, B => 
                           n24789, ZN => n24271);
   U25568 : NAND3_X1 port map( A1 => n28512, A2 => n24269, A3 => n4576, ZN => 
                           n24270);
   U25569 : NAND3_X1 port map( A1 => n24271, A2 => n24270, A3 => n6943, ZN => 
                           n24272);
   U25570 : XNOR2_X1 port map( A => n26095, B => n6653, ZN => n24273);
   U25571 : XNOR2_X1 port map( A => n24274, B => n24273, ZN => n24275);
   U25572 : XNOR2_X1 port map( A => n24276, B => n24275, ZN => n26464);
   U25573 : NOR2_X1 port map( A1 => n24593, A2 => n24278, ZN => n24589);
   U25574 : XNOR2_X1 port map( A => n26011, B => n25820, ZN => n25277);
   U25575 : NAND2_X1 port map( A1 => n24282, A2 => n24280, ZN => n24284);
   U25576 : NAND2_X1 port map( A1 => n22311, A2 => n24602, ZN => n24600);
   U25577 : NAND3_X1 port map( A1 => n24282, A2 => n24736, A3 => n24734, ZN => 
                           n24283);
   U25578 : OAI211_X1 port map( C1 => n22356, C2 => n24284, A => n24600, B => 
                           n24283, ZN => n24286);
   U25580 : XNOR2_X1 port map( A => n25381, B => n25341, ZN => n24287);
   U25581 : XNOR2_X1 port map( A => n24287, B => n25277, ZN => n24302);
   U25582 : AOI22_X1 port map( A1 => n24596, A2 => n24728, B1 => n24730, B2 => 
                           n24729, ZN => n24292);
   U25583 : INV_X1 port map( A => n24598, ZN => n24289);
   U25585 : NAND2_X1 port map( A1 => n4364, A2 => n24295, ZN => n24296);
   U25586 : XNOR2_X1 port map( A => n25760, B => n25890, ZN => n24300);
   U25587 : XNOR2_X1 port map( A => n25179, B => n3423, ZN => n24299);
   U25588 : XNOR2_X1 port map( A => n24300, B => n24299, ZN => n24301);
   U25590 : XNOR2_X1 port map( A => n24306, B => n25782, ZN => n24308);
   U25591 : XNOR2_X1 port map( A => n24308, B => n24307, ZN => n24329);
   U25593 : NAND2_X1 port map( A1 => n29567, A2 => n24310, ZN => n24312);
   U25596 : NOR2_X1 port map( A1 => n24668, A2 => n24383, ZN => n24317);
   U25598 : INV_X1 port map( A => n24383, ZN => n24318);
   U25599 : NAND3_X1 port map( A1 => n24667, A2 => n24669, A3 => n24318, ZN => 
                           n24319);
   U25600 : XNOR2_X1 port map( A => n25386, B => n25780, ZN => n24328);
   U25601 : NOR3_X1 port map( A1 => n29555, A2 => n24677, A3 => n24676, ZN => 
                           n24325);
   U25602 : NOR2_X2 port map( A1 => n24326, A2 => n24325, ZN => n26108);
   U25603 : INV_X1 port map( A => n26108, ZN => n24327);
   U25604 : XNOR2_X1 port map( A => n24328, B => n24327, ZN => n25040);
   U25605 : XNOR2_X1 port map( A => n24329, B => n25040, ZN => n26194);
   U25606 : INV_X1 port map( A => n26194, ZN => n25404);
   U25608 : INV_X1 port map( A => n25375, ZN => n24330);
   U25609 : INV_X1 port map( A => n24772, ZN => n24331);
   U25610 : NOR2_X1 port map( A1 => n24697, A2 => n29624, ZN => n24332);
   U25611 : AOI22_X1 port map( A1 => n24699, A2 => n24768, B1 => n24765, B2 => 
                           n24332, ZN => n24333);
   U25612 : INV_X1 port map( A => n24334, ZN => n24335);
   U25613 : NOR3_X1 port map( A1 => n24337, A2 => n24336, A3 => n24335, ZN => 
                           n24340);
   U25614 : NAND3_X1 port map( A1 => n24341, A2 => n24417, A3 => n29043, ZN => 
                           n24343);
   U25617 : XNOR2_X1 port map( A => n25458, B => n24345, ZN => n24360);
   U25620 : AND3_X2 port map( A1 => n24349, A2 => n24348, A3 => n6945, ZN => 
                           n25535);
   U25621 : XNOR2_X1 port map( A => n24949, B => n25535, ZN => n24358);
   U25622 : NOR2_X1 port map( A1 => n24714, A2 => n24713, ZN => n24350);
   U25623 : MUX2_X1 port map( A => n24351, B => n24350, S => n24712, Z => 
                           n24355);
   U25624 : XNOR2_X1 port map( A => n25149, B => n24356, ZN => n24357);
   U25625 : XNOR2_X1 port map( A => n24358, B => n24357, ZN => n24359);
   U25627 : OAI21_X1 port map( B1 => n25404, B2 => n26469, A => n27394, ZN => 
                           n24361);
   U25628 : OAI211_X1 port map( C1 => n26195, C2 => n25406, A => n24362, B => 
                           n24361, ZN => n27026);
   U25629 : NAND2_X1 port map( A1 => n27032, A2 => n27026, ZN => n24363);
   U25630 : NAND2_X1 port map( A1 => n26705, A2 => n26819, ZN => n24828);
   U25631 : INV_X1 port map( A => n27026, ZN => n26817);
   U25632 : NOR2_X1 port map( A1 => n24366, A2 => n24365, ZN => n24371);
   U25633 : MUX2_X1 port map( A => n25005, B => n24368, S => n24367, Z => 
                           n24370);
   U25635 : NOR2_X1 port map( A1 => n29340, A2 => n24374, ZN => n24379);
   U25636 : XNOR2_X1 port map( A => n25352, B => n25430, ZN => n24389);
   U25637 : MUX2_X1 port map( A => n24667, B => n4605, S => n24669, Z => n24385
                           );
   U25639 : XNOR2_X1 port map( A => n24389, B => n25541, ZN => n24402);
   U25640 : MUX2_X1 port map( A => n466, B => n29471, S => n24390, Z => n24394)
                           ;
   U25641 : INV_X1 port map( A => n24682, ZN => n24392);
   U25642 : INV_X1 port map( A => n24688, ZN => n24681);
   U25644 : OAI21_X1 port map( B1 => n24397, B2 => n24678, A => n24396, ZN => 
                           n24398);
   U25645 : XNOR2_X1 port map( A => n25689, B => n25900, ZN => n25354);
   U25646 : XNOR2_X1 port map( A => n26045, B => n3109, ZN => n24400);
   U25647 : XNOR2_X1 port map( A => n25354, B => n24400, ZN => n24401);
   U25648 : OR2_X1 port map( A1 => n24405, A2 => n24404, ZN => n24406);
   U25649 : NAND2_X1 port map( A1 => n24720, A2 => n24713, ZN => n24414);
   U25651 : XNOR2_X1 port map( A => n25550, B => n25345, ZN => n26091);
   U25652 : NAND2_X1 port map( A1 => n24416, A2 => n24415, ZN => n24419);
   U25653 : AND2_X1 port map( A1 => n24420, A2 => n24514, ZN => n24423);
   U25654 : XNOR2_X1 port map( A => n25737, B => n25864, ZN => n24425);
   U25655 : XNOR2_X1 port map( A => n26091, B => n24425, ZN => n24446);
   U25656 : XNOR2_X1 port map( A => n25867, B => n25708, ZN => n24444);
   U25657 : NOR2_X1 port map( A1 => n24434, A2 => n24433, ZN => n24441);
   U25658 : OR2_X1 port map( A1 => n24435, A2 => n29726, ZN => n24440);
   U25659 : NAND3_X1 port map( A1 => n29726, A2 => n24437, A3 => n29128, ZN => 
                           n24439);
   U25660 : XNOR2_X1 port map( A => n25564, B => n26825, ZN => n24443);
   U25661 : XNOR2_X1 port map( A => n24444, B => n24443, ZN => n24445);
   U25662 : XNOR2_X1 port map( A => n24446, B => n24445, ZN => n26559);
   U25663 : NOR2_X1 port map( A1 => n28385, A2 => n26559, ZN => n24576);
   U25664 : NAND2_X1 port map( A1 => n24449, A2 => n24448, ZN => n24452);
   U25665 : AOI21_X1 port map( B1 => n24757, B2 => n24756, A => n24450, ZN => 
                           n24451);
   U25666 : AOI22_X1 port map( A1 => n24452, A2 => n24451, B1 => n24758, B2 => 
                           n24757, ZN => n25182);
   U25667 : XNOR2_X1 port map( A => n24453, B => n25441, ZN => n24465);
   U25668 : NAND2_X1 port map( A1 => n24780, A2 => n24776, ZN => n24455);
   U25669 : NAND2_X1 port map( A1 => n1426, A2 => n24779, ZN => n24459);
   U25670 : AND3_X1 port map( A1 => n24457, A2 => n24775, A3 => n24779, ZN => 
                           n24458);
   U25671 : NAND2_X1 port map( A1 => n24812, A2 => n24460, ZN => n24464);
   U25672 : NOR2_X1 port map( A1 => n24812, A2 => n24814, ZN => n24498);
   U25673 : OAI21_X1 port map( B1 => n24498, B2 => n24808, A => n24817, ZN => 
                           n24463);
   U25675 : XNOR2_X1 port map( A => n25889, B => n29155, ZN => n25340);
   U25676 : XNOR2_X1 port map( A => n24465, B => n25340, ZN => n24488);
   U25677 : NAND2_X1 port map( A1 => n24583, A2 => n24467, ZN => n24469);
   U25678 : NAND3_X1 port map( A1 => n24471, A2 => n24470, A3 => n24491, ZN => 
                           n24478);
   U25679 : AOI22_X1 port map( A1 => n24473, A2 => n23842, B1 => n24474, B2 => 
                           n24489, ZN => n24477);
   U25680 : NAND2_X1 port map( A1 => n24475, A2 => n24474, ZN => n24476);
   U25681 : NOR2_X1 port map( A1 => n24479, A2 => n24483, ZN => n24481);
   U25683 : XNOR2_X1 port map( A => n24487, B => n26100, ZN => n25529);
   U25684 : AOI21_X1 port map( B1 => n24493, B2 => n24492, A => n24491, ZN => 
                           n24494);
   U25685 : INV_X1 port map( A => n24808, ZN => n24497);
   U25686 : NAND2_X1 port map( A1 => n24498, A2 => n220, ZN => n24501);
   U25687 : NOR2_X1 port map( A1 => n24503, A2 => n24801, ZN => n24504);
   U25688 : NOR2_X1 port map( A1 => n24504, A2 => n24802, ZN => n24505);
   U25689 : XNOR2_X1 port map( A => n25844, B => n25914, ZN => n25330);
   U25690 : AOI21_X1 port map( B1 => n24972, B2 => n24509, A => n24508, ZN => 
                           n24510);
   U25691 : NOR2_X1 port map( A1 => n23467, A2 => n24510, ZN => n24511);
   U25692 : NOR2_X2 port map( A1 => n24512, A2 => n24511, ZN => n26115);
   U25693 : OAI21_X1 port map( B1 => n24518, B2 => n24517, A => n24516, ZN => 
                           n24519);
   U25694 : XNOR2_X1 port map( A => n26115, B => n25909, ZN => n24521);
   U25695 : XNOR2_X1 port map( A => n25330, B => n24521, ZN => n24522);
   U25696 : OAI21_X1 port map( B1 => n24523, B2 => n3061, A => n24653, ZN => 
                           n24525);
   U25697 : NOR2_X1 port map( A1 => n3061, A2 => n28785, ZN => n24527);
   U25698 : NAND2_X1 port map( A1 => n24527, A2 => n24526, ZN => n24528);
   U25699 : XNOR2_X1 port map( A => n24529, B => n26055, ZN => n24549);
   U25700 : NOR2_X1 port map( A1 => n23144, A2 => n24631, ZN => n24893);
   U25701 : NAND2_X1 port map( A1 => n4366, A2 => n24533, ZN => n24628);
   U25702 : INV_X1 port map( A => n24628, ZN => n24534);
   U25703 : NAND2_X1 port map( A1 => n24534, A2 => n24631, ZN => n24535);
   U25705 : AOI21_X1 port map( B1 => n24542, B2 => n24541, A => n23126, ZN => 
                           n24546);
   U25707 : XNOR2_X1 port map( A => n26080, B => n29606, ZN => n25287);
   U25708 : XNOR2_X1 port map( A => n24549, B => n25287, ZN => n24574);
   U25710 : NOR2_X1 port map( A1 => n24559, A2 => n24633, ZN => n24636);
   U25711 : AOI22_X1 port map( A1 => n24561, A2 => n24560, B1 => n24636, B2 => 
                           n465, ZN => n24562);
   U25712 : NOR2_X1 port map( A1 => n24644, A2 => n24564, ZN => n24566);
   U25713 : NOR2_X1 port map( A1 => n24644, A2 => n24638, ZN => n24565);
   U25714 : AOI22_X1 port map( A1 => n24566, A2 => n24642, B1 => n24565, B2 => 
                           n29643, ZN => n24570);
   U25715 : NOR2_X1 port map( A1 => n29643, A2 => n24643, ZN => n24567);
   U25716 : NAND2_X1 port map( A1 => n24568, A2 => n24567, ZN => n24569);
   U25718 : XNOR2_X1 port map( A => n25696, B => n25947, ZN => n24572);
   U25719 : XNOR2_X1 port map( A => n26083, B => n24572, ZN => n24573);
   U25720 : NOR2_X1 port map( A1 => n24578, A2 => n29026, ZN => n24580);
   U25721 : NOR2_X1 port map( A1 => n24583, A2 => n24582, ZN => n24585);
   U25722 : OAI21_X1 port map( B1 => n24586, B2 => n24585, A => n24584, ZN => 
                           n24587);
   U25725 : OAI21_X1 port map( B1 => n24601, B2 => n24602, A => n24744, ZN => 
                           n24606);
   U25726 : AOI22_X1 port map( A1 => n22356, A2 => n24604, B1 => n24603, B2 => 
                           n24602, ZN => n24605);
   U25728 : XNOR2_X1 port map( A => n24608, B => n29518, ZN => n24625);
   U25729 : NOR3_X1 port map( A1 => n459, A2 => n24609, A3 => n5168, ZN => 
                           n24615);
   U25730 : MUX2_X1 port map( A => n24610, B => n29109, S => n24614, Z => 
                           n24611);
   U25731 : AOI21_X1 port map( B1 => n21303, B2 => n2879, A => n24616, ZN => 
                           n24623);
   U25732 : NOR2_X1 port map( A1 => n24618, A2 => n24747, ZN => n24619);
   U25733 : NOR2_X1 port map( A1 => n24620, A2 => n24619, ZN => n24621);
   U25734 : OAI21_X1 port map( B1 => n24623, B2 => n28223, A => n24621, ZN => 
                           n25165);
   U25736 : NOR2_X1 port map( A1 => n26457, A2 => n28578, ZN => n26563);
   U25737 : NAND2_X1 port map( A1 => n26563, A2 => n28385, ZN => n24627);
   U25738 : NOR2_X1 port map( A1 => n26458, A2 => n28578, ZN => n25614);
   U25739 : NAND2_X1 port map( A1 => n25614, A2 => n26559, ZN => n24626);
   U25740 : OAI21_X1 port map( B1 => n24630, B2 => n24629, A => n24628, ZN => 
                           n24632);
   U25741 : INV_X1 port map( A => n29645, ZN => n24640);
   U25742 : OAI22_X1 port map( A1 => n24641, A2 => n24640, B1 => n24639, B2 => 
                           n24638, ZN => n24648);
   U25743 : MUX2_X1 port map( A => n24644, B => n24643, S => n24642, Z => 
                           n24646);
   U25744 : NOR2_X1 port map( A1 => n24646, A2 => n29642, ZN => n24647);
   U25745 : XNOR2_X1 port map( A => n29069, B => n25542, ZN => n25294);
   U25746 : XNOR2_X1 port map( A => n25294, B => n25207, ZN => n24664);
   U25747 : NAND3_X1 port map( A1 => n24649, A2 => n3697, A3 => n3061, ZN => 
                           n24659);
   U25748 : XNOR2_X1 port map( A => n28785, B => n629, ZN => n24654);
   U25749 : NOR2_X1 port map( A1 => n24653, A2 => n3697, ZN => n24652);
   U25750 : AOI22_X1 port map( A1 => n24654, A2 => n24653, B1 => n24652, B2 => 
                           n28481, ZN => n24657);
   U25751 : NAND3_X1 port map( A1 => n24660, A2 => n24659, A3 => n24658, ZN => 
                           n24661);
   U25752 : XNOR2_X1 port map( A => n25352, B => n24661, ZN => n24662);
   U25753 : XNOR2_X1 port map( A => n28576, B => n24662, ZN => n24663);
   U25754 : XNOR2_X2 port map( A => n24664, B => n24663, ZN => n26927);
   U25755 : XNOR2_X1 port map( A => n25215, B => n24671, ZN => n24696);
   U25756 : XNOR2_X1 port map( A => n25345, B => n29534, ZN => n24694);
   U25757 : OAI211_X1 port map( C1 => n24678, C2 => n404, A => n24677, B => 
                           n24676, ZN => n24679);
   U25758 : NAND2_X1 port map( A1 => n24680, A2 => n24679, ZN => n25562);
   U25759 : AOI21_X1 port map( B1 => n24683, B2 => n24682, A => n24681, ZN => 
                           n24693);
   U25760 : NAND4_X1 port map( A1 => n24687, A2 => n24686, A3 => n24685, A4 => 
                           n24684, ZN => n24690);
   U25761 : AOI21_X1 port map( B1 => n24690, B2 => n29471, A => n24688, ZN => 
                           n24692);
   U25762 : OAI21_X1 port map( B1 => n24693, B2 => n24692, A => n24691, ZN => 
                           n25549);
   U25763 : XNOR2_X1 port map( A => n25562, B => n25549, ZN => n25304);
   U25764 : XNOR2_X1 port map( A => n25304, B => n24694, ZN => n24695);
   U25767 : AND2_X1 port map( A1 => n24765, A2 => n24768, ZN => n24701);
   U25768 : XNOR2_X1 port map( A => n25927, B => n25884, ZN => n25298);
   U25769 : XNOR2_X1 port map( A => n25298, B => n24703, ZN => n24723);
   U25770 : MUX2_X1 port map( A => n24712, B => n24714, S => n24711, Z => 
                           n24721);
   U25771 : NAND3_X1 port map( A1 => n24715, A2 => n24714, A3 => n24713, ZN => 
                           n24719);
   U25772 : NAND2_X1 port map( A1 => n28416, A2 => n24716, ZN => n24718);
   U25773 : OAI211_X2 port map( C1 => n24721, C2 => n24720, A => n24719, B => 
                           n24718, ZN => n25885);
   U25774 : XNOR2_X1 port map( A => n25932, B => n25885, ZN => n25486);
   U25775 : XNOR2_X1 port map( A => n25486, B => n25113, ZN => n24722);
   U25776 : XNOR2_X2 port map( A => n24722, B => n24723, ZN => n26933);
   U25777 : NOR2_X1 port map( A1 => n24726, A2 => n24725, ZN => n24727);
   U25778 : NAND2_X1 port map( A1 => n24729, A2 => n24728, ZN => n24731);
   U25779 : AOI21_X1 port map( B1 => n24732, B2 => n24731, A => n24730, ZN => 
                           n24733);
   U25780 : NAND2_X1 port map( A1 => n24740, A2 => n24739, ZN => n24741);
   U25782 : XNOR2_X1 port map( A => n25531, B => n29563, ZN => n25288);
   U25783 : OAI21_X1 port map( B1 => n28550, B2 => n24748, A => n24747, ZN => 
                           n24750);
   U25784 : XNOR2_X1 port map( A => n25288, B => n25479, ZN => n24755);
   U25785 : XNOR2_X1 port map( A => n28630, B => n1187, ZN => n24752);
   U25786 : XNOR2_X1 port map( A => n24753, B => n24752, ZN => n24754);
   U25787 : XNOR2_X1 port map( A => n24755, B => n24754, ZN => n26579);
   U25788 : NAND3_X1 port map( A1 => n26927, A2 => n24788, A3 => n5505, ZN => 
                           n24825);
   U25789 : XNOR2_X1 port map( A => n26115, B => n29614, ZN => n24764);
   U25790 : NAND2_X1 port map( A1 => n24761, A2 => n24760, ZN => n24762);
   U25791 : XNOR2_X1 port map( A => n25251, B => n25810, ZN => n25089);
   U25792 : XNOR2_X1 port map( A => n24764, B => n25089, ZN => n24787);
   U25793 : OAI21_X1 port map( B1 => n24765, B2 => n1856, A => n29624, ZN => 
                           n24766);
   U25794 : OAI21_X1 port map( B1 => n24772, B2 => n24771, A => n24770, ZN => 
                           n24773);
   U25795 : XNOR2_X1 port map( A => n29047, B => n25845, ZN => n24785);
   U25796 : NOR2_X1 port map( A1 => n24777, A2 => n24776, ZN => n24778);
   U25797 : OAI21_X1 port map( B1 => n24778, B2 => n23946, A => n463, ZN => 
                           n24782);
   U25798 : XNOR2_X1 port map( A => n24785, B => n24784, ZN => n24786);
   U25799 : XNOR2_X1 port map( A => n24787, B => n24786, ZN => n25364);
   U25800 : INV_X1 port map( A => n25364, ZN => n26926);
   U25802 : NAND2_X1 port map( A1 => n26929, A2 => n24788, ZN => n24824);
   U25803 : XNOR2_X1 port map( A => n25282, B => n27730, ZN => n24798);
   U25804 : OAI21_X1 port map( B1 => n1955, B2 => n24791, A => n28512, ZN => 
                           n24796);
   U25805 : OAI21_X1 port map( B1 => n24794, B2 => n24793, A => n24792, ZN => 
                           n24795);
   U25806 : XNOR2_X1 port map( A => n24797, B => n25463, ZN => n25753);
   U25807 : XNOR2_X1 port map( A => n24798, B => n25753, ZN => n24822);
   U25808 : OAI21_X1 port map( B1 => n24801, B2 => n24800, A => n28919, ZN => 
                           n24807);
   U25809 : MUX2_X1 port map( A => n24809, B => n24817, S => n24808, Z => 
                           n24811);
   U25810 : XNOR2_X1 port map( A => n25322, B => n25509, ZN => n25153);
   U25811 : XNOR2_X1 port map( A => n24923, B => n25153, ZN => n24821);
   U25812 : XNOR2_X1 port map( A => n24821, B => n24822, ZN => n26581);
   U25813 : XNOR2_X1 port map( A => n24829, B => n622, ZN => Ciphertext(31));
   U25814 : XNOR2_X1 port map( A => n25366, B => n26045, ZN => n25080);
   U25815 : XNOR2_X1 port map( A => n25803, B => n25080, ZN => n24833);
   U25816 : XNOR2_X1 port map( A => n25901, B => n25836, ZN => n24831);
   U25817 : XNOR2_X1 port map( A => n26039, B => n3751, ZN => n24830);
   U25818 : XNOR2_X1 port map( A => n24831, B => n24830, ZN => n24832);
   U25819 : XNOR2_X1 port map( A => n24833, B => n24832, ZN => n26425);
   U25820 : XNOR2_X1 port map( A => n24834, B => n25590, ZN => n24837);
   U25821 : XNOR2_X1 port map( A => n29047, B => n3695, ZN => n24835);
   U25822 : XNOR2_X1 port map( A => n25069, B => n24835, ZN => n24836);
   U25823 : XNOR2_X1 port map( A => n24837, B => n24836, ZN => n26382);
   U25824 : INV_X1 port map( A => n26382, ZN => n26361);
   U25825 : XNOR2_X1 port map( A => n25569, B => n24948, ZN => n24841);
   U25826 : XNOR2_X1 port map( A => n25826, B => n29613, ZN => n24839);
   U25827 : XNOR2_X1 port map( A => n26055, B => n3752, ZN => n24838);
   U25828 : XNOR2_X1 port map( A => n24839, B => n24838, ZN => n24840);
   U25829 : XNOR2_X1 port map( A => n25708, B => n25346, ZN => n26006);
   U25830 : XNOR2_X1 port map( A => n25391, B => n25869, ZN => n24938);
   U25831 : XNOR2_X1 port map( A => n24938, B => n26006, ZN => n24845);
   U25832 : XNOR2_X1 port map( A => n26093, B => n25775, ZN => n24843);
   U25833 : XNOR2_X1 port map( A => n25921, B => n3378, ZN => n24842);
   U25834 : XNOR2_X1 port map( A => n24843, B => n24842, ZN => n24844);
   U25835 : XNOR2_X1 port map( A => n24845, B => n24844, ZN => n26378);
   U25836 : NOR2_X1 port map( A1 => n26426, A2 => n26378, ZN => n24846);
   U25837 : XNOR2_X1 port map( A => n25037, B => n25785, ZN => n24913);
   U25838 : XNOR2_X1 port map( A => n24913, B => n25056, ZN => n24850);
   U25839 : XNOR2_X1 port map( A => n24847, B => n25385, ZN => n24848);
   U25840 : XNOR2_X1 port map( A => n26110, B => n25324, ZN => n26034);
   U25841 : XNOR2_X1 port map( A => n26034, B => n24848, ZN => n24849);
   U25842 : XNOR2_X1 port map( A => n24850, B => n24849, ZN => n26431);
   U25843 : XNOR2_X1 port map( A => n26011, B => n25885, ZN => n24851);
   U25844 : XNOR2_X1 port map( A => n26102, B => n25444, ZN => n25821);
   U25845 : XNOR2_X1 port map( A => n25821, B => n24851, ZN => n24855);
   U25846 : XNOR2_X1 port map( A => n25445, B => n24852, ZN => n25071);
   U25847 : XNOR2_X1 port map( A => n25931, B => n3035, ZN => n24853);
   U25848 : XNOR2_X1 port map( A => n25071, B => n24853, ZN => n24854);
   U25849 : XNOR2_X1 port map( A => n24854, B => n24855, ZN => n26381);
   U25850 : OAI21_X1 port map( B1 => n26380, B2 => n26381, A => n26426, ZN => 
                           n24856);
   U25852 : INV_X1 port map( A => n27646, ZN => n26978);
   U25853 : XNOR2_X1 port map( A => n25913, B => n24858, ZN => n25492);
   U25854 : XNOR2_X1 port map( A => n25492, B => n25330, ZN => n24862);
   U25855 : XNOR2_X1 port map( A => n28771, B => n3787, ZN => n24860);
   U25856 : XNOR2_X1 port map( A => n25808, B => n26118, ZN => n24859);
   U25857 : XNOR2_X1 port map( A => n24860, B => n24859, ZN => n24861);
   U25858 : XNOR2_X1 port map( A => n24862, B => n24861, ZN => n27178);
   U25859 : XNOR2_X1 port map( A => n25165, B => n24984, ZN => n26106);
   U25860 : XNOR2_X1 port map( A => n29518, B => n26106, ZN => n24866);
   U25861 : XNOR2_X1 port map( A => n25577, B => n25509, ZN => n24864);
   U25862 : INV_X1 port map( A => n730, ZN => n27879);
   U25863 : XNOR2_X1 port map( A => n25209, B => n27879, ZN => n24863);
   U25864 : XNOR2_X1 port map( A => n24864, B => n24863, ZN => n24865);
   U25865 : XNOR2_X1 port map( A => n24866, B => n24865, ZN => n26129);
   U25867 : INV_X1 port map( A => n26264, ZN => n27130);
   U25868 : XNOR2_X1 port map( A => n25790, B => n26713, ZN => n24867);
   U25869 : XNOR2_X1 port map( A => n25583, B => n25903, ZN => n25128);
   U25870 : XNOR2_X1 port map( A => n24867, B => n25128, ZN => n24869);
   U25871 : XNOR2_X1 port map( A => n26071, B => n25369, ZN => n25105);
   U25872 : XNOR2_X1 port map( A => n25105, B => n25354, ZN => n24868);
   U25873 : XNOR2_X1 port map( A => n24870, B => n25855, ZN => n25570);
   U25874 : XNOR2_X1 port map( A => n29094, B => n25947, ZN => n24871);
   U25875 : XNOR2_X1 port map( A => n24871, B => n25570, ZN => n24875);
   U25876 : XNOR2_X1 port map( A => n26080, B => n25696, ZN => n24872);
   U25877 : XNOR2_X1 port map( A => n24873, B => n24872, ZN => n24874);
   U25878 : XNOR2_X2 port map( A => n24875, B => n24874, ZN => n27175);
   U25879 : XNOR2_X1 port map( A => n25932, B => n29073, ZN => n25141);
   U25880 : XNOR2_X1 port map( A => n25112, B => n25141, ZN => n24879);
   U25881 : INV_X1 port map( A => n2411, ZN => n27766);
   U25882 : XNOR2_X1 port map( A => n29053, B => n27766, ZN => n24876);
   U25883 : XNOR2_X1 port map( A => n24877, B => n24876, ZN => n24878);
   U25884 : XNOR2_X1 port map( A => n24879, B => n24878, ZN => n27177);
   U25885 : XNOR2_X1 port map( A => n25867, B => n25737, ZN => n25348);
   U25886 : XNOR2_X1 port map( A => n29067, B => n25565, ZN => n25102);
   U25887 : XNOR2_X1 port map( A => n25348, B => n25102, ZN => n24882);
   U25888 : XNOR2_X1 port map( A => n29634, B => n4501, ZN => n24880);
   U25889 : XNOR2_X1 port map( A => n25145, B => n24880, ZN => n24881);
   U25890 : MUX2_X1 port map( A => n27175, B => n27178, S => n26263, Z => 
                           n24883);
   U25891 : NAND2_X1 port map( A1 => n28392, A2 => n24883, ZN => n24884);
   U25892 : XNOR2_X1 port map( A => n25262, B => n25107, ZN => n25791);
   U25893 : XNOR2_X1 port map( A => n24885, B => n25791, ZN => n24889);
   U25894 : XNOR2_X1 port map( A => n25542, B => n25261, ZN => n24887);
   U25895 : XNOR2_X1 port map( A => n25428, B => n6319, ZN => n24886);
   U25896 : XNOR2_X1 port map( A => n24887, B => n24886, ZN => n24888);
   U25897 : XNOR2_X2 port map( A => n24889, B => n24888, ZN => n27193);
   U25898 : AOI22_X1 port map( A1 => n24894, A2 => n24893, B1 => n24892, B2 => 
                           n24891, ZN => n24896);
   U25899 : NAND2_X1 port map( A1 => n24896, A2 => n24895, ZN => n25066);
   U25900 : XNOR2_X1 port map( A => n25251, B => n25066, ZN => n24899);
   U25901 : XNOR2_X1 port map( A => n24899, B => n24898, ZN => n24900);
   U25902 : XNOR2_X1 port map( A => n25549, B => n365, ZN => n24901);
   U25903 : XNOR2_X1 port map( A => n25099, B => n24901, ZN => n24905);
   U25904 : INV_X1 port map( A => n3369, ZN => n24902);
   U25905 : XNOR2_X1 port map( A => n25921, B => n24902, ZN => n24903);
   U25906 : XNOR2_X1 port map( A => n25216, B => n24903, ZN => n24904);
   U25907 : XNOR2_X1 port map( A => n24905, B => n24904, ZN => n27190);
   U25908 : XNOR2_X1 port map( A => n25927, B => n25381, ZN => n24908);
   U25909 : XNOR2_X1 port map( A => n25440, B => n24906, ZN => n24907);
   U25910 : XNOR2_X1 port map( A => n24908, B => n24907, ZN => n24910);
   U25911 : XNOR2_X1 port map( A => n25820, B => n25931, ZN => n25029);
   U25912 : XNOR2_X1 port map( A => n25234, B => n25029, ZN => n24909);
   U25914 : INV_X1 port map( A => n2995, ZN => n27444);
   U25915 : XNOR2_X1 port map( A => n25465, B => n27444, ZN => n24911);
   U25916 : XNOR2_X1 port map( A => n24911, B => n25515, ZN => n24912);
   U25917 : XNOR2_X1 port map( A => n25780, B => n28402, ZN => n25271);
   U25918 : XNOR2_X1 port map( A => n24912, B => n25271, ZN => n24915);
   U25919 : XNOR2_X1 port map( A => n24913, B => n26029, ZN => n24914);
   U25921 : AOI21_X1 port map( B1 => n26140, B2 => n26290, A => n27124, ZN => 
                           n24922);
   U25922 : XNOR2_X1 port map( A => n29103, B => n3372, ZN => n24917);
   U25923 : XNOR2_X1 port map( A => n25375, B => n24916, ZN => n25456);
   U25924 : XNOR2_X1 port map( A => n25456, B => n24917, ZN => n24919);
   U25925 : XNOR2_X1 port map( A => n26054, B => n25826, ZN => n25225);
   U25926 : XNOR2_X1 port map( A => n25943, B => n25149, ZN => n25020);
   U25927 : XNOR2_X1 port map( A => n25225, B => n25020, ZN => n24918);
   U25928 : AOI21_X1 port map( B1 => n24920, B2 => n27191, A => n27193, ZN => 
                           n24921);
   U25929 : NOR2_X2 port map( A1 => n24922, A2 => n24921, ZN => n27641);
   U25930 : AOI21_X1 port map( B1 => n27637, B2 => n28466, A => n27641, ZN => 
                           n27640);
   U25931 : OAI21_X1 port map( B1 => n3606, B2 => n26978, A => n27640, ZN => 
                           n24999);
   U25932 : XNOR2_X1 port map( A => n25786, B => n25714, ZN => n24924);
   U25933 : XNOR2_X1 port map( A => n25751, B => n25385, ZN => n24926);
   U25934 : XNOR2_X1 port map( A => n363, B => n25909, ZN => n24927);
   U25935 : XNOR2_X1 port map( A => n25810, B => n28628, ZN => n25589);
   U25936 : XNOR2_X1 port map( A => n25589, B => n24927, ZN => n24931);
   U25937 : XNOR2_X1 port map( A => n25398, B => n3422, ZN => n24929);
   U25938 : XNOR2_X1 port map( A => n29046, B => n25191, ZN => n24928);
   U25939 : XNOR2_X1 port map( A => n24929, B => n24928, ZN => n24930);
   U25941 : XNOR2_X1 port map( A => n24932, B => n25885, ZN => n24935);
   U25942 : INV_X1 port map( A => n3336, ZN => n24933);
   U25943 : XNOR2_X1 port map( A => n28520, B => n24933, ZN => n24934);
   U25944 : XNOR2_X1 port map( A => n24935, B => n24934, ZN => n24937);
   U25945 : XNOR2_X1 port map( A => n25179, B => n25819, ZN => n24936);
   U25946 : XNOR2_X1 port map( A => n24936, B => n25441, ZN => n25560);
   U25947 : XNOR2_X1 port map( A => n25304, B => n24938, ZN => n24941);
   U25948 : XNOR2_X1 port map( A => n25738, B => n25564, ZN => n25188);
   U25949 : XNOR2_X1 port map( A => n25867, B => n26314, ZN => n24939);
   U25950 : XNOR2_X1 port map( A => n25188, B => n24939, ZN => n24940);
   U25951 : XNOR2_X1 port map( A => n24941, B => n24940, ZN => n27161);
   U25953 : XNOR2_X1 port map( A => n25430, B => n25727, ZN => n25174);
   U25954 : XNOR2_X1 port map( A => n25294, B => n25174, ZN => n24945);
   U25955 : XNOR2_X1 port map( A => n25366, B => n25836, ZN => n24943);
   U25956 : XNOR2_X1 port map( A => n25689, B => n3770, ZN => n24942);
   U25957 : XNOR2_X1 port map( A => n24943, B => n24942, ZN => n24944);
   U25958 : XNOR2_X2 port map( A => n24945, B => n24944, ZN => n27701);
   U25960 : XNOR2_X1 port map( A => n25288, B => n24948, ZN => n24952);
   U25961 : XNOR2_X1 port map( A => n24949, B => n25948, ZN => n25572);
   U25962 : XNOR2_X1 port map( A => n25696, B => n3565, ZN => n24950);
   U25963 : XNOR2_X1 port map( A => n25572, B => n24950, ZN => n24951);
   U25964 : XNOR2_X2 port map( A => n24952, B => n24951, ZN => n27704);
   U25965 : AND2_X1 port map( A1 => n27704, A2 => n27702, ZN => n26128);
   U25966 : INV_X1 port map( A => n27703, ZN => n26350);
   U25967 : NAND2_X1 port map( A1 => n27650, A2 => n27641, ZN => n25001);
   U25968 : INV_X1 port map( A => n25001, ZN => n25004);
   U25969 : INV_X1 port map( A => n25736, ZN => n24954);
   U25970 : XNOR2_X1 port map( A => n25187, B => n24954, ZN => n26008);
   U25971 : XNOR2_X1 port map( A => n29533, B => n29634, ZN => n24955);
   U25972 : XNOR2_X1 port map( A => n25864, B => n2982, ZN => n24956);
   U25973 : XNOR2_X1 port map( A => n24272, B => n25922, ZN => n25547);
   U25974 : XNOR2_X1 port map( A => n24956, B => n25547, ZN => n24957);
   U25975 : INV_X1 port map( A => n26384, ZN => n26387);
   U25976 : XNOR2_X1 port map( A => n25293, B => n26040, ZN => n25172);
   U25977 : XNOR2_X1 port map( A => n25260, B => n25172, ZN => n24962);
   U25978 : XNOR2_X1 port map( A => n26046, B => n24959, ZN => n24960);
   U25979 : INV_X1 port map( A => n25498, ZN => n25351);
   U25980 : XNOR2_X1 port map( A => n25082, B => n24960, ZN => n24961);
   U25981 : XNOR2_X1 port map( A => n25133, B => n25808, ZN => n25254);
   U25982 : XNOR2_X1 port map( A => n25849, B => n24963, ZN => n25521);
   U25983 : XNOR2_X1 port map( A => n25254, B => n25521, ZN => n24967);
   U25984 : XNOR2_X1 port map( A => n25328, B => n25845, ZN => n24965);
   U25985 : INV_X1 port map( A => n3223, ZN => n27263);
   U25986 : XNOR2_X1 port map( A => n25745, B => n27263, ZN => n24964);
   U25987 : XNOR2_X1 port map( A => n24965, B => n24964, ZN => n24966);
   U25988 : XNOR2_X2 port map( A => n24967, B => n24966, ZN => n27165);
   U25989 : MUX2_X1 port map( A => n26387, B => n28572, S => n27165, Z => 
                           n24993);
   U25990 : XNOR2_X1 port map( A => n29094, B => n25535, ZN => n26086);
   U25991 : XNOR2_X1 port map( A => n25532, B => n25534, ZN => n25856);
   U25992 : XNOR2_X1 port map( A => n26086, B => n25856, ZN => n24971);
   U25993 : XNOR2_X1 port map( A => n26059, B => n28630, ZN => n24969);
   U25994 : XNOR2_X1 port map( A => n28465, B => n27324, ZN => n24968);
   U25995 : XNOR2_X1 port map( A => n24969, B => n24968, ZN => n24970);
   U25996 : NAND2_X1 port map( A1 => n24973, A2 => n24972, ZN => n24978);
   U25997 : NOR2_X1 port map( A1 => n24975, A2 => n24974, ZN => n24977);
   U26000 : XNOR2_X1 port map( A => n25341, B => n25884, ZN => n25485);
   U26001 : XNOR2_X1 port map( A => n25411, B => n25485, ZN => n24983);
   U26002 : NAND2_X1 port map( A1 => n28642, A2 => n26386, ZN => n24991);
   U26003 : XNOR2_X1 port map( A => n24984, B => n3244, ZN => n24985);
   U26004 : XNOR2_X1 port map( A => n25386, B => n24985, ZN => n24986);
   U26005 : XNOR2_X1 port map( A => n24986, B => n25516, ZN => n24989);
   U26006 : INV_X1 port map( A => n26028, ZN => n24987);
   U26007 : XNOR2_X1 port map( A => n24987, B => n25282, ZN => n25167);
   U26008 : XNOR2_X1 port map( A => n25508, B => n25876, ZN => n25054);
   U26009 : XNOR2_X1 port map( A => n25167, B => n25054, ZN => n24988);
   U26010 : MUX2_X1 port map( A => n24991, B => n24990, S => n27165, Z => 
                           n24992);
   U26012 : NOR2_X1 port map( A1 => n29532, A2 => n25044, ZN => n25003);
   U26014 : INV_X1 port map( A => n27640, ZN => n24996);
   U26015 : NAND2_X1 port map( A1 => n28466, A2 => n3606, ZN => n25047);
   U26016 : INV_X1 port map( A => n25047, ZN => n24994);
   U26017 : NAND3_X1 port map( A1 => n24994, A2 => n27638, A3 => n29532, ZN => 
                           n24995);
   U26018 : INV_X1 port map( A => n26671, ZN => n27645);
   U26019 : NAND3_X1 port map( A1 => n25001, A2 => n27645, A3 => n25044, ZN => 
                           n25050);
   U26020 : NOR3_X1 port map( A1 => n27637, A2 => n26978, A3 => n27645, ZN => 
                           n25002);
   U26021 : AOI21_X1 port map( B1 => n25004, B2 => n25003, A => n25002, ZN => 
                           n25049);
   U26022 : XNOR2_X1 port map( A => n1514, B => n26119, ZN => n25680);
   U26024 : INV_X1 port map( A => n25134, ZN => n25010);
   U26025 : XNOR2_X1 port map( A => n28565, B => n25010, ZN => n25011);
   U26026 : XNOR2_X1 port map( A => n25680, B => n25011, ZN => n25014);
   U26027 : XNOR2_X1 port map( A => n25910, B => n3180, ZN => n25012);
   U26028 : XNOR2_X1 port map( A => n25449, B => n25012, ZN => n25013);
   U26030 : XNOR2_X1 port map( A => n25081, B => n25015, ZN => n25019);
   U26031 : XNOR2_X1 port map( A => n25352, B => n26046, ZN => n25017);
   U26032 : XNOR2_X1 port map( A => n29129, B => n6016, ZN => n25016);
   U26033 : XNOR2_X1 port map( A => n25017, B => n25016, ZN => n25018);
   U26034 : XNOR2_X1 port map( A => n25019, B => n25018, ZN => n25119);
   U26035 : XNOR2_X1 port map( A => n25020, B => n25533, ZN => n25023);
   U26036 : XNOR2_X1 port map( A => n26059, B => n25361, ZN => n25021);
   U26037 : XNOR2_X1 port map( A => n25697, B => n25372, ZN => n26081);
   U26038 : XNOR2_X1 port map( A => n26081, B => n25021, ZN => n25022);
   U26040 : INV_X1 port map( A => n27181, ZN => n26396);
   U26041 : XNOR2_X1 port map( A => n25345, B => n365, ZN => n25024);
   U26042 : XNOR2_X1 port map( A => n300, B => n25546, ZN => n25711);
   U26043 : XNOR2_X1 port map( A => n25024, B => n25711, ZN => n25028);
   U26044 : XNOR2_X1 port map( A => n26094, B => n25736, ZN => n25026);
   U26045 : XNOR2_X1 port map( A => n25921, B => n3154, ZN => n25025);
   U26046 : XNOR2_X1 port map( A => n25026, B => n25025, ZN => n25027);
   U26047 : XNOR2_X1 port map( A => n25028, B => n25027, ZN => n25034);
   U26048 : INV_X1 port map( A => n25034, ZN => n27183);
   U26049 : XNOR2_X1 port map( A => n25029, B => n26101, ZN => n25033);
   U26050 : XNOR2_X1 port map( A => n25890, B => n25702, ZN => n25031);
   U26051 : XNOR2_X1 port map( A => n25760, B => n1215, ZN => n25030);
   U26052 : XNOR2_X1 port map( A => n25031, B => n25030, ZN => n25032);
   U26053 : XNOR2_X1 port map( A => n25033, B => n25032, ZN => n25124);
   U26055 : NAND2_X1 port map( A1 => n25035, A2 => n25034, ZN => n25043);
   U26056 : INV_X1 port map( A => n3598, ZN => n26814);
   U26057 : XNOR2_X1 port map( A => n25268, B => n26814, ZN => n25036);
   U26058 : XNOR2_X1 port map( A => n26109, B => n25036, ZN => n25039);
   U26059 : XNOR2_X1 port map( A => n25037, B => n25322, ZN => n25038);
   U26060 : XNOR2_X1 port map( A => n25039, B => n25038, ZN => n25041);
   U26061 : XNOR2_X1 port map( A => n25041, B => n25040, ZN => n25120);
   U26062 : INV_X1 port map( A => n25120, ZN => n26356);
   U26063 : NAND3_X1 port map( A1 => n27183, A2 => n28651, A3 => n26356, ZN => 
                           n25042);
   U26064 : INV_X1 port map( A => n27639, ZN => n26980);
   U26065 : NOR3_X1 port map( A1 => n26980, A2 => n28466, A3 => n3606, ZN => 
                           n25046);
   U26066 : NOR2_X1 port map( A1 => n27639, A2 => n25044, ZN => n25045);
   U26067 : OAI21_X1 port map( B1 => n25046, B2 => n25045, A => n29532, ZN => 
                           n25048);
   U26070 : XNOR2_X1 port map( A => n25780, B => n3036, ZN => n25053);
   U26071 : XNOR2_X1 port map( A => n25385, B => n25781, ZN => n25055);
   U26072 : XNOR2_X1 port map( A => n25056, B => n25055, ZN => n25057);
   U26073 : XNOR2_X1 port map( A => n365, B => n300, ZN => n25061);
   U26074 : XNOR2_X1 port map( A => n25391, B => n29111, ZN => n25060);
   U26075 : XNOR2_X1 port map( A => n25708, B => n25864, ZN => n25063);
   U26076 : INV_X1 port map( A => Key(19), ZN => n25991);
   U26077 : XNOR2_X1 port map( A => n26095, B => n25991, ZN => n25062);
   U26078 : XNOR2_X1 port map( A => n25063, B => n25062, ZN => n25064);
   U26079 : NOR2_X1 port map( A1 => n26172, A2 => n26173, ZN => n25079);
   U26080 : XNOR2_X1 port map( A => n26114, B => n25066, ZN => n25068);
   U26081 : XNOR2_X1 port map( A => n25808, B => n3622, ZN => n25067);
   U26082 : XNOR2_X1 port map( A => n25068, B => n25067, ZN => n25070);
   U26083 : INV_X1 port map( A => Key(66), ZN => n27742);
   U26084 : XNOR2_X1 port map( A => n25341, B => n25072, ZN => n26104);
   U26085 : XNOR2_X1 port map( A => n25454, B => n26055, ZN => n25074);
   U26086 : XNOR2_X1 port map( A => n26086, B => n25074, ZN => n25078);
   U26087 : XNOR2_X1 port map( A => n25149, B => n25534, ZN => n25076);
   U26088 : XNOR2_X1 port map( A => n25697, B => n3385, ZN => n25075);
   U26089 : XNOR2_X1 port map( A => n25076, B => n25075, ZN => n25077);
   U26090 : XNOR2_X1 port map( A => n25081, B => n25080, ZN => n25085);
   U26091 : XNOR2_X1 port map( A => n25790, B => n3728, ZN => n25083);
   U26092 : XNOR2_X1 port map( A => n25082, B => n25083, ZN => n25084);
   U26093 : NOR2_X1 port map( A1 => n26917, A2 => n26172, ZN => n26781);
   U26094 : XNOR2_X1 port map( A => n25507, B => n25753, ZN => n25088);
   U26095 : XNOR2_X1 port map( A => n28654, B => n25209, ZN => n25388);
   U26096 : XNOR2_X1 port map( A => n29599, B => n3323, ZN => n25086);
   U26097 : XNOR2_X1 port map( A => n25388, B => n25086, ZN => n25087);
   U26098 : XNOR2_X1 port map( A => n25088, B => n25087, ZN => n26280);
   U26099 : XNOR2_X1 port map( A => n26020, B => n29046, ZN => n25493);
   U26100 : XNOR2_X1 port map( A => n25493, B => n25089, ZN => n25093);
   U26101 : XNOR2_X1 port map( A => n28769, B => n3742, ZN => n25091);
   U26102 : XNOR2_X1 port map( A => n26118, B => n25396, ZN => n25090);
   U26103 : XNOR2_X1 port map( A => n25091, B => n25090, ZN => n25092);
   U26106 : XNOR2_X1 port map( A => n25094, B => n25456, ZN => n25098);
   U26107 : XNOR2_X1 port map( A => n26054, B => n29563, ZN => n25096);
   U26108 : XNOR2_X1 port map( A => n3083, B => n26080, ZN => n25095);
   U26109 : XNOR2_X1 port map( A => n25095, B => n25096, ZN => n25097);
   U26112 : XNOR2_X1 port map( A => n26004, B => n25562, ZN => n25734);
   U26113 : XNOR2_X1 port map( A => n25099, B => n25734, ZN => n25104);
   U26114 : INV_X1 port map( A => n2389, ZN => n25100);
   U26115 : XNOR2_X1 port map( A => n25869, B => n25100, ZN => n25101);
   U26116 : XNOR2_X1 port map( A => n25102, B => n25101, ZN => n25103);
   U26117 : XNOR2_X1 port map( A => n25104, B => n25103, ZN => n26278);
   U26118 : XNOR2_X1 port map( A => n25836, B => n26038, ZN => n25106);
   U26119 : XNOR2_X1 port map( A => n25105, B => n25106, ZN => n25111);
   U26120 : XNOR2_X1 port map( A => n29069, B => n25261, ZN => n25109);
   U26121 : XNOR2_X1 port map( A => n1922, B => n2511, ZN => n25108);
   U26122 : XNOR2_X1 port map( A => n25109, B => n25108, ZN => n25110);
   U26123 : XNOR2_X1 port map( A => n25112, B => n25113, ZN => n25117);
   U26124 : XNOR2_X1 port map( A => n25381, B => n2987, ZN => n25115);
   U26125 : XNOR2_X1 port map( A => n25761, B => n25885, ZN => n25114);
   U26126 : XNOR2_X1 port map( A => n25115, B => n25114, ZN => n25116);
   U26127 : XNOR2_X1 port map( A => n25116, B => n25117, ZN => n26797);
   U26128 : INV_X1 port map( A => n26797, ZN => n26362);
   U26129 : INV_X1 port map( A => n25119, ZN => n26397);
   U26130 : NOR2_X1 port map( A1 => n26397, A2 => n27181, ZN => n25123);
   U26131 : AND2_X1 port map( A1 => n27182, A2 => n28467, ZN => n25122);
   U26132 : NAND2_X1 port map( A1 => n26357, A2 => n25124, ZN => n26399);
   U26133 : INV_X1 port map( A => n27203, ZN => n27538);
   U26134 : XNOR2_X1 port map( A => n26040, B => n25262, ZN => n25126);
   U26135 : XNOR2_X1 port map( A => n25689, B => n25543, ZN => n25839);
   U26136 : XNOR2_X1 port map( A => n25126, B => n25839, ZN => n25130);
   U26137 : XNOR2_X1 port map( A => n25352, B => n28007, ZN => n25127);
   U26138 : XNOR2_X1 port map( A => n25128, B => n25127, ZN => n25129);
   U26140 : XNOR2_X1 port map( A => n28565, B => n363, ZN => n25132);
   U26141 : XNOR2_X1 port map( A => n25132, B => n25492, ZN => n25138);
   U26143 : INV_X1 port map( A => n2946, ZN => n26601);
   U26144 : XNOR2_X1 port map( A => n25328, B => n26601, ZN => n25135);
   U26145 : XNOR2_X1 port map( A => n25136, B => n25135, ZN => n25137);
   U26146 : XNOR2_X1 port map( A => n25889, B => n25820, ZN => n25139);
   U26147 : XNOR2_X1 port map( A => n25411, B => n25139, ZN => n25144);
   U26148 : XNOR2_X1 port map( A => n25140, B => n25928, ZN => n25142);
   U26149 : XNOR2_X1 port map( A => n25142, B => n25141, ZN => n25143);
   U26150 : XNOR2_X1 port map( A => n25143, B => n25144, ZN => n26769);
   U26151 : INV_X1 port map( A => n26769, ZN => n26937);
   U26152 : XNOR2_X1 port map( A => n25922, B => n25345, ZN => n25146);
   U26153 : XNOR2_X1 port map( A => n28496, B => n25146, ZN => n25147);
   U26154 : XNOR2_X1 port map( A => n25148, B => n25147, ZN => n26936);
   U26155 : INV_X1 port map( A => n26772, ZN => n25152);
   U26156 : INV_X1 port map( A => n25696, ZN => n25151);
   U26157 : XNOR2_X1 port map( A => n25151, B => n26083, ZN => n25336);
   U26158 : INV_X1 port map( A => n26935, ZN => n26944);
   U26159 : XNOR2_X1 port map( A => n25516, B => n25714, ZN => n25874);
   U26160 : XNOR2_X1 port map( A => n25874, B => n25153, ZN => n25157);
   U26161 : XNOR2_X1 port map( A => n28534, B => n25577, ZN => n25155);
   U26162 : XNOR2_X1 port map( A => n25780, B => n28294, ZN => n25154);
   U26163 : XNOR2_X1 port map( A => n25155, B => n25154, ZN => n25156);
   U26164 : XNOR2_X1 port map( A => n25157, B => n25156, ZN => n26943);
   U26165 : INV_X1 port map( A => n26943, ZN => n26771);
   U26166 : INV_X1 port map( A => n26436, ZN => n26768);
   U26167 : XNOR2_X1 port map( A => n25531, B => n25947, ZN => n25160);
   U26168 : XNOR2_X1 port map( A => n25160, B => n25572, ZN => n25164);
   U26169 : XNOR2_X1 port map( A => n26080, B => n28630, ZN => n25162);
   U26170 : XNOR2_X1 port map( A => n28465, B => n3276, ZN => n25161);
   U26171 : XNOR2_X1 port map( A => n25162, B => n25161, ZN => n25163);
   U26173 : XNOR2_X1 port map( A => n29599, B => n25751, ZN => n25166);
   U26174 : XNOR2_X1 port map( A => n25167, B => n25166, ZN => n25171);
   U26175 : XNOR2_X1 port map( A => n25754, B => n25515, ZN => n25169);
   U26176 : XNOR2_X1 port map( A => n25169, B => n25168, ZN => n25170);
   U26178 : INV_X1 port map( A => n25172, ZN => n25173);
   U26179 : XNOR2_X1 port map( A => n25173, B => n25174, ZN => n25178);
   U26180 : XNOR2_X1 port map( A => n26071, B => n25900, ZN => n25176);
   U26181 : XNOR2_X1 port map( A => n25542, B => n27231, ZN => n25175);
   U26182 : XNOR2_X1 port map( A => n25176, B => n25175, ZN => n25177);
   U26183 : MUX2_X1 port map( A => n29071, B => n29631, S => n26950, Z => 
                           n25197);
   U26184 : XNOR2_X1 port map( A => n25180, B => n26100, ZN => n25181);
   U26185 : XNOR2_X1 port map( A => n25411, B => n25181, ZN => n25184);
   U26186 : XNOR2_X1 port map( A => n25759, B => n25182, ZN => n25929);
   U26187 : XNOR2_X1 port map( A => n25929, B => n25298, ZN => n25183);
   U26188 : XNOR2_X1 port map( A => n25184, B => n25183, ZN => n26951);
   U26189 : INV_X1 port map( A => n26951, ZN => n26948);
   U26190 : XNOR2_X1 port map( A => n25550, B => n3414, ZN => n25185);
   U26191 : XNOR2_X1 port map( A => n25185, B => n29533, ZN => n25186);
   U26192 : XNOR2_X1 port map( A => n25737, B => n25549, ZN => n25920);
   U26193 : XNOR2_X1 port map( A => n25186, B => n25920, ZN => n25189);
   U26194 : MUX2_X1 port map( A => n26948, B => n28542, S => n29071, Z => 
                           n25196);
   U26195 : XNOR2_X1 port map( A => n25190, B => n25914, ZN => n25744);
   U26196 : XNOR2_X1 port map( A => n25191, B => n25845, ZN => n25312);
   U26197 : XNOR2_X1 port map( A => n25312, B => n25744, ZN => n25195);
   U26198 : XNOR2_X1 port map( A => n25328, B => n25909, ZN => n25193);
   U26199 : XNOR2_X1 port map( A => n26118, B => n27605, ZN => n25192);
   U26200 : XNOR2_X1 port map( A => n25193, B => n25192, ZN => n25194);
   U26201 : XNOR2_X1 port map( A => n25195, B => n25194, ZN => n26440);
   U26203 : INV_X1 port map( A => n26431, ZN => n26275);
   U26204 : NAND3_X1 port map( A1 => n26426, A2 => n26382, A3 => n26381, ZN => 
                           n25198);
   U26205 : OAI21_X1 port map( B1 => n26430, B2 => n26275, A => n25198, ZN => 
                           n25201);
   U26206 : INV_X1 port map( A => n26378, ZN => n26427);
   U26207 : MUX2_X1 port map( A => n26427, B => n26426, S => n26381, Z => 
                           n25199);
   U26208 : NOR2_X1 port map( A1 => n26425, A2 => n25199, ZN => n25200);
   U26209 : AOI22_X1 port map( A1 => n27200, A2 => n27203, B1 => n27199, B2 => 
                           n27547, ZN => n25202);
   U26210 : NAND2_X1 port map( A1 => n25203, A2 => n25202, ZN => n25204);
   U26211 : XNOR2_X1 port map( A => n25204, B => n2912, ZN => Ciphertext(74));
   U26212 : XNOR2_X1 port map( A => n25205, B => n25428, ZN => n25206);
   U26213 : XNOR2_X1 port map( A => n25898, B => n25206, ZN => n25208);
   U26214 : XOR2_X1 port map( A => n25209, B => n25509, Z => n25210);
   U26215 : XNOR2_X1 port map( A => n25876, B => n2446, ZN => n25211);
   U26216 : XNOR2_X1 port map( A => n25864, B => n25565, ZN => n25214);
   U26217 : XNOR2_X1 port map( A => n25564, B => n3191, ZN => n25213);
   U26218 : XNOR2_X1 port map( A => n25214, B => n25213, ZN => n25218);
   U26219 : XNOR2_X1 port map( A => n25216, B => n25215, ZN => n25217);
   U26220 : NOR2_X1 port map( A1 => n26731, A2 => n28560, ZN => n25224);
   U26221 : XNOR2_X1 port map( A => n25681, B => n29614, ZN => n25219);
   U26222 : XNOR2_X1 port map( A => n25493, B => n25219, ZN => n25223);
   U26223 : XNOR2_X1 port map( A => n28771, B => n27225, ZN => n25221);
   U26224 : XNOR2_X1 port map( A => n25849, B => n25909, ZN => n25220);
   U26225 : XNOR2_X1 port map( A => n25220, B => n25221, ZN => n25222);
   U26226 : NOR2_X1 port map( A1 => n25224, A2 => n1622, ZN => n25231);
   U26227 : XNOR2_X1 port map( A => n25225, B => n25479, ZN => n25229);
   U26228 : XNOR2_X1 port map( A => n25944, B => n29606, ZN => n25227);
   U26229 : XNOR2_X1 port map( A => n25948, B => n3321, ZN => n25226);
   U26230 : XNOR2_X1 port map( A => n25227, B => n25226, ZN => n25228);
   U26231 : NOR2_X1 port map( A1 => n25628, A2 => n29579, ZN => n25230);
   U26232 : INV_X1 port map( A => n26729, ZN => n26484);
   U26233 : XNOR2_X1 port map( A => n25441, B => n25891, ZN => n25232);
   U26234 : XNOR2_X1 port map( A => n25486, B => n25232, ZN => n25236);
   U26235 : INV_X1 port map( A => n2381, ZN => n27961);
   U26236 : XNOR2_X1 port map( A => n25933, B => n27961, ZN => n25233);
   U26237 : XNOR2_X1 port map( A => n25234, B => n25233, ZN => n25235);
   U26238 : NOR3_X1 port map( A1 => n26484, A2 => n29501, A3 => n1622, ZN => 
                           n25237);
   U26239 : NOR2_X1 port map( A1 => n26194, A2 => n25406, ZN => n27393);
   U26241 : INV_X1 port map( A => n26466, ZN => n25239);
   U26244 : XNOR2_X1 port map( A => n25532, B => n27669, ZN => n25244);
   U26245 : XNOR2_X1 port map( A => n26055, B => n26053, ZN => n25694);
   U26246 : XNOR2_X1 port map( A => n25245, B => n25694, ZN => n25248);
   U26247 : XNOR2_X1 port map( A => n25246, B => n25149, ZN => n25247);
   U26248 : XNOR2_X1 port map( A => n29612, B => n25247, ZN => n25830);
   U26249 : INV_X1 port map( A => n26754, ZN => n26237);
   U26250 : XNOR2_X1 port map( A => n25249, B => n26019, ZN => n25253);
   U26251 : XNOR2_X1 port map( A => n25251, B => n25250, ZN => n25252);
   U26252 : XNOR2_X1 port map( A => n25253, B => n25252, ZN => n25256);
   U26253 : XNOR2_X1 port map( A => n25806, B => n25254, ZN => n25255);
   U26254 : XNOR2_X1 port map( A => n25255, B => n25256, ZN => n25267);
   U26256 : XNOR2_X1 port map( A => n26041, B => n26045, ZN => n25688);
   U26257 : XNOR2_X1 port map( A => n25260, B => n25688, ZN => n25266);
   U26258 : XNOR2_X1 port map( A => n28475, B => n3586, ZN => n25264);
   U26259 : XNOR2_X1 port map( A => n25261, B => n25262, ZN => n25263);
   U26260 : XNOR2_X1 port map( A => n25264, B => n25263, ZN => n25265);
   U26261 : INV_X1 port map( A => n25267, ZN => n26241);
   U26262 : INV_X1 port map( A => n25268, ZN => n25269);
   U26263 : XNOR2_X1 port map( A => n25270, B => n25269, ZN => n26030);
   U26264 : XNOR2_X1 port map( A => n25271, B => n26030, ZN => n25275);
   U26265 : XNOR2_X1 port map( A => n25324, B => n29247, ZN => n25272);
   U26266 : XNOR2_X1 port map( A => n25272, B => n25781, ZN => n25273);
   U26267 : XNOR2_X1 port map( A => n25273, B => n25516, ZN => n25274);
   U26268 : XNOR2_X1 port map( A => n25274, B => n25275, ZN => n26755);
   U26269 : XNOR2_X1 port map( A => n25412, B => n25277, ZN => n25281);
   U26270 : XNOR2_X1 port map( A => n24852, B => n3374, ZN => n25279);
   U26271 : XNOR2_X1 port map( A => n25702, B => n25440, ZN => n25278);
   U26272 : XNOR2_X1 port map( A => n25279, B => n25278, ZN => n25280);
   U26273 : XNOR2_X1 port map( A => n25281, B => n25280, ZN => n26240);
   U26274 : NAND2_X1 port map( A1 => n26237, A2 => n25603, ZN => n25357);
   U26275 : XNOR2_X1 port map( A => n25517, B => n25875, ZN => n25286);
   U26276 : XNOR2_X1 port map( A => n25786, B => n25515, ZN => n25284);
   U26277 : XNOR2_X1 port map( A => n1871, B => n2916, ZN => n25283);
   U26278 : XNOR2_X1 port map( A => n25284, B => n25283, ZN => n25285);
   U26279 : XNOR2_X1 port map( A => n25287, B => n25288, ZN => n25292);
   U26280 : XNOR2_X1 port map( A => n28630, B => n25855, ZN => n25290);
   U26281 : XNOR2_X1 port map( A => n25372, B => n1927, ZN => n25289);
   U26282 : XNOR2_X1 port map( A => n25290, B => n25289, ZN => n25291);
   U26283 : XNOR2_X1 port map( A => n25583, B => n25293, ZN => n25840);
   U26284 : XNOR2_X1 port map( A => n25294, B => n25840, ZN => n25297);
   U26285 : XNOR2_X1 port map( A => n29129, B => n2894, ZN => n25295);
   U26286 : XNOR2_X1 port map( A => n25541, B => n25295, ZN => n25296);
   U26288 : INV_X1 port map( A => n25659, ZN => n26716);
   U26289 : XNOR2_X1 port map( A => n25298, B => n25408, ZN => n25302);
   U26290 : XNOR2_X1 port map( A => n26100, B => n25819, ZN => n25300);
   U26291 : XNOR2_X1 port map( A => n25891, B => n26531, ZN => n25299);
   U26292 : XNOR2_X1 port map( A => n25300, B => n25299, ZN => n25301);
   U26293 : XNOR2_X1 port map( A => n25302, B => n25301, ZN => n26718);
   U26294 : INV_X1 port map( A => n25868, ZN => n25303);
   U26295 : XNOR2_X1 port map( A => n25303, B => n29533, ZN => n25474);
   U26296 : XNOR2_X1 port map( A => n25304, B => n25474, ZN => n25308);
   U26297 : XNOR2_X1 port map( A => n25864, B => n28485, ZN => n25306);
   U26298 : XNOR2_X1 port map( A => n29067, B => n1062, ZN => n25305);
   U26299 : XNOR2_X1 port map( A => n25306, B => n25305, ZN => n25307);
   U26300 : MUX2_X1 port map( A => n26718, B => n28459, S => n26717, Z => 
                           n25315);
   U26301 : XNOR2_X1 port map( A => n25810, B => n1246, ZN => n25309);
   U26302 : XNOR2_X1 port map( A => n25310, B => n25309, ZN => n25314);
   U26303 : XNOR2_X1 port map( A => n25312, B => n25311, ZN => n25313);
   U26305 : NAND2_X1 port map( A1 => n28503, A2 => n29528, ZN => n25319);
   U26306 : NAND2_X1 port map( A1 => n25666, A2 => n28525, ZN => n25318);
   U26307 : MUX2_X1 port map( A => n25319, B => n25318, S => n28547, Z => 
                           n25320);
   U26308 : XNOR2_X1 port map( A => n26107, B => n29518, ZN => n25327);
   U26309 : XNOR2_X1 port map( A => n1871, B => n26028, ZN => n25717);
   U26310 : XNOR2_X1 port map( A => n25324, B => n2402, ZN => n25325);
   U26311 : XNOR2_X1 port map( A => n25717, B => n25325, ZN => n25326);
   U26312 : XNOR2_X1 port map( A => n26115, B => n25328, ZN => n25329);
   U26313 : XNOR2_X1 port map( A => n25330, B => n25329, ZN => n25334);
   U26314 : XNOR2_X1 port map( A => n28645, B => n29543, ZN => n25332);
   U26315 : XNOR2_X1 port map( A => n26120, B => n27956, ZN => n25331);
   U26316 : XNOR2_X1 port map( A => n25332, B => n25331, ZN => n25333);
   U26317 : XNOR2_X1 port map( A => n25334, B => n25333, ZN => n25344);
   U26318 : INV_X1 port map( A => n25344, ZN => n26235);
   U26319 : XNOR2_X1 port map( A => n25947, B => n29612, ZN => n25335);
   U26320 : XNOR2_X1 port map( A => n25336, B => n25335, ZN => n25339);
   U26321 : XNOR2_X1 port map( A => n25535, B => n3686, ZN => n25337);
   U26322 : XNOR2_X1 port map( A => n25698, B => n25337, ZN => n25338);
   U26323 : XNOR2_X1 port map( A => n25338, B => n25339, ZN => n25654);
   U26325 : XNOR2_X1 port map( A => n26011, B => n3087, ZN => n25342);
   U26326 : INV_X1 port map( A => n25341, ZN => n25526);
   U26327 : XNOR2_X1 port map( A => n25526, B => n25342, ZN => n25343);
   U26329 : NOR2_X1 port map( A1 => n26230, A2 => n26737, ZN => n25349);
   U26330 : XNOR2_X1 port map( A => n26095, B => Key(151), ZN => n25347);
   U26331 : XNOR2_X1 port map( A => n26077, B => n25687, ZN => n25356);
   U26332 : XNOR2_X1 port map( A => n28475, B => n28097, ZN => n25353);
   U26333 : XNOR2_X1 port map( A => n25354, B => n25353, ZN => n25355);
   U26334 : XNOR2_X1 port map( A => n25356, B => n25355, ZN => n25597);
   U26335 : INV_X1 port map( A => n25597, ZN => n26200);
   U26336 : INV_X1 port map( A => n25357, ZN => n25358);
   U26340 : XNOR2_X1 port map( A => n25367, B => n25366, ZN => n25368);
   U26341 : XNOR2_X1 port map( A => n26041, B => n25369, ZN => n25370);
   U26342 : XNOR2_X1 port map( A => n26039, B => n25370, ZN => n25371);
   U26343 : XNOR2_X1 port map( A => n25944, B => n26053, ZN => n25374);
   U26344 : XNOR2_X1 port map( A => n25372, B => n2804, ZN => n25373);
   U26345 : XNOR2_X1 port map( A => n25374, B => n25373, ZN => n25377);
   U26346 : XNOR2_X1 port map( A => n25454, B => n26059, ZN => n25721);
   U26347 : XNOR2_X1 port map( A => n25375, B => n26084, ZN => n25828);
   U26348 : XNOR2_X1 port map( A => n25721, B => n25828, ZN => n25376);
   U26349 : XNOR2_X1 port map( A => n25376, B => n25377, ZN => n26420);
   U26350 : INV_X1 port map( A => n26420, ZN => n26567);
   U26351 : XNOR2_X1 port map( A => n25445, B => n25703, ZN => n25380);
   U26352 : XNOR2_X1 port map( A => n25933, B => n25378, ZN => n25379);
   U26353 : XNOR2_X1 port map( A => n25380, B => n25379, ZN => n25384);
   U26354 : INV_X1 port map( A => n25381, ZN => n25382);
   U26355 : XNOR2_X1 port map( A => n25760, B => n25382, ZN => n25442);
   U26356 : XNOR2_X1 port map( A => n25442, B => n26015, ZN => n25383);
   U26357 : XNOR2_X1 port map( A => n25383, B => n25384, ZN => n26786);
   U26358 : XNOR2_X1 port map( A => n25386, B => n25385, ZN => n25756);
   U26359 : XNOR2_X1 port map( A => n25387, B => n25756, ZN => n25390);
   U26360 : XNOR2_X1 port map( A => n26109, B => n1046, ZN => n25389);
   U26361 : XNOR2_X1 port map( A => n25773, B => n29017, ZN => n25436);
   U26362 : XNOR2_X1 port map( A => n26094, B => n2404, ZN => n25393);
   U26363 : XNOR2_X1 port map( A => n25391, B => n25565, ZN => n25392);
   U26364 : XNOR2_X1 port map( A => n25393, B => n25392, ZN => n25394);
   U26365 : XNOR2_X1 port map( A => n28769, B => n25396, ZN => n25397);
   U26366 : XNOR2_X1 port map( A => n25680, B => n25397, ZN => n25401);
   U26367 : XNOR2_X1 port map( A => n25809, B => n25745, ZN => n26025);
   U26368 : XNOR2_X1 port map( A => n25398, B => n3451, ZN => n25399);
   U26369 : XNOR2_X1 port map( A => n26025, B => n25399, ZN => n25400);
   U26370 : NOR2_X1 port map( A1 => n26912, A2 => n26914, ZN => n26788);
   U26372 : NAND3_X1 port map( A1 => n29617, A2 => n29028, A3 => n25239, ZN => 
                           n25405);
   U26375 : XNOR2_X1 port map( A => n24852, B => n2522, ZN => n25410);
   U26376 : XNOR2_X1 port map( A => n25408, B => n25381, ZN => n25409);
   U26377 : XNOR2_X1 port map( A => n25410, B => n25409, ZN => n25414);
   U26378 : XNOR2_X1 port map( A => n25412, B => n25411, ZN => n25413);
   U26379 : NAND2_X1 port map( A1 => n26179, A2 => n26448, ZN => n26455);
   U26380 : AND2_X1 port map( A1 => n26447, A2 => n26449, ZN => n25416);
   U26382 : NOR2_X1 port map( A1 => n26576, A2 => n28710, ZN => n25419);
   U26383 : INV_X1 port map( A => n26576, ZN => n25421);
   U26384 : NOR3_X1 port map( A1 => n25421, A2 => n29576, A3 => n28711, ZN => 
                           n25422);
   U26386 : NOR2_X1 port map( A1 => n25426, A2 => n25425, ZN => n25427);
   U26387 : XNOR2_X1 port map( A => n25427, B => n3565, ZN => Ciphertext(40));
   U26388 : XNOR2_X1 port map( A => n25428, B => n26070, ZN => n25691);
   U26389 : XNOR2_X1 port map( A => n25429, B => n25691, ZN => n25434);
   U26390 : INV_X1 port map( A => n25430, ZN => n25431);
   U26391 : XNOR2_X1 port map( A => n25431, B => n3164, ZN => n25432);
   U26392 : XNOR2_X2 port map( A => n25434, B => n25433, ZN => n26222);
   U26393 : XNOR2_X1 port map( A => n25564, B => n3501, ZN => n25435);
   U26394 : XNOR2_X1 port map( A => n25436, B => n25435, ZN => n25439);
   U26395 : XNOR2_X1 port map( A => n25775, B => n300, ZN => n25437);
   U26396 : XNOR2_X1 port map( A => n25735, B => n25437, ZN => n25438);
   U26398 : NOR2_X1 port map( A1 => n26222, A2 => n29100, ZN => n25462);
   U26399 : XNOR2_X1 port map( A => n25441, B => n25440, ZN => n25443);
   U26400 : XNOR2_X1 port map( A => n25442, B => n25443, ZN => n25448);
   U26401 : XNOR2_X1 port map( A => n25890, B => n25444, ZN => n25701);
   U26402 : XNOR2_X1 port map( A => n28520, B => n3015, ZN => n25446);
   U26403 : XNOR2_X1 port map( A => n25446, B => n25701, ZN => n25447);
   U26404 : XNOR2_X1 port map( A => n25807, B => n25449, ZN => n25452);
   U26405 : XNOR2_X1 port map( A => n25909, B => n3049, ZN => n25450);
   U26406 : XNOR2_X1 port map( A => n25743, B => n25450, ZN => n25451);
   U26407 : XNOR2_X1 port map( A => n25452, B => n25451, ZN => n26749);
   U26408 : INV_X1 port map( A => n26749, ZN => n25453);
   U26409 : XNOR2_X1 port map( A => n25826, B => n25454, ZN => n25455);
   U26410 : XNOR2_X1 port map( A => n25456, B => n25455, ZN => n25460);
   U26411 : XNOR2_X1 port map( A => n25948, B => n3643, ZN => n25457);
   U26412 : XNOR2_X1 port map( A => n25458, B => n25457, ZN => n25459);
   U26413 : XNOR2_X1 port map( A => n25459, B => n25460, ZN => n26746);
   U26415 : XNOR2_X1 port map( A => n28402, B => n26108, ZN => n25464);
   U26416 : XNOR2_X1 port map( A => n25756, B => n25464, ZN => n25469);
   U26417 : XNOR2_X1 port map( A => n25782, B => n1923, ZN => n25466);
   U26418 : XNOR2_X1 port map( A => n25467, B => n25466, ZN => n25468);
   U26419 : NOR2_X1 port map( A1 => n29159, A2 => n26747, ZN => n25645);
   U26420 : NAND2_X1 port map( A1 => n25645, A2 => n26222, ZN => n25471);
   U26421 : XNOR2_X1 port map( A => n26004, B => n25737, ZN => n25473);
   U26422 : XNOR2_X1 port map( A => n25474, B => n25473, ZN => n25478);
   U26423 : XNOR2_X1 port map( A => n25869, B => n2981, ZN => n25476);
   U26427 : XNOR2_X1 port map( A => n25947, B => n26054, ZN => n25724);
   U26428 : XNOR2_X1 port map( A => n25724, B => n25479, ZN => n25483);
   U26429 : XNOR2_X1 port map( A => n25855, B => n25535, ZN => n25481);
   U26430 : XNOR2_X1 port map( A => n25858, B => n3633, ZN => n25480);
   U26431 : XNOR2_X1 port map( A => n25481, B => n25480, ZN => n25482);
   U26433 : XNOR2_X1 port map( A => n25486, B => n25485, ZN => n25491);
   U26434 : INV_X1 port map( A => n25886, ZN => n25487);
   U26435 : XNOR2_X1 port map( A => n29154, B => n25487, ZN => n25489);
   U26436 : XNOR2_X1 port map( A => n25761, B => n3462, ZN => n25488);
   U26437 : XNOR2_X1 port map( A => n25489, B => n25488, ZN => n25490);
   U26438 : XNOR2_X1 port map( A => n25491, B => n25490, ZN => n27014);
   U26439 : NAND2_X1 port map( A1 => n26623, A2 => n27014, ZN => n25505);
   U26440 : XNOR2_X1 port map( A => n25493, B => n25492, ZN => n25497);
   U26441 : XNOR2_X1 port map( A => n25914, B => n25845, ZN => n25495);
   U26442 : XNOR2_X1 port map( A => n26120, B => n3491, ZN => n25494);
   U26443 : XNOR2_X1 port map( A => n25495, B => n25494, ZN => n25496);
   U26445 : XNOR2_X1 port map( A => n25498, B => n3660, ZN => n25499);
   U26446 : XNOR2_X1 port map( A => n25499, B => n25900, ZN => n25500);
   U26447 : XNOR2_X1 port map( A => n25840, B => n25500, ZN => n25501);
   U26448 : NAND2_X1 port map( A1 => n28639, A2 => n27052, ZN => n25506);
   U26449 : NOR2_X1 port map( A1 => n27052, A2 => n27013, ZN => n25504);
   U26450 : XNOR2_X1 port map( A => n25507, B => n25875, ZN => n25512);
   U26451 : XNOR2_X1 port map( A => n25508, B => n3463, ZN => n25510);
   U26452 : XNOR2_X1 port map( A => n29485, B => n25509, ZN => n25940);
   U26453 : XNOR2_X1 port map( A => n25510, B => n25940, ZN => n25511);
   U26454 : NOR2_X1 port map( A1 => n29160, A2 => n28025, ZN => n28039);
   U26455 : XNOR2_X1 port map( A => n25513, B => n2598, ZN => n25514);
   U26456 : XNOR2_X1 port map( A => n26107, B => n25514, ZN => n25519);
   U26457 : XNOR2_X1 port map( A => n25516, B => n25515, ZN => n25942);
   U26458 : XNOR2_X1 port map( A => n25517, B => n25942, ZN => n25518);
   U26459 : XNOR2_X1 port map( A => n25518, B => n25519, ZN => n27043);
   U26460 : XNOR2_X1 port map( A => n26118, B => n3483, ZN => n25520);
   U26461 : XNOR2_X1 port map( A => n25521, B => n25520, ZN => n25524);
   U26462 : XNOR2_X1 port map( A => n26115, B => n26019, ZN => n25522);
   U26463 : XNOR2_X1 port map( A => n25915, B => n25522, ZN => n25523);
   U26464 : XNOR2_X1 port map( A => n25702, B => n3212, ZN => n25525);
   U26465 : XNOR2_X1 port map( A => n25927, B => n25525, ZN => n25528);
   U26466 : XNOR2_X1 port map( A => n25526, B => n25928, ZN => n25527);
   U26467 : XNOR2_X1 port map( A => n25528, B => n25527, ZN => n25530);
   U26468 : XNOR2_X1 port map( A => n25529, B => n25530, ZN => n27048);
   U26469 : INV_X1 port map( A => n29570, ZN => n27004);
   U26470 : XNOR2_X1 port map( A => n29103, B => n25532, ZN => n25945);
   U26471 : XNOR2_X1 port map( A => n25945, B => n25533, ZN => n25539);
   U26472 : XNOR2_X1 port map( A => n25535, B => n29606, ZN => n25537);
   U26473 : XNOR2_X1 port map( A => n26080, B => n3380, ZN => n25536);
   U26474 : XNOR2_X1 port map( A => n25536, B => n25537, ZN => n25538);
   U26476 : OAI21_X1 port map( B1 => n27001, B2 => n27004, A => n28783, ZN => 
                           n25556);
   U26477 : XNOR2_X1 port map( A => n26041, B => n1123, ZN => n25540);
   U26478 : XNOR2_X1 port map( A => n25541, B => n25540, ZN => n25545);
   U26479 : XNOR2_X1 port map( A => n25542, B => n25543, ZN => n25899);
   U26480 : XNOR2_X1 port map( A => n26077, B => n25899, ZN => n25544);
   U26481 : XNOR2_X1 port map( A => n25546, B => n25345, ZN => n25548);
   U26482 : XNOR2_X1 port map( A => n25548, B => n25547, ZN => n25554);
   U26483 : XNOR2_X1 port map( A => n25864, B => n25549, ZN => n25552);
   U26484 : XNOR2_X1 port map( A => n29067, B => n1175, ZN => n25551);
   U26485 : XNOR2_X1 port map( A => n25552, B => n25551, ZN => n25553);
   U26488 : NOR2_X1 port map( A1 => n28039, A2 => n29031, ZN => n25607);
   U26489 : XNOR2_X1 port map( A => n26102, B => n25931, ZN => n25558);
   U26490 : XNOR2_X1 port map( A => n25559, B => n25558, ZN => n25561);
   U26491 : XNOR2_X1 port map( A => n26093, B => n25562, ZN => n25771);
   U26492 : XNOR2_X1 port map( A => n25771, B => n25563, ZN => n25568);
   U26493 : XNOR2_X1 port map( A => n25565, B => n25564, ZN => n25919);
   U26494 : XNOR2_X1 port map( A => n25868, B => n1248, ZN => n25566);
   U26495 : XNOR2_X1 port map( A => n25919, B => n25566, ZN => n25567);
   U26497 : INV_X1 port map( A => n26998, ZN => n25575);
   U26498 : XNOR2_X1 port map( A => n25569, B => n25570, ZN => n25574);
   U26499 : XNOR2_X1 port map( A => n25825, B => n3457, ZN => n25571);
   U26500 : XNOR2_X1 port map( A => n25572, B => n25571, ZN => n25573);
   U26503 : INV_X1 port map( A => n26997, ZN => n25588);
   U26504 : XNOR2_X1 port map( A => n25939, B => n25576, ZN => n25581);
   U26505 : XNOR2_X1 port map( A => n25786, B => n25577, ZN => n25579);
   U26506 : XNOR2_X1 port map( A => n26110, B => n25751, ZN => n25578);
   U26507 : XNOR2_X1 port map( A => n25579, B => n25578, ZN => n25580);
   U26508 : XNOR2_X1 port map( A => n25581, B => n25580, ZN => n26733);
   U26509 : XNOR2_X1 port map( A => n25901, B => n25727, ZN => n25582);
   U26510 : XNOR2_X1 port map( A => n25898, B => n25582, ZN => n25587);
   U26511 : XNOR2_X1 port map( A => n25729, B => n28540, ZN => n25585);
   U26512 : XNOR2_X1 port map( A => n26039, B => n3710, ZN => n25584);
   U26513 : XNOR2_X1 port map( A => n25585, B => n25584, ZN => n25586);
   U26514 : MUX2_X1 port map( A => n25588, B => n26733, S => n26995, Z => 
                           n25595);
   U26515 : XNOR2_X1 port map( A => n25589, B => n25590, ZN => n25594);
   U26516 : XNOR2_X1 port map( A => n25848, B => n25909, ZN => n25592);
   U26517 : XNOR2_X1 port map( A => n28771, B => n3528, ZN => n25591);
   U26518 : XNOR2_X1 port map( A => n25592, B => n25591, ZN => n25593);
   U26519 : INV_X1 port map( A => n25654, ZN => n26203);
   U26520 : OAI22_X1 port map( A1 => n26204, A2 => n26230, B1 => n26203, B2 => 
                           n26229, ZN => n25598);
   U26521 : INV_X1 port map( A => n26204, ZN => n26228);
   U26522 : AOI22_X1 port map( A1 => n26741, A2 => n26228, B1 => n26230, B2 => 
                           n26200, ZN => n25599);
   U26524 : INV_X1 port map( A => n28038, ZN => n25601);
   U26525 : AOI21_X1 port map( B1 => n26237, B2 => n25603, A => n25602, ZN => 
                           n25605);
   U26526 : NAND2_X1 port map( A1 => n26753, A2 => n26755, ZN => n25604);
   U26527 : OAI21_X1 port map( B1 => n25605, B2 => n26753, A => n25604, ZN => 
                           n25606);
   U26528 : INV_X1 port map( A => n25649, ZN => n26242);
   U26529 : NOR2_X1 port map( A1 => n25606, A2 => n26242, ZN => n26658);
   U26530 : NOR2_X1 port map( A1 => n26760, A2 => n26240, ZN => n26659);
   U26531 : NOR2_X1 port map( A1 => n26658, A2 => n26659, ZN => n26602);
   U26532 : OAI22_X1 port map( A1 => n25607, A2 => n28035, B1 => n26664, B2 => 
                           n26602, ZN => n25608);
   U26533 : XNOR2_X1 port map( A => n25608, B => n2117, ZN => Ciphertext(179));
   U26534 : INV_X1 port map( A => n28547, ZN => n25670);
   U26535 : NAND2_X1 port map( A1 => n26181, A2 => n28503, ZN => n26477);
   U26536 : NOR2_X1 port map( A1 => n25670, A2 => n26477, ZN => n25612);
   U26537 : OAI21_X1 port map( B1 => n26186, B2 => n26185, A => n26476, ZN => 
                           n25609);
   U26538 : AOI21_X1 port map( B1 => n26182, B2 => n28503, A => n25609, ZN => 
                           n25610);
   U26539 : INV_X1 port map( A => n27407, ZN => n27402);
   U26540 : NOR2_X1 port map( A1 => n28476, A2 => n28434, ZN => n25613);
   U26541 : NOR2_X1 port map( A1 => n25614, A2 => n25613, ZN => n26159);
   U26542 : OAI21_X1 port map( B1 => n26560, B2 => n28434, A => n377, ZN => 
                           n25615);
   U26543 : NAND2_X1 port map( A1 => n28385, A2 => n25615, ZN => n25616);
   U26545 : NAND2_X1 port map( A1 => n27402, A2 => n27386, ZN => n27404);
   U26548 : INV_X1 port map( A => n25622, ZN => n25624);
   U26549 : OAI21_X1 port map( B1 => n26448, B2 => n26449, A => n26162, ZN => 
                           n25623);
   U26550 : NOR2_X1 port map( A1 => n25624, A2 => n25623, ZN => n25626);
   U26551 : NOR2_X1 port map( A1 => n26454, A2 => n26448, ZN => n25625);
   U26552 : OAI211_X1 port map( C1 => n27404, C2 => n28607, A => n25627, B => 
                           n1175, ZN => n25634);
   U26553 : NAND2_X1 port map( A1 => n28548, A2 => n29560, ZN => n25665);
   U26554 : INV_X1 port map( A => n26715, ZN => n26209);
   U26556 : INV_X1 port map( A => n26721, ZN => n26208);
   U26557 : INV_X1 port map( A => n26718, ZN => n26215);
   U26558 : OAI21_X1 port map( B1 => n26723, B2 => n26208, A => n26215, ZN => 
                           n25631);
   U26559 : NAND2_X1 port map( A1 => n27402, A2 => n27387, ZN => n25636);
   U26560 : NOR2_X1 port map( A1 => n26960, A2 => n1175, ZN => n25635);
   U26561 : OAI211_X1 port map( C1 => n27410, C2 => n27402, A => n25636, B => 
                           n25635, ZN => n25637);
   U26562 : NAND2_X1 port map( A1 => n25638, A2 => n25637, ZN => n25639);
   U26563 : NOR2_X1 port map( A1 => n25640, A2 => n25639, ZN => Ciphertext(20))
                           ;
   U26564 : NOR2_X1 port map( A1 => n29501, A2 => n28560, ZN => n25641);
   U26565 : NAND2_X1 port map( A1 => n25453, A2 => n26747, ZN => n25647);
   U26566 : NAND2_X1 port map( A1 => n29099, A2 => n26747, ZN => n25642);
   U26567 : NAND2_X1 port map( A1 => n5760, A2 => n25642, ZN => n25643);
   U26568 : OAI21_X1 port map( B1 => n25645, B2 => n25644, A => n25643, ZN => 
                           n25646);
   U26569 : OAI21_X1 port map( B1 => n5035, B2 => n25647, A => n25646, ZN => 
                           n27354);
   U26570 : INV_X1 port map( A => n27354, ZN => n25657);
   U26571 : NOR2_X1 port map( A1 => n27340, A2 => n25657, ZN => n25658);
   U26573 : INV_X1 port map( A => n25650, ZN => n25653);
   U26574 : NOR2_X1 port map( A1 => n26761, A2 => n26237, ZN => n25652);
   U26575 : NAND2_X1 port map( A1 => n26241, A2 => n26755, ZN => n25651);
   U26576 : AOI22_X2 port map( A1 => n25975, A2 => n25653, B1 => n25652, B2 => 
                           n25651, ZN => n27358);
   U26577 : INV_X1 port map( A => n27358, ZN => n27350);
   U26578 : INV_X1 port map( A => n26742, ZN => n25656);
   U26579 : NOR2_X1 port map( A1 => n26204, A2 => n25597, ZN => n26738);
   U26580 : NOR2_X1 port map( A1 => n26203, A2 => n26740, ZN => n25655);
   U26581 : NOR2_X1 port map( A1 => n28473, A2 => n25654, ZN => n26739);
   U26584 : INV_X1 port map( A => n26717, ZN => n26210);
   U26585 : NOR2_X1 port map( A1 => n29560, A2 => n26718, ZN => n25661);
   U26587 : NOR2_X1 port map( A1 => n28548, A2 => n28459, ZN => n25662);
   U26588 : NAND2_X1 port map( A1 => n25662, A2 => n283, ZN => n25663);
   U26589 : NAND3_X1 port map( A1 => n27350, A2 => n29052, A3 => n28549, ZN => 
                           n25672);
   U26590 : OR2_X1 port map( A1 => n27340, A2 => n27352, ZN => n25957);
   U26591 : NOR2_X1 port map( A1 => n26186, A2 => n26182, ZN => n26472);
   U26592 : NOR2_X1 port map( A1 => n25666, A2 => n26185, ZN => n25667);
   U26593 : NOR2_X1 port map( A1 => n26472, A2 => n25667, ZN => n26474);
   U26594 : INV_X1 port map( A => n28561, ZN => n25668);
   U26595 : AOI21_X1 port map( B1 => n26180, B2 => n25668, A => n28525, ZN => 
                           n25669);
   U26597 : INV_X1 port map( A => n1046, ZN => n25674);
   U26598 : XNOR2_X1 port map( A => n25675, B => n25674, ZN => Ciphertext(5));
   U26599 : NOR2_X1 port map( A1 => n27048, A2 => n28130, ZN => n25968);
   U26600 : INV_X1 port map( A => n27044, ZN => n27002);
   U26601 : AOI21_X1 port map( B1 => n28783, B2 => n27002, A => n27048, ZN => 
                           n25677);
   U26602 : OR2_X1 port map( A1 => n25677, A2 => n27041, ZN => n25678);
   U26603 : NAND2_X1 port map( A1 => n25679, A2 => n25678, ZN => n26539);
   U26604 : INV_X1 port map( A => n26539, ZN => n27865);
   U26605 : XNOR2_X1 port map( A => n26021, B => n25680, ZN => n25686);
   U26606 : INV_X1 port map( A => n25681, ZN => n25682);
   U26607 : XNOR2_X1 port map( A => n363, B => n25682, ZN => n25684);
   U26608 : XNOR2_X1 port map( A => n26114, B => n27298, ZN => n25683);
   U26609 : XNOR2_X1 port map( A => n25683, B => n25684, ZN => n25685);
   U26610 : XNOR2_X1 port map( A => n25685, B => n25686, ZN => n26614);
   U26611 : XNOR2_X1 port map( A => n25687, B => n25688, ZN => n25693);
   U26612 : XNOR2_X1 port map( A => n25689, B => n26680, ZN => n25690);
   U26613 : XNOR2_X1 port map( A => n25691, B => n25690, ZN => n25692);
   U26614 : XNOR2_X1 port map( A => n25826, B => n1133, ZN => n25695);
   U26615 : XNOR2_X1 port map( A => n25694, B => n25695, ZN => n25700);
   U26616 : XNOR2_X1 port map( A => n25697, B => n25696, ZN => n25859);
   U26617 : XNOR2_X1 port map( A => n25698, B => n25859, ZN => n25699);
   U26619 : XNOR2_X1 port map( A => n25701, B => n26013, ZN => n25707);
   U26620 : XNOR2_X1 port map( A => n25702, B => n29053, ZN => n25705);
   U26621 : XNOR2_X1 port map( A => n25703, B => n3196, ZN => n25704);
   U26622 : XNOR2_X1 port map( A => n25705, B => n25704, ZN => n25706);
   U26623 : XNOR2_X1 port map( A => n25775, B => n25867, ZN => n25710);
   U26624 : XNOR2_X1 port map( A => n25708, B => n2912, ZN => n25709);
   U26625 : XNOR2_X1 port map( A => n25710, B => n25709, ZN => n25712);
   U26626 : XNOR2_X1 port map( A => n25714, B => n26108, ZN => n25715);
   U26627 : XNOR2_X1 port map( A => n26030, B => n25715, ZN => n25719);
   U26628 : XNOR2_X1 port map( A => n25785, B => n135, ZN => n25716);
   U26629 : XNOR2_X1 port map( A => n25717, B => n25716, ZN => n25718);
   U26631 : NOR2_X1 port map( A1 => n27865, A2 => n27877, ZN => n26594);
   U26632 : XNOR2_X1 port map( A => n25722, B => n25721, ZN => n25726);
   U26633 : XNOR2_X1 port map( A => n29563, B => n3606, ZN => n25723);
   U26634 : XNOR2_X1 port map( A => n25724, B => n25723, ZN => n25725);
   U26635 : XNOR2_X1 port map( A => n25726, B => n25725, ZN => n26988);
   U26636 : INV_X1 port map( A => n26988, ZN => n26991);
   U26637 : XNOR2_X1 port map( A => n25727, B => n26038, ZN => n25728);
   U26638 : XNOR2_X1 port map( A => n25900, B => n440, ZN => n25731);
   U26639 : XNOR2_X1 port map( A => n25729, B => n26046, ZN => n25730);
   U26640 : XNOR2_X1 port map( A => n25730, B => n25731, ZN => n25732);
   U26641 : XNOR2_X2 port map( A => n25733, B => n25732, ZN => n27074);
   U26642 : XNOR2_X1 port map( A => n25735, B => n25734, ZN => n25742);
   U26643 : XNOR2_X1 port map( A => n25737, B => n29017, ZN => n25740);
   U26644 : XNOR2_X1 port map( A => n25738, B => n2505, ZN => n25739);
   U26645 : XNOR2_X1 port map( A => n25740, B => n25739, ZN => n25741);
   U26647 : XNOR2_X1 port map( A => n28593, B => n25810, ZN => n25747);
   U26648 : XNOR2_X1 port map( A => n25745, B => n3662, ZN => n25746);
   U26650 : XNOR2_X1 port map( A => n26029, B => n25751, ZN => n25752);
   U26651 : XNOR2_X1 port map( A => n25752, B => n25753, ZN => n25758);
   U26652 : XNOR2_X1 port map( A => n25754, B => n2510, ZN => n25755);
   U26653 : XNOR2_X1 port map( A => n25756, B => n25755, ZN => n25757);
   U26654 : INV_X1 port map( A => n26322, ZN => n27077);
   U26655 : NOR2_X1 port map( A1 => n27074, A2 => n27077, ZN => n25768);
   U26656 : XNOR2_X1 port map( A => n29155, B => n25819, ZN => n25762);
   U26657 : XNOR2_X1 port map( A => n25760, B => n25761, ZN => n26014);
   U26658 : XNOR2_X1 port map( A => n26014, B => n25762, ZN => n25766);
   U26659 : XNOR2_X1 port map( A => n25445, B => n3673, ZN => n25764);
   U26660 : XNOR2_X1 port map( A => n25763, B => n25764, ZN => n25765);
   U26661 : NOR2_X1 port map( A1 => n26991, A2 => n26989, ZN => n25767);
   U26662 : INV_X1 port map( A => n29623, ZN => n27317);
   U26663 : XNOR2_X1 port map( A => n25772, B => n25771, ZN => n25779);
   U26664 : XNOR2_X1 port map( A => n29634, B => n25773, ZN => n25777);
   U26665 : INV_X1 port map( A => Key(13), ZN => n25774);
   U26666 : XNOR2_X1 port map( A => n25775, B => n25774, ZN => n25776);
   U26667 : XNOR2_X1 port map( A => n25777, B => n25776, ZN => n25778);
   U26668 : XNOR2_X1 port map( A => n25779, B => n25778, ZN => n25815);
   U26669 : XNOR2_X1 port map( A => n25781, B => n25780, ZN => n25784);
   U26670 : XNOR2_X1 port map( A => n25782, B => n1887, ZN => n25783);
   U26671 : XNOR2_X1 port map( A => n25783, B => n25784, ZN => n25789);
   U26672 : XNOR2_X1 port map( A => n25786, B => n25785, ZN => n25787);
   U26673 : XNOR2_X1 port map( A => n26034, B => n25787, ZN => n25788);
   U26674 : XNOR2_X1 port map( A => n25789, B => n25788, ZN => n27018);
   U26676 : XNOR2_X1 port map( A => n25790, B => n26039, ZN => n26076);
   U26677 : XNOR2_X1 port map( A => n26076, B => n25791, ZN => n25805);
   U26678 : INV_X1 port map( A => n25797, ZN => n25792);
   U26679 : NAND2_X1 port map( A1 => n25792, A2 => n3644, ZN => n25801);
   U26680 : INV_X1 port map( A => n25793, ZN => n25796);
   U26681 : NOR2_X1 port map( A1 => n25794, A2 => n3644, ZN => n25795);
   U26682 : NAND2_X1 port map( A1 => n25796, A2 => n25795, ZN => n25799);
   U26683 : INV_X1 port map( A => n3644, ZN => n26257);
   U26684 : NAND2_X1 port map( A1 => n25797, A2 => n26257, ZN => n25798);
   U26685 : OAI211_X1 port map( C1 => n25801, C2 => n25800, A => n25799, B => 
                           n25798, ZN => n25802);
   U26686 : XNOR2_X1 port map( A => n25803, B => n25802, ZN => n25804);
   U26687 : MUX2_X1 port map( A => n25815, B => n28640, S => n26841, Z => 
                           n25814);
   U26688 : XNOR2_X1 port map( A => n25806, B => n25807, ZN => n25813);
   U26689 : XNOR2_X1 port map( A => n25809, B => n25808, ZN => n26116);
   U26690 : XNOR2_X1 port map( A => n25810, B => n3317, ZN => n25811);
   U26691 : XNOR2_X1 port map( A => n26116, B => n25811, ZN => n25812);
   U26692 : NOR2_X1 port map( A1 => n26841, A2 => n27086, ZN => n25833);
   U26693 : XNOR2_X1 port map( A => n26011, B => n2541, ZN => n25818);
   U26694 : XNOR2_X1 port map( A => n25818, B => n25817, ZN => n25824);
   U26695 : XNOR2_X1 port map( A => n25820, B => n25819, ZN => n25822);
   U26696 : XNOR2_X1 port map( A => n25821, B => n25822, ZN => n25823);
   U26697 : NOR2_X1 port map( A1 => n26507, A2 => n26840, ZN => n25832);
   U26698 : XNOR2_X1 port map( A => n25825, B => n26909, ZN => n25827);
   U26699 : XNOR2_X1 port map( A => n25826, B => n25827, ZN => n25829);
   U26700 : XNOR2_X1 port map( A => n25829, B => n25828, ZN => n25831);
   U26701 : XNOR2_X1 port map( A => n25831, B => n25830, ZN => n27081);
   U26702 : INV_X1 port map( A => n27081, ZN => n26842);
   U26703 : XNOR2_X1 port map( A => n26070, B => n25836, ZN => n25838);
   U26704 : XNOR2_X1 port map( A => n25838, B => n25837, ZN => n25842);
   U26705 : XNOR2_X1 port map( A => n25839, B => n25840, ZN => n25841);
   U26706 : XNOR2_X1 port map( A => n25133, B => n363, ZN => n25847);
   U26707 : XNOR2_X1 port map( A => n26114, B => n25845, ZN => n25846);
   U26708 : XNOR2_X1 port map( A => n25846, B => n25847, ZN => n25854);
   U26709 : XNOR2_X1 port map( A => n25849, B => n25848, ZN => n25852);
   U26710 : XNOR2_X1 port map( A => n29046, B => n72, ZN => n25851);
   U26711 : XNOR2_X1 port map( A => n25852, B => n25851, ZN => n25853);
   U26712 : NOR2_X1 port map( A1 => n27120, A2 => n26837, ZN => n26516);
   U26713 : XNOR2_X1 port map( A => n25856, B => n25857, ZN => n25862);
   U26714 : XNOR2_X1 port map( A => n25858, B => n3554, ZN => n25860);
   U26715 : XNOR2_X1 port map( A => n25859, B => n25860, ZN => n25861);
   U26717 : XNOR2_X1 port map( A => n29534, B => n300, ZN => n25866);
   U26718 : XNOR2_X1 port map( A => n25864, B => n25922, ZN => n25865);
   U26719 : XNOR2_X1 port map( A => n25866, B => n25865, ZN => n25873);
   U26720 : XNOR2_X1 port map( A => n25868, B => n25867, ZN => n25871);
   U26721 : XNOR2_X1 port map( A => n25869, B => n27643, ZN => n25870);
   U26722 : XNOR2_X1 port map( A => n25871, B => n25870, ZN => n25872);
   U26723 : XNOR2_X1 port map( A => n25873, B => n25872, ZN => n26835);
   U26724 : XNOR2_X1 port map( A => n25875, B => n25874, ZN => n25880);
   U26725 : XNOR2_X1 port map( A => n25876, B => n3386, ZN => n25878);
   U26726 : XNOR2_X1 port map( A => n25878, B => n25877, ZN => n25879);
   U26727 : XNOR2_X1 port map( A => n25880, B => n25879, ZN => n27121);
   U26728 : NAND2_X1 port map( A1 => n6951, A2 => n27121, ZN => n25883);
   U26729 : NAND2_X1 port map( A1 => n28631, A2 => n28437, ZN => n25881);
   U26730 : INV_X1 port map( A => n27121, ZN => n26334);
   U26731 : NAND2_X1 port map( A1 => n25881, A2 => n26334, ZN => n25882);
   U26732 : OAI21_X1 port map( B1 => n26516, B2 => n25883, A => n25882, ZN => 
                           n25896);
   U26733 : XNOR2_X1 port map( A => n25928, B => n25884, ZN => n25888);
   U26734 : XNOR2_X1 port map( A => n29073, B => n25885, ZN => n25887);
   U26735 : XNOR2_X1 port map( A => n25888, B => n25887, ZN => n25895);
   U26736 : XNOR2_X1 port map( A => n25890, B => n29053, ZN => n25893);
   U26737 : XNOR2_X1 port map( A => n25891, B => n2403, ZN => n25892);
   U26738 : XNOR2_X1 port map( A => n25893, B => n25892, ZN => n25894);
   U26739 : XNOR2_X1 port map( A => n25895, B => n25894, ZN => n26512);
   U26740 : NAND2_X1 port map( A1 => n27118, A2 => n26512, ZN => n26302);
   U26741 : NAND2_X1 port map( A1 => n25896, A2 => n26302, ZN => n27862);
   U26742 : XNOR2_X1 port map( A => n25898, B => n25899, ZN => n25907);
   U26743 : XNOR2_X1 port map( A => n25901, B => n25900, ZN => n25905);
   U26744 : XNOR2_X1 port map( A => n25903, B => n25902, ZN => n25904);
   U26745 : XNOR2_X1 port map( A => n25905, B => n25904, ZN => n25906);
   U26746 : XNOR2_X1 port map( A => n28771, B => n3219, ZN => n25912);
   U26747 : XNOR2_X1 port map( A => n25910, B => n25909, ZN => n25911);
   U26748 : XNOR2_X1 port map( A => n25912, B => n25911, ZN => n25918);
   U26749 : XNOR2_X1 port map( A => n29039, B => n25914, ZN => n25916);
   U26750 : XNOR2_X1 port map( A => n25915, B => n25916, ZN => n25917);
   U26751 : XNOR2_X1 port map( A => n25920, B => n25919, ZN => n25926);
   U26752 : XNOR2_X1 port map( A => n25921, B => n27462, ZN => n25924);
   U26753 : XNOR2_X1 port map( A => n25924, B => n25923, ZN => n25925);
   U26754 : XNOR2_X1 port map( A => n25926, B => n25925, ZN => n26848);
   U26755 : XNOR2_X1 port map( A => n25927, B => n25928, ZN => n25930);
   U26756 : XNOR2_X1 port map( A => n25929, B => n25930, ZN => n25937);
   U26757 : XNOR2_X1 port map( A => n25932, B => n25931, ZN => n25935);
   U26758 : XNOR2_X1 port map( A => n25933, B => n3650, ZN => n25934);
   U26759 : XNOR2_X1 port map( A => n25935, B => n25934, ZN => n25936);
   U26760 : AOI22_X1 port map( A1 => n26510, A2 => n26849, B1 => n26848, B2 => 
                           n27056, ZN => n26301);
   U26761 : INV_X1 port map( A => n26850, ZN => n27898);
   U26762 : XNOR2_X1 port map( A => n25939, B => n25938, ZN => n25941);
   U26763 : XNOR2_X1 port map( A => n25943, B => n25944, ZN => n25946);
   U26764 : XNOR2_X1 port map( A => n25946, B => n25945, ZN => n25952);
   U26765 : INV_X1 port map( A => n2527, ZN => n27915);
   U26766 : XNOR2_X1 port map( A => n25948, B => n27915, ZN => n25949);
   U26767 : XNOR2_X1 port map( A => n25950, B => n25949, ZN => n25951);
   U26768 : XNOR2_X2 port map( A => n25952, B => n25951, ZN => n27902);
   U26770 : OAI21_X1 port map( B1 => n26849, B2 => n29536, A => n26852, ZN => 
                           n25953);
   U26771 : MUX2_X1 port map( A => n27865, B => n27872, S => n27871, Z => 
                           n25954);
   U26772 : XNOR2_X1 port map( A => n25955, B => n6016, ZN => Ciphertext(147));
   U26773 : OAI21_X1 port map( B1 => n27358, B2 => n27354, A => n29052, ZN => 
                           n25956);
   U26774 : NAND2_X1 port map( A1 => n27355, A2 => n27354, ZN => n27330);
   U26775 : MUX2_X1 port map( A => n27357, B => n25956, S => n27330, Z => 
                           n25959);
   U26776 : NOR2_X1 port map( A1 => n27340, A2 => n27357, ZN => n27328);
   U26777 : NAND2_X1 port map( A1 => n25959, A2 => n25958, ZN => n25961);
   U26778 : INV_X1 port map( A => n3081, ZN => n25960);
   U26779 : XNOR2_X1 port map( A => n25961, B => n25960, ZN => Ciphertext(4));
   U26780 : NAND2_X1 port map( A1 => n27066, A2 => n25963, ZN => n25966);
   U26781 : NOR2_X1 port map( A1 => n922, A2 => n28452, ZN => n25964);
   U26782 : OR2_X1 port map( A1 => n25964, A2 => n29520, ZN => n25965);
   U26784 : OAI211_X1 port map( C1 => n29524, C2 => n29058, A => n28130, B => 
                           n398, ZN => n25969);
   U26785 : NAND2_X1 port map( A1 => n25970, A2 => n25969, ZN => n28017);
   U26786 : INV_X1 port map( A => n28017, ZN => n28001);
   U26787 : NOR2_X1 port map( A1 => n29482, A2 => n26733, ZN => n26734);
   U26788 : NOR2_X1 port map( A1 => n26997, A2 => n26998, ZN => n28099);
   U26790 : INV_X1 port map( A => n26755, ZN => n26236);
   U26791 : OR2_X1 port map( A1 => n29479, A2 => n28575, ZN => n25973);
   U26792 : AOI21_X1 port map( B1 => n25973, B2 => n25603, A => n26753, ZN => 
                           n25974);
   U26794 : NOR2_X1 port map( A1 => n29099, A2 => n26748, ZN => n25977);
   U26795 : NOR2_X1 port map( A1 => n5035, A2 => n25977, ZN => n25982);
   U26796 : INV_X1 port map( A => n26747, ZN => n26223);
   U26797 : AOI21_X1 port map( B1 => n26223, B2 => n29159, A => n26222, ZN => 
                           n25981);
   U26798 : AOI22_X1 port map( A1 => n26222, A2 => n25979, B1 => n25453, B2 => 
                           n25978, ZN => n25980);
   U26799 : OAI21_X1 port map( B1 => n25982, B2 => n25981, A => n25980, ZN => 
                           n28021);
   U26800 : NOR2_X1 port map( A1 => n26984, A2 => n28021, ZN => n27034);
   U26801 : MUX2_X1 port map( A => n27014, B => n26623, S => n29062, Z => 
                           n25986);
   U26802 : INV_X1 port map( A => n29062, ZN => n25983);
   U26803 : INV_X1 port map( A => n27010, ZN => n27053);
   U26804 : NOR2_X1 port map( A1 => n28446, A2 => n27053, ZN => n25984);
   U26805 : NOR2_X1 port map( A1 => n27017, A2 => n25984, ZN => n25985);
   U26806 : NAND2_X1 port map( A1 => n27034, A2 => n28019, ZN => n25989);
   U26807 : NOR2_X1 port map( A1 => n28019, A2 => n28411, ZN => n25987);
   U26808 : NAND2_X1 port map( A1 => n25987, A2 => n28003, ZN => n25988);
   U26809 : NAND3_X1 port map( A1 => n25990, A2 => n25989, A3 => n25988, ZN => 
                           n25993);
   U26810 : XNOR2_X1 port map( A => n25993, B => n25992, ZN => Ciphertext(170))
                           ;
   U26811 : INV_X1 port map( A => n27371, ZN => n26497);
   U26812 : INV_X1 port map( A => n26808, ZN => n25994);
   U26813 : XNOR2_X1 port map( A => n25996, B => n857, ZN => Ciphertext(7));
   U26814 : NOR2_X1 port map( A1 => n29538, A2 => n28562, ZN => n25999);
   U26815 : NOR2_X1 port map( A1 => n25994, A2 => n27371, ZN => n27365);
   U26816 : AOI22_X1 port map( A1 => n25999, A2 => n27362, B1 => n27365, B2 => 
                           n27368, ZN => n26001);
   U26817 : NAND2_X1 port map( A1 => n27366, A2 => n27368, ZN => n26000);
   U26818 : INV_X1 port map( A => n3622, ZN => n26003);
   U26819 : XNOR2_X1 port map( A => n26004, B => n26214, ZN => n26005);
   U26820 : XNOR2_X1 port map( A => n26006, B => n26005, ZN => n26010);
   U26821 : INV_X1 port map( A => n27155, ZN => n26018);
   U26822 : XNOR2_X1 port map( A => n26011, B => n4029, ZN => n26012);
   U26823 : XNOR2_X1 port map( A => n26013, B => n26012, ZN => n26017);
   U26824 : XNOR2_X1 port map( A => n26014, B => n26015, ZN => n26016);
   U26825 : XNOR2_X1 port map( A => n26016, B => n26017, ZN => n26867);
   U26826 : INV_X1 port map( A => n26867, ZN => n27153);
   U26827 : NOR2_X1 port map( A1 => n26018, A2 => n27153, ZN => n26052);
   U26828 : XNOR2_X1 port map( A => n26020, B => n26019, ZN => n26022);
   U26829 : XNOR2_X1 port map( A => n26021, B => n26022, ZN => n26027);
   U26830 : XNOR2_X1 port map( A => n26023, B => n27452, ZN => n26024);
   U26831 : XNOR2_X1 port map( A => n26025, B => n26024, ZN => n26026);
   U26832 : XNOR2_X1 port map( A => n28534, B => n26029, ZN => n26031);
   U26833 : XNOR2_X1 port map( A => n26030, B => n26031, ZN => n26037);
   U26834 : XNOR2_X1 port map( A => n25386, B => n26032, ZN => n26035);
   U26835 : XNOR2_X1 port map( A => n26034, B => n26035, ZN => n26036);
   U26836 : XNOR2_X1 port map( A => n26037, B => n26036, ZN => n26868);
   U26838 : XNOR2_X1 port map( A => n26039, B => n26038, ZN => n26043);
   U26839 : XNOR2_X1 port map( A => n26041, B => n26040, ZN => n26042);
   U26841 : XNOR2_X1 port map( A => n28475, B => n3003, ZN => n26048);
   U26842 : XNOR2_X1 port map( A => n26046, B => n26045, ZN => n26047);
   U26843 : XNOR2_X1 port map( A => n26047, B => n26048, ZN => n26049);
   U26845 : XNOR2_X1 port map( A => n26054, B => n26053, ZN => n26058);
   U26846 : XNOR2_X1 port map( A => n29613, B => n26055, ZN => n26057);
   U26847 : XNOR2_X1 port map( A => n26057, B => n26058, ZN => n26064);
   U26848 : XNOR2_X1 port map( A => n26084, B => n26059, ZN => n26062);
   U26849 : XNOR2_X1 port map( A => n26060, B => n2889, ZN => n26061);
   U26850 : XNOR2_X1 port map( A => n26062, B => n26061, ZN => n26063);
   U26852 : NOR2_X1 port map( A1 => n29474, A2 => n29048, ZN => n26066);
   U26856 : NOR2_X1 port map( A1 => n26067, A2 => n26867, ZN => n26068);
   U26857 : INV_X1 port map( A => n27728, ZN => n26126);
   U26858 : XNOR2_X1 port map( A => n26071, B => n26070, ZN => n26075);
   U26859 : INV_X1 port map( A => n28693, ZN => n26072);
   U26860 : XNOR2_X1 port map( A => n29129, B => n26072, ZN => n26074);
   U26861 : XNOR2_X1 port map( A => n26075, B => n26074, ZN => n26079);
   U26862 : XNOR2_X1 port map( A => n26080, B => n3482, ZN => n26082);
   U26863 : XNOR2_X1 port map( A => n26082, B => n26081, ZN => n26088);
   U26864 : XNOR2_X1 port map( A => n26084, B => n26083, ZN => n26085);
   U26865 : XNOR2_X1 port map( A => n26086, B => n26085, ZN => n26087);
   U26866 : XNOR2_X1 port map( A => n300, B => n26089, ZN => n26092);
   U26867 : XNOR2_X1 port map( A => n26091, B => n26092, ZN => n26099);
   U26868 : XNOR2_X1 port map( A => n26094, B => n26093, ZN => n26097);
   U26869 : INV_X1 port map( A => n2385, ZN => n27887);
   U26870 : XNOR2_X1 port map( A => n26095, B => n27887, ZN => n26096);
   U26871 : XNOR2_X1 port map( A => n26097, B => n26096, ZN => n26098);
   U26872 : INV_X1 port map( A => n27137, ZN => n26858);
   U26874 : XNOR2_X1 port map( A => n26105, B => n26104, ZN => n26518);
   U26875 : XNOR2_X1 port map( A => n1871, B => n26108, ZN => n26112);
   U26876 : XNOR2_X1 port map( A => n26110, B => n27788, ZN => n26111);
   U26877 : XNOR2_X1 port map( A => n26112, B => n26111, ZN => n26113);
   U26878 : XNOR2_X1 port map( A => n26114, B => n26115, ZN => n26117);
   U26879 : XNOR2_X1 port map( A => n26117, B => n26116, ZN => n26124);
   U26880 : XNOR2_X1 port map( A => n29543, B => n26118, ZN => n26122);
   U26881 : INV_X1 port map( A => n2465, ZN => n28050);
   U26882 : XNOR2_X1 port map( A => n26120, B => n28050, ZN => n26121);
   U26883 : XNOR2_X1 port map( A => n26122, B => n26121, ZN => n26123);
   U26885 : INV_X1 port map( A => n26518, ZN => n27142);
   U26886 : NOR2_X1 port map( A1 => n26350, A2 => n27704, ZN => n26127);
   U26888 : NOR2_X1 port map( A1 => n27691, A2 => n27707, ZN => n27727);
   U26889 : NAND2_X1 port map( A1 => n6953, A2 => n27727, ZN => n26148);
   U26890 : INV_X1 port map( A => n27178, ZN => n27129);
   U26891 : NOR2_X1 port map( A1 => n27175, A2 => n28536, ZN => n26130);
   U26892 : OAI21_X1 port map( B1 => n26130, B2 => n28392, A => n27178, ZN => 
                           n26131);
   U26893 : INV_X1 port map( A => n26386, ZN => n26132);
   U26894 : NOR2_X1 port map( A1 => n26260, A2 => n26133, ZN => n26137);
   U26896 : AND2_X1 port map( A1 => n26384, A2 => n1907, ZN => n26135);
   U26897 : OAI21_X1 port map( B1 => n27171, B2 => n26135, A => n28535, ZN => 
                           n26136);
   U26899 : NAND2_X1 port map( A1 => n27193, A2 => n28595, ZN => n26139);
   U26900 : MUX2_X1 port map( A => n26139, B => n26138, S => n27123, Z => 
                           n26144);
   U26901 : NOR3_X1 port map( A1 => n27193, A2 => n4109, A3 => n27124, ZN => 
                           n26142);
   U26902 : NOR2_X1 port map( A1 => n26140, A2 => n28595, ZN => n26141);
   U26906 : NOR2_X1 port map( A1 => n26576, A2 => n26789, ZN => n26924);
   U26907 : NAND2_X1 port map( A1 => n26924, A2 => n26791, ZN => n26154);
   U26911 : INV_X1 port map( A => n26458, ZN => n26461);
   U26912 : NOR2_X1 port map( A1 => n26461, A2 => n28578, ZN => n26562);
   U26913 : NAND2_X1 port map( A1 => n28578, A2 => n26457, ZN => n26157);
   U26914 : NAND3_X1 port map( A1 => n26157, A2 => n26560, A3 => n28434, ZN => 
                           n26158);
   U26916 : INV_X1 port map( A => n27460, ZN => n27467);
   U26917 : INV_X1 port map( A => n26455, ZN => n26161);
   U26919 : INV_X1 port map( A => n26454, ZN => n26177);
   U26920 : NOR2_X1 port map( A1 => n29105, A2 => n26454, ZN => n26163);
   U26921 : OAI21_X1 port map( B1 => n26163, B2 => n26162, A => n29467, ZN => 
                           n26164);
   U26922 : OAI21_X1 port map( B1 => n27465, B2 => n27467, A => n29468, ZN => 
                           n26170);
   U26923 : AND2_X1 port map( A1 => n28435, A2 => n27463, ZN => n27236);
   U26924 : INV_X1 port map( A => n26914, ZN => n26568);
   U26925 : MUX2_X1 port map( A => n29610, B => n26568, S => n26567, Z => 
                           n26169);
   U26926 : NOR2_X1 port map( A1 => n5625, A2 => n26786, ZN => n26168);
   U26927 : INV_X1 port map( A => n27457, ZN => n27235);
   U26928 : AOI22_X1 port map( A1 => n26170, A2 => n27458, B1 => n27236, B2 => 
                           n27235, ZN => n26175);
   U26929 : NAND2_X1 port map( A1 => n26920, A2 => n4820, ZN => n26171);
   U26930 : INV_X1 port map( A => n26782, ZN => n26174);
   U26931 : NOR2_X1 port map( A1 => n27457, A2 => n27447, ZN => n26606);
   U26932 : NOR2_X1 port map( A1 => n26180, A2 => n26476, ZN => n26184);
   U26933 : NOR2_X1 port map( A1 => n26181, A2 => n28503, ZN => n26183);
   U26934 : MUX2_X1 port map( A => n26184, B => n26183, S => n28547, Z => 
                           n26190);
   U26936 : NAND3_X1 port map( A1 => n28561, A2 => n28503, A3 => n28525, ZN => 
                           n26187);
   U26937 : OAI21_X1 port map( B1 => n29596, B2 => n26475, A => n26187, ZN => 
                           n26189);
   U26938 : NAND2_X1 port map( A1 => n26464, A2 => n26191, ZN => n26193);
   U26939 : AOI21_X1 port map( B1 => n26193, B2 => n26192, A => n27395, ZN => 
                           n26197);
   U26940 : AND3_X1 port map( A1 => n28908, A2 => n280, A3 => n26469, ZN => 
                           n26196);
   U26941 : MUX2_X1 port map( A => n28560, B => n26728, S => n26729, Z => 
                           n26198);
   U26942 : NAND2_X1 port map( A1 => n26198, A2 => n1622, ZN => n26199);
   U26943 : NAND3_X1 port map( A1 => n26200, A2 => n26204, A3 => n26737, ZN => 
                           n26207);
   U26944 : NOR2_X1 port map( A1 => n26204, A2 => n26235, ZN => n26201);
   U26945 : NAND2_X1 port map( A1 => n26201, A2 => n1874, ZN => n26206);
   U26946 : NAND2_X1 port map( A1 => n28473, A2 => n1874, ZN => n26234);
   U26947 : NAND3_X1 port map( A1 => n26204, A2 => n26203, A3 => n26740, ZN => 
                           n26205);
   U26948 : AND4_X1 port map( A1 => n26207, A2 => n26206, A3 => n26234, A4 => 
                           n26205, ZN => n27379);
   U26949 : INV_X1 port map( A => n26217, ZN => n26213);
   U26950 : AND2_X1 port map( A1 => n26715, A2 => n26718, ZN => n26216);
   U26951 : NAND2_X1 port map( A1 => n26216, A2 => n26208, ZN => n26212);
   U26953 : AOI21_X1 port map( B1 => n283, B2 => n28459, A => n26215, ZN => 
                           n26219);
   U26955 : NOR2_X1 port map( A1 => n26222, A2 => n5760, ZN => n26221);
   U26956 : AOI21_X1 port map( B1 => n26223, B2 => n26222, A => n26221, ZN => 
                           n26226);
   U26957 : INV_X1 port map( A => n29100, ZN => n26224);
   U26959 : INV_X1 port map( A => n28069, ZN => n26227);
   U26960 : NAND2_X1 port map( A1 => n26231, A2 => n26234, ZN => n26232);
   U26961 : NAND2_X1 port map( A1 => n26236, A2 => n26757, ZN => n26239);
   U26962 : MUX2_X1 port map( A => n26239, B => n26238, S => n26753, Z => 
                           n26244);
   U26963 : AND2_X1 port map( A1 => n28575, A2 => n26240, ZN => n26758);
   U26964 : AOI22_X1 port map( A1 => n26242, A2 => n26761, B1 => n26758, B2 => 
                           n26241, ZN => n26243);
   U26965 : INV_X1 port map( A => n27014, ZN => n27049);
   U26966 : NAND2_X1 port map( A1 => n29062, A2 => n27049, ZN => n26245);
   U26967 : NAND2_X1 port map( A1 => n26246, A2 => n26245, ZN => n26249);
   U26968 : OAI21_X1 port map( B1 => n27053, B2 => n399, A => n28639, ZN => 
                           n26248);
   U26969 : NOR2_X1 port map( A1 => n27010, A2 => n27050, ZN => n26247);
   U26970 : NOR3_X1 port map( A1 => n28543, A2 => n28065, A3 => n28063, ZN => 
                           n26250);
   U26971 : AOI21_X1 port map( B1 => n28055, B2 => n28067, A => n26250, ZN => 
                           n26256);
   U26972 : NAND2_X1 port map( A1 => n26632, A2 => n26998, ZN => n26251);
   U26973 : OAI21_X1 port map( B1 => n29481, B2 => n5389, A => n28099, ZN => 
                           n26252);
   U26974 : INV_X1 port map( A => n28066, ZN => n28044);
   U26975 : OAI21_X1 port map( B1 => n28044, B2 => n28063, A => n28069, ZN => 
                           n26254);
   U26976 : NOR2_X1 port map( A1 => n28543, A2 => n28066, ZN => n28053);
   U26977 : NAND2_X1 port map( A1 => n26256, A2 => n26255, ZN => n26258);
   U26978 : XNOR2_X1 port map( A => n26258, B => n26257, ZN => Ciphertext(183))
                           ;
   U26979 : NOR2_X1 port map( A1 => n28535, A2 => n28572, ZN => n26261);
   U26980 : INV_X1 port map( A => n27165, ZN => n27168);
   U26981 : INV_X1 port map( A => n26129, ZN => n27131);
   U26982 : MUX2_X1 port map( A => n29071, B => n26950, S => n26949, Z => 
                           n26269);
   U26983 : MUX2_X1 port map( A => n26267, B => n26948, S => n26952, Z => 
                           n26268);
   U26985 : AOI21_X1 port map( B1 => n1901, B2 => n27585, A => n28179, ZN => 
                           n26286);
   U26986 : OAI21_X1 port map( B1 => n28650, B2 => n27183, A => n26270, ZN => 
                           n26271);
   U26987 : NAND2_X1 port map( A1 => n26271, A2 => n26397, ZN => n26274);
   U26988 : AND3_X1 port map( A1 => n28651, A2 => n27181, A3 => n25124, ZN => 
                           n26272);
   U26989 : AOI21_X1 port map( B1 => n28652, B2 => n26357, A => n26272, ZN => 
                           n26273);
   U26990 : MUX2_X2 port map( A => n26277, B => n26276, S => n26361, Z => 
                           n27596);
   U26991 : NAND2_X1 port map( A1 => n26798, A2 => n26362, ZN => n26804);
   U26992 : INV_X1 port map( A => n26392, ZN => n26279);
   U26994 : AOI22_X1 port map( A1 => n26279, A2 => n28470, B1 => n26800, B2 => 
                           n29573, ZN => n26282);
   U26995 : OR3_X1 port map( A1 => n26798, A2 => n26280, A3 => n26799, ZN => 
                           n26281);
   U26996 : OAI211_X1 port map( C1 => n29573, C2 => n26804, A => n26282, B => 
                           n26281, ZN => n27590);
   U26997 : INV_X1 port map( A => n27590, ZN => n26284);
   U26998 : NOR2_X1 port map( A1 => n26284, A2 => n27586, ZN => n26285);
   U26999 : INV_X1 port map( A => n2598, ZN => n26288);
   U27000 : MUX2_X1 port map( A => n28487, B => n29621, S => n27137, Z => 
                           n26289);
   U27001 : AND2_X1 port map( A1 => n29621, A2 => n27141, ZN => n26326);
   U27002 : INV_X1 port map( A => n26290, ZN => n26291);
   U27003 : INV_X1 port map( A => n26292, ZN => n26293);
   U27004 : NOR2_X1 port map( A1 => n29070, A2 => n27768, ZN => n27782);
   U27005 : NAND2_X1 port map( A1 => n27700, A2 => n27702, ZN => n26297);
   U27006 : NAND2_X1 port map( A1 => n26350, A2 => n27704, ZN => n26296);
   U27007 : INV_X1 port map( A => n27161, ZN => n26352);
   U27008 : OAI21_X1 port map( B1 => n400, B2 => n26352, A => n455, ZN => 
                           n26295);
   U27009 : NOR2_X1 port map( A1 => n27782, A2 => n26298, ZN => n26315);
   U27011 : AOI21_X1 port map( B1 => n27902, B2 => n26848, A => n28600, ZN => 
                           n26300);
   U27012 : NAND2_X1 port map( A1 => n26315, A2 => n29537, ZN => n26313);
   U27013 : INV_X1 port map( A => n26302, ZN => n26305);
   U27014 : INV_X1 port map( A => n27120, ZN => n26303);
   U27015 : NOR2_X1 port map( A1 => n26303, A2 => n27121, ZN => n26304);
   U27016 : MUX2_X1 port map( A => n26305, B => n26304, S => n26837, Z => 
                           n26308);
   U27017 : INV_X1 port map( A => n26512, ZN => n27117);
   U27018 : MUX2_X1 port map( A => n28631, B => n402, S => n27117, Z => n26306)
                           ;
   U27019 : NOR2_X1 port map( A1 => n26306, A2 => n29016, ZN => n26307);
   U27020 : NOR2_X1 port map( A1 => n26308, A2 => n26307, ZN => n27762);
   U27021 : INV_X1 port map( A => n27111, ZN => n27154);
   U27022 : AOI21_X1 port map( B1 => n27110, B2 => n27154, A => n26865, ZN => 
                           n26311);
   U27023 : NOR2_X1 port map( A1 => n27762, A2 => n27777, ZN => n27771);
   U27025 : OAI21_X1 port map( B1 => n26317, B2 => n2441, A => n26316, ZN => 
                           n26318);
   U27026 : NOR2_X1 port map( A1 => n26319, A2 => n26318, ZN => Ciphertext(122)
                           );
   U27027 : INV_X1 port map( A => n27074, ZN => n26321);
   U27028 : INV_X1 port map( A => n26989, ZN => n26320);
   U27029 : MUX2_X1 port map( A => n26989, B => n26323, S => n27074, Z => 
                           n26324);
   U27031 : INV_X1 port map( A => n27140, ZN => n26855);
   U27032 : NOR2_X1 port map( A1 => n29621, A2 => n27137, ZN => n26325);
   U27033 : NAND2_X1 port map( A1 => n27136, A2 => n26326, ZN => n26327);
   U27034 : NOR2_X1 port map( A1 => n29232, A2 => n27807, ZN => n26339);
   U27035 : INV_X1 port map( A => n27902, ZN => n27836);
   U27036 : AND2_X1 port map( A1 => n27902, A2 => n27898, ZN => n26511);
   U27037 : AOI21_X1 port map( B1 => n26510, B2 => n27836, A => n26511, ZN => 
                           n26329);
   U27038 : NOR2_X1 port map( A1 => n29497, A2 => n26848, ZN => n26328);
   U27042 : NOR2_X1 port map( A1 => n27155, A2 => n26867, ZN => n27151);
   U27043 : NAND2_X1 port map( A1 => n27154, A2 => n27155, ZN => n27109);
   U27044 : NOR2_X1 port map( A1 => n29060, A2 => n26865, ZN => n26332);
   U27046 : INV_X1 port map( A => n27118, ZN => n26836);
   U27047 : AND2_X1 port map( A1 => n26837, A2 => n27117, ZN => n26333);
   U27048 : NAND2_X1 port map( A1 => n26516, A2 => n26334, ZN => n26335);
   U27049 : AOI22_X1 port map( A1 => n26339, A2 => n27800, B1 => n27819, B2 => 
                           n27812, ZN => n26341);
   U27051 : OAI21_X1 port map( B1 => n27795, B2 => n29469, A => n27818, ZN => 
                           n26338);
   U27052 : INV_X1 port map( A => n27807, ZN => n27821);
   U27053 : INV_X1 port map( A => n27791, ZN => n26344);
   U27054 : NAND2_X1 port map( A1 => n27800, A2 => n28403, ZN => n26343);
   U27055 : AND2_X1 port map( A1 => n27819, A2 => n27818, ZN => n26342);
   U27056 : AOI22_X1 port map( A1 => n27823, A2 => n26344, B1 => n26343, B2 => 
                           n26342, ZN => n26345);
   U27057 : XNOR2_X1 port map( A => n26345, B => n3673, ZN => Ciphertext(127));
   U27058 : MUX2_X1 port map( A => n27597, B => n26346, S => n27596, Z => 
                           n26348);
   U27059 : NOR2_X1 port map( A1 => n27582, A2 => n27594, ZN => n27265);
   U27060 : AND2_X1 port map( A1 => n27582, A2 => n27590, ZN => n27593);
   U27061 : NOR2_X1 port map( A1 => n27265, A2 => n27593, ZN => n26347);
   U27063 : XNOR2_X1 port map( A => n26349, B => n1079, ZN => Ciphertext(86));
   U27066 : NAND2_X1 port map( A1 => n26397, A2 => n27181, ZN => n26401);
   U27067 : NAND2_X1 port map( A1 => n26357, A2 => n26356, ZN => n27188);
   U27069 : MUX2_X1 port map( A => n27183, B => n25124, S => n27181, Z => 
                           n26359);
   U27070 : INV_X1 port map( A => n28650, ZN => n26358);
   U27071 : INV_X1 port map( A => n27630, ZN => n27619);
   U27072 : AND2_X1 port map( A1 => n26427, A2 => n26381, ZN => n26432);
   U27073 : MUX2_X1 port map( A => n26798, B => n26362, S => n26799, Z => 
                           n26365);
   U27075 : OR2_X1 port map( A1 => n26799, A2 => n26280, ZN => n26363);
   U27076 : OAI22_X1 port map( A1 => n27626, A2 => n27619, B1 => n27627, B2 => 
                           n27632, ZN => n27610);
   U27077 : NAND2_X1 port map( A1 => n27175, A2 => n27177, ZN => n27134);
   U27078 : NAND2_X1 port map( A1 => n27129, A2 => n29132, ZN => n26366);
   U27080 : AOI21_X1 port map( B1 => n27165, B2 => n26384, A => n28572, ZN => 
                           n26367);
   U27081 : INV_X1 port map( A => n26367, ZN => n26369);
   U27082 : NOR2_X1 port map( A1 => n26385, A2 => n27168, ZN => n26368);
   U27083 : INV_X1 port map( A => n27625, ZN => n27613);
   U27084 : OAI21_X1 port map( B1 => n27627, B2 => n27613, A => n3366, ZN => 
                           n26370);
   U27085 : AOI22_X1 port map( A1 => n27610, A2 => n27628, B1 => n26370, B2 => 
                           n27619, ZN => n26371);
   U27086 : XNOR2_X1 port map( A => n26371, B => n3232, ZN => Ciphertext(95));
   U27087 : NOR2_X1 port map( A1 => n28646, A2 => n26775, ZN => n26373);
   U27088 : AOI21_X1 port map( B1 => n26949, B2 => n26440, A => n26952, ZN => 
                           n26372);
   U27090 : INV_X1 port map( A => n27571, ZN => n27552);
   U27091 : NAND2_X1 port map( A1 => n26935, A2 => n26936, ZN => n26376);
   U27092 : AOI21_X1 port map( B1 => n26772, B2 => n26376, A => n26943, ZN => 
                           n26377);
   U27093 : MUX2_X1 port map( A => n26382, B => n26426, S => n26378, Z => 
                           n26379);
   U27095 : OAI21_X1 port map( B1 => n28573, B2 => n27165, A => n27166, ZN => 
                           n26390);
   U27096 : OAI21_X1 port map( B1 => n26387, B2 => n1907, A => n26385, ZN => 
                           n26389);
   U27097 : AOI22_X2 port map( A1 => n27169, A2 => n26390, B1 => n26389, B2 => 
                           n28573, ZN => n27562);
   U27098 : OAI21_X1 port map( B1 => n28470, B2 => n26797, A => n29573, ZN => 
                           n26410);
   U27099 : NAND2_X1 port map( A1 => n26392, A2 => n26799, ZN => n26394);
   U27100 : NOR2_X1 port map( A1 => n26800, A2 => n29573, ZN => n26413);
   U27101 : MUX2_X1 port map( A => n26394, B => n26280, S => n26413, Z => 
                           n26395);
   U27102 : AOI21_X1 port map( B1 => n28651, B2 => n26396, A => n25124, ZN => 
                           n26402);
   U27103 : NAND3_X1 port map( A1 => n26397, A2 => n28650, A3 => n27182, ZN => 
                           n26398);
   U27104 : OAI21_X1 port map( B1 => n26399, B2 => n25034, A => n26398, ZN => 
                           n26400);
   U27105 : NAND2_X1 port map( A1 => n27561, A2 => n27562, ZN => n27567);
   U27106 : NAND2_X1 port map( A1 => n27572, A2 => n27567, ZN => n26403);
   U27107 : OAI21_X1 port map( B1 => n27149, B2 => n29085, A => n26403, ZN => 
                           n26404);
   U27109 : XNOR2_X1 port map( A => n26406, B => n1062, ZN => Ciphertext(80));
   U27110 : NAND2_X1 port map( A1 => n28035, A2 => n28038, ZN => n28037);
   U27111 : NOR2_X1 port map( A1 => n29161, A2 => n29032, ZN => n28028);
   U27112 : INV_X1 port map( A => n28028, ZN => n26408);
   U27113 : INV_X1 port map( A => n3372, ZN => n26409);
   U27114 : INV_X1 port map( A => n26410, ZN => n26414);
   U27115 : AND2_X1 port map( A1 => n26280, A2 => n29330, ZN => n26412);
   U27116 : NOR3_X1 port map( A1 => n26414, A2 => n26413, A3 => n26412, ZN => 
                           n26417);
   U27117 : MUX2_X1 port map( A => n26799, B => n26798, S => n26797, Z => 
                           n26415);
   U27118 : NOR2_X1 port map( A1 => n26415, A2 => n26800, ZN => n26416);
   U27120 : NAND2_X1 port map( A1 => n26565, A2 => n26420, ZN => n26418);
   U27121 : OAI21_X1 port map( B1 => n29610, B2 => n1872, A => n26418, ZN => 
                           n26419);
   U27122 : NOR2_X1 port map( A1 => n26419, A2 => n26914, ZN => n27305);
   U27123 : NOR2_X1 port map( A1 => n26565, A2 => n26911, ZN => n26421);
   U27124 : NOR2_X2 port map( A1 => n27305, A2 => n27304, ZN => n27308);
   U27125 : INV_X1 port map( A => n26920, ZN => n26422);
   U27126 : OAI21_X1 port map( B1 => n26172, B2 => n26919, A => n26422, ZN => 
                           n26424);
   U27127 : NAND2_X1 port map( A1 => n26782, A2 => n454, ZN => n26423);
   U27128 : MUX2_X1 port map( A => n26424, B => n26423, S => n4820, Z => n27302
                           );
   U27129 : NAND2_X1 port map( A1 => n26917, A2 => n26919, ZN => n27303);
   U27130 : NAND2_X1 port map( A1 => n27302, A2 => n27303, ZN => n26879);
   U27132 : NAND2_X1 port map( A1 => n26430, A2 => n26429, ZN => n26434);
   U27133 : NAND2_X1 port map( A1 => n26432, A2 => n4679, ZN => n26433);
   U27134 : INV_X1 port map( A => n26936, ZN => n26435);
   U27135 : NAND3_X1 port map( A1 => n28541, A2 => n26943, A3 => n26768, ZN => 
                           n26437);
   U27136 : OAI22_X1 port map( A1 => n27308, A2 => n28510, B1 => n29493, B2 => 
                           n27301, ZN => n26887);
   U27137 : INV_X1 port map( A => n26952, ZN => n26439);
   U27138 : MUX2_X1 port map( A => n26439, B => n26440, S => n28542, Z => 
                           n26444);
   U27139 : NAND2_X1 port map( A1 => n28646, A2 => n26439, ZN => n26441);
   U27140 : MUX2_X1 port map( A => n26442, B => n26441, S => n26440, Z => 
                           n26443);
   U27144 : XNOR2_X1 port map( A => n26446, B => n3386, ZN => Ciphertext(71));
   U27145 : NAND2_X1 port map( A1 => n29105, A2 => n26451, ZN => n26453);
   U27146 : NOR2_X1 port map( A1 => n28385, A2 => n26457, ZN => n26460);
   U27147 : NAND2_X1 port map( A1 => n26464, A2 => n26466, ZN => n26465);
   U27148 : OAI21_X1 port map( B1 => n28908, B2 => n280, A => n26465, ZN => 
                           n26468);
   U27149 : INV_X1 port map( A => n26468, ZN => n26470);
   U27150 : MUX2_X2 port map( A => n26471, B => n26470, S => n26469, Z => 
                           n27429);
   U27151 : MUX2_X1 port map( A => n29542, B => n27426, S => n27429, Z => 
                           n26494);
   U27152 : NOR2_X1 port map( A1 => n26472, A2 => n28503, ZN => n26473);
   U27153 : NOR2_X1 port map( A1 => n26474, A2 => n26473, ZN => n26479);
   U27154 : AND3_X1 port map( A1 => n28561, A2 => n26477, A3 => n26475, ZN => 
                           n26478);
   U27155 : NOR2_X2 port map( A1 => n26479, A2 => n26478, ZN => n27428);
   U27156 : NAND3_X1 port map( A1 => n26482, A2 => n28560, A3 => n26480, ZN => 
                           n26488);
   U27157 : NOR2_X1 port map( A1 => n26482, A2 => n26727, ZN => n26483);
   U27158 : NOR2_X1 port map( A1 => n26927, A2 => n25364, ZN => n26582);
   U27159 : NOR2_X1 port map( A1 => n26489, A2 => n26933, ZN => n26490);
   U27160 : NOR2_X1 port map( A1 => n26582, A2 => n26490, ZN => n26493);
   U27161 : OAI21_X1 port map( B1 => n26928, B2 => n26933, A => n26927, ZN => 
                           n26492);
   U27162 : NOR2_X1 port map( A1 => n28477, A2 => n26933, ZN => n26491);
   U27163 : OAI22_X2 port map( A1 => n26493, A2 => n26581, B1 => n26492, B2 => 
                           n26491, ZN => n27425);
   U27164 : XNOR2_X1 port map( A => n26495, B => n3191, ZN => Ciphertext(26));
   U27165 : NOR2_X1 port map( A1 => n27366, A2 => n29541, ZN => n26498);
   U27168 : NAND2_X1 port map( A1 => n29075, A2 => n27063, ZN => n26501);
   U27169 : INV_X1 port map( A => n27088, ZN => n26506);
   U27171 : NOR2_X1 port map( A1 => n28458, A2 => n27085, ZN => n26504);
   U27172 : NOR2_X1 port map( A1 => n27086, A2 => n26840, ZN => n26503);
   U27173 : NOR2_X1 port map( A1 => n26504, A2 => n26503, ZN => n26505);
   U27174 : NOR2_X1 port map( A1 => n26841, A2 => n28640, ZN => n26509);
   U27175 : AND2_X1 port map( A1 => n27085, A2 => n26840, ZN => n26508);
   U27176 : NOR3_X1 port map( A1 => n27852, A2 => n26638, A3 => n26639, ZN => 
                           n27849);
   U27178 : NAND2_X1 port map( A1 => n27849, A2 => n447, ZN => n26525);
   U27179 : NOR2_X1 port map( A1 => n402, A2 => n28631, ZN => n26513);
   U27180 : OAI21_X1 port map( B1 => n26334, B2 => n28437, A => n26513, ZN => 
                           n26515);
   U27181 : NOR2_X1 port map( A1 => n27136, A2 => n29621, ZN => n26857);
   U27182 : AND2_X1 port map( A1 => n27137, A2 => n27141, ZN => n26517);
   U27183 : OAI21_X1 port map( B1 => n26857, B2 => n26517, A => n27147, ZN => 
                           n26521);
   U27184 : OAI21_X1 port map( B1 => n26519, B2 => n27138, A => n27139, ZN => 
                           n26520);
   U27185 : INV_X1 port map( A => n26641, ZN => n27851);
   U27186 : AOI21_X1 port map( B1 => n27855, B2 => n27851, A => n27847, ZN => 
                           n26522);
   U27187 : OAI21_X1 port map( B1 => n27855, B2 => n5295, A => n26522, ZN => 
                           n26524);
   U27188 : NAND2_X1 port map( A1 => n27855, A2 => n6907, ZN => n26523);
   U27189 : INV_X1 port map( A => n27425, ZN => n27418);
   U27192 : INV_X1 port map( A => n26669, ZN => n26529);
   U27193 : INV_X1 port map( A => n26531, ZN => n26528);
   U27194 : INV_X1 port map( A => n27426, ZN => n26668);
   U27195 : AND2_X1 port map( A1 => n27424, A2 => n27428, ZN => n26530);
   U27196 : OAI21_X1 port map( B1 => n26668, B2 => n27425, A => n26530, ZN => 
                           n26532);
   U27197 : AND3_X1 port map( A1 => n26529, A2 => n26528, A3 => n26532, ZN => 
                           n26536);
   U27198 : NAND2_X1 port map( A1 => n27429, A2 => n27425, ZN => n27417);
   U27202 : OAI21_X1 port map( B1 => n27875, B2 => n27866, A => n3378, ZN => 
                           n26538);
   U27203 : INV_X1 port map( A => n26538, ZN => n26543);
   U27205 : INV_X1 port map( A => n27864, ZN => n26540);
   U27206 : NAND3_X1 port map( A1 => n27875, A2 => n27872, A3 => n26540, ZN => 
                           n26542);
   U27207 : NAND3_X1 port map( A1 => n27872, A2 => n27873, A3 => n27864, ZN => 
                           n26541);
   U27208 : NAND4_X1 port map( A1 => n26544, A2 => n26543, A3 => n26542, A4 => 
                           n26541, ZN => n26551);
   U27209 : AOI22_X1 port map( A1 => n27317, A2 => n27313, B1 => n27864, B2 => 
                           n27862, ZN => n26548);
   U27210 : INV_X1 port map( A => n27872, ZN => n26595);
   U27211 : AOI21_X1 port map( B1 => n26595, B2 => n27875, A => n3378, ZN => 
                           n26547);
   U27212 : INV_X1 port map( A => n27327, ZN => n26546);
   U27213 : NAND3_X1 port map( A1 => n26548, A2 => n26547, A3 => n26546, ZN => 
                           n26549);
   U27214 : AND3_X1 port map( A1 => n26551, A2 => n26550, A3 => n26549, ZN => 
                           Ciphertext(146));
   U27215 : AND2_X1 port map( A1 => n26920, A2 => n26782, ZN => n26554);
   U27216 : MUX2_X1 port map( A => n26554, B => n26553, S => n454, Z => n26557)
                           ;
   U27217 : MUX2_X1 port map( A => n4820, B => n26920, S => n26782, Z => n26555
                           );
   U27218 : NOR2_X1 port map( A1 => n26917, A2 => n26555, ZN => n26556);
   U27219 : NOR2_X2 port map( A1 => n26557, A2 => n26556, ZN => n27492);
   U27220 : AND2_X1 port map( A1 => n26560, A2 => n26559, ZN => n26561);
   U27221 : OAI21_X1 port map( B1 => n26563, B2 => n377, A => n28482, ZN => 
                           n26564);
   U27222 : NAND2_X1 port map( A1 => n26568, A2 => n1872, ZN => n26566);
   U27223 : NOR3_X1 port map( A1 => n26568, A2 => n26567, A3 => n26786, ZN => 
                           n26569);
   U27224 : AOI21_X1 port map( B1 => n26788, B2 => n5625, A => n26569, ZN => 
                           n26570);
   U27227 : OR2_X1 port map( A1 => n26791, A2 => n26575, ZN => n26922);
   U27228 : NOR2_X1 port map( A1 => n29552, A2 => n26922, ZN => n26577);
   U27229 : NAND3_X1 port map( A1 => n27492, A2 => n29093, A3 => n27497, ZN => 
                           n26589);
   U27230 : NAND2_X1 port map( A1 => n26928, A2 => n29054, ZN => n26586);
   U27231 : NOR2_X1 port map( A1 => n28477, A2 => n26928, ZN => n26584);
   U27232 : NAND2_X1 port map( A1 => n26581, A2 => n29054, ZN => n26583);
   U27233 : AOI21_X1 port map( B1 => n26584, B2 => n26583, A => n26582, ZN => 
                           n26585);
   U27234 : OAI21_X1 port map( B1 => n26933, B2 => n26586, A => n26585, ZN => 
                           n27493);
   U27235 : INV_X1 port map( A => n27493, ZN => n26965);
   U27236 : NOR2_X1 port map( A1 => n29522, A2 => n26965, ZN => n26587);
   U27237 : NAND2_X1 port map( A1 => n27492, A2 => n26587, ZN => n26588);
   U27238 : INV_X1 port map( A => n3483, ZN => n26590);
   U27239 : INV_X1 port map( A => n2404, ZN => n26592);
   U27240 : XNOR2_X1 port map( A => n26593, B => n26592, ZN => Ciphertext(32));
   U27241 : NOR2_X1 port map( A1 => n27873, A2 => n27872, ZN => n27311);
   U27242 : INV_X1 port map( A => n27311, ZN => n26600);
   U27243 : NAND3_X1 port map( A1 => n27872, A2 => n27877, A3 => n27863, ZN => 
                           n26599);
   U27244 : NAND2_X1 port map( A1 => n26595, A2 => n26594, ZN => n26598);
   U27245 : INV_X1 port map( A => n27877, ZN => n26596);
   U27247 : NOR2_X1 port map( A1 => n28035, A2 => n29032, ZN => n28026);
   U27248 : INV_X1 port map( A => n26602, ZN => n28030);
   U27249 : MUX2_X1 port map( A => n29032, B => n29160, S => n28025, Z => 
                           n26603);
   U27250 : INV_X1 port map( A => n3770, ZN => n26604);
   U27251 : MUX2_X1 port map( A => n27465, B => n27447, S => n28435, Z => 
                           n26608);
   U27254 : XNOR2_X1 port map( A => n26609, B => n440, ZN => Ciphertext(45));
   U27255 : INV_X1 port map( A => n27379, ZN => n27377);
   U27256 : OAI21_X1 port map( B1 => n27209, B2 => n28393, A => n27377, ZN => 
                           n26613);
   U27257 : OAI21_X1 port map( B1 => n5581, B2 => n446, A => n27379, ZN => 
                           n26612);
   U27258 : NOR2_X1 port map( A1 => n295, A2 => n27382, ZN => n26611);
   U27259 : NOR2_X1 port map( A1 => n26614, A2 => n28452, ZN => n26615);
   U27260 : NAND2_X1 port map( A1 => n26616, A2 => n26615, ZN => n26619);
   U27261 : NOR2_X1 port map( A1 => n28545, A2 => n29520, ZN => n26617);
   U27262 : NAND2_X1 port map( A1 => n26617, A2 => n27066, ZN => n26618);
   U27263 : MUX2_X1 port map( A => n26841, B => n27085, S => n27018, Z => 
                           n26622);
   U27264 : NOR2_X1 port map( A1 => n27018, A2 => n25815, ZN => n26620);
   U27265 : MUX2_X1 port map( A => n26840, B => n26620, S => n26842, Z => 
                           n26621);
   U27266 : NOR2_X1 port map( A1 => n27050, A2 => n27014, ZN => n26625);
   U27268 : MUX2_X1 port map( A => n26995, B => n29481, S => n28532, Z => 
                           n26631);
   U27270 : NOR2_X1 port map( A1 => n26632, A2 => n26998, ZN => n26628);
   U27274 : INV_X1 port map( A => n29095, ZN => n26640);
   U27275 : NAND2_X1 port map( A1 => n6907, A2 => n26640, ZN => n26644);
   U27276 : XNOR2_X1 port map( A => n26645, B => n2804, ZN => Ciphertext(142));
   U27277 : OR2_X1 port map( A1 => n29095, A2 => n27847, ZN => n27858);
   U27278 : NAND2_X1 port map( A1 => n27851, A2 => n27854, ZN => n26646);
   U27279 : AOI21_X1 port map( B1 => n27636, B2 => n27641, A => n27639, ZN => 
                           n26649);
   U27280 : OAI22_X1 port map( A1 => n29532, A2 => n27641, B1 => n26978, B2 => 
                           n26980, ZN => n27649);
   U27281 : INV_X1 port map( A => n27641, ZN => n26648);
   U27282 : AOI22_X1 port map( A1 => n26649, A2 => n27637, B1 => n27649, B2 => 
                           n26979, ZN => n26650);
   U27283 : XNOR2_X1 port map( A => n26650, B => n3256, ZN => Ciphertext(97));
   U27284 : NOR2_X1 port map( A1 => n27202, A2 => n27203, ZN => n26651);
   U27285 : AOI21_X1 port map( B1 => n27539, B2 => n27202, A => n26651, ZN => 
                           n26655);
   U27286 : NOR2_X1 port map( A1 => n27549, A2 => n27203, ZN => n27541);
   U27287 : NOR2_X1 port map( A1 => n27539, A2 => n28468, ZN => n26653);
   U27288 : OAI21_X1 port map( B1 => n26655, B2 => n27547, A => n26654, ZN => 
                           n26657);
   U27289 : XNOR2_X1 port map( A => n26657, B => n26656, ZN => Ciphertext(75));
   U27290 : INV_X1 port map( A => n26658, ZN => n26662);
   U27291 : INV_X1 port map( A => n26659, ZN => n26660);
   U27292 : AND2_X1 port map( A1 => n28038, A2 => n26660, ZN => n26661);
   U27293 : NAND3_X1 port map( A1 => n28036, A2 => n29160, A3 => n28025, ZN => 
                           n26663);
   U27294 : OAI21_X1 port map( B1 => n26664, B2 => n28026, A => n26663, ZN => 
                           n26666);
   U27295 : XNOR2_X1 port map( A => n26666, B => n630, ZN => Ciphertext(175));
   U27296 : INV_X1 port map( A => n27427, ZN => n27430);
   U27297 : OAI21_X1 port map( B1 => n27428, B2 => n29542, A => n27430, ZN => 
                           n26667);
   U27298 : AOI22_X1 port map( A1 => n26669, A2 => n26668, B1 => n27429, B2 => 
                           n26667, ZN => n26670);
   U27299 : XNOR2_X1 port map( A => n26670, B => n2996, ZN => Ciphertext(29));
   U27300 : NAND2_X1 port map( A1 => n26978, A2 => n27641, ZN => n26673);
   U27301 : OAI22_X1 port map( A1 => n26979, A2 => n27636, B1 => n26673, B2 => 
                           n27638, ZN => n26674);
   U27302 : NOR2_X1 port map( A1 => n26675, A2 => n26674, ZN => n26676);
   U27303 : XNOR2_X1 port map( A => n26676, B => n2577, ZN => Ciphertext(99));
   U27305 : INV_X1 port map( A => n27818, ZN => n27790);
   U27306 : INV_X1 port map( A => n27800, ZN => n27822);
   U27307 : INV_X1 port map( A => n26680, ZN => n26681);
   U27308 : INV_X1 port map( A => n26830, ZN => n27438);
   U27309 : INV_X1 port map( A => n27442, ZN => n26831);
   U27310 : OAI21_X1 port map( B1 => n27442, B2 => n26710, A => n25417, ZN => 
                           n26683);
   U27311 : NAND2_X1 port map( A1 => n26683, A2 => n27439, ZN => n26684);
   U27312 : XNOR2_X1 port map( A => n26685, B => n633, ZN => Ciphertext(36));
   U27313 : NOR2_X1 port map( A1 => n27308, A2 => n27300, ZN => n27310);
   U27314 : NOR2_X1 port map( A1 => n27310, A2 => n29493, ZN => n26687);
   U27315 : NAND2_X1 port map( A1 => n26687, A2 => n26686, ZN => n26688);
   U27316 : OAI21_X1 port map( B1 => n26689, B2 => n26880, A => n26688, ZN => 
                           n26690);
   U27317 : XNOR2_X1 port map( A => n26690, B => n3369, ZN => Ciphertext(68));
   U27318 : NAND2_X1 port map( A1 => n27025, A2 => n29588, ZN => n26691);
   U27319 : NOR2_X1 port map( A1 => n26692, A2 => n27025, ZN => n26693);
   U27320 : NOR2_X1 port map( A1 => n26694, A2 => n26693, ZN => n26695);
   U27321 : XNOR2_X1 port map( A => n26695, B => n3607, ZN => Ciphertext(30));
   U27322 : NOR2_X1 port map( A1 => n27859, A2 => n27847, ZN => n26697);
   U27323 : AOI21_X1 port map( B1 => n29095, B2 => n26697, A => n26696, ZN => 
                           n26700);
   U27324 : NAND3_X1 port map( A1 => n27855, A2 => n29095, A3 => n27854, ZN => 
                           n26699);
   U27325 : OAI211_X1 port map( C1 => n27855, C2 => n27858, A => n26700, B => 
                           n26699, ZN => n26702);
   U27326 : XNOR2_X1 port map( A => n26702, B => n26701, ZN => Ciphertext(138))
                           ;
   U27327 : NAND2_X1 port map( A1 => n29093, A2 => n27497, ZN => n27478);
   U27328 : INV_X1 port map( A => n3586, ZN => n26703);
   U27329 : XNOR2_X1 port map( A => n26704, B => n26703, ZN => Ciphertext(51));
   U27330 : OAI21_X1 port map( B1 => n27025, B2 => n26817, A => n27032, ZN => 
                           n26706);
   U27332 : NOR2_X1 port map( A1 => n27439, A2 => n26708, ZN => n26709);
   U27333 : AOI21_X1 port map( B1 => n26830, B2 => n27439, A => n26709, ZN => 
                           n27435);
   U27334 : NOR2_X1 port map( A1 => n27433, A2 => n26710, ZN => n26828);
   U27335 : AOI22_X1 port map( A1 => n26831, A2 => n26833, B1 => n26828, B2 => 
                           n27438, ZN => n26711);
   U27336 : OAI21_X1 port map( B1 => n26712, B2 => n27435, A => n26711, ZN => 
                           n26714);
   U27337 : XNOR2_X1 port map( A => n26714, B => n26713, ZN => Ciphertext(39));
   U27338 : NOR2_X1 port map( A1 => n26716, A2 => n28459, ZN => n26720);
   U27340 : NOR3_X1 port map( A1 => n26723, A2 => n28548, A3 => n29560, ZN => 
                           n26724);
   U27342 : OAI21_X1 port map( B1 => n29579, B2 => n26727, A => n26726, ZN => 
                           n26732);
   U27343 : NOR2_X1 port map( A1 => n28115, A2 => n28794, ZN => n28094);
   U27345 : MUX2_X1 port map( A => n26742, B => n26741, S => n26740, Z => 
                           n26743);
   U27348 : AOI21_X1 port map( B1 => n29159, B2 => n26747, A => n28563, ZN => 
                           n26752);
   U27349 : AND2_X1 port map( A1 => n29159, A2 => n26748, ZN => n26751);
   U27350 : MUX2_X1 port map( A => n26752, B => n26751, S => n29099, Z => 
                           n28103);
   U27351 : INV_X1 port map( A => n28089, ZN => n28112);
   U27352 : AOI21_X1 port map( B1 => n28591, B2 => n28112, A => n29056, ZN => 
                           n26763);
   U27353 : NAND2_X1 port map( A1 => n26758, A2 => n26757, ZN => n26759);
   U27355 : NAND3_X1 port map( A1 => n28107, A2 => n28590, A3 => n29121, ZN => 
                           n26762);
   U27356 : OAI21_X1 port map( B1 => n26764, B2 => n26763, A => n26762, ZN => 
                           n26766);
   U27357 : INV_X1 port map( A => n3491, ZN => n26765);
   U27358 : XNOR2_X1 port map( A => n26766, B => n26765, ZN => Ciphertext(186))
                           ;
   U27359 : MUX2_X1 port map( A => n26935, B => n26768, S => n26936, Z => 
                           n26767);
   U27360 : NOR2_X1 port map( A1 => n26767, A2 => n28541, ZN => n26774);
   U27363 : NOR2_X2 port map( A1 => n26774, A2 => n26773, ZN => n27275);
   U27364 : MUX2_X1 port map( A => n26950, B => n26775, S => n29071, Z => 
                           n26779);
   U27365 : NOR2_X1 port map( A1 => n26949, A2 => n26775, ZN => n26777);
   U27366 : NOR2_X1 port map( A1 => n26948, A2 => n28542, ZN => n26776);
   U27367 : MUX2_X1 port map( A => n26777, B => n26776, S => n26950, Z => 
                           n26778);
   U27368 : AOI21_X2 port map( B1 => n26948, B2 => n26779, A => n26778, ZN => 
                           n27291);
   U27369 : NOR2_X1 port map( A1 => n457, A2 => n26920, ZN => n26780);
   U27370 : NOR2_X1 port map( A1 => n26781, A2 => n26780, ZN => n26784);
   U27371 : MUX2_X1 port map( A => n26782, B => n4820, S => n26920, Z => n26783
                           );
   U27372 : MUX2_X1 port map( A => n27275, B => n27291, S => n27282, Z => 
                           n26806);
   U27373 : NAND2_X1 port map( A1 => n28471, A2 => n26911, ZN => n26785);
   U27374 : AND3_X1 port map( A1 => n26914, A2 => n5625, A3 => n26786, ZN => 
                           n26787);
   U27375 : NOR2_X1 port map( A1 => n25418, A2 => n26789, ZN => n26790);
   U27379 : MUX2_X1 port map( A => n27286, B => n27287, S => n27275, Z => 
                           n26805);
   U27383 : XNOR2_X1 port map( A => n26807, B => n3414, ZN => Ciphertext(62));
   U27384 : XNOR2_X1 port map( A => n26810, B => n3244, ZN => Ciphertext(11));
   U27385 : INV_X1 port map( A => n27277, ZN => n27288);
   U27386 : NOR2_X1 port map( A1 => n27282, A2 => n27288, ZN => n26812);
   U27388 : NOR2_X1 port map( A1 => n26812, A2 => n26811, ZN => n26897);
   U27389 : INV_X1 port map( A => n27275, ZN => n27290);
   U27390 : AOI21_X1 port map( B1 => n27280, B2 => n27290, A => n27287, ZN => 
                           n26813);
   U27391 : OAI22_X1 port map( A1 => n26897, A2 => n27291, B1 => n27278, B2 => 
                           n26813, ZN => n26815);
   U27392 : XNOR2_X1 port map( A => n26815, B => n26814, ZN => Ciphertext(65));
   U27393 : NOR2_X1 port map( A1 => n27032, A2 => n306, ZN => n26818);
   U27394 : NAND2_X1 port map( A1 => n27025, A2 => n26818, ZN => n26820);
   U27395 : INV_X1 port map( A => n3728, ZN => n26821);
   U27396 : MUX2_X1 port map( A => n27354, B => n29052, S => n27357, Z => 
                           n26824);
   U27397 : NAND2_X1 port map( A1 => n27358, A2 => n28549, ZN => n26822);
   U27398 : MUX2_X1 port map( A => n26822, B => n27348, S => n27357, Z => 
                           n26823);
   U27399 : OAI21_X1 port map( B1 => n26824, B2 => n27355, A => n26823, ZN => 
                           n26826);
   U27400 : XNOR2_X1 port map( A => n26826, B => n26825, ZN => Ciphertext(2));
   U27401 : NOR2_X1 port map( A1 => n25417, A2 => n26830, ZN => n26827);
   U27402 : NOR2_X1 port map( A1 => n26828, A2 => n26827, ZN => n27443);
   U27403 : OAI211_X1 port map( C1 => n26831, C2 => n27434, A => n26830, B => 
                           n26829, ZN => n26832);
   U27405 : XNOR2_X1 port map( A => n26834, B => n5892, ZN => Ciphertext(37));
   U27406 : MUX2_X1 port map( A => n27117, B => n26835, S => n28631, Z => 
                           n26839);
   U27407 : MUX2_X1 port map( A => n27121, B => n26836, S => n27120, Z => 
                           n26838);
   U27408 : INV_X1 port map( A => n27843, ZN => n26846);
   U27409 : OAI21_X1 port map( B1 => n26842, B2 => n25815, A => n26840, ZN => 
                           n26843);
   U27410 : NAND2_X1 port map( A1 => n26843, A2 => n27088, ZN => n26844);
   U27412 : OAI21_X1 port map( B1 => n26849, B2 => n29575, A => n29497, ZN => 
                           n26853);
   U27413 : OAI21_X1 port map( B1 => n26853, B2 => n26852, A => n26851, ZN => 
                           n26854);
   U27414 : AOI21_X1 port map( B1 => n27137, B2 => n27138, A => n26855, ZN => 
                           n26856);
   U27415 : NOR2_X1 port map( A1 => n26857, A2 => n26856, ZN => n27830);
   U27416 : NAND2_X1 port map( A1 => n28487, A2 => n26858, ZN => n26859);
   U27417 : NOR2_X1 port map( A1 => n26860, A2 => n26859, ZN => n27829);
   U27418 : MUX2_X1 port map( A => n27074, B => n27076, S => n26991, Z => 
                           n26864);
   U27419 : NAND2_X1 port map( A1 => n26992, A2 => n27076, ZN => n26861);
   U27420 : MUX2_X1 port map( A => n26862, B => n26861, S => n27074, Z => 
                           n26863);
   U27421 : OAI21_X1 port map( B1 => n26864, B2 => n28521, A => n26863, ZN => 
                           n27826);
   U27422 : NAND2_X1 port map( A1 => n26866, A2 => n26865, ZN => n27834);
   U27423 : NAND2_X1 port map( A1 => n26867, A2 => n29048, ZN => n26871);
   U27424 : INV_X1 port map( A => n26868, ZN => n27159);
   U27426 : OAI21_X1 port map( B1 => n27155, B2 => n29060, A => n27154, ZN => 
                           n26869);
   U27427 : OAI21_X1 port map( B1 => n26871, B2 => n26870, A => n26869, ZN => 
                           n27831);
   U27428 : NAND2_X1 port map( A1 => n27834, A2 => n27831, ZN => n27841);
   U27429 : AOI21_X1 port map( B1 => n27826, B2 => n27827, A => n27841, ZN => 
                           n26872);
   U27430 : XNOR2_X1 port map( A => n26873, B => n625, ZN => Ciphertext(132));
   U27431 : MUX2_X1 port map( A => n27825, B => n27101, S => n27100, Z => 
                           n26876);
   U27432 : NAND2_X1 port map( A1 => n26902, A2 => n27826, ZN => n26874);
   U27433 : OAI211_X1 port map( C1 => n26876, C2 => n27828, A => n26875, B => 
                           n26874, ZN => n26878);
   U27434 : XNOR2_X1 port map( A => n26878, B => n26877, ZN => Ciphertext(135))
                           ;
   U27435 : NOR2_X1 port map( A1 => n27300, A2 => n26879, ZN => n26886);
   U27436 : OAI21_X1 port map( B1 => n26880, B2 => n28510, A => n444, ZN => 
                           n26883);
   U27437 : OAI211_X1 port map( C1 => n26886, C2 => n26883, A => n26882, B => 
                           n26881, ZN => n26884);
   U27438 : XNOR2_X1 port map( A => n26884, B => n6174, ZN => Ciphertext(69));
   U27439 : NAND2_X1 port map( A1 => n29493, A2 => n27255, ZN => n26885);
   U27440 : XNOR2_X1 port map( A => n26888, B => n3336, ZN => Ciphertext(67));
   U27441 : INV_X1 port map( A => n27727, ZN => n26894);
   U27442 : INV_X1 port map( A => n326, ZN => n27715);
   U27443 : OAI21_X1 port map( B1 => n27714, B2 => n27715, A => n26889, ZN => 
                           n26893);
   U27444 : NOR2_X1 port map( A1 => n324, A2 => n27728, ZN => n27681);
   U27445 : NOR2_X1 port map( A1 => n27725, A2 => n27711, ZN => n26890);
   U27446 : AOI22_X1 port map( A1 => n27691, A2 => n27681, B1 => n325, B2 => 
                           n26890, ZN => n26892);
   U27447 : NAND2_X1 port map( A1 => n27681, A2 => n27707, ZN => n26891);
   U27448 : NAND2_X1 port map( A1 => n27282, A2 => n27277, ZN => n27285);
   U27449 : INV_X1 port map( A => n27285, ZN => n26898);
   U27450 : INV_X1 port map( A => n27291, ZN => n26895);
   U27451 : OAI211_X1 port map( C1 => n26895, C2 => n27277, A => n27275, B => 
                           n27286, ZN => n26896);
   U27452 : OAI21_X1 port map( B1 => n26898, B2 => n26897, A => n26896, ZN => 
                           n26900);
   U27453 : XNOR2_X1 port map( A => n26900, B => n26899, ZN => Ciphertext(61));
   U27454 : INV_X1 port map( A => n27841, ZN => n26901);
   U27455 : INV_X1 port map( A => n26902, ZN => n26905);
   U27456 : AND2_X1 port map( A1 => n27101, A2 => n27100, ZN => n26904);
   U27457 : NOR2_X1 port map( A1 => n27826, A2 => n27827, ZN => n27102);
   U27458 : INV_X1 port map( A => n27102, ZN => n26903);
   U27459 : AOI22_X1 port map( A1 => n26905, A2 => n27249, B1 => n26904, B2 => 
                           n26903, ZN => n26906);
   U27460 : XNOR2_X1 port map( A => n26906, B => n3374, ZN => Ciphertext(133));
   U27461 : NAND2_X1 port map( A1 => n27235, A2 => n27447, ZN => n26908);
   U27462 : INV_X1 port map( A => n27447, ZN => n27472);
   U27463 : INV_X1 port map( A => n26909, ZN => n26910);
   U27464 : MUX2_X1 port map( A => n26911, B => n28423, S => n28471, Z => 
                           n26916);
   U27465 : INV_X1 port map( A => n27531, ZN => n27506);
   U27466 : NAND2_X1 port map( A1 => n26922, A2 => n26921, ZN => n26923);
   U27467 : OAI21_X1 port map( B1 => n26925, B2 => n26924, A => n26923, ZN => 
                           n27528);
   U27468 : INV_X1 port map( A => n27528, ZN => n27502);
   U27469 : AOI22_X1 port map( A1 => n26928, A2 => n5505, B1 => n26927, B2 => 
                           n1279, ZN => n26932);
   U27470 : INV_X1 port map( A => n26929, ZN => n26931);
   U27471 : MUX2_X1 port map( A => n26932, B => n26931, S => n26930, Z => 
                           n26934);
   U27472 : OAI21_X1 port map( B1 => n27520, B2 => n27502, A => n27527, ZN => 
                           n26958);
   U27473 : AND2_X1 port map( A1 => n6768, A2 => n26935, ZN => n26939);
   U27474 : NOR2_X1 port map( A1 => n6768, A2 => n26936, ZN => n26938);
   U27475 : OAI21_X1 port map( B1 => n26939, B2 => n26938, A => n28541, ZN => 
                           n26946);
   U27476 : NOR2_X1 port map( A1 => n28541, A2 => n26940, ZN => n26942);
   U27478 : INV_X1 port map( A => n26950, ZN => n26954);
   U27479 : AOI21_X1 port map( B1 => n29071, B2 => n28542, A => n28646, ZN => 
                           n26953);
   U27481 : NAND3_X1 port map( A1 => n27527, A2 => n27528, A3 => n27525, ZN => 
                           n26956);
   U27482 : OAI21_X1 port map( B1 => n27506, B2 => n27221, A => n26956, ZN => 
                           n26957);
   U27483 : AOI21_X1 port map( B1 => n27506, B2 => n26958, A => n26957, ZN => 
                           n26959);
   U27484 : XNOR2_X1 port map( A => n26959, B => n2544, ZN => Ciphertext(59));
   U27485 : OAI21_X1 port map( B1 => n27386, B2 => n27410, A => n28177, ZN => 
                           n26962);
   U27486 : OAI21_X1 port map( B1 => n27400, B2 => n27387, A => n27390, ZN => 
                           n26961);
   U27488 : NAND2_X1 port map( A1 => n27496, A2 => n27493, ZN => n26964);
   U27489 : OAI21_X1 port map( B1 => n27494, B2 => n27480, A => n26964, ZN => 
                           n27477);
   U27490 : INV_X1 port map( A => n27498, ZN => n27487);
   U27491 : OAI21_X1 port map( B1 => n27487, B2 => n26965, A => n27496, ZN => 
                           n26966);
   U27492 : AOI22_X1 port map( A1 => n5368, A2 => n27477, B1 => n26966, B2 => 
                           n29093, ZN => n26967);
   U27493 : XNOR2_X1 port map( A => n26967, B => n2916, ZN => Ciphertext(53));
   U27494 : OAI21_X1 port map( B1 => n27417, B2 => n27426, A => n26968, ZN => 
                           n26971);
   U27496 : NAND2_X1 port map( A1 => n29529, A2 => n27425, ZN => n26969);
   U27497 : INV_X1 port map( A => n27424, ZN => n27420);
   U27498 : NOR2_X1 port map( A1 => n26971, A2 => n26970, ZN => n26972);
   U27500 : INV_X1 port map( A => n27629, ZN => n26973);
   U27501 : OAI21_X1 port map( B1 => n26973, B2 => n27627, A => n27630, ZN => 
                           n26974);
   U27502 : NOR2_X1 port map( A1 => n27614, A2 => n27625, ZN => n27609);
   U27503 : NAND2_X1 port map( A1 => n1912, A2 => n27632, ZN => n27601);
   U27504 : OAI22_X1 port map( A1 => n26974, A2 => n27609, B1 => n27601, B2 => 
                           n27625, ZN => n26976);
   U27505 : NOR2_X1 port map( A1 => n1912, A2 => n27630, ZN => n27607);
   U27506 : AND2_X1 port map( A1 => n27607, A2 => n27628, ZN => n26975);
   U27507 : NOR2_X1 port map( A1 => n26976, A2 => n26975, ZN => n26977);
   U27508 : XNOR2_X1 port map( A => n26977, B => n2973, ZN => Ciphertext(93));
   U27509 : OAI21_X1 port map( B1 => n27636, B2 => n27641, A => n26978, ZN => 
                           n26982);
   U27510 : OAI21_X1 port map( B1 => n26980, B2 => n27638, A => n26979, ZN => 
                           n26981);
   U27512 : XNOR2_X1 port map( A => n26983, B => Key(173), ZN => Ciphertext(96)
                           );
   U27515 : INV_X1 port map( A => n28021, ZN => n28006);
   U27516 : OAI21_X1 port map( B1 => n28006, B2 => n28003, A => n28015, ZN => 
                           n26985);
   U27517 : AOI22_X1 port map( A1 => n26986, A2 => n28006, B1 => n28411, B2 => 
                           n26985, ZN => n26987);
   U27518 : XNOR2_X1 port map( A => n26987, B => n1919, ZN => Ciphertext(168));
   U27520 : INV_X1 port map( A => n27944, ZN => n27927);
   U27521 : MUX2_X1 port map( A => n29500, B => n27069, S => n28660, Z => 
                           n27000);
   U27522 : MUX2_X1 port map( A => n28452, B => n29076, S => n28545, Z => 
                           n26999);
   U27523 : MUX2_X1 port map( A => n27000, B => n26999, S => n29520, Z => 
                           n27925);
   U27524 : NOR2_X1 port map( A1 => n27004, A2 => n29058, ZN => n27005);
   U27525 : NAND2_X1 port map( A1 => n27005, A2 => n398, ZN => n27008);
   U27526 : AND2_X1 port map( A1 => n28783, A2 => n28130, ZN => n27006);
   U27527 : NAND2_X1 port map( A1 => n27041, A2 => n27006, ZN => n27007);
   U27529 : NOR2_X1 port map( A1 => n26623, A2 => n27014, ZN => n27012);
   U27530 : NOR2_X1 port map( A1 => n27010, A2 => n28639, ZN => n27011);
   U27531 : NAND2_X1 port map( A1 => n29062, A2 => n27013, ZN => n27015);
   U27532 : NAND2_X1 port map( A1 => n27015, A2 => n27014, ZN => n27016);
   U27533 : NOR2_X1 port map( A1 => n26507, A2 => n27018, ZN => n27089);
   U27534 : NOR3_X1 port map( A1 => n27089, A2 => n27086, A3 => n27085, ZN => 
                           n27019);
   U27535 : AOI21_X1 port map( B1 => n27927, B2 => n27023, A => n27022, ZN => 
                           n27024);
   U27536 : XNOR2_X1 port map( A => n27024, B => n3643, ZN => Ciphertext(160));
   U27537 : NOR2_X1 port map( A1 => n27032, A2 => n29588, ZN => n27027);
   U27538 : NAND2_X1 port map( A1 => n27027, A2 => n28592, ZN => n27031);
   U27539 : NOR2_X1 port map( A1 => n6568, A2 => n306, ZN => n27030);
   U27540 : INV_X1 port map( A => n27034, ZN => n27035);
   U27541 : AOI22_X1 port map( A1 => n27035, A2 => n28000, B1 => n28005, B2 => 
                           n28022, ZN => n27036);
   U27542 : XNOR2_X1 port map( A => n27036, B => n2353, ZN => Ciphertext(169));
   U27543 : OAI21_X1 port map( B1 => n27382, B2 => n28393, A => n27379, ZN => 
                           n27037);
   U27544 : XNOR2_X1 port map( A => n27039, B => n3787, ZN => Ciphertext(12));
   U27545 : NAND2_X1 port map( A1 => n27048, A2 => n28130, ZN => n27046);
   U27546 : MUX2_X1 port map( A => n4497, B => n27046, S => n27045, Z => n27047
                           );
   U27548 : AOI21_X1 port map( B1 => n29062, B2 => n26623, A => n27049, ZN => 
                           n27051);
   U27549 : OR2_X1 port map( A1 => n29536, A2 => n27898, ZN => n27058);
   U27550 : OAI211_X1 port map( C1 => n29536, C2 => n27056, A => n27902, B => 
                           n27055, ZN => n27057);
   U27551 : OAI21_X1 port map( B1 => n29497, B2 => n27058, A => n27057, ZN => 
                           n27062);
   U27552 : NOR2_X1 port map( A1 => n27902, A2 => n29575, ZN => n27903);
   U27553 : AND2_X1 port map( A1 => n27903, A2 => n27060, ZN => n27061);
   U27554 : NOR2_X1 port map( A1 => n922, A2 => n27063, ZN => n27064);
   U27555 : NOR2_X1 port map( A1 => n27065, A2 => n27064, ZN => n27073);
   U27556 : INV_X1 port map( A => n27066, ZN => n27072);
   U27557 : NOR2_X1 port map( A1 => n28228, A2 => n28545, ZN => n27071);
   U27558 : NOR2_X1 port map( A1 => n27069, A2 => n29076, ZN => n27070);
   U27559 : OAI211_X1 port map( C1 => n27092, C2 => n27908, A => n27905, B => 
                           n27080, ZN => n27094);
   U27560 : NAND2_X1 port map( A1 => n27077, A2 => n27076, ZN => n27078);
   U27561 : AND2_X1 port map( A1 => n27079, A2 => n27078, ZN => n27899);
   U27563 : INV_X1 port map( A => n28453, ZN => n27918);
   U27564 : OAI21_X1 port map( B1 => n27919, B2 => n27920, A => n27918, ZN => 
                           n27093);
   U27565 : AOI21_X1 port map( B1 => n27084, B2 => n28458, A => n27081, ZN => 
                           n27083);
   U27566 : OAI21_X1 port map( B1 => n27088, B2 => n27084, A => n27083, ZN => 
                           n27091);
   U27567 : OAI21_X1 port map( B1 => n27087, B2 => n27086, A => n27085, ZN => 
                           n27090);
   U27568 : INV_X1 port map( A => n27271, ZN => n27913);
   U27569 : AOI22_X1 port map( A1 => n27094, A2 => n27093, B1 => n27889, B2 => 
                           n27092, ZN => n27095);
   U27570 : XNOR2_X1 port map( A => n27095, B => n3422, ZN => Ciphertext(150));
   U27571 : OAI21_X1 port map( B1 => n27520, B2 => n27528, A => n27096, ZN => 
                           n27097);
   U27572 : XNOR2_X1 port map( A => n27098, B => n3109, ZN => Ciphertext(57));
   U27573 : NAND2_X1 port map( A1 => n27825, A2 => n27099, ZN => n27104);
   U27574 : NAND2_X1 port map( A1 => n27102, A2 => n27828, ZN => n27103);
   U27575 : NAND2_X1 port map( A1 => n27703, A2 => n27161, ZN => n27106);
   U27577 : INV_X1 port map( A => n27755, ZN => n27745);
   U27578 : AOI21_X1 port map( B1 => n27155, B2 => n29474, A => n27152, ZN => 
                           n27116);
   U27579 : INV_X1 port map( A => n27109, ZN => n27115);
   U27580 : NOR2_X1 port map( A1 => n29474, A2 => n27159, ZN => n27113);
   U27581 : NOR2_X1 port map( A1 => n27153, A2 => n29048, ZN => n27112);
   U27583 : NAND2_X1 port map( A1 => n27745, A2 => n29049, ZN => n27227);
   U27584 : AOI21_X1 port map( B1 => n28631, B2 => n402, A => n27117, ZN => 
                           n27119);
   U27585 : INV_X1 port map( A => n27128, ZN => n27732);
   U27586 : MUX2_X1 port map( A => n27124, B => n27123, S => n27193, Z => 
                           n27127);
   U27587 : NAND2_X1 port map( A1 => n27130, A2 => n27175, ZN => n27133);
   U27588 : NAND3_X1 port map( A1 => n27173, A2 => n27131, A3 => n28536, ZN => 
                           n27132);
   U27589 : AOI21_X1 port map( B1 => n27137, B2 => n27142, A => n27136, ZN => 
                           n27145);
   U27590 : NAND2_X1 port map( A1 => n27139, A2 => n27138, ZN => n27144);
   U27591 : NOR3_X1 port map( A1 => n27142, A2 => n28487, A3 => n29621, ZN => 
                           n27143);
   U27592 : AOI21_X1 port map( B1 => n27145, B2 => n27144, A => n27143, ZN => 
                           n27146);
   U27593 : OAI21_X1 port map( B1 => n27690, B2 => n27147, A => n27146, ZN => 
                           n27739);
   U27594 : INV_X1 port map( A => n27739, ZN => n27757);
   U27595 : NOR2_X1 port map( A1 => n27551, A2 => n29085, ZN => n27148);
   U27596 : NOR2_X1 port map( A1 => n27572, A2 => n27562, ZN => n27576);
   U27597 : MUX2_X1 port map( A => n27148, B => n27576, S => n27552, Z => 
                           n27150);
   U27598 : NOR2_X1 port map( A1 => n27561, A2 => n27562, ZN => n27554);
   U27599 : OAI21_X1 port map( B1 => n27155, B2 => n27154, A => n27153, ZN => 
                           n27156);
   U27601 : OR2_X1 port map( A1 => n27704, A2 => n27703, ZN => n27162);
   U27602 : OAI21_X1 port map( B1 => n27169, B2 => n27168, A => n27167, ZN => 
                           n27170);
   U27603 : NOR2_X1 port map( A1 => n28392, A2 => n29132, ZN => n27172);
   U27604 : AOI21_X1 port map( B1 => n28392, B2 => n27173, A => n27172, ZN => 
                           n27180);
   U27605 : MUX2_X1 port map( A => n27177, B => n28536, S => n27175, Z => 
                           n27179);
   U27606 : INV_X1 port map( A => n27661, ZN => n27674);
   U27607 : NAND2_X1 port map( A1 => n26396, A2 => n25124, ZN => n27185);
   U27608 : OAI21_X1 port map( B1 => n27183, B2 => n27182, A => n27181, ZN => 
                           n27184);
   U27609 : OAI21_X1 port map( B1 => n28652, B2 => n27185, A => n27184, ZN => 
                           n27187);
   U27610 : OAI21_X1 port map( B1 => n28650, B2 => n27188, A => n27187, ZN => 
                           n27671);
   U27612 : NOR2_X1 port map( A1 => n27652, A2 => n27676, ZN => n27194);
   U27613 : AOI211_X1 port map( C1 => n27196, C2 => n27674, A => n27195, B => 
                           n27194, ZN => n27197);
   U27614 : XNOR2_X1 port map( A => n27197, B => n3164, ZN => Ciphertext(105));
   U27615 : NAND2_X1 port map( A1 => n27537, A2 => n27202, ZN => n27198);
   U27617 : OAI21_X1 port map( B1 => n27537, B2 => n27538, A => n28386, ZN => 
                           n27201);
   U27618 : NOR2_X1 port map( A1 => n27201, A2 => n27200, ZN => n27207);
   U27619 : NAND2_X1 port map( A1 => n27547, A2 => n27548, ZN => n27205);
   U27621 : NAND2_X1 port map( A1 => n394, A2 => n27203, ZN => n27204);
   U27623 : NOR2_X1 port map( A1 => n295, A2 => n446, ZN => n27211);
   U27624 : AND2_X1 port map( A1 => n27208, A2 => n27379, ZN => n27210);
   U27626 : XNOR2_X1 port map( A => n27215, B => n28693, ZN => Ciphertext(15));
   U27627 : NOR2_X1 port map( A1 => n27572, A2 => n27561, ZN => n27216);
   U27629 : XNOR2_X1 port map( A => n27220, B => n2986, ZN => Ciphertext(82));
   U27630 : NOR3_X1 port map( A1 => n27531, A2 => n27505, A3 => n29556, ZN => 
                           n27224);
   U27631 : INV_X1 port map( A => n27527, ZN => n27222);
   U27632 : NAND2_X1 port map( A1 => n27755, A2 => n397, ZN => n27226);
   U27633 : INV_X1 port map( A => n27759, ZN => n27749);
   U27634 : AOI21_X1 port map( B1 => n27227, B2 => n27226, A => n27749, ZN => 
                           n27230);
   U27636 : NAND2_X1 port map( A1 => n28445, A2 => n27732, ZN => n27228);
   U27637 : XNOR2_X1 port map( A => n27232, B => n27231, ZN => Ciphertext(117))
                           ;
   U27638 : AOI21_X1 port map( B1 => n27762, B2 => n27777, A => n6419, ZN => 
                           n27233);
   U27639 : XNOR2_X1 port map( A => n27234, B => n3180, ZN => Ciphertext(120));
   U27640 : OAI211_X1 port map( C1 => n27235, C2 => n27472, A => n27465, B => 
                           n27467, ZN => n27238);
   U27641 : NAND2_X1 port map( A1 => n27447, A2 => n27236, ZN => n27237);
   U27642 : OAI211_X1 port map( C1 => n27458, C2 => n27447, A => n27238, B => 
                           n27237, ZN => n27240);
   U27643 : INV_X1 port map( A => n2403, ZN => n27239);
   U27644 : XNOR2_X1 port map( A => n27240, B => n27239, ZN => Ciphertext(43));
   U27645 : OAI21_X1 port map( B1 => n27400, B2 => n27386, A => n27241, ZN => 
                           n27243);
   U27646 : INV_X1 port map( A => n27387, ZN => n27242);
   U27647 : MUX2_X1 port map( A => n27246, B => n27245, S => n28441, Z => 
                           n27247);
   U27648 : XNOR2_X1 port map( A => n27247, B => n2981, ZN => Ciphertext(158));
   U27649 : NAND2_X1 port map( A1 => n27248, A2 => n27841, ZN => n27250);
   U27652 : AOI21_X1 port map( B1 => n27278, B2 => n27253, A => n27252, ZN => 
                           n27254);
   U27653 : XNOR2_X1 port map( A => n27254, B => n2511, ZN => Ciphertext(63));
   U27655 : OAI21_X1 port map( B1 => n6910, B2 => n395, A => n29619, ZN => 
                           n27262);
   U27656 : NOR2_X1 port map( A1 => n28510, A2 => n27300, ZN => n27260);
   U27657 : OAI21_X1 port map( B1 => n27260, B2 => n27259, A => n27255, ZN => 
                           n27261);
   U27658 : NAND2_X1 port map( A1 => n27262, A2 => n27261, ZN => n27264);
   U27659 : XNOR2_X1 port map( A => n27264, B => n27263, ZN => Ciphertext(66));
   U27660 : INV_X1 port map( A => n27265, ZN => n27266);
   U27661 : INV_X1 port map( A => n27596, ZN => n27588);
   U27662 : NOR3_X1 port map( A1 => n27588, A2 => n27597, A3 => n27585, ZN => 
                           n27268);
   U27663 : NOR3_X1 port map( A1 => n27596, A2 => n28429, A3 => n28179, ZN => 
                           n27267);
   U27664 : NOR3_X1 port map( A1 => n27269, A2 => n27268, A3 => n27267, ZN => 
                           n27270);
   U27665 : XNOR2_X1 port map( A => n27270, B => n3385, ZN => Ciphertext(88));
   U27666 : INV_X1 port map( A => n27889, ZN => n27273);
   U27667 : OAI22_X1 port map( A1 => n27919, A2 => n27905, B1 => n27923, B2 => 
                           n27908, ZN => n27921);
   U27668 : INV_X1 port map( A => n27919, ZN => n27272);
   U27669 : NOR2_X1 port map( A1 => n27272, A2 => n27080, ZN => n27893);
   U27670 : AOI22_X1 port map( A1 => n27273, A2 => n27921, B1 => n27883, B2 => 
                           n27893, ZN => n27274);
   U27671 : XNOR2_X1 port map( A => n27274, B => Key(126), ZN => 
                           Ciphertext(151));
   U27672 : MUX2_X1 port map( A => n27277, B => n27282, S => n27275, Z => 
                           n27276);
   U27673 : NAND2_X1 port map( A1 => n27276, A2 => n27281, ZN => n27284);
   U27674 : NOR2_X1 port map( A1 => n27291, A2 => n27277, ZN => n27279);
   U27675 : NAND2_X1 port map( A1 => n27279, A2 => n27278, ZN => n27283);
   U27676 : OAI21_X1 port map( B1 => n27286, B2 => n27290, A => n27285, ZN => 
                           n27292);
   U27677 : OAI21_X1 port map( B1 => n27291, B2 => n2438, A => n27287, ZN => 
                           n27289);
   U27678 : AOI22_X1 port map( A1 => n27292, A2 => n27291, B1 => n27290, B2 => 
                           n27289, ZN => n27293);
   U27679 : XNOR2_X1 port map( A => n27293, B => n3451, ZN => Ciphertext(60));
   U27680 : NAND2_X1 port map( A1 => n28655, A2 => n27663, ZN => n27295);
   U27681 : AOI21_X1 port map( B1 => n27676, B2 => n27672, A => n27673, ZN => 
                           n27294);
   U27682 : AOI21_X1 port map( B1 => n29091, B2 => n27295, A => n27294, ZN => 
                           n27297);
   U27683 : INV_X1 port map( A => n27664, ZN => n27668);
   U27684 : NOR2_X1 port map( A1 => n27652, A2 => n28655, ZN => n27296);
   U27685 : NOR3_X1 port map( A1 => n27297, A2 => n27668, A3 => n27296, ZN => 
                           n27299);
   U27686 : XNOR2_X1 port map( A => n27299, B => n27298, ZN => Ciphertext(102))
                           ;
   U27687 : INV_X1 port map( A => n27303, ZN => n27306);
   U27688 : NOR2_X1 port map( A1 => n27317, A2 => n27324, ZN => n27314);
   U27689 : INV_X1 port map( A => n27313, ZN => n27319);
   U27690 : NOR2_X1 port map( A1 => n27875, A2 => n27324, ZN => n27316);
   U27691 : AOI22_X1 port map( A1 => n27314, A2 => n27319, B1 => n27311, B2 => 
                           n27316, ZN => n27326);
   U27692 : NOR3_X1 port map( A1 => n27875, A2 => n3537, A3 => n27871, ZN => 
                           n27312);
   U27693 : NOR2_X1 port map( A1 => n27875, A2 => n27872, ZN => n27315);
   U27694 : OAI21_X1 port map( B1 => n27315, B2 => n3537, A => n27862, ZN => 
                           n27322);
   U27695 : NAND2_X1 port map( A1 => n27316, A2 => n29504, ZN => n27321);
   U27696 : NOR2_X1 port map( A1 => n27317, A2 => n3537, ZN => n27318);
   U27697 : NAND2_X1 port map( A1 => n27319, A2 => n27318, ZN => n27320);
   U27699 : INV_X1 port map( A => n27328, ZN => n27332);
   U27700 : OAI22_X1 port map( A1 => n5421, A2 => n27357, B1 => n27358, B2 => 
                           n27355, ZN => n27329);
   U27701 : NAND2_X1 port map( A1 => n27329, A2 => n27340, ZN => n27331);
   U27702 : OAI211_X1 port map( C1 => n27332, C2 => n27353, A => n27331, B => 
                           n27330, ZN => n27334);
   U27703 : XNOR2_X1 port map( A => n27334, B => n27333, ZN => Ciphertext(0));
   U27704 : AND2_X1 port map( A1 => n27358, A2 => n2522, ZN => n27343);
   U27705 : XNOR2_X1 port map( A => n27354, B => n2522, ZN => n27335);
   U27706 : OAI21_X1 port map( B1 => n27335, B2 => n27358, A => n27357, ZN => 
                           n27336);
   U27707 : AOI21_X1 port map( B1 => n27340, B2 => n27343, A => n27336, ZN => 
                           n27347);
   U27708 : INV_X1 port map( A => n2522, ZN => n27337);
   U27709 : OAI21_X1 port map( B1 => n27358, B2 => n27337, A => n27351, ZN => 
                           n27339);
   U27710 : OR2_X1 port map( A1 => n27351, A2 => n27337, ZN => n27338);
   U27711 : AOI21_X1 port map( B1 => n27339, B2 => n27338, A => n27357, ZN => 
                           n27346);
   U27712 : INV_X1 port map( A => n27340, ZN => n27342);
   U27713 : INV_X1 port map( A => n27357, ZN => n27349);
   U27714 : NOR3_X1 port map( A1 => n27350, A2 => n2522, A3 => n28549, ZN => 
                           n27341);
   U27715 : OAI21_X1 port map( B1 => n27342, B2 => n27349, A => n27341, ZN => 
                           n27345);
   U27716 : OAI211_X1 port map( C1 => n27351, C2 => n27357, A => n27343, B => 
                           n28549, ZN => n27344);
   U27717 : OAI211_X1 port map( C1 => n27347, C2 => n27346, A => n27345, B => 
                           n27344, ZN => Ciphertext(1));
   U27718 : INV_X1 port map( A => n27348, ZN => n27360);
   U27719 : OAI21_X1 port map( B1 => n27351, B2 => n27350, A => n27349, ZN => 
                           n27359);
   U27720 : NOR2_X1 port map( A1 => n27354, A2 => n28549, ZN => n27356);
   U27721 : XNOR2_X1 port map( A => n27361, B => n629, ZN => Ciphertext(3));
   U27722 : AOI211_X1 port map( C1 => n29541, C2 => n27362, A => n3751, B => 
                           n27364, ZN => n27367);
   U27723 : NAND2_X1 port map( A1 => n27365, A2 => n27364, ZN => n27375);
   U27725 : NAND2_X1 port map( A1 => n27368, A2 => n27370, ZN => n27369);
   U27726 : NAND3_X1 port map( A1 => n28494, A2 => n27372, A3 => n29541, ZN => 
                           n27374);
   U27728 : OAI21_X1 port map( B1 => n27380, B2 => n27379, A => n295, ZN => 
                           n27381);
   U27730 : XNOR2_X1 port map( A => n27385, B => n27384, ZN => Ciphertext(17));
   U27731 : OAI22_X1 port map( A1 => n27400, A2 => n28177, B1 => n27386, B2 => 
                           n342, ZN => n27411);
   U27732 : NOR2_X1 port map( A1 => n25629, A2 => n27387, ZN => n27389);
   U27733 : AOI22_X1 port map( A1 => n27411, A2 => n27390, B1 => n27389, B2 => 
                           n27388, ZN => n27391);
   U27734 : XNOR2_X1 port map( A => n27391, B => n3196, ZN => Ciphertext(19));
   U27735 : NOR2_X1 port map( A1 => n27408, A2 => n27392, ZN => n27399);
   U27736 : INV_X1 port map( A => n27393, ZN => n27397);
   U27737 : MUX2_X1 port map( A => n27397, B => n27396, S => n27395, Z => 
                           n27398);
   U27738 : AOI22_X1 port map( A1 => n27400, A2 => n28177, B1 => n27399, B2 => 
                           n27398, ZN => n27401);
   U27739 : OAI222_X1 port map( A1 => n27404, A2 => n27410, B1 => n27403, B2 =>
                           n28177, C1 => n27402, C2 => n27401, ZN => n27406);
   U27740 : INV_X1 port map( A => n3457, ZN => n27405);
   U27741 : XNOR2_X1 port map( A => n27406, B => n27405, ZN => Ciphertext(22));
   U27742 : OAI21_X1 port map( B1 => n27409, B2 => n28177, A => n342, ZN => 
                           n27413);
   U27743 : NAND2_X1 port map( A1 => n27411, A2 => n4922, ZN => n27412);
   U27744 : NAND2_X1 port map( A1 => n27413, A2 => n27412, ZN => n27414);
   U27745 : XNOR2_X1 port map( A => n27414, B => n4222, ZN => Ciphertext(23));
   U27748 : OAI21_X1 port map( B1 => n27426, B2 => n6738, A => n27427, ZN => 
                           n27419);
   U27749 : AOI22_X1 port map( A1 => n27421, A2 => n27426, B1 => n27420, B2 => 
                           n27419, ZN => n27423);
   U27750 : XNOR2_X1 port map( A => n27423, B => n27422, ZN => Ciphertext(24));
   U27752 : INV_X1 port map( A => n2982, ZN => n27436);
   U27753 : XNOR2_X1 port map( A => n27437, B => n27436, ZN => Ciphertext(38));
   U27754 : AOI21_X1 port map( B1 => n27439, B2 => n27438, A => n25417, ZN => 
                           n27440);
   U27755 : OAI22_X1 port map( A1 => n27443, A2 => n27442, B1 => n27441, B2 => 
                           n27440, ZN => n27445);
   U27756 : XNOR2_X1 port map( A => n27445, B => n27444, ZN => Ciphertext(41));
   U27757 : NAND3_X1 port map( A1 => n27458, A2 => n27457, A3 => n27472, ZN => 
                           n27451);
   U27758 : INV_X1 port map( A => n27446, ZN => n27450);
   U27759 : OR3_X1 port map( A1 => n27465, A2 => n27447, A3 => n27457, ZN => 
                           n27449);
   U27760 : NAND3_X1 port map( A1 => n27457, A2 => n27465, A3 => n28435, ZN => 
                           n27448);
   U27761 : INV_X1 port map( A => n27452, ZN => n27453);
   U27762 : INV_X1 port map( A => n27462, ZN => n27466);
   U27763 : NOR2_X1 port map( A1 => n27465, A2 => n27466, ZN => n27461);
   U27764 : AND2_X1 port map( A1 => n27465, A2 => n27466, ZN => n27454);
   U27765 : NOR2_X1 port map( A1 => n27461, A2 => n27454, ZN => n27456);
   U27767 : AOI21_X1 port map( B1 => n27456, B2 => n4823, A => n27472, ZN => 
                           n27474);
   U27768 : XNOR2_X1 port map( A => n27457, B => n27462, ZN => n27459);
   U27769 : NAND2_X1 port map( A1 => n27459, A2 => n27458, ZN => n27473);
   U27770 : NAND2_X1 port map( A1 => n27461, A2 => n28435, ZN => n27470);
   U27771 : XNOR2_X1 port map( A => n27463, B => n27462, ZN => n27464);
   U27772 : NAND2_X1 port map( A1 => n27464, A2 => n27465, ZN => n27469);
   U27773 : NAND3_X1 port map( A1 => n449, A2 => n27467, A3 => n27466, ZN => 
                           n27468);
   U27774 : NAND3_X1 port map( A1 => n27470, A2 => n27469, A3 => n27468, ZN => 
                           n27471);
   U27775 : AOI22_X1 port map( A1 => n27474, A2 => n27473, B1 => n27472, B2 => 
                           n27471, ZN => Ciphertext(44));
   U27777 : AOI22_X1 port map( A1 => n27478, A2 => n27477, B1 => n27476, B2 => 
                           n27475, ZN => n27479);
   U27778 : XNOR2_X1 port map( A => n27479, B => n1225, ZN => Ciphertext(49));
   U27779 : XNOR2_X1 port map( A => n27492, B => n3501, ZN => n27484);
   U27780 : NAND2_X1 port map( A1 => n29093, A2 => n27480, ZN => n27483);
   U27781 : XNOR2_X1 port map( A => n29523, B => n5513, ZN => n27482);
   U27782 : OR2_X1 port map( A1 => n29093, A2 => n27497, ZN => n27481);
   U27783 : OAI22_X1 port map( A1 => n27484, A2 => n27483, B1 => n27482, B2 => 
                           n27481, ZN => n27491);
   U27784 : XNOR2_X1 port map( A => n27496, B => n3501, ZN => n27485);
   U27785 : OAI21_X1 port map( B1 => n27485, B2 => n29522, A => n27497, ZN => 
                           n27489);
   U27786 : XNOR2_X1 port map( A => n27493, B => n3501, ZN => n27486);
   U27787 : NOR2_X1 port map( A1 => n27487, A2 => n27486, ZN => n27488);
   U27788 : NOR2_X1 port map( A1 => n27489, A2 => n27488, ZN => n27490);
   U27789 : NOR2_X1 port map( A1 => n27491, A2 => n27490, ZN => Ciphertext(50))
                           ;
   U27791 : NOR2_X1 port map( A1 => n27496, A2 => n27493, ZN => n27495);
   U27792 : NAND3_X1 port map( A1 => n29522, A2 => n27497, A3 => n27496, ZN => 
                           n27499);
   U27793 : XNOR2_X1 port map( A => n27501, B => n628, ZN => Ciphertext(52));
   U27794 : NAND3_X1 port map( A1 => n27520, A2 => n27502, A3 => n27510, ZN => 
                           n27504);
   U27795 : NAND3_X1 port map( A1 => n27527, A2 => n27526, A3 => n27528, ZN => 
                           n27503);
   U27796 : OAI211_X1 port map( C1 => n27506, C2 => n27505, A => n27504, B => 
                           n27503, ZN => n27507);
   U27797 : XNOR2_X1 port map( A => n27507, B => n632, ZN => Ciphertext(55));
   U27798 : INV_X1 port map( A => n27509, ZN => n27512);
   U27799 : AOI21_X1 port map( B1 => n27531, B2 => n27512, A => n27511, ZN => 
                           n27514);
   U27800 : NOR3_X1 port map( A1 => n27526, A2 => n27520, A3 => n27528, ZN => 
                           n27516);
   U27801 : NAND2_X1 port map( A1 => n27516, A2 => n27515, ZN => n27517);
   U27802 : AND3_X1 port map( A1 => n27518, A2 => n27519, A3 => n27517, ZN => 
                           Ciphertext(56));
   U27803 : INV_X1 port map( A => n27531, ZN => n27521);
   U27804 : AOI21_X1 port map( B1 => n27524, B2 => n27523, A => n27522, ZN => 
                           n27533);
   U27805 : AND2_X1 port map( A1 => n27526, A2 => n27525, ZN => n27530);
   U27806 : NOR3_X1 port map( A1 => n27531, A2 => n27528, A3 => n27527, ZN => 
                           n27529);
   U27807 : AOI21_X1 port map( B1 => n27531, B2 => n27530, A => n27529, ZN => 
                           n27532);
   U27810 : OAI21_X1 port map( B1 => n27541, B2 => n28386, A => n27539, ZN => 
                           n27542);
   U27811 : OAI21_X1 port map( B1 => n27543, B2 => n394, A => n27542, ZN => 
                           n27544);
   U27812 : XNOR2_X1 port map( A => n27544, B => n621, ZN => Ciphertext(72));
   U27813 : INV_X1 port map( A => n3114, ZN => n27550);
   U27814 : AOI22_X1 port map( A1 => n27551, A2 => n27552, B1 => n29085, B2 => 
                           n2433, ZN => n27556);
   U27815 : INV_X1 port map( A => n27561, ZN => n27575);
   U27816 : NOR2_X1 port map( A1 => n27554, A2 => n27553, ZN => n27555);
   U27817 : OAI22_X1 port map( A1 => n27556, A2 => n27575, B1 => n27551, B2 => 
                           n27555, ZN => n27558);
   U27818 : INV_X1 port map( A => n3049, ZN => n27557);
   U27819 : XNOR2_X1 port map( A => n27558, B => n27557, ZN => Ciphertext(78));
   U27820 : AOI21_X1 port map( B1 => n27571, B2 => n27551, A => n27576, ZN => 
                           n27566);
   U27821 : NOR2_X1 port map( A1 => n27571, A2 => n27573, ZN => n27577);
   U27822 : AOI21_X1 port map( B1 => n27577, B2 => n29158, A => n3087, ZN => 
                           n27559);
   U27823 : NAND2_X1 port map( A1 => n27566, A2 => n27559, ZN => n27570);
   U27824 : AND3_X1 port map( A1 => n27562, A2 => n27561, A3 => n27560, ZN => 
                           n27565);
   U27825 : NAND2_X1 port map( A1 => n27562, A2 => n3087, ZN => n27563);
   U27826 : NAND2_X1 port map( A1 => n27577, A2 => n27563, ZN => n27564);
   U27827 : OAI21_X1 port map( B1 => n27577, B2 => n27565, A => n27564, ZN => 
                           n27569);
   U27828 : INV_X1 port map( A => n27566, ZN => n27568);
   U27829 : NOR2_X1 port map( A1 => n27551, A2 => n27571, ZN => n27574);
   U27830 : OAI21_X1 port map( B1 => n27574, B2 => n29578, A => n29085, ZN => 
                           n27579);
   U27831 : OAI21_X1 port map( B1 => n27577, B2 => n27576, A => n27575, ZN => 
                           n27578);
   U27832 : NAND2_X1 port map( A1 => n27578, A2 => n27579, ZN => n27581);
   U27833 : INV_X1 port map( A => n2602, ZN => n27580);
   U27834 : XNOR2_X1 port map( A => n27581, B => n27580, ZN => Ciphertext(83));
   U27835 : OAI21_X1 port map( B1 => n1901, B2 => n27585, A => n27589, ZN => 
                           n27583);
   U27836 : OAI21_X1 port map( B1 => n27598, B2 => n27592, A => n27583, ZN => 
                           n27584);
   U27837 : XNOR2_X1 port map( A => n27584, B => n22534, ZN => Ciphertext(85));
   U27838 : NOR2_X1 port map( A1 => n930, A2 => n27593, ZN => n27595);
   U27839 : OAI22_X1 port map( A1 => n27598, A2 => n27597, B1 => n27596, B2 => 
                           n27595, ZN => n27600);
   U27840 : INV_X1 port map( A => n28294, ZN => n27599);
   U27841 : XNOR2_X1 port map( A => n27600, B => n27599, ZN => Ciphertext(89));
   U27842 : NAND2_X1 port map( A1 => n27601, A2 => n27625, ZN => n27604);
   U27843 : NOR2_X1 port map( A1 => n27628, A2 => n3366, ZN => n27603);
   U27844 : NOR2_X1 port map( A1 => n27627, A2 => n27625, ZN => n27602);
   U27845 : XNOR2_X1 port map( A => n27606, B => n27605, ZN => Ciphertext(90));
   U27847 : NAND2_X1 port map( A1 => n27626, A2 => n27617, ZN => n27608);
   U27848 : AOI22_X1 port map( A1 => n27610, A2 => n28505, B1 => n27609, B2 => 
                           n27608, ZN => n27612);
   U27849 : XNOR2_X1 port map( A => n27612, B => n3035, ZN => Ciphertext(91));
   U27850 : MUX2_X1 port map( A => n27614, B => n3366, S => n27613, Z => n27615
                           );
   U27852 : XNOR2_X1 port map( A => n27625, B => n28213, ZN => n27616);
   U27853 : NAND3_X1 port map( A1 => n27619, A2 => n27617, A3 => n3154, ZN => 
                           n27621);
   U27854 : NAND3_X1 port map( A1 => n27619, A2 => n28213, A3 => n27628, ZN => 
                           n27620);
   U27855 : NOR3_X1 port map( A1 => n27624, A2 => n27623, A3 => n27622, ZN => 
                           Ciphertext(92));
   U27856 : NAND2_X1 port map( A1 => n1912, A2 => n27628, ZN => n27631);
   U27857 : INV_X1 port map( A => n3334, ZN => n27633);
   U27858 : XNOR2_X1 port map( A => n27634, B => n27633, ZN => Ciphertext(94));
   U27859 : MUX2_X1 port map( A => n27637, B => n27636, S => n29532, Z => 
                           n27642);
   U27860 : NAND2_X1 port map( A1 => n27639, A2 => n27638, ZN => n27647);
   U27863 : AOI21_X1 port map( B1 => n27647, B2 => n28466, A => n27645, ZN => 
                           n27648);
   U27864 : AOI21_X1 port map( B1 => n27650, B2 => n27649, A => n27648, ZN => 
                           n27651);
   U27865 : XNOR2_X1 port map( A => n27651, B => n1887, ZN => Ciphertext(101));
   U27866 : INV_X1 port map( A => n27652, ZN => n27655);
   U27867 : AOI22_X1 port map( A1 => n27674, A2 => n27663, B1 => n27672, B2 => 
                           n27671, ZN => n27677);
   U27868 : INV_X1 port map( A => n29091, ZN => n27653);
   U27869 : OAI21_X1 port map( B1 => n27655, B2 => n27677, A => n27654, ZN => 
                           n27657);
   U27870 : XNOR2_X1 port map( A => n27657, B => n27656, ZN => Ciphertext(103))
                           ;
   U27871 : MUX2_X1 port map( A => n29091, B => n28655, S => n27661, Z => 
                           n27659);
   U27872 : MUX2_X1 port map( A => n27659, B => n27658, S => n27663, Z => 
                           n27660);
   U27873 : XNOR2_X1 port map( A => n27660, B => n4503, ZN => Ciphertext(104));
   U27877 : XNOR2_X1 port map( A => n27670, B => n27669, ZN => Ciphertext(106))
                           ;
   U27878 : AOI21_X1 port map( B1 => n29090, B2 => n27672, A => n85, ZN => 
                           n27675);
   U27879 : OAI22_X1 port map( A1 => n27677, A2 => n27676, B1 => n27675, B2 => 
                           n27674, ZN => n27679);
   U27880 : XNOR2_X1 port map( A => n27679, B => n27678, ZN => Ciphertext(107))
                           ;
   U27882 : NOR2_X1 port map( A1 => n27714, A2 => n27725, ZN => n27680);
   U27883 : NAND2_X1 port map( A1 => n1826, A2 => n27680, ZN => n27683);
   U27884 : OAI21_X1 port map( B1 => n27681, B2 => n27711, A => n27725, ZN => 
                           n27682);
   U27885 : OAI211_X1 port map( C1 => n27727, C2 => n27684, A => n27683, B => 
                           n27682, ZN => n27686);
   U27886 : INV_X1 port map( A => n1246, ZN => n27685);
   U27887 : XNOR2_X1 port map( A => n27686, B => n27685, ZN => Ciphertext(108))
                           ;
   U27888 : INV_X1 port map( A => n27707, ZN => n27689);
   U27889 : NAND2_X1 port map( A1 => n27689, A2 => n27687, ZN => n27693);
   U27890 : NAND3_X1 port map( A1 => n27690, A2 => n27689, A3 => n27688, ZN => 
                           n27692);
   U27891 : AOI21_X1 port map( B1 => n27693, B2 => n27692, A => n27691, ZN => 
                           n27695);
   U27892 : INV_X1 port map( A => n27711, ZN => n27723);
   U27893 : NOR2_X1 port map( A1 => n27695, A2 => n27694, ZN => n27729);
   U27894 : NOR2_X1 port map( A1 => n27727, A2 => n326, ZN => n27697);
   U27895 : OAI21_X1 port map( B1 => n28396, B2 => n27697, A => n27696, ZN => 
                           n27698);
   U27896 : XNOR2_X1 port map( A => n27698, B => n22755, ZN => Ciphertext(109))
                           ;
   U27897 : NOR2_X1 port map( A1 => n27701, A2 => n27704, ZN => n27699);
   U27898 : AOI211_X1 port map( C1 => n27701, C2 => n27700, A => n27702, B => 
                           n27699, ZN => n27709);
   U27899 : NAND2_X1 port map( A1 => n27703, A2 => n27702, ZN => n27705);
   U27900 : NOR2_X1 port map( A1 => n27705, A2 => n27704, ZN => n27706);
   U27901 : OR2_X1 port map( A1 => n27707, A2 => n27706, ZN => n27708);
   U27902 : NOR2_X1 port map( A1 => n27709, A2 => n27708, ZN => n27716);
   U27905 : INV_X1 port map( A => n27725, ZN => n27712);
   U27906 : NAND2_X1 port map( A1 => n27713, A2 => n27712, ZN => n27721);
   U27907 : NAND3_X1 port map( A1 => n27715, A2 => n27714, A3 => n27725, ZN => 
                           n27720);
   U27908 : INV_X1 port map( A => n27716, ZN => n27717);
   U27909 : NAND3_X1 port map( A1 => n1826, A2 => n324, A3 => n27717, ZN => 
                           n27719);
   U27911 : XNOR2_X1 port map( A => n27722, B => n3062, ZN => Ciphertext(110));
   U27912 : AOI21_X1 port map( B1 => n27725, B2 => n27724, A => n27723, ZN => 
                           n27726);
   U27913 : OAI22_X1 port map( A1 => n27729, A2 => n1826, B1 => n27727, B2 => 
                           n27726, ZN => n27731);
   U27914 : XNOR2_X1 port map( A => n27731, B => n27730, ZN => Ciphertext(113))
                           ;
   U27915 : INV_X1 port map( A => n29049, ZN => n27746);
   U27916 : AOI21_X1 port map( B1 => n27739, B2 => n28430, A => n27744, ZN => 
                           n27736);
   U27917 : NOR2_X1 port map( A1 => n27745, A2 => n29049, ZN => n27734);
   U27918 : NOR2_X1 port map( A1 => n27739, A2 => n27732, ZN => n27733);
   U27919 : XNOR2_X1 port map( A => n27738, B => n27737, ZN => Ciphertext(114))
                           ;
   U27920 : OR2_X1 port map( A1 => n29049, A2 => n27755, ZN => n27741);
   U27921 : NOR2_X1 port map( A1 => n27739, A2 => n28430, ZN => n27740);
   U27922 : AOI22_X1 port map( A1 => n27755, A2 => n27744, B1 => n27759, B2 => 
                           n397, ZN => n27758);
   U27923 : XNOR2_X1 port map( A => n27743, B => n27742, ZN => Ciphertext(115))
                           ;
   U27924 : NOR2_X1 port map( A1 => n27745, A2 => n27744, ZN => n27747);
   U27925 : OAI22_X1 port map( A1 => n27747, A2 => n27759, B1 => n27746, B2 => 
                           n28445, ZN => n27752);
   U27926 : NOR3_X1 port map( A1 => n27757, A2 => n27749, A3 => n397, ZN => 
                           n27751);
   U27927 : NOR2_X1 port map( A1 => n28445, A2 => n397, ZN => n27748);
   U27928 : OAI211_X1 port map( C1 => n27757, C2 => n27749, A => n27748, B => 
                           n29049, ZN => n27750);
   U27931 : AOI21_X1 port map( B1 => n29049, B2 => n27755, A => n28445, ZN => 
                           n27760);
   U27932 : OAI22_X1 port map( A1 => n27760, A2 => n27759, B1 => n27758, B2 => 
                           n27757, ZN => n27761);
   U27933 : XNOR2_X1 port map( A => n27761, B => n4882, ZN => Ciphertext(119));
   U27935 : OAI211_X1 port map( C1 => n29027, C2 => n29537, A => n29070, B => 
                           n29118, ZN => n27765);
   U27936 : INV_X1 port map( A => n27784, ZN => n27764);
   U27937 : NOR2_X1 port map( A1 => n28414, A2 => n29117, ZN => n27785);
   U27938 : XNOR2_X1 port map( A => n27767, B => n27766, ZN => Ciphertext(121))
                           ;
   U27939 : OAI211_X1 port map( C1 => n27777, C2 => n27776, A => n27775, B => 
                           n27774, ZN => n27779);
   U27940 : XNOR2_X1 port map( A => n27779, B => n27778, ZN => Ciphertext(124))
                           ;
   U27941 : OAI21_X1 port map( B1 => n27782, B2 => n28414, A => n27780, ZN => 
                           n27787);
   U27942 : OAI21_X1 port map( B1 => n27785, B2 => n27784, A => n29027, ZN => 
                           n27786);
   U27943 : NAND2_X1 port map( A1 => n27787, A2 => n27786, ZN => n27789);
   U27944 : XNOR2_X1 port map( A => n27789, B => n27788, ZN => Ciphertext(125))
                           ;
   U27946 : NAND2_X1 port map( A1 => n27790, A2 => n27817, ZN => n27793);
   U27947 : OAI211_X1 port map( C1 => n27800, C2 => n29535, A => n27793, B => 
                           n27792, ZN => n27794);
   U27948 : XNOR2_X1 port map( A => n27794, B => n4070, ZN => Ciphertext(126));
   U27949 : NAND2_X1 port map( A1 => n28403, A2 => n3380, ZN => n27799);
   U27950 : AND2_X1 port map( A1 => n27817, A2 => n3380, ZN => n27806);
   U27951 : OAI21_X1 port map( B1 => n27795, B2 => n3380, A => n27807, ZN => 
                           n27796);
   U27952 : AOI21_X1 port map( B1 => n27812, B2 => n27806, A => n27796, ZN => 
                           n27798);
   U27953 : NAND2_X1 port map( A1 => n27800, A2 => n27811, ZN => n27797);
   U27954 : OAI211_X1 port map( C1 => n27800, C2 => n27799, A => n27798, B => 
                           n27797, ZN => n27816);
   U27955 : NAND2_X1 port map( A1 => n29469, A2 => n27811, ZN => n27805);
   U27956 : AOI21_X1 port map( B1 => n27819, B2 => n3380, A => n27807, ZN => 
                           n27804);
   U27957 : NAND2_X1 port map( A1 => n27818, A2 => n27811, ZN => n27802);
   U27958 : NAND2_X1 port map( A1 => n27802, A2 => n27817, ZN => n27803);
   U27959 : OAI211_X1 port map( C1 => n27819, C2 => n27805, A => n27804, B => 
                           n27803, ZN => n27815);
   U27960 : INV_X1 port map( A => n27806, ZN => n27808);
   U27961 : NOR3_X1 port map( A1 => n27808, A2 => n27818, A3 => n27807, ZN => 
                           n27809);
   U27962 : NAND2_X1 port map( A1 => n29535, A2 => n27809, ZN => n27814);
   U27963 : NAND3_X1 port map( A1 => n27812, A2 => n27811, A3 => n27817, ZN => 
                           n27813);
   U27964 : NAND4_X1 port map( A1 => n27816, A2 => n27815, A3 => n27814, A4 => 
                           n27813, ZN => Ciphertext(130));
   U27965 : OAI21_X1 port map( B1 => n27819, B2 => n27818, A => n27817, ZN => 
                           n27820);
   U27966 : AOI22_X1 port map( A1 => n27823, A2 => n27822, B1 => n27821, B2 => 
                           n27820, ZN => n27824);
   U27967 : XNOR2_X1 port map( A => n27824, B => n3463, ZN => Ciphertext(131));
   U27968 : INV_X1 port map( A => n27829, ZN => n27833);
   U27969 : INV_X1 port map( A => n27830, ZN => n27832);
   U27970 : NAND4_X1 port map( A1 => n27834, A2 => n27833, A3 => n27832, A4 => 
                           n27831, ZN => n27845);
   U27971 : MUX2_X1 port map( A => n27898, B => n27836, S => n29575, Z => 
                           n27837);
   U27972 : NOR2_X1 port map( A1 => n27837, A2 => n5299, ZN => n27840);
   U27973 : NOR3_X1 port map( A1 => n27840, A2 => n27839, A3 => n27838, ZN => 
                           n27842);
   U27974 : NAND2_X1 port map( A1 => n27842, A2 => n27841, ZN => n27844);
   U27975 : AOI21_X1 port map( B1 => n27845, B2 => n27844, A => n27843, ZN => 
                           n27846);
   U27976 : NOR2_X1 port map( A1 => n27851, A2 => n27852, ZN => n27853);
   U27977 : AOI22_X1 port map( A1 => n27855, A2 => n27853, B1 => n27859, B2 => 
                           n6949, ZN => n27857);
   U27978 : OAI211_X1 port map( C1 => n27859, C2 => n27858, A => n27857, B => 
                           n27856, ZN => n27861);
   U27979 : INV_X1 port map( A => n3527, ZN => n27860);
   U27980 : XNOR2_X1 port map( A => n27861, B => n27860, ZN => Ciphertext(141))
                           ;
   U27981 : AOI22_X1 port map( A1 => n27875, A2 => n27864, B1 => n27862, B2 => 
                           n27863, ZN => n27878);
   U27982 : NOR2_X1 port map( A1 => n27875, A2 => n26540, ZN => n27868);
   U27983 : NAND3_X1 port map( A1 => n27872, A2 => n27871, A3 => n27866, ZN => 
                           n27867);
   U27984 : OAI21_X1 port map( B1 => n27878, B2 => n27868, A => n27867, ZN => 
                           n27870);
   U27985 : INV_X1 port map( A => n2987, ZN => n27869);
   U27986 : XNOR2_X1 port map( A => n27870, B => n27869, ZN => Ciphertext(145))
                           ;
   U27987 : NOR2_X1 port map( A1 => n27872, A2 => n27871, ZN => n27874);
   U27988 : NOR2_X1 port map( A1 => n27874, A2 => n27873, ZN => n27876);
   U27989 : OAI22_X1 port map( A1 => n27878, A2 => n27877, B1 => n27876, B2 => 
                           n27875, ZN => n27880);
   U27990 : XNOR2_X1 port map( A => n27880, B => n27879, ZN => Ciphertext(149))
                           ;
   U27991 : NAND2_X1 port map( A1 => n27919, A2 => n27080, ZN => n27882);
   U27992 : OAI21_X1 port map( B1 => n27905, B2 => n27908, A => n27918, ZN => 
                           n27881);
   U27993 : OAI21_X1 port map( B1 => n27882, B2 => n27908, A => n27881, ZN => 
                           n27886);
   U27994 : NAND2_X1 port map( A1 => n27908, A2 => n27923, ZN => n27885);
   U27995 : INV_X1 port map( A => n27883, ZN => n27884);
   U27996 : XNOR2_X1 port map( A => n27888, B => n27887, ZN => Ciphertext(152))
                           ;
   U27997 : INV_X1 port map( A => n27908, ZN => n27909);
   U27998 : OAI21_X1 port map( B1 => n27919, B2 => n27909, A => n1843, ZN => 
                           n27892);
   U27999 : NAND3_X1 port map( A1 => n27918, A2 => n27908, A3 => n27905, ZN => 
                           n27891);
   U28000 : NAND2_X1 port map( A1 => n27889, A2 => n27920, ZN => n27890);
   U28004 : OAI21_X1 port map( B1 => n27060, B2 => n27898, A => n28600, ZN => 
                           n27901);
   U28005 : AOI211_X1 port map( C1 => n27902, C2 => n27901, A => n27900, B => 
                           n27899, ZN => n27907);
   U28006 : OAI21_X1 port map( B1 => n27904, B2 => n27903, A => n27060, ZN => 
                           n27906);
   U28007 : INV_X1 port map( A => n27905, ZN => n27917);
   U28008 : NAND3_X1 port map( A1 => n27920, A2 => n27908, A3 => n1843, ZN => 
                           n27912);
   U28009 : NAND3_X1 port map( A1 => n27080, A2 => n27909, A3 => n27917, ZN => 
                           n27911);
   U28010 : OAI211_X1 port map( C1 => n27914, C2 => n1843, A => n27912, B => 
                           n27911, ZN => n27916);
   U28011 : XNOR2_X1 port map( A => n27916, B => n27915, ZN => Ciphertext(154))
                           ;
   U28012 : OAI21_X1 port map( B1 => n27919, B2 => n27918, A => n27917, ZN => 
                           n27922);
   U28013 : AOI22_X1 port map( A1 => n27923, A2 => n27922, B1 => n27921, B2 => 
                           n27920, ZN => n27924);
   U28014 : XNOR2_X1 port map( A => n27924, B => n2510, ZN => Ciphertext(155));
   U28015 : INV_X1 port map( A => n27925, ZN => n27950);
   U28016 : INV_X1 port map( A => n27934, ZN => n27942);
   U28018 : OAI21_X1 port map( B1 => n27948, B2 => n27927, A => n27926, ZN => 
                           n27929);
   U28019 : OAI211_X1 port map( C1 => n27942, C2 => n28451, A => n27929, B => 
                           n27928, ZN => n27931);
   U28020 : INV_X1 port map( A => n3317, ZN => n27930);
   U28021 : XNOR2_X1 port map( A => n27931, B => n27930, ZN => Ciphertext(156))
                           ;
   U28022 : NOR2_X1 port map( A1 => n27944, A2 => n27938, ZN => n27947);
   U28023 : NOR2_X1 port map( A1 => n27244, A2 => n27947, ZN => n27935);
   U28024 : NAND2_X1 port map( A1 => n27941, A2 => n28441, ZN => n27932);
   U28025 : OAI21_X1 port map( B1 => n27935, B2 => n27934, A => n27933, ZN => 
                           n27937);
   U28026 : XNOR2_X1 port map( A => n27937, B => n27936, ZN => Ciphertext(157))
                           ;
   U28027 : XNOR2_X1 port map( A => n27943, B => n5802, ZN => Ciphertext(159));
   U28028 : AOI21_X1 port map( B1 => n27926, B2 => n4998, A => n27944, ZN => 
                           n27951);
   U28029 : AOI22_X1 port map( A1 => n27948, A2 => n27950, B1 => n27947, B2 => 
                           n28451, ZN => n27949);
   U28030 : OAI21_X1 port map( B1 => n27951, B2 => n27950, A => n27949, ZN => 
                           n27953);
   U28031 : XNOR2_X1 port map( A => n27953, B => n27952, ZN => Ciphertext(161))
                           ;
   U28032 : NOR2_X1 port map( A1 => n27972, A2 => n27996, ZN => n27965);
   U28034 : AND2_X1 port map( A1 => n29021, A2 => n27977, ZN => n27954);
   U28035 : INV_X1 port map( A => n27956, ZN => n27957);
   U28038 : INV_X1 port map( A => n27997, ZN => n27964);
   U28040 : OAI211_X1 port map( C1 => n27964, C2 => n29092, A => n27977, B => 
                           n27979, ZN => n27960);
   U28041 : OAI21_X1 port map( B1 => n27998, B2 => n27965, A => n27960, ZN => 
                           n27962);
   U28042 : XNOR2_X1 port map( A => n27962, B => n27961, ZN => Ciphertext(163))
                           ;
   U28043 : MUX2_X1 port map( A => n27970, B => n27977, S => n27979, Z => 
                           n27967);
   U28044 : INV_X1 port map( A => n27996, ZN => n27983);
   U28045 : AND2_X1 port map( A1 => n27977, A2 => n27972, ZN => n27963);
   U28046 : AOI22_X1 port map( A1 => n27965, A2 => n27964, B1 => n27963, B2 => 
                           n28456, ZN => n27966);
   U28047 : OAI21_X1 port map( B1 => n27967, B2 => n27983, A => n27966, ZN => 
                           n27969);
   U28048 : INV_X1 port map( A => n3211, ZN => n27968);
   U28049 : XNOR2_X1 port map( A => n27969, B => n27968, ZN => Ciphertext(165))
                           ;
   U28050 : NOR2_X1 port map( A1 => n28456, A2 => n27977, ZN => n27987);
   U28051 : INV_X1 port map( A => n27987, ZN => n27971);
   U28052 : NOR2_X1 port map( A1 => n27971, A2 => n27970, ZN => n27991);
   U28053 : AND2_X1 port map( A1 => n27972, A2 => n3722, ZN => n27976);
   U28054 : INV_X1 port map( A => n27976, ZN => n27975);
   U28055 : AOI21_X1 port map( B1 => n28636, B2 => n27978, A => n27983, ZN => 
                           n27974);
   U28056 : NAND2_X1 port map( A1 => n29092, A2 => n27978, ZN => n27985);
   U28057 : OAI211_X1 port map( C1 => n28636, C2 => n27975, A => n27974, B => 
                           n27985, ZN => n27990);
   U28058 : AND2_X1 port map( A1 => n27987, A2 => n27976, ZN => n27984);
   U28059 : NAND2_X1 port map( A1 => n27977, A2 => n27978, ZN => n27982);
   U28060 : XNOR2_X1 port map( A => n27979, B => n27978, ZN => n27980);
   U28061 : INV_X1 port map( A => n27985, ZN => n27986);
   U28062 : NAND2_X1 port map( A1 => n27987, A2 => n27986, ZN => n27988);
   U28063 : OAI211_X1 port map( C1 => n27991, C2 => n27990, A => n27989, B => 
                           n27988, ZN => Ciphertext(166));
   U28064 : AOI21_X1 port map( B1 => n29021, B2 => n29063, A => n28456, ZN => 
                           n27995);
   U28065 : OAI22_X1 port map( A1 => n27998, A2 => n28636, B1 => n27996, B2 => 
                           n27995, ZN => n27999);
   U28066 : XNOR2_X1 port map( A => n27999, B => n635, ZN => Ciphertext(167));
   U28067 : NAND3_X1 port map( A1 => n445, A2 => n28003, A3 => n28015, ZN => 
                           n28004);
   U28068 : INV_X1 port map( A => n28015, ZN => n28008);
   U28069 : NAND3_X1 port map( A1 => n28411, A2 => n28008, A3 => n26984, ZN => 
                           n28011);
   U28070 : NAND2_X1 port map( A1 => n6955, A2 => n443, ZN => n28010);
   U28071 : XNOR2_X1 port map( A => n28014, B => n28013, ZN => Ciphertext(172))
                           ;
   U28072 : NAND2_X1 port map( A1 => n28017, A2 => n28016, ZN => n28018);
   U28073 : NAND2_X1 port map( A1 => n28008, A2 => n28018, ZN => n28020);
   U28074 : AOI22_X1 port map( A1 => n28022, A2 => n28021, B1 => n28020, B2 => 
                           n28019, ZN => n28023);
   U28075 : XNOR2_X1 port map( A => n28023, B => n3323, ZN => Ciphertext(173));
   U28076 : AOI22_X1 port map( A1 => n28030, A2 => n28028, B1 => n28034, B2 => 
                           n28027, ZN => n28029);
   U28077 : OAI21_X1 port map( B1 => n28031, B2 => n28030, A => n28029, ZN => 
                           n28033);
   U28078 : INV_X1 port map( A => n3695, ZN => n28032);
   U28079 : XNOR2_X1 port map( A => n28033, B => n28032, ZN => Ciphertext(174))
                           ;
   U28080 : NOR3_X1 port map( A1 => n28040, A2 => n28039, A3 => n28038, ZN => 
                           n28041);
   U28081 : NOR2_X1 port map( A1 => n28042, A2 => n28041, ZN => n28043);
   U28082 : XNOR2_X1 port map( A => n28043, B => n4501, ZN => Ciphertext(176));
   U28083 : NOR2_X1 port map( A1 => n28044, A2 => n28543, ZN => n28046);
   U28084 : INV_X1 port map( A => n28067, ZN => n28045);
   U28085 : OAI21_X1 port map( B1 => n28055, B2 => n28046, A => n28045, ZN => 
                           n28049);
   U28086 : OAI21_X1 port map( B1 => n28047, B2 => n28065, A => n28543, ZN => 
                           n28048);
   U28087 : NAND2_X1 port map( A1 => n28049, A2 => n28048, ZN => n28051);
   U28088 : XNOR2_X1 port map( A => n28051, B => n28050, ZN => Ciphertext(180))
                           ;
   U28089 : NOR2_X1 port map( A1 => n28052, A2 => n28063, ZN => n28056);
   U28090 : OAI21_X1 port map( B1 => n28067, B2 => n28063, A => n28053, ZN => 
                           n28054);
   U28091 : OAI21_X1 port map( B1 => n28056, B2 => n28055, A => n28054, ZN => 
                           n28058);
   U28092 : INV_X1 port map( A => n3650, ZN => n28057);
   U28093 : XNOR2_X1 port map( A => n28058, B => n28057, ZN => Ciphertext(181))
                           ;
   U28094 : MUX2_X1 port map( A => n28067, B => n28543, S => n28069, Z => 
                           n28060);
   U28095 : MUX2_X1 port map( A => n28060, B => n28059, S => n28063, Z => 
                           n28062);
   U28096 : INV_X1 port map( A => n2505, ZN => n28061);
   U28097 : XNOR2_X1 port map( A => n28062, B => n28061, ZN => Ciphertext(182))
                           ;
   U28098 : INV_X1 port map( A => n28063, ZN => n28068);
   U28099 : MUX2_X1 port map( A => n28069, B => n28068, S => n28543, Z => 
                           n28072);
   U28100 : OR2_X1 port map( A1 => n28066, A2 => n28065, ZN => n28070);
   U28101 : XNOR2_X1 port map( A => n28074, B => n28073, ZN => Ciphertext(184))
                           ;
   U28103 : INV_X1 port map( A => n28115, ZN => n28075);
   U28104 : OAI211_X1 port map( C1 => n28075, C2 => n29121, A => n28089, B => 
                           n28090, ZN => n28076);
   U28106 : INV_X1 port map( A => n3015, ZN => n28078);
   U28107 : XNOR2_X1 port map( A => n28079, B => n28078, ZN => Ciphertext(187))
                           ;
   U28109 : NAND2_X1 port map( A1 => n28590, A2 => n28794, ZN => n28081);
   U28111 : OAI21_X1 port map( B1 => n29480, B2 => n28081, A => n28080, ZN => 
                           n28087);
   U28112 : NAND2_X1 port map( A1 => n28090, A2 => n28794, ZN => n28084);
   U28113 : NAND3_X1 port map( A1 => n28111, A2 => n28090, A3 => n29121, ZN => 
                           n28083);
   U28114 : OAI211_X1 port map( C1 => n28107, C2 => n28084, A => n1928, B => 
                           n28083, ZN => n28086);
   U28115 : NOR2_X1 port map( A1 => n28111, A2 => n28794, ZN => n28105);
   U28116 : AND2_X1 port map( A1 => n28087, A2 => n4359, ZN => n28088);
   U28117 : NAND2_X1 port map( A1 => n29056, A2 => n28089, ZN => n28096);
   U28118 : NOR3_X1 port map( A1 => n28107, A2 => n28089, A3 => n28794, ZN => 
                           n28093);
   U28119 : AND3_X1 port map( A1 => n28111, A2 => n28794, A3 => n28090, ZN => 
                           n28092);
   U28120 : NOR2_X1 port map( A1 => n28093, A2 => n28092, ZN => n28095);
   U28122 : AOI21_X1 port map( B1 => n29056, B2 => n28112, A => n28111, ZN => 
                           n28114);
   U28123 : INV_X1 port map( A => n2446, ZN => n28116);
   U6151 : NAND2_X2 port map( A1 => n5663, A2 => n5665, ZN => n22434);
   U3467 : XNOR2_X2 port map( A => Key(105), B => Plaintext(105), ZN => n8231);
   U2036 : OAI21_X2 port map( B1 => n6976, B2 => n8231, A => n6975, ZN => n5945
                           );
   U1808 : BUF_X1 port map( A => n7560, Z => n8044);
   U5612 : NOR2_X2 port map( A1 => n26355, A2 => n26354, ZN => n1912);
   U14802 : INV_X1 port map( A => n7198, ZN => n8281);
   U3188 : XNOR2_X2 port map( A => n9769, B => n9768, ZN => n3441);
   U1772 : OAI211_X2 port map( C1 => n20932, C2 => n20931, A => n20930, B => 
                           n20929, ZN => n22094);
   U14624 : XNOR2_X2 port map( A => n7077, B => Key(185), ZN => n7093);
   U775 : BUF_X1 port map( A => n24205, Z => n24814);
   U1023 : XNOR2_X1 port map( A => n15043, B => n15044, ZN => n337);
   U10135 : NOR2_X1 port map( A1 => n3991, A2 => n10050, ZN => n11855);
   U2015 : XNOR2_X2 port map( A => n4506, B => n4505, ZN => n11209);
   U2541 : AND2_X2 port map( A1 => n20402, A2 => n5871, ZN => n21539);
   U1999 : NOR2_X2 port map( A1 => n11405, A2 => n11403, ZN => n11848);
   U1253 : OAI21_X1 port map( B1 => n11952, B2 => n11665, A => n5901, ZN => 
                           n11668);
   U3263 : NAND3_X2 port map( A1 => n3296, A2 => n8406, A3 => n8405, ZN => 
                           n10128);
   U2202 : NAND3_X2 port map( A1 => n24884, A2 => n2615, A3 => n1995, ZN => 
                           n27638);
   U462 : OAI21_X1 port map( B1 => n11784, B2 => n666, A => n667, ZN => n12542)
                           ;
   U2363 : OAI21_X2 port map( B1 => n23574, B2 => n23573, A => n23572, ZN => 
                           n24760);
   U1864 : AND3_X2 port map( A1 => n873, A2 => n5350, A3 => n5348, ZN => n25681
                           );
   U21 : NAND2_X2 port map( A1 => n24090, A2 => n24091, ZN => n24471);
   U27204 : BUF_X1 port map( A => n26539, Z => n27864);
   U1879 : MUX2_X2 port map( A => n23249, B => n23248, S => n23247, Z => n24367
                           );
   U248 : XNOR2_X1 port map( A => n24301, B => n24302, ZN => n26191);
   U4391 : XNOR2_X2 port map( A => n19204, B => n19205, ZN => n20349);
   U445 : INV_X1 port map( A => n17780, ZN => n18168);
   U20591 : XNOR2_X2 port map( A => n16276, B => n16275, ZN => n17148);
   U2038 : BUF_X1 port map( A => n7371, Z => n8222);
   U12034 : XNOR2_X1 port map( A => n4753, B => n16342, ZN => n17179);
   U219 : AOI22_X1 port map( A1 => n28807, A2 => n125, B1 => n11611, B2 => 
                           n11767, ZN => n12548);
   U2052 : CLKBUF_X1 port map( A => Key(92), Z => n3164);
   U3493 : CLKBUF_X1 port map( A => Key(158), Z => n3644);
   U3450 : CLKBUF_X1 port map( A => Key(111), Z => n26909);
   U113 : CLKBUF_X1 port map( A => Key(125), Z => n2946);
   U821 : XNOR2_X1 port map( A => Key(28), B => Plaintext(28), ZN => n8151);
   U642 : CLKBUF_X1 port map( A => Key(138), Z => n2403);
   U1045 : CLKBUF_X1 port map( A => Key(152), Z => n3527);
   U3483 : CLKBUF_X1 port map( A => Key(77), Z => n2961);
   U228 : CLKBUF_X1 port map( A => Key(99), Z => n2527);
   U115 : CLKBUF_X1 port map( A => Key(95), Z => n72);
   U14797 : XNOR2_X1 port map( A => Key(138), B => Plaintext(138), ZN => n8275)
                           ;
   U846 : AND2_X1 port map( A1 => n7857, A2 => n7858, ZN => n9015);
   U3381 : NAND3_X1 port map( A1 => n7323, A2 => n7280, A3 => n2716, ZN => 
                           n8889);
   U6648 : OAI211_X1 port map( C1 => n5559, C2 => n5558, A => n7305, B => n7304
                           , ZN => n9421);
   U8556 : NAND2_X1 port map( A1 => n7246, A2 => n2470, ZN => n8749);
   U1321 : OAI211_X1 port map( C1 => n7967, C2 => n7188, A => n7962, B => n5470
                           , ZN => n8809);
   U4350 : OAI211_X1 port map( C1 => n4939, C2 => n1700, A => n1404, B => n7091
                           , ZN => n8586);
   U423 : NAND2_X1 port map( A1 => n7078, A2 => n2507, ZN => n8521);
   U6673 : INV_X1 port map( A => n8589, ZN => n8594);
   U2032 : NAND2_X1 port map( A1 => n6382, A2 => n6381, ZN => n8610);
   U391 : NAND2_X1 port map( A1 => n2388, A2 => n2080, ZN => n9202);
   U1191 : OR2_X1 port map( A1 => n8439, A2 => n8720, ZN => n224);
   U715 : BUF_X1 port map( A => n8230, Z => n8961);
   U16085 : BUF_X1 port map( A => n9306, Z => n9725);
   U889 : AND3_X1 port map( A1 => n9365, A2 => n3273, A3 => n3272, ZN => n10352
                           );
   U3264 : NAND3_X1 port map( A1 => n1118, A2 => n9048, A3 => n1117, ZN => 
                           n10435);
   U3258 : NAND2_X1 port map( A1 => n8083, A2 => n8082, ZN => n10289);
   U3233 : XNOR2_X1 port map( A => n10262, B => n10261, ZN => n10876);
   U10153 : XNOR2_X1 port map( A => n9554, B => n9553, ZN => n11275);
   U4315 : XNOR2_X1 port map( A => n5185, B => n10058, ZN => n11154);
   U15875 : XNOR2_X1 port map( A => n8922, B => n8923, ZN => n10810);
   U469 : NAND4_X1 port map( A1 => n4146, A2 => n10527, A3 => n10526, A4 => 
                           n10838, ZN => n11747);
   U940 : AND3_X1 port map( A1 => n11080, A2 => n11079, A3 => n11078, ZN => 
                           n12270);
   U408 : AOI21_X1 port map( B1 => n10807, B2 => n7814, A => n6347, ZN => 
                           n12145);
   U783 : NAND2_X1 port map( A1 => n139, A2 => n5902, ZN => n11951);
   U2007 : INV_X1 port map( A => n11473, ZN => n431);
   U3073 : OR2_X1 port map( A1 => n12148, A2 => n5636, ZN => n12559);
   U233 : XNOR2_X1 port map( A => n12854, B => n13484, ZN => n13347);
   U18835 : XNOR2_X1 port map( A => n13477, B => n13476, ZN => n13719);
   U3028 : XNOR2_X1 port map( A => n11511, B => n11510, ZN => n14240);
   U17990 : XNOR2_X1 port map( A => n12393, B => n12392, ZN => n14406);
   U282 : INV_X1 port map( A => n12607, ZN => n14294);
   U854 : OR2_X1 port map( A1 => n14165, A2 => n14484, ZN => n14483);
   U404 : NOR2_X1 port map( A1 => n14483, A2 => n14164, ZN => n14660);
   U10190 : NOR2_X1 port map( A1 => n14290, A2 => n14289, ZN => n15054);
   U2968 : NAND3_X1 port map( A1 => n6234, A2 => n6235, A3 => n6233, ZN => 
                           n15370);
   U836 : BUF_X1 port map( A => n14600, Z => n14845);
   U1347 : MUX2_X1 port map( A => n13940, B => n13939, S => n14253, Z => n15300
                           );
   U5630 : AOI22_X1 port map( A1 => n13960, A2 => n13959, B1 => n13961, B2 => 
                           n14437, ZN => n15323);
   U186 : NAND3_X1 port map( A1 => n2742, A2 => n2745, A3 => n2743, ZN => 
                           n15790);
   U342 : AND3_X1 port map( A1 => n36, A2 => n5093, A3 => n5092, ZN => n16393);
   U973 : XNOR2_X1 port map( A => n15604, B => n15603, ZN => n17386);
   U474 : XNOR2_X1 port map( A => n4215, B => n15614, ZN => n16878);
   U10808 : XNOR2_X1 port map( A => n3677, B => n5828, ZN => n17261);
   U19212 : XNOR2_X1 port map( A => n14028, B => n14027, ZN => n17428);
   U567 : XNOR2_X1 port map( A => n15573, B => n15574, ZN => n17155);
   U511 : BUF_X1 port map( A => n17255, Z => n1880);
   U241 : AND3_X2 port map( A1 => n6800, A2 => n6799, A3 => n5986, ZN => n18506
                           );
   U14303 : CLKBUF_X1 port map( A => n16693, Z => n17948);
   U2735 : BUF_X2 port map( A => n16685, Z => n514);
   U904 : BUF_X1 port map( A => n15810, Z => n18064);
   U1090 : NAND3_X1 port map( A1 => n1480, A2 => n4244, A3 => n4191, ZN => 
                           n19534);
   U40 : AND3_X1 port map( A1 => n1170, A2 => n3933, A3 => n3931, ZN => n19243)
                           ;
   U8922 : AOI22_X1 port map( A1 => n17748, A2 => n3239, B1 => n17747, B2 => 
                           n18195, ZN => n18856);
   U5418 : OAI211_X1 port map( C1 => n1759, C2 => n1758, A => n17247, B => 
                           n4761, ZN => n19246);
   U9607 : NAND4_X1 port map( A1 => n17578, A2 => n3086, A3 => n3085, A4 => 
                           n3084, ZN => n19373);
   U609 : AOI22_X1 port map( A1 => n18103, A2 => n18104, B1 => n1143, B2 => 
                           n106, ZN => n19004);
   U1323 : NAND2_X1 port map( A1 => n6342, A2 => n16873, ZN => n19686);
   U2639 : AND2_X1 port map( A1 => n5492, A2 => n19172, ZN => n19692);
   U2652 : INV_X1 port map( A => n19245, ZN => n19348);
   U1563 : XNOR2_X1 port map( A => n4339, B => n18086, ZN => n20205);
   U1149 : AOI21_X1 port map( B1 => n6261, B2 => n20546, A => n19958, ZN => 
                           n20392);
   U1550 : NAND2_X1 port map( A1 => n3473, A2 => n19821, ZN => n21495);
   U1289 : AOI21_X1 port map( B1 => n20195, B2 => n20821, A => n20824, ZN => 
                           n21677);
   U1381 : AND2_X1 port map( A1 => n20891, A2 => n20890, ZN => n21087);
   U2542 : OR2_X1 port map( A1 => n2529, A2 => n2528, ZN => n20688);
   U12584 : NAND3_X1 port map( A1 => n5252, A2 => n19881, A3 => n5253, ZN => 
                           n21713);
   U883 : OAI22_X1 port map( A1 => n28797, A2 => n21039, B1 => n21038, B2 => 
                           n21037, ZN => n21903);
   U2485 : AND3_X1 port map( A1 => n1940, A2 => n2041, A3 => n1948, ZN => 
                           n22194);
   U881 : AND3_X1 port map( A1 => n658, A2 => n5128, A3 => n656, ZN => n22898);
   U6159 : XNOR2_X1 port map( A => n22643, B => n22898, ZN => n22481);
   U1669 : XNOR2_X1 port map( A => n20708, B => n20709, ZN => n23351);
   U197 : OAI21_X1 port map( B1 => n23401, B2 => n23402, A => n23400, ZN => 
                           n24077);
   U14074 : MUX2_X1 port map( A => n24158, B => n24157, S => n28512, Z => 
                           n26041);
   U12962 : AND3_X1 port map( A1 => n5654, A2 => n5655, A3 => n5653, ZN => 
                           n25714);
   U519 : XNOR2_X1 port map( A => n5755, B => n5754, ZN => n27700);
   U13844 : XNOR2_X1 port map( A => n25058, B => n25057, ZN => n26172);
   U5574 : BUF_X1 port map( A => n26436, Z => n26940);
   U8458 : NAND4_X1 port map( A1 => n27135, A2 => n27134, A3 => n27133, A4 => 
                           n27132, ZN => n27744);
   U1358 : AND2_X1 port map( A1 => n26521, A2 => n26520, ZN => n26641);
   U1384 : AND2_X1 port map( A1 => n3376, A2 => n3397, ZN => n27591);
   U970 : AND3_X1 port map( A1 => n26486, A2 => n26488, A3 => n26487, ZN => 
                           n27427);
   U853 : NOR2_X1 port map( A1 => n27877, A2 => n26539, ZN => n27313);
   U3484 : CLKBUF_X1 port map( A => Key(1), Z => n27462);
   U3456 : CLKBUF_X1 port map( A => Key(117), Z => n3385);
   U760 : CLKBUF_X1 port map( A => Key(166), Z => n135);
   U5163 : NOR2_X1 port map( A1 => n9184, A2 => n9007, ZN => n2250);
   U3364 : INV_X1 port map( A => n9425, ZN => n604);
   U661 : AND2_X1 port map( A1 => n8109, A2 => n9041, ZN => n9042);
   U8339 : AND2_X1 port map( A1 => n7490, A2 => n9084, ZN => n8724);
   U999 : NAND2_X1 port map( A1 => n8483, A2 => n8484, ZN => n10250);
   U3239 : INV_X1 port map( A => n11000, ZN => n592);
   U2014 : INV_X1 port map( A => n10687, ZN => n10959);
   U1106 : CLKBUF_X1 port map( A => n10668, Z => n11048);
   U10428 : AND2_X1 port map( A1 => n11881, A2 => n11875, ZN => n11883);
   U1362 : AOI22_X1 port map( A1 => n2430, A2 => n10870, B1 => n1630, B2 => 
                           n11883, ZN => n13195);
   U4337 : NAND3_X1 port map( A1 => n3020, A2 => n3021, A3 => n11513, ZN => 
                           n13137);
   U19201 : INV_X1 port map( A => n14132, ZN => n14341);
   U11243 : INV_X1 port map( A => n5584, ZN => n14411);
   U13346 : INV_X1 port map( A => n13920, ZN => n14033);
   U612 : BUF_X1 port map( A => n13677, Z => n14466);
   U1457 : OAI21_X1 port map( B1 => n13813, B2 => n14411, A => n5542, ZN => 
                           n14904);
   U744 : NAND3_X1 port map( A1 => n6433, A2 => n13712, A3 => n13713, ZN => 
                           n15135);
   U1963 : INV_X1 port map( A => n17389, ZN => n424);
   U20851 : BUF_X1 port map( A => n16712, Z => n17379);
   U10285 : NOR2_X1 port map( A1 => n16803, A2 => n17474, ZN => n17475);
   U536 : AND3_X1 port map( A1 => n16972, A2 => n16971, A3 => n17267, ZN => 
                           n18285);
   U6061 : INV_X1 port map( A => n18476, ZN => n18480);
   U4403 : OAI211_X1 port map( C1 => n17950, C2 => n17906, A => n17949, B => 
                           n6387, ZN => n19622);
   U2670 : OAI211_X1 port map( C1 => n18423, C2 => n18044, A => n5496, B => 
                           n5495, ZN => n19389);
   U2492 : OR2_X1 port map( A1 => n21227, A2 => n21632, ZN => n21036);
   U8131 : INV_X1 port map( A => n23789, ZN => n23792);
   U1118 : OR2_X1 port map( A1 => n23375, A2 => n24072, ZN => n205);
   U155 : OR2_X1 port map( A1 => n23916, A2 => n23917, ZN => n985);
   U26486 : XNOR2_X1 port map( A => n25554, B => n25553, ZN => n27044);
   U4317 : XNOR2_X1 port map( A => n25496, B => n25497, ZN => n27013);
   U14388 : NAND2_X1 port map( A1 => n26623, A2 => n27013, ZN => n26624);
   U26586 : AOI22_X1 port map( A1 => n26217, A2 => n28459, B1 => n26210, B2 => 
                           n25661, ZN => n25664);
   U11169 : AND2_X2 port map( A1 => n3928, A2 => n3927, ZN => n15343);
   U9574 : OR2_X2 port map( A1 => n7699, A2 => n7698, ZN => n9034);
   U4450 : AND3_X2 port map( A1 => n3709, A2 => n3823, A3 => n3825, ZN => 
                           n19228);
   U3816 : OR2_X2 port map( A1 => n24336, A2 => n24337, ZN => n24341);
   U624 : BUF_X2 port map( A => n14061, Z => n14064);
   U708 : OR2_X2 port map( A1 => n8172, A2 => n8171, ZN => n8984);
   U2251 : BUF_X2 port map( A => n26518, Z => n27138);
   U1333 : MUX2_X2 port map( A => n15450, B => n15449, S => n15448, Z => n16557
                           );
   U779 : OR2_X2 port map( A1 => n19918, A2 => n19917, ZN => n21875);
   U543 : AND2_X2 port map( A1 => n4209, A2 => n3402, ZN => n18913);
   U11200 : AND3_X2 port map( A1 => n3956, A2 => n3960, A3 => n3955, ZN => 
                           n13175);
   U11407 : OAI21_X2 port map( B1 => n10862, B2 => n11512, A => n4140, ZN => 
                           n12566);
   U13213 : AND3_X2 port map( A1 => n5906, A2 => n5908, A3 => n5907, ZN => 
                           n19251);
   U17368 : AOI21_X2 port map( B1 => n11327, B2 => n11328, A => n11326, ZN => 
                           n11801);
   U4110 : XNOR2_X2 port map( A => n19515, B => n19514, ZN => n20299);
   U72 : OAI211_X2 port map( C1 => n15507, C2 => n15506, A => n15505, B => 
                           n15504, ZN => n16607);
   U1105 : AND3_X2 port map( A1 => n14130, A2 => n14129, A3 => n14128, ZN => 
                           n14752);
   U8465 : XNOR2_X2 port map( A => Key(111), B => Plaintext(111), ZN => n7626);
   U8079 : AND3_X2 port map( A1 => n2049, A2 => n20984, A3 => n21812, ZN => 
                           n22713);
   U4045 : NAND2_X2 port map( A1 => n910, A2 => n5547, ZN => n23467);
   U3426 : BUF_X1 port map( A => n7017, Z => n8245);
   U1101 : OR2_X2 port map( A1 => n8684, A2 => n8683, ZN => n9949);
   U1697 : NAND2_X2 port map( A1 => n6444, A2 => n6443, ZN => n19025);
   U2035 : MUX2_X2 port map( A => n7820, B => n7819, S => n8243, Z => n9016);
   U938 : OR2_X2 port map( A1 => n17585, A2 => n1376, ZN => n19245);
   U849 : AND2_X2 port map( A1 => n17705, A2 => n17704, ZN => n19603);
   U10806 : NAND3_X2 port map( A1 => n3676, A2 => n3675, A3 => n7227, ZN => 
                           n9971);
   U9935 : MUX2_X2 port map( A => n7081, B => n7080, S => n8812, Z => n10037);
   U1437 : NAND2_X2 port map( A1 => n5034, A2 => n5033, ZN => n21932);
   U348 : NAND2_X2 port map( A1 => n2678, A2 => n10857, ZN => n12241);
   U10408 : MUX2_X2 port map( A => n26839, B => n26838, S => n26837, Z => 
                           n27843);
   U24797 : OR2_X2 port map( A1 => n22983, A2 => n22982, ZN => n24433);
   U1533 : BUF_X2 port map( A => n8847, Z => n12205);
   U2465 : AND3_X2 port map( A1 => n20796, A2 => n20795, A3 => n20794, ZN => 
                           n22790);
   U12 : MUX2_X2 port map( A => n24371, B => n24370, S => n24369, Z => n25430);
   U4745 : NAND3_X2 port map( A1 => n23439, A2 => n1228, A3 => n23438, ZN => 
                           n24256);
   U1568 : BUF_X1 port map( A => n20224, Z => n296);
   U684 : NAND2_X2 port map( A1 => n11296, A2 => n3556, ZN => n12841);
   U11437 : NAND2_X2 port map( A1 => n26934, A2 => n6950, ZN => n27527);
   U2043 : XNOR2_X2 port map( A => n7138, B => Key(48), ZN => n8013);
   U10033 : NAND2_X2 port map( A1 => n24333, A2 => n3696, ZN => n26059);
   U3215 : XNOR2_X2 port map( A => n9804, B => n9803, ZN => n10992);
   U22792 : MUX2_X2 port map( A => n19862, B => n19861, S => n385, Z => n20744)
                           ;
   U19927 : OAI211_X2 port map( C1 => n15495, C2 => n15494, A => n15493, B => 
                           n15492, ZN => n16309);
   U9185 : OAI21_X2 port map( B1 => n8743, B2 => n8742, A => n2859, ZN => 
                           n10265);
   U8068 : NOR2_X1 port map( A1 => n7569, A2 => n8326, ZN => n8581);
   U1548 : AOI21_X2 port map( B1 => n9145, B2 => n9144, A => n9143, ZN => 
                           n10159);
   U3202 : BUF_X1 port map( A => n10482, Z => n11258);
   U5280 : AND2_X1 port map( A1 => n1663, A2 => n11974, ZN => n1664);
   U1754 : BUF_X1 port map( A => n18522, Z => n374);
   U2570 : OAI21_X1 port map( B1 => n20694, B2 => n6730, A => n20693, ZN => 
                           n21810);
   U5902 : BUF_X1 port map( A => n23702, Z => n23387);
   U4140 : NAND3_X1 port map( A1 => n24342, A2 => n2460, A3 => n24343, ZN => 
                           n25697);
   U47 : XNOR2_X1 port map( A => n6447, B => n16080, ZN => n16812);
   U77 : BUF_X1 port map( A => n8151, Z => n28149);
   U118 : NAND3_X2 port map( A1 => n28306, A2 => n15038, A3 => n28305, ZN => 
                           n15989);
   U126 : NAND3_X2 port map( A1 => n4550, A2 => n4551, A3 => n7826, ZN => n9012
                           );
   U135 : NAND3_X2 port map( A1 => n28707, A2 => n3499, A3 => n5387, ZN => 
                           n24697);
   U194 : OAI21_X2 port map( B1 => n19857, B2 => n20556, A => n19856, ZN => 
                           n21481);
   U216 : BUF_X1 port map( A => n1308, Z => n28407);
   U235 : OR2_X2 port map( A1 => n14269, A2 => n14270, ZN => n15260);
   U293 : XNOR2_X1 port map( A => n26064, B => n26063, ZN => n27111);
   U307 : OAI21_X2 port map( B1 => n4351, B2 => n10871, A => n4350, ZN => 
                           n12236);
   U323 : AND3_X2 port map( A1 => n3023, A2 => n4045, A3 => n4171, ZN => n11430
                           );
   U335 : XNOR2_X1 port map( A => n12458, B => n12457, ZN => n14416);
   U353 : NOR2_X1 port map( A1 => n14036, A2 => n13719, ZN => n28121);
   U378 : XOR2_X1 port map( A => n21492, B => n21491, Z => n28122);
   U383 : XNOR2_X2 port map( A => n24522, B => n4643, ZN => n28578);
   U396 : INV_X1 port map( A => n17696, ZN => n16898);
   U429 : XNOR2_X1 port map( A => n19432, B => n19431, ZN => n21355);
   U444 : NAND2_X2 port map( A1 => n4609, A2 => n4608, ZN => n14733);
   U471 : XNOR2_X2 port map( A => n4764, B => n25928, ZN => n25412);
   U500 : NOR2_X2 port map( A1 => n20596, A2 => n20595, ZN => n21801);
   U507 : OAI21_X2 port map( B1 => n7578, B2 => n7577, A => n7576, ZN => n8717)
                           ;
   U525 : BUF_X2 port map( A => n21356, Z => n28133);
   U527 : XNOR2_X1 port map( A => n19437, B => n19436, ZN => n21356);
   U551 : XNOR2_X2 port map( A => n25098, B => n25097, ZN => n26799);
   U562 : XNOR2_X2 port map( A => n9093, B => n9092, ZN => n11192);
   U566 : XNOR2_X2 port map( A => n15628, B => n15627, ZN => n17359);
   U587 : XNOR2_X1 port map( A => n22049, B => n22048, ZN => n23250);
   U592 : NOR2_X2 port map( A1 => n13313, A2 => n13312, ZN => n16346);
   U601 : XNOR2_X2 port map( A => n6074, B => n21757, ZN => n23036);
   U608 : OAI21_X2 port map( B1 => n17778, B2 => n17980, A => n6264, ZN => 
                           n19685);
   U623 : AOI21_X2 port map( B1 => n26249, B2 => n26248, A => n26247, ZN => 
                           n28065);
   U634 : OAI211_X2 port map( C1 => n21187, C2 => n22288, A => n1694, B => 
                           n1692, ZN => n22690);
   U636 : OR2_X2 port map( A1 => n3486, A2 => n21592, ZN => n21998);
   U670 : OAI21_X2 port map( B1 => n18627, B2 => n20381, A => n18626, ZN => 
                           n21218);
   U695 : NOR2_X2 port map( A1 => n20898, A2 => n20897, ZN => n1925);
   U697 : XNOR2_X2 port map( A => n13047, B => n13046, ZN => n14354);
   U718 : XNOR2_X2 port map( A => n15820, B => n15821, ZN => n17555);
   U721 : OAI21_X2 port map( B1 => n7923, B2 => n8234, A => n7922, ZN => n9108)
                           ;
   U735 : OR2_X2 port map( A1 => n20138, A2 => n20139, ZN => n21425);
   U746 : NOR2_X1 port map( A1 => n17010, A2 => n17011, ZN => n18601);
   U753 : INV_X1 port map( A => n13842, ZN => n14345);
   U756 : NOR2_X1 port map( A1 => n18543, A2 => n28339, ZN => n19556);
   U757 : AND2_X2 port map( A1 => n11134, A2 => n11775, ZN => n11551);
   U766 : BUF_X2 port map( A => n20354, Z => n383);
   U778 : XNOR2_X2 port map( A => n13515, B => n13514, ZN => n13587);
   U785 : NOR2_X2 port map( A1 => n3243, A2 => n19975, ZN => n21956);
   U794 : CLKBUF_X1 port map( A => n11275, Z => n28147);
   U831 : XNOR2_X2 port map( A => n4747, B => n4745, ZN => n20494);
   U857 : AND3_X2 port map( A1 => n23379, A2 => n23381, A3 => n23380, ZN => 
                           n25933);
   U882 : XNOR2_X2 port map( A => n25286, B => n25285, ZN => n26723);
   U896 : XNOR2_X2 port map( A => n7105, B => Key(186), ZN => n7312);
   U905 : INV_X1 port map( A => n10544, ZN => n10742);
   U911 : AND3_X2 port map( A1 => n1105, A2 => n19919, A3 => n4658, ZN => 
                           n20658);
   U964 : XNOR2_X2 port map( A => n6980, B => Key(96), ZN => n7828);
   U968 : XNOR2_X2 port map( A => n23861, B => n23860, ZN => n25418);
   U1058 : XNOR2_X2 port map( A => n7003, B => Key(72), ZN => n7250);
   U1067 : NAND2_X2 port map( A1 => n5619, A2 => n5618, ZN => n24408);
   U1077 : OAI211_X2 port map( C1 => n8823, C2 => n7529, A => n8475, B => n7528
                           , ZN => n10395);
   U1091 : BUF_X2 port map( A => n21565, Z => n28155);
   U1096 : OAI211_X1 port map( C1 => n19792, C2 => n20488, A => n5208, B => 
                           n2383, ZN => n21565);
   U1143 : CLKBUF_X1 port map( A => n7141, Z => n28161);
   U1155 : AOI22_X2 port map( A1 => n2220, A2 => n11750, B1 => n28698, B2 => 
                           n11501, ZN => n12965);
   U1183 : NOR3_X1 port map( A1 => n20428, A2 => n20427, A3 => n20426, ZN => 
                           n22765);
   U1203 : XNOR2_X2 port map( A => n15540, B => n15539, ZN => n17025);
   U1207 : AND3_X2 port map( A1 => n17468, A2 => n3981, A3 => n3980, ZN => 
                           n18500);
   U1228 : AND2_X2 port map( A1 => n1539, A2 => n1542, ZN => n22522);
   U1281 : INV_X1 port map( A => n10830, ZN => n11338);
   U1305 : NOR2_X2 port map( A1 => n24026, A2 => n24025, ZN => n4764);
   U1324 : AND2_X2 port map( A1 => n4177, A2 => n3204, ZN => n24405);
   U1325 : OAI211_X2 port map( C1 => n12587, C2 => n13711, A => n12586, B => 
                           n12585, ZN => n15094);
   U1326 : OAI211_X2 port map( C1 => n3880, C2 => n1581, A => n3878, B => n3879
                           , ZN => n18421);
   U1342 : AND2_X2 port map( A1 => n2942, A2 => n2941, ZN => n9140);
   U1348 : AOI21_X2 port map( B1 => n21234, B2 => n21389, A => n21233, ZN => 
                           n22195);
   U1353 : XNOR2_X2 port map( A => n19471, B => n19470, ZN => n20443);
   U1364 : OAI21_X2 port map( B1 => n5863, B2 => n24146, A => n24145, ZN => 
                           n25391);
   U1391 : XNOR2_X2 port map( A => n4430, B => n5184, ZN => n4086);
   U1393 : OAI22_X2 port map( A1 => n4661, A2 => n4660, B1 => n14580, B2 => 
                           n15095, ZN => n16494);
   U1394 : XNOR2_X2 port map( A => n9288, B => n9287, ZN => n10942);
   U1415 : XNOR2_X2 port map( A => n12530, B => n12531, ZN => n13872);
   U1422 : AOI21_X2 port map( B1 => n792, B2 => n17226, A => n4763, ZN => 
                           n18431);
   U1488 : BUF_X2 port map( A => n24074, Z => n24072);
   U1529 : AND2_X1 port map( A1 => n17423, A2 => n17421, ZN => n28739);
   U1530 : BUF_X1 port map( A => n17452, Z => n28193);
   U1532 : BUF_X1 port map( A => n15980, Z => n17275);
   U1545 : INV_X1 port map( A => n13730, ZN => n28171);
   U1559 : INV_X1 port map( A => n10957, ZN => n28173);
   U1572 : INV_X1 port map( A => n11045, ZN => n28174);
   U1573 : INV_X1 port map( A => n11158, ZN => n28175);
   U1574 : INV_X1 port map( A => n10703, ZN => n28176);
   U1579 : AND2_X1 port map( A1 => n9196, A2 => n9197, ZN => n231);
   U1608 : AND3_X1 port map( A1 => n2432, A2 => n28341, A3 => n2434, ZN => 
                           n27220);
   U1609 : AOI22_X1 port map( A1 => n29021, A2 => n27958, B1 => n29092, B2 => 
                           n27996, ZN => n27998);
   U1611 : NAND3_X1 port map( A1 => n27009, A2 => n27008, A3 => n27007, ZN => 
                           n27926);
   U1613 : OAI21_X1 port map( B1 => n24857, B2 => n4679, A => n24856, ZN => 
                           n28466);
   U1625 : AND3_X1 port map( A1 => n28216, A2 => n28238, A3 => n28237, ZN => 
                           n27800);
   U1632 : INV_X1 port map( A => n27594, ZN => n28179);
   U1634 : OR3_X1 port map( A1 => n26129, A2 => n28392, A3 => n27129, ZN => 
                           n27135);
   U1644 : XNOR2_X1 port map( A => n25478, B => n28230, ZN => n26623);
   U1645 : INV_X1 port map( A => n29474, ZN => n28180);
   U1657 : AND2_X1 port map( A1 => n24102, A2 => n24101, ZN => n28256);
   U1658 : NOR2_X1 port map( A1 => n22177, A2 => n24468, ZN => n22178);
   U1659 : OR2_X1 port map( A1 => n24583, A2 => n24584, ZN => n28315);
   U1663 : BUF_X1 port map( A => n24790, Z => n28512);
   U1673 : OR2_X1 port map( A1 => n29567, A2 => n24391, ZN => n2648);
   U1676 : CLKBUF_X1 port map( A => n24717, Z => n28416);
   U1679 : AND4_X1 port map( A1 => n6154, A2 => n4234, A3 => n4233, A4 => n6153
                           , ZN => n28509);
   U1680 : AND2_X1 port map( A1 => n23783, A2 => n23787, ZN => n21769);
   U1684 : OR2_X1 port map( A1 => n23772, A2 => n23771, ZN => n23021);
   U1692 : INV_X1 port map( A => n22566, ZN => n28181);
   U1698 : XNOR2_X1 port map( A => n22850, B => n22849, ZN => n28609);
   U1699 : OR2_X1 port map( A1 => n23769, A2 => n23763, ZN => n28354);
   U1702 : INV_X1 port map( A => n23725, ZN => n28183);
   U1717 : AOI22_X1 port map( A1 => n28750, A2 => n28749, B1 => n22012, B2 => 
                           n20537, ZN => n20798);
   U1718 : INV_X1 port map( A => n21068, ZN => n28301);
   U1719 : INV_X1 port map( A => n20853, ZN => n20852);
   U1723 : OR2_X1 port map( A1 => n21581, A2 => n21481, ZN => n28723);
   U1729 : BUF_X1 port map( A => n21343, Z => n28440);
   U1730 : INV_X1 port map( A => n20663, ZN => n28184);
   U1734 : INV_X1 port map( A => n21541, ZN => n28185);
   U1736 : OAI21_X1 port map( B1 => n2715, B2 => n18831, A => n19773, ZN => 
                           n28326);
   U1738 : INV_X1 port map( A => n20162, ZN => n28187);
   U1742 : INV_X1 port map( A => n20099, ZN => n28188);
   U1746 : XNOR2_X1 port map( A => n6157, B => n19135, ZN => n20506);
   U1755 : INV_X1 port map( A => n19413, ZN => n18628);
   U1764 : NOR2_X1 port map( A1 => n17724, A2 => n373, ZN => n19659);
   U1765 : OR2_X1 port map( A1 => n18291, A2 => n18292, ZN => n3768);
   U1767 : INV_X1 port map( A => n18493, ZN => n18487);
   U1777 : OR2_X1 port map( A1 => n18387, A2 => n18393, ZN => n686);
   U1787 : OR2_X1 port map( A1 => n4732, A2 => n526, ZN => n17330);
   U1794 : OR2_X1 port map( A1 => n18193, A2 => n16718, ZN => n1025);
   U1796 : NAND2_X1 port map( A1 => n1592, A2 => n1591, ZN => n18493);
   U1801 : OR2_X1 port map( A1 => n526, A2 => n18144, ZN => n193);
   U1803 : INV_X1 port map( A => n17762, ZN => n28191);
   U1848 : OR2_X1 port map( A1 => n28323, A2 => n4270, ZN => n2858);
   U1880 : AND2_X1 port map( A1 => n17355, A2 => n17357, ZN => n16713);
   U1889 : XNOR2_X1 port map( A => n15699, B => n15700, ZN => n17368);
   U1893 : INV_X1 port map( A => n17426, ZN => n28194);
   U1947 : INV_X1 port map( A => n14942, ZN => n28195);
   U1991 : AND2_X1 port map( A1 => n12414, A2 => n12415, ZN => n14906);
   U2008 : INV_X1 port map( A => n15060, ZN => n28197);
   U2021 : INV_X1 port map( A => n14695, ZN => n28198);
   U2031 : OR2_X1 port map( A1 => n28569, A2 => n13587, ZN => n28257);
   U2104 : INV_X1 port map( A => n13703, ZN => n28199);
   U2144 : INV_X1 port map( A => n14438, ZN => n28200);
   U2148 : INV_X1 port map( A => n12696, ZN => n12861);
   U2174 : NAND3_X1 port map( A1 => n28682, A2 => n3987, A3 => n11391, ZN => 
                           n4474);
   U2201 : OR2_X1 port map( A1 => n12081, A2 => n3558, ZN => n28703);
   U2249 : INV_X1 port map( A => n12232, ZN => n28201);
   U2255 : INV_X1 port map( A => n12211, ZN => n28203);
   U2258 : AND2_X1 port map( A1 => n4352, A2 => n10666, ZN => n28363);
   U2259 : INV_X1 port map( A => n10668, ZN => n28204);
   U2263 : INV_X1 port map( A => n11113, ZN => n28205);
   U2281 : INV_X1 port map( A => n11145, ZN => n28206);
   U2286 : XNOR2_X1 port map( A => n6891, B => n9309, ZN => n28608);
   U2307 : INV_X1 port map( A => n10467, ZN => n28208);
   U2345 : AND3_X1 port map( A1 => n1045, A2 => n28352, A3 => n5130, ZN => 
                           n9323);
   U2357 : AOI21_X1 port map( B1 => n9419, B2 => n604, A => n9420, ZN => n2290)
                           ;
   U2414 : INV_X1 port map( A => n9028, ZN => n28210);
   U2422 : INV_X1 port map( A => n8109, ZN => n28211);
   U2442 : INV_X1 port map( A => n9075, ZN => n28212);
   U2446 : OR2_X1 port map( A1 => n6988, A2 => n7822, ZN => n7426);
   U2452 : OR2_X1 port map( A1 => n7935, A2 => n7933, ZN => n7616);
   U2466 : INV_X1 port map( A => n3154, ZN => n28213);
   U2467 : CLKBUF_X1 port map( A => Key(172), Z => n28294);
   U2503 : INV_X1 port map( A => n7822, ZN => n3821);
   U2526 : INV_X1 port map( A => n441, ZN => n7870);
   U2544 : OAI21_X1 port map( B1 => n627, B2 => n8217, A => n7925, ZN => n6961)
                           ;
   U2557 : BUF_X1 port map( A => n7093, Z => n7309);
   U2565 : OR2_X1 port map( A1 => n9009, A2 => n9007, ZN => n9189);
   U2585 : INV_X1 port map( A => n8440, ZN => n28743);
   U2590 : OR2_X1 port map( A1 => n7952, A2 => n8258, ZN => n117);
   U2603 : AND3_X1 port map( A1 => n1418, A2 => n1417, A3 => n7574, ZN => 
                           n28281);
   U2605 : OR2_X1 port map( A1 => n8351, A2 => n8353, ZN => n238);
   U2620 : BUF_X1 port map( A => n7665, Z => n8265);
   U2656 : NAND2_X1 port map( A1 => n4673, A2 => n4674, ZN => n8192);
   U2657 : OR2_X1 port map( A1 => n8976, A2 => n8819, ZN => n142);
   U2660 : OR2_X1 port map( A1 => n10406, A2 => n3787, ZN => n2891);
   U2674 : OR2_X1 port map( A1 => n8575, A2 => n9421, ZN => n28352);
   U2684 : OR2_X1 port map( A1 => n9139, A2 => n8185, ZN => n8187);
   U2710 : AOI21_X1 port map( B1 => n8738, B2 => n8731, A => n8730, ZN => n8374
                           );
   U2717 : AND2_X1 port map( A1 => n8702, A2 => n8700, ZN => n105);
   U2747 : INV_X1 port map( A => n8077, ZN => n8431);
   U2756 : NOR2_X1 port map( A1 => n8491, A2 => n8666, ZN => n8495);
   U2792 : OR2_X1 port map( A1 => n8598, A2 => n9062, ZN => n8402);
   U2799 : XNOR2_X1 port map( A => n9635, B => n9634, ZN => n11047);
   U2822 : OR2_X1 port map( A1 => n10942, A2 => n10703, ZN => n28310);
   U2831 : MUX2_X1 port map( A => n11034, B => n10671, S => n28147, Z => n10672
                           );
   U2836 : NOR2_X1 port map( A1 => n11106, A2 => n10871, ZN => n10280);
   U2855 : INV_X1 port map( A => n10482, ZN => n4296);
   U2886 : NOR2_X1 port map( A1 => n4389, A2 => n10741, ZN => n4390);
   U2900 : XNOR2_X1 port map( A => n2662, B => n1988, ZN => n10930);
   U2927 : AND2_X1 port map( A1 => n6703, A2 => n2063, ZN => n28336);
   U2932 : AND2_X1 port map( A1 => n11888, A2 => n12328, ZN => n28260);
   U2934 : OR2_X1 port map( A1 => n349, A2 => n11933, ZN => n11594);
   U2935 : INV_X1 port map( A => n11377, ZN => n12167);
   U2959 : OAI211_X1 port map( C1 => n11799, C2 => n12289, A => n11798, B => 
                           n11797, ZN => n12734);
   U2975 : INV_X1 port map( A => n12589, ZN => n13539);
   U2981 : AND2_X1 port map( A1 => n14295, A2 => n14293, ZN => n28322);
   U2983 : AND2_X1 port map( A1 => n14304, A2 => n5341, ZN => n28273);
   U2986 : XNOR2_X1 port map( A => n11866, B => n11865, ZN => n14252);
   U3037 : OAI21_X1 port map( B1 => n12122, B2 => n12121, A => n14487, ZN => 
                           n141);
   U3044 : NAND2_X1 port map( A1 => n1389, A2 => n57, ZN => n14971);
   U3085 : OR2_X1 port map( A1 => n14583, A2 => n14971, ZN => n14886);
   U3098 : OAI211_X1 port map( C1 => n13651, C2 => n14302, A => n13650, B => 
                           n13649, ZN => n15117);
   U3116 : OR2_X1 port map( A1 => n15351, A2 => n15343, ZN => n150);
   U3147 : CLKBUF_X1 port map( A => n14826, Z => n15030);
   U3163 : AND2_X1 port map( A1 => n15009, A2 => n15370, ZN => n15376);
   U3170 : OAI21_X1 port map( B1 => n1662, B2 => n15376, A => n15371, ZN => n5)
                           ;
   U3191 : XNOR2_X1 port map( A => n6080, B => n16494, ZN => n15903);
   U3214 : AND2_X1 port map( A1 => n5714, A2 => n17304, ZN => n28233);
   U3228 : NOR2_X1 port map( A1 => n28233, A2 => n16968, ZN => n28232);
   U3265 : OR2_X1 port map( A1 => n17139, A2 => n16887, ZN => n17135);
   U3279 : NOR2_X1 port map( A1 => n16706, A2 => n16884, ZN => n16430);
   U3303 : AND2_X1 port map( A1 => n18181, A2 => n18180, ZN => n17738);
   U3342 : OR2_X1 port map( A1 => n517, A2 => n17762, ZN => n66);
   U3412 : OR2_X1 port map( A1 => n1384, A2 => n18467, ZN => n17917);
   U3420 : AND2_X1 port map( A1 => n18458, A2 => n18106, ZN => n28241);
   U3496 : OR2_X1 port map( A1 => n2853, A2 => n18430, ZN => n18147);
   U3502 : BUF_X1 port map( A => n18708, Z => n28558);
   U3507 : OR2_X1 port map( A1 => n17814, A2 => n420, ZN => n17247);
   U3518 : INV_X1 port map( A => n18423, ZN => n512);
   U3519 : OR2_X1 port map( A1 => n5203, A2 => n18171, ZN => n17785);
   U3532 : XNOR2_X1 port map( A => n18737, B => n19475, ZN => n19040);
   U3541 : OR2_X1 port map( A1 => n18019, A2 => n28370, ZN => n3070);
   U3570 : XNOR2_X1 port map( A => n18926, B => n18925, ZN => n28479);
   U3578 : AND2_X1 port map( A1 => n21088, A2 => n628, ZN => n28275);
   U3584 : NOR2_X1 port map( A1 => n20382, A2 => n28508, ZN => n20385);
   U3593 : OR2_X1 port map( A1 => n21227, A2 => n21392, ZN => n3418);
   U3615 : AND2_X1 port map( A1 => n21171, A2 => n21047, ZN => n28287);
   U3616 : OR2_X1 port map( A1 => n21144, A2 => n21118, ZN => n20853);
   U3641 : XNOR2_X1 port map( A => n1859, B => n5803, ZN => n22058);
   U3642 : OR2_X1 port map( A1 => n4104, A2 => n43, ZN => n4203);
   U3655 : AND3_X1 port map( A1 => n20532, A2 => n20933, A3 => n20533, ZN => 
                           n20426);
   U3682 : INV_X1 port map( A => n4872, ZN => n23150);
   U3701 : OR2_X1 port map( A1 => n23712, A2 => n22174, ZN => n22163);
   U3716 : NOR2_X1 port map( A1 => n23629, A2 => n23630, ZN => n23555);
   U3723 : XNOR2_X1 port map( A => n22115, B => n22114, ZN => n23726);
   U3729 : OR2_X1 port map( A1 => n23647, A2 => n2779, ZN => n640);
   U3739 : XNOR2_X1 port map( A => n22083, B => n22082, ZN => n23386);
   U3745 : XNOR2_X1 port map( A => n21104, B => n21105, ZN => n23360);
   U3760 : AND2_X1 port map( A1 => n23147, A2 => n23461, ZN => n4872);
   U3772 : OR2_X1 port map( A1 => n23465, A2 => n22926, ZN => n28317);
   U3850 : OR2_X1 port map( A1 => n23388, A2 => n23704, ZN => n28695);
   U3856 : OR2_X1 port map( A1 => n22867, A2 => n22866, ZN => n28519);
   U3866 : OR2_X1 port map( A1 => n23373, A2 => n24316, ZN => n28681);
   U3871 : NOR2_X1 port map( A1 => n24816, A2 => n24461, ZN => n28678);
   U3893 : AND2_X1 port map( A1 => n23590, A2 => n24447, ZN => n28330);
   U3906 : XNOR2_X1 port map( A => n25693, B => n25692, ZN => n28545);
   U3912 : BUF_X1 port map( A => n26941, Z => n28541);
   U3943 : AOI21_X1 port map( B1 => n28289, B2 => n28288, A => n26352, ZN => 
                           n26354);
   U3994 : XNOR2_X1 port map( A => n25854, B => n25853, ZN => n26837);
   U4001 : NOR2_X1 port map( A1 => n25814, A2 => n27087, ZN => n28249);
   U4032 : NOR2_X1 port map( A1 => n27038, A2 => n27379, ZN => n26610);
   U4118 : AND3_X1 port map( A1 => n3390, A2 => n6634, A3 => n6633, ZN => 
                           n27548);
   U4131 : INV_X1 port map( A => n26696, ZN => n28248);
   U4135 : NAND3_X1 port map( A1 => n6755, A2 => n5391, A3 => n5390, ZN => 
                           n27244);
   U4144 : CLKBUF_X1 port map( A => Key(151), Z => n27105);
   U4146 : CLKBUF_X1 port map( A => Key(154), Z => n2510);
   U4151 : AND2_X1 port map( A1 => n29537, A2 => n26314, ZN => n28214);
   U4160 : NAND3_X1 port map( A1 => n29644, A2 => n20191, A3 => n20541, ZN => 
                           n28215);
   U4162 : OR3_X1 port map( A1 => n5299, A2 => n27060, A3 => n26849, ZN => 
                           n28216);
   U4190 : OR2_X1 port map( A1 => n28228, A2 => n29076, ZN => n28217);
   U4198 : INV_X1 port map( A => n7424, ZN => n28721);
   U4201 : AND2_X1 port map( A1 => n7837, A2 => n7700, ZN => n28218);
   U4202 : AND2_X1 port map( A1 => n7492, A2 => n8850, ZN => n28219);
   U4229 : INV_X1 port map( A => n10929, ZN => n10927);
   U4247 : INV_X1 port map( A => n12042, ZN => n28726);
   U4265 : AND2_X1 port map( A1 => n14455, A2 => n14200, ZN => n28220);
   U4266 : INV_X1 port map( A => n14696, ZN => n15288);
   U4268 : OR2_X1 port map( A1 => n15081, A2 => n15082, ZN => n28221);
   U4279 : NOR2_X1 port map( A1 => n14763, A2 => n15260, ZN => n28222);
   U4281 : INV_X1 port map( A => n17294, ZN => n28729);
   U4282 : INV_X1 port map( A => n15691, ZN => n28666);
   U4308 : INV_X1 port map( A => n18020, ZN => n28370);
   U4323 : NAND4_X2 port map( A1 => n4189, A2 => n4190, A3 => n6410, A4 => 
                           n6409, ZN => n22290);
   U4335 : OR2_X1 port map( A1 => n20657, A2 => n20656, ZN => n28223);
   U4351 : NAND3_X1 port map( A1 => n23326, A2 => n23034, A3 => n23760, ZN => 
                           n28224);
   U4360 : XOR2_X1 port map( A => n22191, B => n22190, Z => n28225);
   U4387 : XOR2_X1 port map( A => n24962, B => n24961, Z => n28226);
   U4393 : AND2_X1 port map( A1 => n24668, A2 => n24665, ZN => n28227);
   U4394 : XOR2_X1 port map( A => n25719, B => n25718, Z => n28228);
   U4421 : INV_X1 port map( A => n23862, ZN => n28710);
   U4423 : AND2_X1 port map( A1 => n29060, A2 => n29474, ZN => n28229);
   U4428 : XOR2_X1 port map( A => n25476, B => n25475, Z => n28230);
   U4511 : NAND2_X1 port map( A1 => n4543, A2 => n6053, ZN => n4542);
   U4550 : NAND2_X1 port map( A1 => n28232, A2 => n28231, ZN => n6224);
   U4551 : NAND2_X1 port map( A1 => n28768, A2 => n1738, ZN => n28231);
   U4572 : NAND2_X1 port map( A1 => n20377, A2 => n20371, ZN => n28235);
   U4583 : NAND2_X1 port map( A1 => n20376, A2 => n351, ZN => n28236);
   U4593 : NAND2_X1 port map( A1 => n26328, A2 => n28600, ZN => n28237);
   U4597 : NAND2_X1 port map( A1 => n26329, A2 => n27056, ZN => n28238);
   U4603 : NAND2_X1 port map( A1 => n6931, A2 => n19951, ZN => n28244);
   U4616 : NAND2_X1 port map( A1 => n28240, A2 => n20192, ZN => n3016);
   U4642 : NOR2_X1 port map( A1 => n503, A2 => n20416, ZN => n28240);
   U4651 : NAND3_X1 port map( A1 => n4033, A2 => n28393, A3 => n4236, ZN => 
                           n4032);
   U4664 : NAND2_X1 port map( A1 => n17729, A2 => n18109, ZN => n3849);
   U4710 : NAND2_X1 port map( A1 => n28242, A2 => n5822, ZN => n5820);
   U4733 : NAND2_X1 port map( A1 => n5804, A2 => n13935, ZN => n28242);
   U4741 : NAND2_X1 port map( A1 => n28243, A2 => n5943, ZN => n21581);
   U4742 : NAND3_X1 port map( A1 => n19839, A2 => n5100, A3 => n5099, ZN => 
                           n28243);
   U4764 : NOR2_X1 port map( A1 => n19953, A2 => n28244, ZN => n21729);
   U4767 : NAND3_X1 port map( A1 => n28641, A2 => n27862, A3 => n27324, ZN => 
                           n27325);
   U4778 : NAND2_X1 port map( A1 => n24241, A2 => n24559, ZN => n5332);
   U4786 : AOI21_X1 port map( B1 => n15267, B2 => n15266, A => n15506, ZN => 
                           n28245);
   U4925 : NAND2_X1 port map( A1 => n1483, A2 => n24780, ZN => n24781);
   U4945 : NAND2_X1 port map( A1 => n28246, A2 => n8204, ZN => n8206);
   U4977 : NOR2_X2 port map( A1 => n5289, A2 => n28247, ZN => n4384);
   U4996 : NOR2_X1 port map( A1 => n24058, A2 => n459, ZN => n28247);
   U4998 : OR2_X1 port map( A1 => n20381, A2 => n20573, ZN => n19834);
   U4999 : NAND3_X1 port map( A1 => n447, A2 => n3681, A3 => n28248, ZN => 
                           n26643);
   U5011 : NOR2_X2 port map( A1 => n25834, A2 => n28249, ZN => n27872);
   U5049 : NOR2_X2 port map( A1 => n28251, A2 => n28250, ZN => n18802);
   U5063 : OAI22_X1 port map( A1 => n18013, A2 => n18480, B1 => n18012, B2 => 
                           n18011, ZN => n28250);
   U5067 : NAND2_X1 port map( A1 => n6574, A2 => n6575, ZN => n28251);
   U5113 : NAND2_X1 port map( A1 => n28894, A2 => n20430, ZN => n28252);
   U5118 : NAND2_X1 port map( A1 => n24590, A2 => n831, ZN => n4692);
   U5131 : NAND2_X2 port map( A1 => n28317, A2 => n5269, ZN => n831);
   U5149 : OAI21_X2 port map( B1 => n12310, B2 => n28253, A => n12309, ZN => 
                           n13419);
   U5153 : NOR2_X1 port map( A1 => n12299, A2 => n12303, ZN => n28253);
   U5154 : NAND3_X1 port map( A1 => n26930, A2 => n26927, A3 => n26926, ZN => 
                           n1277);
   U5180 : NAND2_X1 port map( A1 => n1561, A2 => n18172, ZN => n28254);
   U5183 : NAND2_X1 port map( A1 => n24099, A2 => n53, ZN => n28255);
   U5195 : OAI21_X1 port map( B1 => n14976, B2 => n14974, A => n14973, ZN => 
                           n14975);
   U5196 : NAND2_X1 port map( A1 => n14971, A2 => n13789, ZN => n14974);
   U5244 : NAND2_X1 port map( A1 => n21440, A2 => n6275, ZN => n28258);
   U5246 : NAND2_X1 port map( A1 => n20244, A2 => n21661, ZN => n28259);
   U5254 : AOI21_X1 port map( B1 => n12333, B2 => n12332, A => n28260, ZN => 
                           n11748);
   U5299 : OAI21_X1 port map( B1 => n6097, B2 => n24493, A => n28261, ZN => 
                           n690);
   U5300 : NAND3_X1 port map( A1 => n24470, A2 => n23942, A3 => n29033, ZN => 
                           n28261);
   U5301 : NAND2_X1 port map( A1 => n26573, A2 => n29576, ZN => n28284);
   U5318 : NAND2_X1 port map( A1 => n28263, A2 => n28262, ZN => n24393);
   U5320 : NAND2_X1 port map( A1 => n24392, A2 => n29471, ZN => n28263);
   U5376 : NAND3_X2 port map( A1 => n11620, A2 => n28265, A3 => n28264, ZN => 
                           n13055);
   U5379 : NAND2_X1 port map( A1 => n11618, A2 => n5637, ZN => n28264);
   U5388 : INV_X1 port map( A => n11989, ZN => n28265);
   U5425 : NAND2_X1 port map( A1 => n28268, A2 => n28266, ZN => n8815);
   U5441 : NAND2_X1 port map( A1 => n8814, A2 => n28267, ZN => n28266);
   U5465 : INV_X1 port map( A => n8812, ZN => n28267);
   U5483 : NAND2_X1 port map( A1 => n8681, A2 => n8810, ZN => n8814);
   U5498 : NAND2_X1 port map( A1 => n8813, A2 => n8812, ZN => n28268);
   U5503 : AOI21_X1 port map( B1 => n10569, B2 => n4101, A => n28270, ZN => 
                           n28269);
   U5511 : INV_X1 port map( A => n10795, ZN => n28270);
   U5523 : NAND2_X1 port map( A1 => n17833, A2 => n17832, ZN => n17838);
   U5524 : XNOR2_X1 port map( A => n28271, B => n26214, ZN => Ciphertext(14));
   U5540 : NAND2_X1 port map( A1 => n4032, A2 => n4034, ZN => n28271);
   U5555 : NAND3_X1 port map( A1 => n27721, A2 => n27719, A3 => n27720, ZN => 
                           n27722);
   U5584 : OAI21_X2 port map( B1 => n11209, B2 => n10656, A => n10655, ZN => 
                           n375);
   U5597 : NAND2_X1 port map( A1 => n2196, A2 => n8359, ZN => n9948);
   U5598 : OAI21_X2 port map( B1 => n20116, B2 => n20117, A => n20115, ZN => 
                           n21424);
   U5626 : NAND2_X1 port map( A1 => n1422, A2 => n1426, ZN => n28274);
   U5632 : NAND2_X1 port map( A1 => n1420, A2 => n23946, ZN => n1425);
   U5677 : NAND2_X1 port map( A1 => n11220, A2 => n11223, ZN => n11106);
   U5681 : NAND2_X1 port map( A1 => n3237, A2 => n28275, ZN => n1267);
   U5711 : NAND3_X1 port map( A1 => n28276, A2 => n1606, A3 => n7354, ZN => 
                           n9139);
   U5740 : NAND2_X1 port map( A1 => n1608, A2 => n7353, ZN => n28276);
   U5743 : NAND2_X1 port map( A1 => n13829, A2 => n14360, ZN => n14075);
   U5764 : XNOR2_X1 port map( A => n28277, B => n27643, ZN => Ciphertext(98));
   U5797 : AOI22_X1 port map( A1 => n27642, A2 => n27641, B1 => n27647, B2 => 
                           n27640, ZN => n28277);
   U5810 : OAI21_X1 port map( B1 => n20078, B2 => n20079, A => n20077, ZN => 
                           n20086);
   U5828 : NOR2_X1 port map( A1 => n7454, A2 => n28278, ZN => n7461);
   U5831 : INV_X1 port map( A => n7984, ZN => n28278);
   U5839 : NAND2_X1 port map( A1 => n7643, A2 => n7456, ZN => n7984);
   U5867 : INV_X1 port map( A => n9575, ZN => n8715);
   U5939 : NAND2_X1 port map( A1 => n1251, A2 => n3121, ZN => n24154);
   U5942 : OR2_X1 port map( A1 => n7164, A2 => n7320, ZN => n3167);
   U5983 : NAND2_X1 port map( A1 => n3809, A2 => n3808, ZN => n19962);
   U5984 : NAND2_X1 port map( A1 => n28279, A2 => n28737, ZN => n23842);
   U5991 : NOR2_X1 port map( A1 => n23822, A2 => n23821, ZN => n28279);
   U5997 : OR2_X1 port map( A1 => n5918, A2 => n14039, ZN => n59);
   U6024 : NAND3_X1 port map( A1 => n16940, A2 => n211, A3 => n16939, ZN => n42
                           );
   U6037 : OAI22_X1 port map( A1 => n8268, A2 => n8267, B1 => n341, B2 => n8270
                           , ZN => n8272);
   U6180 : XNOR2_X1 port map( A => n28280, B => n26681, ZN => Ciphertext(129));
   U6192 : NAND3_X1 port map( A1 => n3561, A2 => n26678, A3 => n6902, ZN => 
                           n28280);
   U6230 : NAND2_X1 port map( A1 => n1355, A2 => n28281, ZN => n1884);
   U6271 : NAND3_X1 port map( A1 => n24422, A2 => n24421, A3 => n24517, ZN => 
                           n903);
   U6394 : NAND2_X1 port map( A1 => n11774, A2 => n10497, ZN => n28282);
   U6411 : INV_X1 port map( A => n10716, ZN => n28283);
   U6463 : NAND2_X1 port map( A1 => n26574, A2 => n28286, ZN => n28285);
   U6484 : INV_X1 port map( A => n26575, ZN => n28286);
   U6524 : NAND2_X1 port map( A1 => n3803, A2 => n3802, ZN => n3800);
   U6526 : NAND2_X1 port map( A1 => n8438, A2 => n224, ZN => n8441);
   U6536 : NAND2_X1 port map( A1 => n28184, A2 => n28287, ZN => n5477);
   U6559 : NAND2_X1 port map( A1 => n400, A2 => n27703, ZN => n28288);
   U6561 : NAND2_X1 port map( A1 => n27701, A2 => n27704, ZN => n28289);
   U6579 : NAND2_X1 port map( A1 => n5651, A2 => n5652, ZN => n5650);
   U6590 : NAND2_X1 port map( A1 => n7932, A2 => n7613, ZN => n8310);
   U6604 : NAND3_X1 port map( A1 => n28290, A2 => n20901, A3 => n5830, ZN => 
                           n5014);
   U6684 : NAND2_X1 port map( A1 => n20896, A2 => n21426, ZN => n28290);
   U6718 : NAND2_X1 port map( A1 => n28291, A2 => n15288, ZN => n1392);
   U6766 : NAND2_X1 port map( A1 => n1394, A2 => n756, ZN => n28291);
   U6795 : NAND2_X1 port map( A1 => n29023, A2 => n17592, ZN => n28292);
   U6830 : AOI22_X1 port map( A1 => n26981, A2 => n27636, B1 => n26982, B2 => 
                           n27638, ZN => n26983);
   U6852 : NAND2_X1 port map( A1 => n8271, A2 => n8270, ZN => n7210);
   U6855 : NAND2_X1 port map( A1 => n18490, A2 => n18488, ZN => n18291);
   U6872 : NAND2_X1 port map( A1 => n52, A2 => n54, ZN => n51);
   U7082 : XNOR2_X1 port map( A => n21817, B => n22882, ZN => n21979);
   U7162 : NAND2_X1 port map( A1 => n2250, A2 => n8784, ZN => n1566);
   U7243 : INV_X1 port map( A => n7775, ZN => n28692);
   U7251 : OAI22_X1 port map( A1 => n27418, A2 => n27429, B1 => n27428, B2 => 
                           n27427, ZN => n26669);
   U7254 : XNOR2_X1 port map( A => n13432, B => n12919, ZN => n12921);
   U7340 : OAI21_X2 port map( B1 => n11748, B2 => n6432, A => n3281, ZN => 
                           n13432);
   U7353 : NOR2_X1 port map( A1 => n20251, A2 => n20252, ZN => n28295);
   U7389 : INV_X1 port map( A => n11271, ZN => n652);
   U7400 : NAND2_X1 port map( A1 => n279, A2 => n11038, ZN => n11271);
   U7433 : OAI21_X1 port map( B1 => n8720, B2 => n8718, A => n28296, ZN => 
                           n8413);
   U7458 : NAND2_X1 port map( A1 => n8718, A2 => n8788, ZN => n28296);
   U7468 : OAI21_X1 port map( B1 => n28298, B2 => n28532, A => n28297, ZN => 
                           n25596);
   U7470 : NAND2_X1 port map( A1 => n25575, A2 => n28532, ZN => n28297);
   U7520 : INV_X1 port map( A => n26996, ZN => n28298);
   U7521 : NAND2_X1 port map( A1 => n11574, A2 => n12264, ZN => n5963);
   U7546 : AND3_X2 port map( A1 => n11041, A2 => n11040, A3 => n11042, ZN => 
                           n11574);
   U7579 : NAND3_X1 port map( A1 => n21069, A2 => n22403, A3 => n28299, ZN => 
                           n22830);
   U7605 : NAND2_X1 port map( A1 => n28301, A2 => n28300, ZN => n28299);
   U7635 : NOR2_X1 port map( A1 => n22402, A2 => n22404, ZN => n28300);
   U7637 : NAND2_X1 port map( A1 => n27715, A2 => n1826, ZN => n27684);
   U7645 : NAND4_X2 port map( A1 => n28302, A2 => n3512, A3 => n1522, A4 => 
                           n3514, ZN => n26011);
   U7678 : NAND2_X1 port map( A1 => n28419, A2 => n24368, ZN => n28302);
   U7684 : XNOR2_X1 port map( A => n2813, B => n28303, ZN => n26230);
   U7702 : INV_X1 port map( A => n2812, ZN => n28303);
   U7711 : NAND2_X1 port map( A1 => n27977, A2 => n28456, ZN => n28355);
   U7756 : NAND2_X1 port map( A1 => n18433, A2 => n18430, ZN => n17815);
   U7779 : OAI21_X2 port map( B1 => n17218, B2 => n17217, A => n17216, ZN => 
                           n18430);
   U7782 : NAND2_X1 port map( A1 => n2576, A2 => n6023, ZN => n14936);
   U7817 : BUF_X1 port map( A => n22991, Z => n23180);
   U7837 : NAND2_X1 port map( A1 => n15040, A2 => n14517, ZN => n28305);
   U7852 : NAND3_X1 port map( A1 => n5811, A2 => n14971, A3 => n14793, ZN => 
                           n5810);
   U7871 : NOR2_X2 port map( A1 => n28307, A2 => n5201, ZN => n18114);
   U7916 : OAI21_X1 port map( B1 => n1708, B2 => n5203, A => n853, ZN => n28307
                           );
   U7920 : NAND2_X1 port map( A1 => n4419, A2 => n4420, ZN => n28308);
   U7973 : OAI21_X1 port map( B1 => n27711, B2 => n27714, A => n26146, ZN => 
                           n26145);
   U8011 : NAND2_X1 port map( A1 => n27725, A2 => n27711, ZN => n26146);
   U8018 : AND2_X1 port map( A1 => n14400, A2 => n29628, ZN => n13962);
   U8019 : OAI21_X1 port map( B1 => n6128, B2 => n16790, A => n28309, ZN => 
                           n6126);
   U8027 : NAND3_X1 port map( A1 => n28768, A2 => n17421, A3 => n17012, ZN => 
                           n28309);
   U8052 : NOR2_X1 port map( A1 => n15222, A2 => n15223, ZN => n5238);
   U8060 : NAND2_X1 port map( A1 => n10940, A2 => n10942, ZN => n10702);
   U8073 : XNOR2_X1 port map( A => n13442, B => n13443, ZN => n28311);
   U8074 : NOR2_X1 port map( A1 => n21349, A2 => n28312, ZN => n21351);
   U8080 : NAND2_X1 port map( A1 => n21346, A2 => n21347, ZN => n28312);
   U8094 : NAND2_X1 port map( A1 => n6314, A2 => n21698, ZN => n21347);
   U8095 : NAND2_X1 port map( A1 => n14677, A2 => n3315, ZN => n6681);
   U8101 : NAND2_X1 port map( A1 => n14902, A2 => n15097, ZN => n14677);
   U8103 : NAND2_X1 port map( A1 => n28313, A2 => n18078, ZN => n18080);
   U8106 : OAI22_X1 port map( A1 => n18076, A2 => n18075, B1 => n18074, B2 => 
                           n5814, ZN => n28313);
   U8110 : NAND2_X1 port map( A1 => n24557, A2 => n24633, ZN => n24558);
   U8111 : NAND2_X1 port map( A1 => n24461, A2 => n28314, ZN => n24462);
   U8112 : AND2_X1 port map( A1 => n24812, A2 => n24809, ZN => n28314);
   U8123 : BUF_X2 port map( A => n21729, Z => n1930);
   U8143 : AND3_X2 port map( A1 => n6518, A2 => n6519, A3 => n11542, ZN => 
                           n13273);
   U8164 : NAND2_X1 port map( A1 => n28316, A2 => n28315, ZN => n23921);
   U8187 : NAND2_X1 port map( A1 => n6740, A2 => n24583, ZN => n28316);
   U8223 : NAND2_X1 port map( A1 => n24592, A2 => n831, ZN => n24142);
   U8282 : OAI21_X1 port map( B1 => n4370, B2 => n7977, A => n7976, ZN => n7978
                           );
   U8297 : NAND2_X1 port map( A1 => n28320, A2 => n28319, ZN => n26069);
   U8298 : NAND2_X1 port map( A1 => n401, A2 => n28229, ZN => n28319);
   U8326 : NAND2_X1 port map( A1 => n26052, A2 => n28180, ZN => n28320);
   U8349 : XNOR2_X1 port map( A => n28321, B => n22841, ZN => n23289);
   U8351 : XNOR2_X1 port map( A => n22839, B => n22838, ZN => n28321);
   U8376 : NAND2_X1 port map( A1 => n28322, A2 => n14294, ZN => n14296);
   U8403 : NAND3_X1 port map( A1 => n5198, A2 => n15154, A3 => n5199, ZN => 
                           n5197);
   U8427 : INV_X1 port map( A => n520, ZN => n5690);
   U8429 : NAND2_X1 port map( A1 => n28324, A2 => n2938, ZN => n2442);
   U8431 : NAND2_X1 port map( A1 => n2937, A2 => n23655, ZN => n28324);
   U8475 : NAND3_X1 port map( A1 => n772, A2 => n1458, A3 => n770, ZN => n25205
                           );
   U8481 : OR2_X1 port map( A1 => n2096, A2 => n20170, ZN => n4640);
   U8514 : NAND3_X1 port map( A1 => n27621, A2 => n27620, A3 => n1912, ZN => 
                           n1186);
   U8516 : NAND3_X1 port map( A1 => n29126, A2 => n23619, A3 => n23270, ZN => 
                           n23271);
   U8523 : NAND3_X1 port map( A1 => n7939, A2 => n7657, A3 => n8301, ZN => 
                           n7658);
   U8538 : NAND2_X1 port map( A1 => n24484, A2 => n24483, ZN => n967);
   U8598 : NAND2_X1 port map( A1 => n2283, A2 => n28329, ZN => n10270);
   U8604 : NAND2_X1 port map( A1 => n10872, A2 => n11219, ZN => n28329);
   U8608 : AOI21_X2 port map( B1 => n28331, B2 => n23591, A => n28330, ZN => 
                           n25785);
   U8609 : NAND2_X1 port map( A1 => n23575, A2 => n2079, ZN => n28331);
   U8610 : NAND3_X1 port map( A1 => n14379, A2 => n14005, A3 => n14007, ZN => 
                           n6106);
   U8616 : XNOR2_X2 port map( A => n12247, B => n12248, ZN => n14259);
   U8658 : NAND2_X1 port map( A1 => n28333, A2 => n11338, ZN => n28332);
   U8710 : NAND2_X1 port map( A1 => n11336, A2 => n11176, ZN => n28333);
   U8714 : NAND2_X1 port map( A1 => n11178, A2 => n10830, ZN => n28334);
   U8716 : NAND2_X1 port map( A1 => n14550, A2 => n14549, ZN => n15476);
   U8744 : AND2_X2 port map( A1 => n28335, A2 => n87, ZN => n9233);
   U8758 : NAND2_X1 port map( A1 => n6963, A2 => n6962, ZN => n28335);
   U8771 : NAND2_X1 port map( A1 => n471, A2 => n24972, ZN => n1251);
   U8775 : NAND2_X1 port map( A1 => n10694, A2 => n10985, ZN => n10695);
   U8821 : NAND2_X1 port map( A1 => n6704, A2 => n28336, ZN => n11599);
   U8822 : NAND2_X1 port map( A1 => n8064, A2 => n582, ZN => n6704);
   U8907 : NAND2_X1 port map( A1 => n17379, A2 => n17179, ZN => n17177);
   U8921 : NOR2_X1 port map( A1 => n26953, A2 => n26954, ZN => n28337);
   U8927 : OR2_X1 port map( A1 => n7145, A2 => n7146, ZN => n28674);
   U8941 : NAND2_X1 port map( A1 => n6284, A2 => n6285, ZN => n28339);
   U8959 : NOR2_X1 port map( A1 => n28094, A2 => n28340, ZN => n26764);
   U8972 : NAND2_X1 port map( A1 => n29056, A2 => n28111, ZN => n28340);
   U9030 : NAND2_X1 port map( A1 => n27219, A2 => n27572, ZN => n28341);
   U9065 : XNOR2_X2 port map( A => n12617, B => n12618, ZN => n14295);
   U9125 : NAND2_X1 port map( A1 => n5624, A2 => n28343, ZN => n26682);
   U9184 : AOI21_X1 port map( B1 => n26788, B2 => n1872, A => n28344, ZN => 
                           n28343);
   U9195 : AND2_X1 port map( A1 => n26912, A2 => n28423, ZN => n28344);
   U9225 : NAND2_X1 port map( A1 => n14487, A2 => n14481, ZN => n14169);
   U9237 : OAI211_X1 port map( C1 => n3976, C2 => n14761, A => n15055, B => 
                           n28345, ZN => n3979);
   U9246 : NAND2_X1 port map( A1 => n4162, A2 => n14761, ZN => n28345);
   U9309 : NAND2_X1 port map( A1 => n507, A2 => n20133, ZN => n19903);
   U9401 : NAND2_X1 port map( A1 => n85, A2 => n27672, ZN => n28347);
   U9405 : NAND2_X1 port map( A1 => n28348, A2 => n18658, ZN => n20966);
   U9435 : OAI21_X1 port map( B1 => n20559, B2 => n18650, A => n20563, ZN => 
                           n28348);
   U9453 : AND2_X1 port map( A1 => n9421, A2 => n8327, ZN => n1386);
   U9487 : NAND3_X1 port map( A1 => n24261, A2 => n24503, A3 => n24801, ZN => 
                           n24262);
   U9527 : AND2_X2 port map( A1 => n7259, A2 => n3683, ZN => n9562);
   U9597 : INV_X1 port map( A => n12512, ZN => n28349);
   U9609 : NOR2_X2 port map( A1 => n2655, A2 => n10102, ZN => n12512);
   U9686 : NAND2_X1 port map( A1 => n14299, A2 => n13816, ZN => n28351);
   U9740 : OR2_X1 port map( A1 => n430, A2 => n12991, ZN => n28677);
   U9743 : NAND2_X1 port map( A1 => n24814, A2 => n24812, ZN => n2246);
   U9784 : NAND3_X1 port map( A1 => n23332, A2 => n23768, A3 => n28354, ZN => 
                           n28353);
   U9799 : OAI21_X1 port map( B1 => n21012, B2 => n21443, A => n20833, ZN => 
                           n20836);
   U9815 : OAI21_X1 port map( B1 => n27977, B2 => n29021, A => n28355, ZN => 
                           n26637);
   U9829 : OR2_X2 port map( A1 => n6060, A2 => n28357, ZN => n9073);
   U9833 : AOI21_X1 port map( B1 => n7430, B2 => n7431, A => n8234, ZN => 
                           n28357);
   U9924 : XNOR2_X1 port map( A => n28359, B => n18579, ZN => n18834);
   U9971 : XNOR2_X1 port map( A => n18576, B => n19693, ZN => n28359);
   U9982 : OAI21_X1 port map( B1 => n4819, B2 => n26174, A => n28360, ZN => 
                           n4817);
   U10020 : NAND3_X1 port map( A1 => n26172, A2 => n26917, A3 => n26919, ZN => 
                           n28360);
   U10062 : NAND3_X1 port map( A1 => n24422, A2 => n24515, A3 => n24421, ZN => 
                           n28361);
   U10126 : NAND3_X1 port map( A1 => n23871, A2 => n23870, A3 => n24514, ZN => 
                           n28362);
   U10141 : MUX2_X1 port map( A => n12280, B => n11357, S => n12404, Z => 
                           n11358);
   U10147 : NAND2_X1 port map( A1 => n12281, A2 => n12407, ZN => n12404);
   U10193 : OR2_X1 port map( A1 => n10667, A2 => n11077, ZN => n28364);
   U10198 : NAND2_X1 port map( A1 => n28722, A2 => n14109, ZN => n14517);
   U10199 : NAND2_X1 port map( A1 => n28218, A2 => n439, ZN => n28365);
   U10235 : NAND4_X2 port map( A1 => n24319, A2 => n28369, A3 => n28368, A4 => 
                           n28367, ZN => n25780);
   U10255 : NAND2_X1 port map( A1 => n24317, A2 => n24316, ZN => n28367);
   U10259 : NAND2_X1 port map( A1 => n28227, A2 => n24072, ZN => n28368);
   U10296 : NAND2_X1 port map( A1 => n24315, A2 => n24669, ZN => n28369);
   U10299 : NAND2_X1 port map( A1 => n17771, A2 => n17772, ZN => n18019);
   U10300 : NAND2_X1 port map( A1 => n9124, A2 => n8899, ZN => n1651);
   U10311 : NAND3_X1 port map( A1 => n618, A2 => n7521, A3 => n8030, ZN => 
                           n8031);
   U10335 : NAND3_X1 port map( A1 => n149, A2 => n2940, A3 => n2939, ZN => n851
                           );
   U10347 : NAND2_X1 port map( A1 => n28371, A2 => n485, ZN => n1676);
   U10360 : OAI22_X1 port map( A1 => n28626, A2 => n23417, B1 => n480, B2 => 
                           n23416, ZN => n28371);
   U10424 : NAND2_X1 port map( A1 => n8008, A2 => n8504, ZN => n28372);
   U10504 : AND2_X1 port map( A1 => n19827, A2 => n20311, ZN => n5826);
   U10526 : NAND2_X1 port map( A1 => n6752, A2 => n21495, ZN => n21127);
   U10586 : NAND2_X1 port map( A1 => n28377, A2 => n28376, ZN => n27214);
   U10587 : NAND2_X1 port map( A1 => n27209, A2 => n27210, ZN => n28376);
   U10601 : NAND2_X1 port map( A1 => n27211, A2 => n27038, ZN => n28377);
   U10602 : INV_X1 port map( A => n27209, ZN => n28378);
   U10665 : NAND2_X1 port map( A1 => n28381, A2 => n28379, ZN => n10218);
   U10704 : INV_X1 port map( A => n28380, ZN => n28379);
   U10711 : OAI21_X1 port map( B1 => n9000, B2 => n329, A => n9001, ZN => 
                           n28380);
   U10728 : OAI211_X1 port map( C1 => n329, C2 => n9202, A => n8779, B => 
                           n28862, ZN => n28381);
   U10812 : NAND2_X1 port map( A1 => n25470, A2 => n25471, ZN => n28670);
   U10852 : NAND2_X1 port map( A1 => n18835, A2 => n29582, ZN => n28383);
   U10859 : NAND2_X1 port map( A1 => n18836, A2 => n29315, ZN => n28384);
   U10862 : NAND2_X1 port map( A1 => n4672, A2 => n23835, ZN => n6557);
   U10889 : INV_X1 port map( A => n10844, ZN => n1812);
   U10895 : NAND2_X1 port map( A1 => n11272, A2 => n11269, ZN => n10844);
   U10911 : XNOR2_X1 port map( A => n24402, B => n24401, ZN => n28385);
   U10968 : NAND3_X1 port map( A1 => n3390, A2 => n6634, A3 => n6633, ZN => 
                           n28386);
   U10969 : NAND2_X1 port map( A1 => n21262, A2 => n3318, ZN => n28387);
   U10970 : XNOR2_X1 port map( A => n28388, B => n22562, ZN => n22564);
   U10981 : XOR2_X1 port map( A => n22561, B => n22690, Z => n28388);
   U10991 : NAND2_X1 port map( A1 => n21262, A2 => n3318, ZN => n22561);
   U11015 : XOR2_X1 port map( A => n10306, B => n8477, Z => n8479);
   U11031 : NAND2_X1 port map( A1 => n23972, A2 => n24209, ZN => n4754);
   U11051 : XNOR2_X1 port map( A => n22231, B => n22230, ZN => n28390);
   U11088 : INV_X1 port map( A => n23193, ZN => n28391);
   U11105 : XNOR2_X1 port map( A => n24868, B => n24869, ZN => n28392);
   U11127 : AND2_X1 port map( A1 => n6125, A2 => n6124, ZN => n28393);
   U11191 : AND2_X1 port map( A1 => n6125, A2 => n6124, ZN => n28394);
   U11229 : AND2_X1 port map( A1 => n6125, A2 => n6124, ZN => n27208);
   U11267 : OAI21_X1 port map( B1 => n14888, B2 => n14889, A => n14887, ZN => 
                           n28395);
   U11276 : XOR2_X1 port map( A => n16555, B => n16026, Z => n16030);
   U11295 : OAI21_X1 port map( B1 => n14888, B2 => n14889, A => n14887, ZN => 
                           n3792);
   U11307 : AOI21_X1 port map( B1 => n18346, B2 => n514, A => n18344, ZN => 
                           n17950);
   U11343 : NOR2_X1 port map( A1 => n27695, A2 => n27694, ZN => n28396);
   U11363 : XOR2_X1 port map( A => n28397, B => n3321, Z => Ciphertext(136));
   U11377 : NAND3_X1 port map( A1 => n2765, A2 => n2764, A3 => n2763, ZN => 
                           n28397);
   U11388 : MUX2_X1 port map( A => n28399, B => n28400, S => n27701, Z => 
                           n28398);
   U11434 : OR2_X1 port map( A1 => n27702, A2 => n27700, ZN => n28399);
   U11441 : OR2_X1 port map( A1 => n27703, A2 => n27161, ZN => n28400);
   U11459 : NOR2_X1 port map( A1 => n6277, A2 => n6278, ZN => n28401);
   U11478 : NOR2_X1 port map( A1 => n24116, A2 => n24115, ZN => n28402);
   U11498 : NOR2_X1 port map( A1 => n1008, A2 => n26324, ZN => n28403);
   U11499 : NOR2_X1 port map( A1 => n24116, A2 => n24115, ZN => n25463);
   U11509 : OR2_X1 port map( A1 => n3283, A2 => n18376, ZN => n28404);
   U11510 : XOR2_X1 port map( A => n13420, B => n13067, Z => n12943);
   U11532 : XNOR2_X1 port map( A => n9394, B => n9395, ZN => n11004);
   U11593 : XNOR2_X1 port map( A => n9408, B => n9407, ZN => n1308);
   U11628 : XNOR2_X1 port map( A => n19282, B => n19281, ZN => n28408);
   U11658 : NAND2_X1 port map( A1 => n3758, A2 => n1050, ZN => n28409);
   U11699 : NAND2_X1 port map( A1 => n3758, A2 => n1050, ZN => n22887);
   U11716 : NAND3_X1 port map( A1 => n664, A2 => n25971, A3 => n663, ZN => 
                           n28411);
   U11724 : NAND3_X1 port map( A1 => n664, A2 => n25971, A3 => n663, ZN => 
                           n28016);
   U11729 : CLKBUF_X1 port map( A => Key(44), Z => n27894);
   U11761 : NAND2_X1 port map( A1 => n28412, A2 => n28413, ZN => n994);
   U11837 : OR2_X1 port map( A1 => n17659, A2 => n18467, ZN => n28412);
   U11874 : OR2_X1 port map( A1 => n18464, A2 => n1383, ZN => n28413);
   U11875 : BUF_X1 port map( A => n11739, Z => n11742);
   U11902 : AND2_X1 port map( A1 => n6025, A2 => n6024, ZN => n28414);
   U11908 : XOR2_X1 port map( A => n19269, B => n18858, Z => n18861);
   U11971 : AOI22_X1 port map( A1 => n456, A2 => n26436, B1 => n26937, B2 => 
                           n26936, ZN => n5546);
   U12005 : OAI21_X1 port map( B1 => n6091, B2 => n23419, A => n23063, ZN => 
                           n24717);
   U12012 : XNOR2_X1 port map( A => n19545, B => n19544, ZN => n28417);
   U12023 : XNOR2_X1 port map( A => n6846, B => n6847, ZN => n23280);
   U12025 : NOR2_X1 port map( A1 => n24369, A2 => n23897, ZN => n28419);
   U12026 : NAND2_X1 port map( A1 => n20605, A2 => n20606, ZN => n21599);
   U12029 : XNOR2_X1 port map( A => n25862, B => n25861, ZN => n28631);
   U12038 : AND2_X1 port map( A1 => n28420, A2 => n23211, ZN => n21978);
   U12041 : OR2_X1 port map( A1 => n23577, A2 => n23603, ZN => n28420);
   U12046 : INV_X1 port map( A => n26937, ZN => n28421);
   U12076 : AND2_X1 port map( A1 => n25159, A2 => n25158, ZN => n28422);
   U12101 : XOR2_X1 port map( A => n25383, B => n25384, Z => n28423);
   U12105 : MUX2_X1 port map( A => n26805, B => n26806, S => n2438, Z => n26807
                           );
   U12134 : OAI21_X1 port map( B1 => n480, B2 => n22808, A => n22807, ZN => 
                           n24556);
   U12149 : INV_X1 port map( A => n24382, ZN => n28424);
   U12150 : XNOR2_X1 port map( A => n28425, B => n28426, ZN => n5306);
   U12169 : XNOR2_X1 port map( A => n25743, B => n25744, ZN => n28425);
   U12192 : XOR2_X1 port map( A => n25747, B => n25746, Z => n28426);
   U12222 : OAI21_X1 port map( B1 => n23350, B2 => n4429, A => n23349, ZN => 
                           n24665);
   U12318 : XNOR2_X1 port map( A => n22070, B => n22071, ZN => n23700);
   U12397 : BUF_X1 port map( A => n27590, Z => n28429);
   U12418 : INV_X1 port map( A => n27732, ZN => n28430);
   U12444 : XOR2_X1 port map( A => n9648, B => n9899, Z => n10156);
   U12477 : XOR2_X1 port map( A => n13565, B => n12834, Z => n12381);
   U12482 : XOR2_X1 port map( A => n22070, B => n22071, Z => n28431);
   U12483 : OR2_X1 port map( A1 => n24560, A2 => n23990, ZN => n28687);
   U12515 : XOR2_X1 port map( A => n22093, B => n28387, Z => n28432);
   U12518 : AOI21_X1 port map( B1 => n219, B2 => n28679, A => n28678, ZN => 
                           n28433);
   U12519 : AOI21_X1 port map( B1 => n219, B2 => n28679, A => n28678, ZN => 
                           n4263);
   U12520 : XOR2_X1 port map( A => n24446, B => n24445, Z => n28434);
   U12525 : BUF_X1 port map( A => n27460, Z => n28435);
   U12527 : OAI21_X1 port map( B1 => n26159, B2 => n26562, A => n26158, ZN => 
                           n27460);
   U12548 : BUF_X1 port map( A => n11787, Z => n28436);
   U12551 : XOR2_X1 port map( A => n25854, B => n25853, Z => n28437);
   U12558 : OAI21_X1 port map( B1 => n10729, B2 => n10730, A => n10728, ZN => 
                           n11787);
   U12574 : MUX2_X2 port map( A => n26783, B => n26784, S => n454, Z => n27282)
                           ;
   U12604 : AND3_X1 port map( A1 => n27009, A2 => n27008, A3 => n27007, ZN => 
                           n28438);
   U12605 : AND3_X1 port map( A1 => n27009, A2 => n27008, A3 => n27007, ZN => 
                           n28439);
   U12620 : AOI22_X1 port map( A1 => n18546, A2 => n19967, B1 => n18547, B2 => 
                           n20123, ZN => n21343);
   U12634 : AND3_X1 port map( A1 => n6755, A2 => n5391, A3 => n5390, ZN => 
                           n28441);
   U12641 : NAND2_X1 port map( A1 => n5779, A2 => n5780, ZN => n28442);
   U12708 : XOR2_X1 port map( A => n12383, B => n12087, Z => n12119);
   U12714 : XNOR2_X1 port map( A => n21882, B => n21883, ZN => n28444);
   U12740 : AND4_X1 port map( A1 => n27135, A2 => n27134, A3 => n27133, A4 => 
                           n27132, ZN => n28445);
   U12759 : XNOR2_X1 port map( A => n21882, B => n21883, ZN => n23687);
   U12786 : XNOR2_X1 port map( A => n25502, B => n25501, ZN => n27052);
   U12804 : CLKBUF_X1 port map( A => n22205, Z => n28514);
   U12832 : NOR2_X1 port map( A1 => n17817, A2 => n17816, ZN => n28447);
   U12847 : INV_X1 port map( A => n20049, ZN => n28448);
   U12848 : XNOR2_X1 port map( A => n22053, B => n22052, ZN => n22600);
   U12858 : XNOR2_X1 port map( A => n25823, B => n25824, ZN => n26840);
   U12864 : NAND3_X1 port map( A1 => n2299, A2 => n19803, A3 => n4225, ZN => 
                           n28449);
   U12952 : BUF_X1 port map( A => n1534, Z => n28451);
   U12959 : NAND2_X1 port map( A1 => n25001, A2 => n25003, ZN => n894);
   U12997 : XNOR2_X1 port map( A => n25719, B => n25718, ZN => n28452);
   U12999 : OAI211_X1 port map( C1 => n27073, C2 => n27072, A => n3786, B => 
                           n3785, ZN => n28453);
   U13018 : INV_X1 port map( A => n16693, ZN => n18343);
   U13067 : XNOR2_X1 port map( A => n15786, B => n15785, ZN => n17541);
   U13070 : OAI211_X1 port map( C1 => n29126, C2 => n23626, A => n5554, B => 
                           n5556, ZN => n28455);
   U13110 : OAI211_X1 port map( C1 => n29126, C2 => n23626, A => n5554, B => 
                           n5556, ZN => n23655);
   U13133 : XNOR2_X1 port map( A => n20872, B => n20873, ZN => n28457);
   U13142 : XOR2_X1 port map( A => n25823, B => n25824, Z => n28458);
   U13143 : XNOR2_X1 port map( A => n20872, B => n20873, ZN => n23686);
   U13148 : XNOR2_X1 port map( A => n25308, B => n25307, ZN => n28459);
   U13187 : XNOR2_X1 port map( A => n25308, B => n25307, ZN => n26715);
   U13188 : INV_X1 port map( A => n7298, ZN => n8162);
   U13189 : AOI22_X1 port map( A1 => n25632, A2 => n26723, B1 => n26717, B2 => 
                           n25631, ZN => n27408);
   U13202 : BUF_X1 port map( A => n22232, Z => n28461);
   U13234 : OAI22_X1 port map( A1 => n20719, A2 => n28602, B1 => n5622, B2 => 
                           n20899, ZN => n22232);
   U13262 : AOI21_X1 port map( B1 => n3950, B2 => n14345, A => n3947, ZN => 
                           n28462);
   U13289 : AOI21_X1 port map( B1 => n3950, B2 => n14345, A => n3947, ZN => 
                           n15175);
   U13290 : OR2_X1 port map( A1 => n10828, A2 => n11337, ZN => n1190);
   U13345 : OR2_X1 port map( A1 => n24056, A2 => n5507, ZN => n24916);
   U13376 : NAND2_X1 port map( A1 => n23915, A2 => n985, ZN => n28465);
   U13385 : NAND2_X1 port map( A1 => n985, A2 => n23915, ZN => n26060);
   U13398 : OAI21_X1 port map( B1 => n24857, B2 => n4679, A => n24856, ZN => 
                           n27646);
   U13400 : XOR2_X1 port map( A => n25697, B => n26059, Z => n25458);
   U13417 : XOR2_X1 port map( A => n22218, B => n22219, Z => n22712);
   U13418 : XNOR2_X1 port map( A => n1502, B => n1055, ZN => n23370);
   U13442 : XOR2_X1 port map( A => n25033, B => n25032, Z => n28467);
   U13466 : INV_X1 port map( A => n27203, ZN => n28468);
   U13547 : XOR2_X1 port map( A => n25098, B => n25097, Z => n28470);
   U13548 : XNOR2_X1 port map( A => n25376, B => n25377, ZN => n28471);
   U13567 : OAI211_X1 port map( C1 => n21011, C2 => n21010, A => n21009, B => 
                           n2343, ZN => n28472);
   U13598 : OAI211_X1 port map( C1 => n21011, C2 => n21010, A => n21009, B => 
                           n2343, ZN => n22910);
   U13647 : XNOR2_X1 port map( A => n2813, B => n2812, ZN => n28473);
   U13676 : OR2_X1 port map( A1 => n11322, A2 => n29316, ZN => n22);
   U13682 : INV_X1 port map( A => n29157, ZN => n28474);
   U13696 : NOR2_X1 port map( A1 => n22178, A2 => n22179, ZN => n28475);
   U13704 : NOR2_X1 port map( A1 => n22178, A2 => n22179, ZN => n26044);
   U13710 : XNOR2_X1 port map( A => n3596, B => n25258, ZN => n26447);
   U13718 : XNOR2_X1 port map( A => n13276, B => n13275, ZN => n28478);
   U13719 : XNOR2_X1 port map( A => n18926, B => n18925, ZN => n21095);
   U13729 : XOR2_X1 port map( A => n24879, B => n24878, Z => n28480);
   U13874 : OAI21_X1 port map( B1 => n23232, B2 => n1862, A => n23231, ZN => 
                           n28481);
   U13875 : XOR2_X1 port map( A => n24574, B => n24573, Z => n28482);
   U13879 : AND2_X1 port map( A1 => n9207, A2 => n41, ZN => n9437);
   U13898 : NAND4_X1 port map( A1 => n6425, A2 => n6427, A3 => n6426, A4 => 
                           n20216, ZN => n28483);
   U13917 : NAND4_X1 port map( A1 => n6425, A2 => n6427, A3 => n6426, A4 => 
                           n20216, ZN => n22568);
   U13925 : NOR2_X1 port map( A1 => n23967, A2 => n23966, ZN => n28485);
   U13935 : XNOR2_X1 port map( A => n22121, B => n22120, ZN => n23725);
   U13936 : NOR2_X1 port map( A1 => n23967, A2 => n23966, ZN => n26094);
   U13969 : NOR2_X1 port map( A1 => n21112, A2 => n4755, ZN => n28486);
   U13970 : XOR2_X1 port map( A => n22159, B => n21836, Z => n21840);
   U13973 : NOR2_X1 port map( A1 => n21112, A2 => n4755, ZN => n22756);
   U13977 : XNOR2_X1 port map( A => n26087, B => n26088, ZN => n28487);
   U13980 : XNOR2_X1 port map( A => n26087, B => n26088, ZN => n27141);
   U13982 : XNOR2_X1 port map( A => n25561, B => n25560, ZN => n26632);
   U14077 : BUF_X1 port map( A => n27972, Z => n27970);
   U14098 : INV_X1 port map( A => n4950, ZN => n28738);
   U14099 : OR2_X1 port map( A1 => n15787, A2 => n17542, ZN => n16940);
   U14107 : OAI211_X1 port map( C1 => n9167, C2 => n9163, A => n8317, B => 
                           n8316, ZN => n9921);
   U14130 : NAND2_X1 port map( A1 => n1810, A2 => n20276, ZN => n28492);
   U14274 : OR2_X1 port map( A1 => n17415, A2 => n17413, ZN => n17301);
   U14306 : AND2_X1 port map( A1 => n25359, A2 => n25357, ZN => n28494);
   U14316 : XNOR2_X1 port map( A => n9270, B => n9269, ZN => n28495);
   U14322 : CLKBUF_X1 port map( A => n25187, Z => n28496);
   U14340 : XNOR2_X1 port map( A => n9270, B => n9269, ZN => n10941);
   U14423 : NOR2_X1 port map( A1 => n4466, A2 => n4465, ZN => n28499);
   U14510 : NAND2_X1 port map( A1 => n7482, A2 => n7483, ZN => n9080);
   U14511 : XNOR2_X1 port map( A => n16871, B => n16870, ZN => n28501);
   U14537 : XNOR2_X1 port map( A => n24088, B => n24089, ZN => n28503);
   U14625 : NAND2_X1 port map( A1 => n23293, A2 => n4175, ZN => n3797);
   U14633 : NAND3_X1 port map( A1 => n5427, A2 => n24030, A3 => n24031, ZN => 
                           n25703);
   U14666 : XOR2_X1 port map( A => n24931, B => n24930, Z => n28504);
   U14747 : OR2_X1 port map( A1 => n1912, A2 => n27630, ZN => n28505);
   U14786 : MUX2_X2 port map( A => n26360, B => n26359, S => n26358, Z => 
                           n27630);
   U14843 : XOR2_X1 port map( A => n5702, B => n5703, Z => n28506);
   U14848 : INV_X1 port map( A => n14358, ZN => n28507);
   U14907 : OR2_X1 port map( A1 => n29037, A2 => n13672, ZN => n2965);
   U15011 : XNOR2_X1 port map( A => n5703, B => n5702, ZN => n23801);
   U15032 : CLKBUF_X1 port map( A => n20573, Z => n28508);
   U15033 : XNOR2_X1 port map( A => n18609, B => n19683, ZN => n20573);
   U15037 : AND2_X1 port map( A1 => n27302, A2 => n27303, ZN => n28510);
   U15073 : MUX2_X2 port map( A => n25316, B => n25315, S => n29560, Z => 
                           n27364);
   U15128 : XNOR2_X1 port map( A => n24918, B => n24919, ZN => n28513);
   U15131 : AOI22_X1 port map( A1 => n23608, A2 => n23607, B1 => n23605, B2 => 
                           n23606, ZN => n24790);
   U15132 : CLKBUF_X1 port map( A => n20333, Z => n28515);
   U15138 : XNOR2_X1 port map( A => n19288, B => n19287, ZN => n20333);
   U15238 : OAI22_X1 port map( A1 => n23108, A2 => n23107, B1 => n23106, B2 => 
                           n486, ZN => n24211);
   U15286 : OAI21_X1 port map( B1 => n14004, B2 => n13575, A => n13574, ZN => 
                           n28518);
   U15305 : OAI21_X1 port map( B1 => n14004, B2 => n13575, A => n13574, ZN => 
                           n14942);
   U15309 : AOI21_X1 port map( B1 => n24177, B2 => n24178, A => n24176, ZN => 
                           n28520);
   U15315 : XNOR2_X1 port map( A => n25766, B => n25765, ZN => n28521);
   U15373 : AOI21_X1 port map( B1 => n24177, B2 => n24178, A => n24176, ZN => 
                           n25445);
   U15492 : XNOR2_X2 port map( A => n24841, B => n24840, ZN => n26426);
   U15493 : NOR2_X1 port map( A1 => n6599, A2 => n23797, ZN => n28522);
   U15508 : NOR2_X1 port map( A1 => n6599, A2 => n23797, ZN => n28523);
   U15511 : NOR2_X1 port map( A1 => n6599, A2 => n23797, ZN => n24803);
   U15516 : OAI211_X1 port map( C1 => n23694, C2 => n23135, A => n6442, B => 
                           n6441, ZN => n24409);
   U15528 : XNOR2_X1 port map( A => n24198, B => n24199, ZN => n28525);
   U15535 : XNOR2_X1 port map( A => n24198, B => n24199, ZN => n26185);
   U15572 : XNOR2_X1 port map( A => n22022, B => n22021, ZN => n28527);
   U15617 : OR2_X1 port map( A1 => n5320, A2 => n23255, ZN => n28528);
   U15620 : XNOR2_X1 port map( A => n22022, B => n22021, ZN => n23406);
   U15625 : XNOR2_X2 port map( A => n24625, B => n24624, ZN => n26457);
   U15640 : NOR2_X1 port map( A1 => n4803, A2 => n174, ZN => n28530);
   U15722 : NOR2_X1 port map( A1 => n4803, A2 => n174, ZN => n19636);
   U15759 : INV_X1 port map( A => n24697, ZN => n28531);
   U15779 : XNOR2_X1 port map( A => n25574, B => n25573, ZN => n28532);
   U15804 : XNOR2_X1 port map( A => n25574, B => n25573, ZN => n26997);
   U15828 : XNOR2_X1 port map( A => n24882, B => n24881, ZN => n28536);
   U15995 : XNOR2_X1 port map( A => n19416, B => n19415, ZN => n28538);
   U15996 : XNOR2_X1 port map( A => n19416, B => n19415, ZN => n20634);
   U16017 : XNOR2_X1 port map( A => n22210, B => n22209, ZN => n23562);
   U16066 : OAI211_X1 port map( C1 => n17897, C2 => n18268, A => n1718, B => 
                           n1716, ZN => n18928);
   U16088 : OAI22_X1 port map( A1 => n23889, A2 => n23888, B1 => n23887, B2 => 
                           n24434, ZN => n28540);
   U16159 : OAI22_X1 port map( A1 => n23889, A2 => n23888, B1 => n23887, B2 => 
                           n24434, ZN => n25583);
   U16245 : XNOR2_X1 port map( A => n25129, B => n25130, ZN => n26941);
   U16380 : XNOR2_X1 port map( A => n25189, B => n6789, ZN => n28542);
   U16535 : XNOR2_X1 port map( A => n25189, B => n6789, ZN => n26266);
   U16536 : XOR2_X1 port map( A => n16566, B => n15256, Z => n15257);
   U16829 : NAND2_X1 port map( A1 => n26243, A2 => n26244, ZN => n28064);
   U16831 : INV_X1 port map( A => n4599, ZN => n28544);
   U16952 : XNOR2_X1 port map( A => n25693, B => n25692, ZN => n27067);
   U16961 : XNOR2_X1 port map( A => n24170, B => n24169, ZN => n28547);
   U16965 : XNOR2_X1 port map( A => n24170, B => n24169, ZN => n26182);
   U17022 : XNOR2_X1 port map( A => n25296, B => n25297, ZN => n28548);
   U17039 : NAND3_X1 port map( A1 => n25664, A2 => n6288, A3 => n25663, ZN => 
                           n28549);
   U17040 : NAND3_X1 port map( A1 => n25664, A2 => n6288, A3 => n25663, ZN => 
                           n27355);
   U17051 : XOR2_X1 port map( A => n25901, B => n26038, Z => n24885);
   U17098 : CLKBUF_X3 port map( A => n26537, Z => n27875);
   U17103 : XNOR2_X1 port map( A => n25171, B => n25170, ZN => n26949);
   U17208 : XOR2_X1 port map( A => n22466, B => n22465, Z => n28551);
   U17328 : XNOR2_X1 port map( A => n19524, B => n19523, ZN => n28552);
   U17523 : XOR2_X1 port map( A => n19713, B => n19712, Z => n28555);
   U17611 : OAI211_X1 port map( C1 => n24743, C2 => n24744, A => n24742, B => 
                           n24741, ZN => n25825);
   U17664 : AOI22_X1 port map( A1 => n14114, A2 => n15116, B1 => n13668, B2 => 
                           n1001, ZN => n28557);
   U17689 : AOI22_X1 port map( A1 => n14114, A2 => n15116, B1 => n13668, B2 => 
                           n1001, ZN => n16039);
   U17776 : AOI22_X1 port map( A1 => n17380, A2 => n4295, B1 => n17378, B2 => 
                           n17379, ZN => n18708);
   U17840 : CLKBUF_X1 port map( A => n10556, Z => n28559);
   U17841 : BUF_X1 port map( A => n26481, Z => n28560);
   U17844 : XNOR2_X1 port map( A => n25217, B => n25218, ZN => n26481);
   U17856 : OR2_X1 port map( A1 => n7164, A2 => n7770, ZN => n7323);
   U17893 : XNOR2_X1 port map( A => n24063, B => n24062, ZN => n28561);
   U17939 : BUF_X1 port map( A => n26808, Z => n28562);
   U17944 : XNOR2_X1 port map( A => n24063, B => n24062, ZN => n26476);
   U17980 : OAI21_X1 port map( B1 => n25321, B2 => n28525, A => n25320, ZN => 
                           n26808);
   U17981 : OR3_X1 port map( A1 => n17259, A2 => n17260, A3 => n17262, ZN => 
                           n3587);
   U18075 : XNOR2_X1 port map( A => n15564, B => n6929, ZN => n28564);
   U18110 : OR2_X1 port map( A1 => n24512, A2 => n24511, ZN => n28565);
   U18211 : XOR2_X1 port map( A => n6212, B => n21728, Z => n28566);
   U18328 : OR2_X1 port map( A1 => n22948, A2 => n22947, ZN => n28567);
   U18329 : NOR2_X2 port map( A1 => n24648, A2 => n24647, ZN => n25542);
   U18438 : XNOR2_X1 port map( A => n9714, B => n6916, ZN => n28568);
   U18458 : XNOR2_X1 port map( A => n19282, B => n19281, ZN => n20598);
   U18477 : OR2_X1 port map( A1 => n23683, A2 => n23686, ZN => n3434);
   U18854 : XNOR2_X1 port map( A => n13483, B => n6651, ZN => n28569);
   U18911 : XNOR2_X1 port map( A => n21419, B => n21418, ZN => n28570);
   U18915 : XNOR2_X1 port map( A => n13483, B => n6651, ZN => n14039);
   U18959 : XNOR2_X1 port map( A => n21419, B => n21418, ZN => n23343);
   U18983 : INV_X1 port map( A => n17012, ZN => n16968);
   U18984 : NAND2_X1 port map( A1 => n5228, A2 => n17863, ZN => n28571);
   U19007 : NAND2_X1 port map( A1 => n5228, A2 => n17863, ZN => n19725);
   U19010 : XNOR2_X1 port map( A => n24962, B => n24961, ZN => n28572);
   U19044 : XNOR2_X1 port map( A => n24962, B => n24961, ZN => n28573);
   U19059 : NOR2_X1 port map( A1 => n28226, A2 => n27165, ZN => n27171);
   U19065 : XOR2_X1 port map( A => n6870, B => n6869, Z => n28574);
   U19131 : XNOR2_X1 port map( A => n25830, B => n25248, ZN => n28575);
   U19284 : OR2_X1 port map( A1 => n20494, A2 => n20493, ZN => n19867);
   U19386 : XOR2_X1 port map( A => n21689, B => n21688, Z => n28577);
   U19419 : NAND2_X1 port map( A1 => n3344, A2 => n13988, ZN => n28579);
   U19477 : NAND2_X1 port map( A1 => n3967, A2 => n19798, ZN => n28580);
   U19672 : XNOR2_X1 port map( A => n22191, B => n22190, ZN => n28581);
   U19699 : XNOR2_X1 port map( A => n22191, B => n22190, ZN => n28582);
   U19726 : XOR2_X1 port map( A => n25448, B => n25447, Z => n28583);
   U19728 : XOR2_X1 port map( A => n22698, B => n22699, Z => n22701);
   U19805 : BUF_X1 port map( A => n13566, Z => n28587);
   U19826 : XOR2_X1 port map( A => n11866, B => n11865, Z => n28588);
   U19866 : OAI21_X1 port map( B1 => n11863, B2 => n11862, A => n1526, ZN => 
                           n13566);
   U19871 : NAND2_X1 port map( A1 => n3531, A2 => n3530, ZN => n28589);
   U19942 : NAND2_X1 port map( A1 => n3531, A2 => n3530, ZN => n22762);
   U20053 : NOR2_X1 port map( A1 => n26725, A2 => n26724, ZN => n28591);
   U20146 : OAI21_X1 port map( B1 => n24038, B2 => n24039, A => n24037, ZN => 
                           n27029);
   U20172 : XNOR2_X1 port map( A => n19379, B => n19378, ZN => n19641);
   U20226 : NAND2_X1 port map( A1 => n6513, A2 => n1223, ZN => n28593);
   U20358 : XOR2_X1 port map( A => n22598, B => n22597, Z => n28594);
   U20400 : XOR2_X1 port map( A => n24905, B => n24904, Z => n28595);
   U20423 : NOR2_X1 port map( A1 => n23083, A2 => n23082, ZN => n28596);
   U20425 : OAI21_X1 port map( B1 => n14669, B2 => n15304, A => n14668, ZN => 
                           n28597);
   U20426 : INV_X1 port map( A => n24426, ZN => n28598);
   U20645 : OAI21_X1 port map( B1 => n14669, B2 => n15304, A => n14668, ZN => 
                           n16470);
   U20745 : OAI21_X1 port map( B1 => n23535, B2 => n23534, A => n6942, ZN => 
                           n24767);
   U20809 : NAND2_X1 port map( A1 => n6513, A2 => n1223, ZN => n26020);
   U20853 : XOR2_X1 port map( A => n25937, B => n25936, Z => n28600);
   U20908 : XOR2_X1 port map( A => n12773, B => n12772, Z => n28601);
   U20940 : BUF_X1 port map( A => n1925, Z => n28602);
   U20944 : NOR2_X1 port map( A1 => n12185, A2 => n12184, ZN => n28603);
   U21033 : XNOR2_X1 port map( A => n21300, B => n21299, ZN => n28604);
   U21048 : XNOR2_X1 port map( A => n21300, B => n21299, ZN => n23676);
   U21119 : OR2_X1 port map( A1 => n29629, A2 => n7257, ZN => n7512);
   U21125 : XNOR2_X1 port map( A => n6977, B => Key(101), ZN => n28605);
   U21158 : OR2_X1 port map( A1 => n20480, A2 => n19995, ZN => n20230);
   U21159 : NOR2_X1 port map( A1 => n20357, A2 => n20356, ZN => n20782);
   U21237 : INV_X1 port map( A => n27242, ZN => n28607);
   U21290 : NOR2_X1 port map( A1 => n3445, A2 => n155, ZN => n9081);
   U21318 : XNOR2_X1 port map( A => n6891, B => n9309, ZN => n10948);
   U21330 : XOR2_X1 port map( A => n19444, B => n19443, Z => n28610);
   U21334 : INV_X1 port map( A => n20393, ZN => n28611);
   U21376 : XOR2_X1 port map( A => n9527, B => n9526, Z => n28612);
   U21395 : XOR2_X1 port map( A => n22326, B => n22414, Z => n28613);
   U21419 : MUX2_X1 port map( A => n7616, B => n7615, S => n29135, Z => n7617);
   U21424 : XNOR2_X1 port map( A => n7219, B => Key(128), ZN => n28614);
   U21440 : XNOR2_X1 port map( A => n7219, B => Key(128), ZN => n28615);
   U21463 : XNOR2_X1 port map( A => n7219, B => Key(128), ZN => n8256);
   U21495 : AND2_X1 port map( A1 => n20573, A2 => n19838, ZN => n19833);
   U21498 : OR2_X1 port map( A1 => n12057, A2 => n12320, ZN => n28747);
   U21514 : XNOR2_X1 port map( A => n7220, B => Key(129), ZN => n28617);
   U21549 : XNOR2_X1 port map( A => n7220, B => Key(129), ZN => n28618);
   U21550 : AOI22_X1 port map( A1 => n20387, A2 => n20386, B1 => n20385, B2 => 
                           n20384, ZN => n28619);
   U21554 : XNOR2_X1 port map( A => n7220, B => Key(129), ZN => n8263);
   U21784 : AOI22_X1 port map( A1 => n20387, A2 => n20386, B1 => n20385, B2 => 
                           n20384, ZN => n21501);
   U21803 : XNOR2_X1 port map( A => n19080, B => n19081, ZN => n28620);
   U21817 : XNOR2_X1 port map( A => n19081, B => n19080, ZN => n20485);
   U21819 : XOR2_X1 port map( A => n19121, B => n19120, Z => n28621);
   U21900 : NOR2_X1 port map( A1 => n2205, A2 => n24559, ZN => n24561);
   U21910 : NOR2_X1 port map( A1 => n19656, A2 => n19659, ZN => n28623);
   U22058 : XNOR2_X1 port map( A => n10125, B => n10124, ZN => n28624);
   U22085 : XNOR2_X1 port map( A => n10124, B => n10125, ZN => n11210);
   U22105 : XOR2_X1 port map( A => n12897, B => n12898, Z => n28625);
   U22116 : XNOR2_X1 port map( A => n22775, B => n22774, ZN => n28626);
   U22120 : XNOR2_X1 port map( A => n22775, B => n22774, ZN => n2452);
   U22305 : XNOR2_X1 port map( A => n7811, B => n7812, ZN => n28627);
   U22412 : XNOR2_X1 port map( A => n7811, B => n7812, ZN => n11145);
   U22413 : OAI21_X1 port map( B1 => n1777, B2 => n1828, A => n23094, ZN => 
                           n25190);
   U22509 : OAI211_X1 port map( C1 => n23857, C2 => n23856, A => n841, B => 
                           n840, ZN => n28630);
   U22513 : OAI211_X1 port map( C1 => n23857, C2 => n23856, A => n841, B => 
                           n840, ZN => n25858);
   U22671 : XNOR2_X1 port map( A => n25862, B => n25861, ZN => n27118);
   U22715 : BUF_X1 port map( A => n18492, Z => n28633);
   U22737 : AOI22_X1 port map( A1 => n16878, A2 => n15616, B1 => n15615, B2 => 
                           n424, ZN => n18492);
   U22764 : OAI211_X1 port map( C1 => n9106, C2 => n8512, A => n9105, B => 
                           n8072, ZN => n28634);
   U22883 : OAI211_X1 port map( C1 => n9106, C2 => n8512, A => n9105, B => 
                           n8072, ZN => n10145);
   U23009 : AOI21_X1 port map( B1 => n26632, B2 => n26631, A => n26630, ZN => 
                           n27997);
   U23010 : XNOR2_X1 port map( A => n18586, B => n18585, ZN => n28637);
   U23015 : XNOR2_X1 port map( A => n18586, B => n18585, ZN => n19836);
   U23016 : XNOR2_X1 port map( A => n8520, B => n8519, ZN => n28638);
   U23067 : XOR2_X1 port map( A => n25496, B => n25497, Z => n28639);
   U23076 : XNOR2_X1 port map( A => n8520, B => n8519, ZN => n10814);
   U23077 : XOR2_X1 port map( A => n25789, B => n25788, Z => n28640);
   U23081 : INV_X1 port map( A => n26546, ZN => n28641);
   U23091 : NOR2_X1 port map( A1 => n27865, A2 => n27872, ZN => n27327);
   U23105 : XNOR2_X1 port map( A => n24982, B => n24983, ZN => n28642);
   U23106 : OAI21_X1 port map( B1 => n7161, B2 => n7160, A => n7159, ZN => 
                           n28643);
   U23122 : CLKBUF_X1 port map( A => n23631, Z => n28644);
   U23158 : OAI21_X1 port map( B1 => n22970, B2 => n22969, A => n22968, ZN => 
                           n28645);
   U23159 : BUF_X1 port map( A => n26951, Z => n28646);
   U23175 : XNOR2_X1 port map( A => n12480, B => n12479, ZN => n28647);
   U23205 : XNOR2_X1 port map( A => n12480, B => n12479, ZN => n28648);
   U23259 : INV_X1 port map( A => n4044, ZN => n28649);
   U23318 : XNOR2_X1 port map( A => n12480, B => n12479, ZN => n14444);
   U23368 : NOR2_X1 port map( A1 => n17781, A2 => n17782, ZN => n18174);
   U23377 : OR2_X1 port map( A1 => n14845, A2 => n15284, ZN => n14849);
   U23418 : XNOR2_X1 port map( A => n25014, B => n25013, ZN => n28650);
   U23428 : XNOR2_X1 port map( A => n25014, B => n25013, ZN => n28651);
   U23433 : NOR2_X1 port map( A1 => n26356, A2 => n28650, ZN => n28652);
   U23552 : XNOR2_X1 port map( A => n22604, B => n22603, ZN => n28653);
   U23614 : AOI21_X1 port map( B1 => n24376, B2 => n23999, A => n23998, ZN => 
                           n28654);
   U23625 : XNOR2_X1 port map( A => n22604, B => n22603, ZN => n23809);
   U23634 : AOI21_X1 port map( B1 => n24376, B2 => n23999, A => n23998, ZN => 
                           n25465);
   U23651 : OAI211_X1 port map( C1 => n27192, C2 => n27193, A => n4108, B => 
                           n4110, ZN => n28655);
   U23669 : OAI211_X1 port map( C1 => n27192, C2 => n27193, A => n4108, B => 
                           n4110, ZN => n27662);
   U23671 : BUF_X1 port map( A => n17872, Z => n28656);
   U23703 : BUF_X1 port map( A => n20282, Z => n28657);
   U23736 : XOR2_X1 port map( A => n18568, B => n18567, Z => n28658);
   U23838 : XNOR2_X1 port map( A => n21492, B => n21491, ZN => n28659);
   U23857 : XNOR2_X1 port map( A => n25699, B => n25700, ZN => n28660);
   U23922 : XNOR2_X1 port map( A => n19128, B => n19127, ZN => n20225);
   U23977 : NOR2_X1 port map( A1 => n20583, A2 => n20582, ZN => n28661);
   U24006 : NAND2_X1 port map( A1 => n2372, A2 => n2371, ZN => n28662);
   U24054 : AOI21_X1 port map( B1 => n28663, B2 => n3771, A => n5263, ZN => 
                           n1008);
   U24064 : NAND2_X1 port map( A1 => n26320, A2 => n26992, ZN => n28663);
   U24097 : OAI21_X2 port map( B1 => n8122, B2 => n8351, A => n8121, ZN => 
                           n10088);
   U24133 : OR2_X1 port map( A1 => n20248, A2 => n20033, ZN => n20641);
   U24179 : OAI21_X1 port map( B1 => n15689, B2 => n28666, A => n28665, ZN => 
                           n15693);
   U24213 : NAND2_X1 port map( A1 => n15689, A2 => n15690, ZN => n28665);
   U24219 : NOR2_X1 port map( A1 => n20044, A2 => n20158, ZN => n19982);
   U24220 : NAND2_X1 port map( A1 => n17762, A2 => n17942, ZN => n17761);
   U24408 : NAND2_X1 port map( A1 => n15388, A2 => n15144, ZN => n15390);
   U24475 : NAND2_X1 port map( A1 => n27107, A2 => n28667, ZN => n27755);
   U24547 : NAND2_X1 port map( A1 => n4794, A2 => n23370, ZN => n2119);
   U24549 : XNOR2_X1 port map( A => n28668, B => n3083, ZN => Ciphertext(118));
   U24573 : OAI21_X1 port map( B1 => n27752, B2 => n27751, A => n27750, ZN => 
                           n28668);
   U24698 : OAI21_X1 port map( B1 => n20362, B2 => n21520, A => n21180, ZN => 
                           n20363);
   U24748 : NOR2_X1 port map( A1 => n8509, A2 => n8510, ZN => n9431);
   U24752 : NAND2_X1 port map( A1 => n28671, A2 => n17849, ZN => n6444);
   U24779 : NAND2_X1 port map( A1 => n2719, A2 => n17845, ZN => n28671);
   U24923 : NAND3_X1 port map( A1 => n11661, A2 => n2142, A3 => n12163, ZN => 
                           n12104);
   U24993 : NAND2_X1 port map( A1 => n12167, A2 => n11376, ZN => n11381);
   U24995 : NAND2_X1 port map( A1 => n5234, A2 => n18388, ZN => n28672);
   U24998 : AND4_X2 port map( A1 => n1556, A2 => n1555, A3 => n4994, A4 => 
                           n1558, ZN => n24633);
   U25074 : NAND2_X1 port map( A1 => n24460, A2 => n24808, ZN => n24816);
   U25166 : INV_X1 port map( A => n5759, ZN => n5245);
   U25171 : NAND2_X1 port map( A1 => n5758, A2 => n5756, ZN => n5759);
   U25174 : INV_X1 port map( A => n21634, ZN => n21635);
   U25283 : NAND2_X1 port map( A1 => n12149, A2 => n12991, ZN => n28676);
   U25328 : NAND2_X1 port map( A1 => n24811, A2 => n24810, ZN => n28679);
   U25348 : NAND2_X1 port map( A1 => n21013, A2 => n2639, ZN => n22053);
   U25376 : NAND2_X1 port map( A1 => n25966, A2 => n25965, ZN => n28680);
   U25377 : NAND3_X1 port map( A1 => n8630, A2 => n8627, A3 => n8664, ZN => 
                           n8629);
   U25397 : NAND3_X1 port map( A1 => n24372, A2 => n23994, A3 => n23995, ZN => 
                           n28717);
   U25423 : NAND2_X1 port map( A1 => n7968, A2 => n1938, ZN => n7970);
   U25432 : NAND2_X1 port map( A1 => n20948, A2 => n21499, ZN => n20949);
   U25434 : OAI21_X1 port map( B1 => n24073, B2 => n23372, A => n28681, ZN => 
                           n23374);
   U25505 : NAND2_X1 port map( A1 => n3989, A2 => n11548, ZN => n28682);
   U25517 : OAI211_X2 port map( C1 => n14511, C2 => n14512, A => n14509, B => 
                           n28683, ZN => n16023);
   U25527 : NAND2_X1 port map( A1 => n14512, A2 => n15251, ZN => n28683);
   U25592 : NAND3_X1 port map( A1 => n12278, A2 => n11801, A3 => n12280, ZN => 
                           n2288);
   U25595 : AOI21_X2 port map( B1 => n8118, B2 => n8653, A => n5819, ZN => 
                           n10087);
   U25615 : NAND2_X1 port map( A1 => n981, A2 => n28685, ZN => n28684);
   U25616 : NOR2_X1 port map( A1 => n14204, A2 => n28220, ZN => n28685);
   U25643 : NAND3_X2 port map( A1 => n28687, A2 => n23201, A3 => n28686, ZN => 
                           n25775);
   U25650 : INV_X1 port map( A => n24561, ZN => n28686);
   U25674 : NAND2_X1 port map( A1 => n6046, A2 => n3881, ZN => n6044);
   U25682 : OAI21_X1 port map( B1 => n29547, B2 => n18410, A => n28688, ZN => 
                           n17820);
   U25709 : NAND2_X1 port map( A1 => n18028, A2 => n18410, ZN => n28688);
   U25735 : NAND2_X1 port map( A1 => n7755, A2 => n887, ZN => n28689);
   U25781 : NAND2_X1 port map( A1 => n28690, A2 => n23751, ZN => n2818);
   U25851 : NAND2_X1 port map( A1 => n23747, A2 => n409, ZN => n28690);
   U25940 : OAI21_X1 port map( B1 => n28692, B2 => n7890, A => n28691, ZN => 
                           n7090);
   U25952 : NAND2_X1 port map( A1 => n7315, A2 => n7890, ZN => n28691);
   U26013 : NAND2_X1 port map( A1 => n11114, A2 => n10490, ZN => n10547);
   U26023 : NAND2_X1 port map( A1 => n22971, A2 => n6728, ZN => n4233);
   U26029 : NAND2_X1 port map( A1 => n24712, A2 => n28524, ZN => n24410);
   U26054 : NAND2_X1 port map( A1 => n15362, A2 => n15363, ZN => n15364);
   U26139 : NAND2_X1 port map( A1 => n28694, A2 => n27417, ZN => n27421);
   U26304 : NAND2_X1 port map( A1 => n29529, A2 => n29542, ZN => n28694);
   U26371 : NAND3_X1 port map( A1 => n7293, A2 => n8156, A3 => n7781, ZN => 
                           n28696);
   U26424 : INV_X1 port map( A => n19881, ZN => n20604);
   U26425 : NAND2_X1 port map( A1 => n20598, A2 => n4569, ZN => n19881);
   U26426 : NAND2_X1 port map( A1 => n14885, A2 => n14972, ZN => n14582);
   U26444 : NAND2_X1 port map( A1 => n14971, A2 => n14969, ZN => n14885);
   U26501 : NAND2_X1 port map( A1 => n390, A2 => n11751, ZN => n28698);
   U26502 : NAND2_X1 port map( A1 => n12219, A2 => n12218, ZN => n12222);
   U26630 : OAI21_X1 port map( B1 => n8718, B2 => n8717, A => n28699, ZN => 
                           n8442);
   U26646 : NAND2_X1 port map( A1 => n8718, A2 => n8719, ZN => n28699);
   U26789 : NAND2_X1 port map( A1 => n28702, A2 => n10717, ZN => n28701);
   U26793 : INV_X1 port map( A => n11793, ZN => n28702);
   U26837 : NAND2_X1 port map( A1 => n21698, A2 => n21696, ZN => n21695);
   U26844 : NAND3_X1 port map( A1 => n3016, A2 => n2019, A3 => n17754, ZN => 
                           n21698);
   U26851 : NAND3_X2 port map( A1 => n5543, A2 => n28704, A3 => n28703, ZN => 
                           n13447);
   U26895 : NAND2_X1 port map( A1 => n12083, A2 => n12289, ZN => n28704);
   U26898 : NAND2_X1 port map( A1 => n7591, A2 => n441, ZN => n5483);
   U26915 : AND2_X1 port map( A1 => n21503, A2 => n21539, ZN => n20947);
   U26952 : NAND3_X1 port map( A1 => n28706, A2 => n29552, A3 => n26151, ZN => 
                           n26153);
   U26954 : NAND2_X1 port map( A1 => n28710, A2 => n26789, ZN => n28706);
   U26984 : NAND2_X1 port map( A1 => n3459, A2 => n23779, ZN => n28707);
   U26993 : OAI21_X1 port map( B1 => n26792, B2 => n28709, A => n28708, ZN => 
                           n26795);
   U27010 : NAND2_X1 port map( A1 => n26792, A2 => n26793, ZN => n28708);
   U27039 : INV_X1 port map( A => n26791, ZN => n28711);
   U27045 : NAND2_X1 port map( A1 => n1764, A2 => n1763, ZN => n28712);
   U27065 : NAND2_X1 port map( A1 => n28714, A2 => n28713, ZN => n26796);
   U27131 : NAND2_X1 port map( A1 => n26790, A2 => n26791, ZN => n28713);
   U27170 : NAND2_X1 port map( A1 => n26924, A2 => n28711, ZN => n28714);
   U27191 : NAND2_X1 port map( A1 => n28715, A2 => n8176, ZN => n2659);
   U27201 : NAND2_X1 port map( A1 => n7763, A2 => n7347, ZN => n28715);
   U27226 : AOI21_X1 port map( B1 => n28716, B2 => n7313, A => n7176, ZN => 
                           n7112);
   U27267 : NAND2_X1 port map( A1 => n7896, A2 => n7895, ZN => n28716);
   U27341 : OAI21_X1 port map( B1 => n1828, B2 => n23997, A => n28717, ZN => 
                           n23998);
   U27346 : NAND2_X1 port map( A1 => n23819, A2 => n23820, ZN => n23090);
   U27376 : NAND2_X1 port map( A1 => n17316, A2 => n4220, ZN => n16836);
   U27377 : AOI22_X1 port map( A1 => n28718, A2 => n27382, B1 => n27037, B2 => 
                           n28378, ZN => n27039);
   U27382 : NAND2_X1 port map( A1 => n27212, A2 => n5312, ZN => n28718);
   U27477 : XNOR2_X1 port map( A => n12861, B => n3871, ZN => n253);
   U27480 : NAND2_X1 port map( A1 => n11569, A2 => n11568, ZN => n28719);
   U27511 : NAND2_X1 port map( A1 => n11570, A2 => n4341, ZN => n28720);
   U27528 : NAND2_X1 port map( A1 => n28721, A2 => n7822, ZN => n7823);
   U27562 : NAND3_X1 port map( A1 => n16804, A2 => n16802, A3 => n16801, ZN => 
                           n17780);
   U27576 : NAND3_X1 port map( A1 => n26, A2 => n11469, A3 => n11468, ZN => n25
                           );
   U27616 : NAND2_X1 port map( A1 => n14104, A2 => n14103, ZN => n28722);
   U27620 : NOR2_X1 port map( A1 => n21484, A2 => n28723, ZN => n19859);
   U27625 : NAND2_X1 port map( A1 => n1528, A2 => n1529, ZN => n1527);
   U27628 : NAND2_X1 port map( A1 => n18111, A2 => n17902, ZN => n17905);
   U27654 : NAND2_X1 port map( A1 => n11965, A2 => n28726, ZN => n28725);
   U27698 : NAND2_X1 port map( A1 => n17487, A2 => n17076, ZN => n17486);
   U27724 : OR2_X1 port map( A1 => n14947, A2 => n6855, ZN => n28727);
   U27766 : OR2_X1 port map( A1 => n20577, A2 => n20580, ZN => n5545);
   U27851 : NAND3_X1 port map( A1 => n28730, A2 => n9244, A3 => n9410, ZN => 
                           n9251);
   U27861 : NAND2_X1 port map( A1 => n28211, A2 => n9243, ZN => n28730);
   U27862 : NAND2_X1 port map( A1 => n17804, A2 => n16898, ZN => n28);
   U27876 : OR2_X1 port map( A1 => n7266, A2 => n7265, ZN => n8029);
   U27881 : NAND2_X1 port map( A1 => n2170, A2 => n4129, ZN => n7259);
   U27903 : NAND2_X1 port map( A1 => n342, A2 => n26960, ZN => n27390);
   U27929 : NAND2_X1 port map( A1 => n28732, A2 => n2954, ZN => n11058);
   U27930 : OAI21_X1 port map( B1 => n11030, B2 => n11031, A => n11283, ZN => 
                           n28732);
   U28002 : NAND3_X1 port map( A1 => n28404, A2 => n18349, A3 => n17646, ZN => 
                           n28733);
   U28003 : INV_X1 port map( A => n13857, ZN => n13856);
   U28017 : NAND2_X1 port map( A1 => n13673, A2 => n13855, ZN => n13857);
   U28037 : NAND2_X1 port map( A1 => n28734, A2 => n6465, ZN => n16667);
   U28039 : OAI21_X1 port map( B1 => n17277, B2 => n17278, A => n16844, ZN => 
                           n28734);
   U28121 : NAND3_X2 port map( A1 => n2645, A2 => n14700, A3 => n2642, ZN => 
                           n16216);
   U28126 : NAND2_X1 port map( A1 => n6097, A2 => n6098, ZN => n23878);
   U28127 : OAI21_X1 port map( B1 => n7964, B2 => n7963, A => n28736, ZN => 
                           n7578);
   U28128 : NAND2_X1 port map( A1 => n7964, A2 => n7965, ZN => n28736);
   U28129 : XNOR2_X1 port map( A => n22681, B => n22903, ZN => n22495);
   U28130 : OAI21_X1 port map( B1 => n23817, B2 => n23818, A => n28738, ZN => 
                           n28737);
   U28131 : INV_X1 port map( A => n15617, ZN => n15106);
   U28133 : NOR2_X1 port map( A1 => n16965, A2 => n28739, ZN => n16966);
   U28135 : AOI22_X2 port map( A1 => n5407, A2 => n14780, B1 => n14683, B2 => 
                           n14684, ZN => n15909);
   U28138 : NAND2_X1 port map( A1 => n28741, A2 => n26946, ZN => n27525);
   U28139 : AOI22_X1 port map( A1 => n6948, A2 => n26944, B1 => n26942, B2 => 
                           n26943, ZN => n28741);
   U28140 : NAND2_X1 port map( A1 => n28744, A2 => n28742, ZN => n9916);
   U28141 : NAND2_X1 port map( A1 => n8442, A2 => n28743, ZN => n28742);
   U28142 : NAND2_X1 port map( A1 => n8441, A2 => n8440, ZN => n28744);
   U28143 : INV_X1 port map( A => n18292, ZN => n28745);
   U28144 : NOR2_X1 port map( A1 => n1630, A2 => n567, ZN => n2542);
   U28145 : OAI211_X2 port map( C1 => n13781, C2 => n14254, A => n13779, B => 
                           n28746, ZN => n15208);
   U28146 : NAND3_X1 port map( A1 => n14253, A2 => n14254, A3 => n29312, ZN => 
                           n28746);
   U28147 : NAND2_X1 port map( A1 => n307, A2 => n27029, ZN => n26819);
   U28148 : NAND3_X2 port map( A1 => n14726, A2 => n3605, A3 => n14727, ZN => 
                           n16280);
   U28149 : NAND3_X1 port map( A1 => n6678, A2 => n6680, A3 => n28747, ZN => 
                           n12589);
   U28150 : NAND2_X1 port map( A1 => n28748, A2 => n5889, ZN => n3781);
   U28151 : NAND2_X1 port map( A1 => n9025, A2 => n9024, ZN => n28748);
   U28152 : NAND2_X1 port map( A1 => n697, A2 => n18322, ZN => n17714);
   U28155 : NAND2_X1 port map( A1 => n20535, A2 => n20934, ZN => n28749);
   U28156 : NAND2_X1 port map( A1 => n20534, A2 => n21078, ZN => n28750);
   U28157 : NAND2_X1 port map( A1 => n2697, A2 => n405, ZN => n4686);
   U28158 : INV_X1 port map( A => n28752, ZN => n28751);
   U28159 : OAI21_X1 port map( B1 => n7423, B2 => n370, A => n7422, ZN => 
                           n28752);
   U28162 : NAND2_X1 port map( A1 => n28121, A2 => n58, ZN => n28753);
   U28163 : OR2_X1 port map( A1 => n13898, A2 => n58, ZN => n28754);
   U28165 : NAND3_X2 port map( A1 => n1463, A2 => n1468, A3 => n17448, ZN => 
                           n18942);
   U28167 : OAI211_X1 port map( C1 => n28015, C2 => n28411, A => n26984, B => 
                           n28018, ZN => n25990);
   U28168 : NAND3_X1 port map( A1 => n1802, A2 => n1800, A3 => n1801, ZN => 
                           n1798);
   U28170 : NAND3_X1 port map( A1 => n17803, A2 => n3994, A3 => n18277, ZN => 
                           n27);
   U28171 : NAND2_X1 port map( A1 => n416, A2 => n19946, ZN => n3809);
   U28172 : NAND2_X1 port map( A1 => n17106, A2 => n17470, ZN => n17515);
   U28174 : XNOR2_X2 port map( A => n12086, B => n12085, ZN => n14484);
   U28175 : NAND2_X1 port map( A1 => n26315, A2 => n28214, ZN => n26316);
   U28178 : NAND3_X1 port map( A1 => n7464, A2 => n7618, A3 => n7463, ZN => 
                           n7469);
   U28179 : NAND2_X1 port map( A1 => n8246, A2 => n7690, ZN => n3510);
   U28181 : NAND2_X1 port map( A1 => n3658, A2 => n698, ZN => n22835);
   U28182 : NAND2_X1 port map( A1 => n4048, A2 => n4050, ZN => n15047);
   U28183 : NAND2_X1 port map( A1 => n693, A2 => n695, ZN => n15341);
   U28184 : NAND2_X1 port map( A1 => n18500, A2 => n520, ZN => n4707);
   U28185 : NAND2_X1 port map( A1 => n12079, A2 => n12058, ZN => n5543);
   U28186 : OAI22_X1 port map( A1 => n12291, A2 => n12080, B1 => n29324, B2 => 
                           n11795, ZN => n12079);
   U28188 : NAND3_X1 port map( A1 => n15205, A2 => n15203, A3 => n15204, ZN => 
                           n28756);
   U28191 : NAND3_X1 port map( A1 => n28757, A2 => n217, A3 => n15509, ZN => 
                           n4708);
   U28192 : NAND2_X1 port map( A1 => n2347, A2 => n15515, ZN => n28757);
   U28194 : NAND3_X1 port map( A1 => n18509, A2 => n510, A3 => n18510, ZN => 
                           n6255);
   U28195 : NAND3_X1 port map( A1 => n28759, A2 => n3690, A3 => n2463, ZN => 
                           n1688);
   U28196 : OAI21_X1 port map( B1 => n1691, B2 => n1690, A => n28107, ZN => 
                           n28759);
   U28198 : OR3_X1 port map( A1 => n16992, A2 => n29299, A3 => n17263, ZN => 
                           n16771);
   U28200 : NAND2_X1 port map( A1 => n4892, A2 => n4872, ZN => n4871);
   U28201 : OAI22_X1 port map( A1 => n27113, A2 => n401, B1 => n26865, B2 => 
                           n27112, ZN => n27114);
   U28202 : OAI211_X2 port map( C1 => n8738, C2 => n8739, A => n8737, B => 
                           n8736, ZN => n9931);
   U28203 : AND2_X1 port map( A1 => n1876, A2 => n14432, ZN => n28761);
   U28204 : AND2_X1 port map( A1 => n15374, A2 => n14863, ZN => n28762);
   U28206 : NAND2_X1 port map( A1 => n18506, A2 => n18213, ZN => n28763);
   U28207 : CLKBUF_X1 port map( A => n20425, Z => n22012);
   U28208 : OAI211_X2 port map( C1 => n5826, C2 => n6914, A => n19828, B => 
                           n1972, ZN => n21496);
   U28209 : OR2_X1 port map( A1 => n23194, A2 => n23647, ZN => n28764);
   U28210 : NAND2_X2 port map( A1 => n5309, A2 => n1162, ZN => n6348);
   U28212 : OR2_X1 port map( A1 => n23183, A2 => n23641, ZN => n28765);
   U28215 : OR2_X2 port map( A1 => n26190, A2 => n26189, ZN => n27038);
   U1524 : OR2_X2 port map( A1 => n28308, A2 => n17893, ZN => n18691);
   U627 : XNOR2_X2 port map( A => n22917, B => n22916, ZN => n23460);
   U2310 : XNOR2_X2 port map( A => n10155, B => n10154, ZN => n11086);
   U932 : MUX2_X2 port map( A => n8660, B => n8659, S => n8658, Z => n9915);
   U1752 : AND2_X2 port map( A1 => n669, A2 => n670, ZN => n19331);
   U1204 : AND2_X2 port map( A1 => n5791, A2 => n5792, ZN => n18471);
   U12394 : OAI21_X2 port map( B1 => n22939, B2 => n23449, A => n22938, ZN => 
                           n24591);
   U4286 : AND2_X2 port map( A1 => n1189, A2 => n1188, ZN => n21657);
   U5085 : OAI21_X2 port map( B1 => n23111, B2 => n29295, A => n1498, ZN => 
                           n24479);
   U9238 : NAND2_X2 port map( A1 => n3850, A2 => n14208, ZN => n15334);
   U18658 : XNOR2_X2 port map( A => n13188, B => n13187, ZN => n14031);
   U11500 : OR2_X2 port map( A1 => n17817, A2 => n17816, ZN => n19500);
   U1453 : AND2_X2 port map( A1 => n9865, A2 => n12194, ZN => n2483);
   U2217 : NAND2_X2 port map( A1 => n11693, A2 => n11694, ZN => n12219);
   U1269 : MUX2_X2 port map( A => n8435, B => n8434, S => n9034, Z => n10295);
   U2252 : AND3_X2 port map( A1 => n6373, A2 => n10112, A3 => n10111, ZN => 
                           n10863);
   U19384 : BUF_X1 port map( A => n25293, Z => n28576);
   U3435 : XNOR2_X2 port map( A => n7140, B => Key(49), ZN => n7743);
   U907 : BUF_X2 port map( A => n12166, Z => n1931);
   U8002 : AND2_X2 port map( A1 => n20095, A2 => n20094, ZN => n21078);
   U2344 : BUF_X1 port map( A => n23599, Z => n24973);
   U930 : MUX2_X2 port map( A => n8070, B => n8069, S => n8501, Z => n10219);
   U9983 : OR2_X2 port map( A1 => n6516, A2 => n6514, ZN => n12233);
   U231 : NAND2_X2 port map( A1 => n3574, A2 => n3577, ZN => n16416);
   U22399 : XNOR2_X2 port map( A => n19266, B => n19265, ZN => n19271);
   U292 : AND2_X2 port map( A1 => n6103, A2 => n6101, ZN => n19584);
   U10925 : OR2_X2 port map( A1 => n8728, A2 => n8727, ZN => n10264);
   U3427 : BUF_X1 port map( A => n7377, Z => n7818);
   U17446 : OAI211_X2 port map( C1 => n12334, C2 => n12327, A => n11452, B => 
                           n11451, ZN => n13278);
   U1237 : OR2_X1 port map( A1 => n6034, A2 => n23167, ZN => n23681);
   U754 : BUF_X1 port map( A => n19556, Z => n28143);
   U1199 : BUF_X1 port map( A => n27718, Z => n324);
   U685 : OR2_X2 port map( A1 => n21437, A2 => n5274, ZN => n20833);
   U3463 : INV_X2 port map( A => n18469, ZN => n6079);
   U60 : MUX2_X2 port map( A => n16228, B => n16227, S => n17138, Z => n18469);
   U4047 : NAND3_X2 port map( A1 => n4127, A2 => n1525, A3 => n4128, ZN => 
                           n11867);
   U3087 : OAI211_X2 port map( C1 => n11883, C2 => n11882, A => n2349, B => 
                           n2348, ZN => n13478);
   U15571 : OAI211_X2 port map( C1 => n22404, C2 => n21018, A => n1720, B => 
                           n21017, ZN => n22735);
   U5769 : NAND4_X2 port map( A1 => n7683, A2 => n7682, A3 => n7680, A4 => 
                           n7681, ZN => n10322);
   U1110 : AND3_X2 port map( A1 => n20884, A2 => n20883, A3 => n20882, ZN => 
                           n21994);
   U1933 : MUX2_X2 port map( A => n16493, B => n16492, S => n18464, Z => n18912
                           );
   U9665 : MUX2_X2 port map( A => n9091, B => n9090, S => n2320, Z => n10344);
   U1894 : OAI211_X2 port map( C1 => n15288, C2 => n14849, A => n14848, B => 
                           n14847, ZN => n16017);
   U3359 : OAI21_X2 port map( B1 => n7677, B2 => n7678, A => n6540, ZN => n9434
                           );
   U12642 : OAI211_X2 port map( C1 => n21138, C2 => n21605, A => n21604, B => 
                           n5719, ZN => n22500);
   U13340 : AOI22_X1 port map( A1 => n24580, A2 => n24581, B1 => n6056, B2 => 
                           n24467, ZN => n6055);
   U12485 : XNOR2_X1 port map( A => n23125, B => n23124, ZN => n26789);
   U5199 : OAI21_X1 port map( B1 => n1596, B2 => n16951, A => n16950, ZN => 
                           n18538);
   U5477 : AOI22_X1 port map( A1 => n20271, A2 => n20270, B1 => n20269, B2 => 
                           n21665, ZN => n1810);
   U2671 : MUX2_X2 port map( A => n17821, B => n17820, S => n18418, Z => n19706
                           );
   U1294 : OAI21_X1 port map( B1 => n24297, B2 => n24894, A => n24296, ZN => 
                           n24298);
   U6738 : MUX2_X2 port map( A => n3863, B => n10463, S => n11137, Z => n10766)
                           ;
   U4670 : AOI22_X1 port map( A1 => n21021, A2 => n22023, B1 => n21053, B2 => 
                           n22026, ZN => n21917);
   U23577 : AND3_X2 port map( A1 => n21176, A2 => n21175, A3 => n21174, ZN => 
                           n22678);
   U8743 : XNOR2_X1 port map( A => n9276, B => n9275, ZN => n10703);
   U1214 : MUX2_X2 port map( A => n12046, B => n12045, S => n12219, Z => n13525
                           );
   U4815 : AND2_X2 port map( A1 => n4153, A2 => n1282, ZN => n25322);
   U3948 : BUF_X1 port map( A => n26125, Z => n27147);
   U2559 : NAND4_X2 port map( A1 => n20030, A2 => n20029, A3 => n4933, A4 => 
                           n4567, ZN => n21392);
   U2918 : AND4_X2 port map( A1 => n2068, A2 => n5848, A3 => n5886, A4 => n5845
                           , ZN => n14810);
   U22015 : OAI21_X1 port map( B1 => n21220, B2 => n21215, A => n18786, ZN => 
                           n18787);
   U232 : NAND2_X1 port map( A1 => n3030, A2 => n7247, ZN => n8941);
   U5741 : XNOR2_X1 port map( A => n22213, B => n21905, ZN => n23790);
   U20810 : XNOR2_X1 port map( A => n4453, B => n4452, ZN => n17271);
   U164 : MUX2_X2 port map( A => n21944, B => n21943, S => n24729, Z => n26038)
                           ;
   U1957 : XNOR2_X1 port map( A => n3938, B => n3937, ZN => n16879);
   U563 : OAI21_X2 port map( B1 => n23207, B2 => n24550, A => n23206, ZN => 
                           n25565);
   U1635 : BUF_X1 port map( A => n27718, Z => n325);
   U2842 : XNOR2_X2 port map( A => n16466, B => n16465, ZN => n17506);
   U23512 : INV_X1 port map( A => n23686, ZN => n23516);
   U2668 : NAND2_X2 port map( A1 => n18112, A2 => n3074, ZN => n19700);
   U279 : MUX2_X1 port map( A => n19926, B => n19925, S => n5935, Z => n21748);
   U2125 : CLKBUF_X1 port map( A => Key(150), Z => n3673);
   U1597 : CLKBUF_X1 port map( A => Key(112), Z => n2916);
   U1589 : CLKBUF_X1 port map( A => Key(4), Z => n3598);
   U1817 : CLKBUF_X1 port map( A => Key(105), Z => n3081);
   U2127 : CLKBUF_X1 port map( A => Key(29), Z => n3483);
   U76 : CLKBUF_X1 port map( A => Key(116), Z => n3654);
   U1826 : CLKBUF_X1 port map( A => Key(47), Z => n3695);
   U14714 : XNOR2_X1 port map( A => n7139, B => Key(52), ZN => n7533);
   U6646 : BUF_X1 port map( A => n7191, Z => n7642);
   U512 : NAND3_X1 port map( A1 => n7918, A2 => n2569, A3 => n2568, ZN => n9116
                           );
   U9155 : OAI211_X1 port map( C1 => n8039, C2 => n8038, A => n8037, B => n2841
                           , ZN => n9123);
   U3349 : AND2_X1 port map( A1 => n7567, A2 => n7566, ZN => n9064);
   U192 : AND2_X1 port map( A1 => n7277, A2 => n7276, ZN => n8886);
   U902 : INV_X1 port map( A => n9245, ZN => n9410);
   U3367 : NAND3_X1 port map( A1 => n3034, A2 => n7602, A3 => n7603, ZN => 
                           n8787);
   U302 : OAI211_X1 port map( C1 => n7297, C2 => n8159, A => n7158, B => n7296,
                           ZN => n9243);
   U371 : NAND2_X1 port map( A1 => n1033, A2 => n1032, ZN => n8977);
   U4523 : NAND2_X1 port map( A1 => n1139, A2 => n5989, ZN => n8873);
   U249 : INV_X1 port map( A => n8635, ZN => n8653);
   U15171 : INV_X1 port map( A => n7679, ZN => n9438);
   U2030 : INV_X1 port map( A => n8735, ZN => n8731);
   U768 : AND2_X1 port map( A1 => n7066, A2 => n7065, ZN => n2238);
   U201 : AOI21_X1 port map( B1 => n7860, B2 => n7859, A => n1614, ZN => n10353
                           );
   U3283 : AND3_X1 port map( A1 => n9251, A2 => n9250, A3 => n9249, ZN => n9785
                           );
   U3284 : OAI21_X1 port map( B1 => n9174, B2 => n9173, A => n9172, ZN => 
                           n10391);
   U3286 : AND3_X1 port map( A1 => n3718, A2 => n4932, A3 => n1047, ZN => n9446
                           );
   U4464 : OAI21_X1 port map( B1 => n9174, B2 => n8963, A => n8470, ZN => 
                           n10263);
   U1317 : NAND2_X1 port map( A1 => n3101, A2 => n240, ZN => n10202);
   U8678 : MUX2_X1 port map( A => n8668, B => n8667, S => n8666, Z => n10133);
   U3260 : OR2_X1 port map( A1 => n8633, A2 => n8632, ZN => n9986);
   U5590 : OR2_X1 port map( A1 => n8374, A2 => n8373, ZN => n1895);
   U9241 : NAND2_X1 port map( A1 => n8815, A2 => n2899, ZN => n9852);
   U3247 : XNOR2_X1 port map( A => n748, B => n10064, ZN => n10332);
   U3252 : NAND2_X1 port map( A1 => n8571, A2 => n9378, ZN => n10311);
   U11328 : XNOR2_X1 port map( A => n10341, B => n10340, ZN => n11282);
   U16033 : XNOR2_X1 port map( A => n9263, B => n9264, ZN => n10592);
   U11514 : XNOR2_X1 port map( A => n9394, B => n9395, ZN => n28405);
   U3211 : CLKBUF_X1 port map( A => n9608, Z => n10476);
   U683 : BUF_X2 port map( A => n10522, Z => n10523);
   U14235 : OR2_X1 port map( A1 => n11127, A2 => n11123, ZN => n10760);
   U8939 : OR2_X1 port map( A1 => n28204, A2 => n11045, ZN => n11262);
   U311 : AND2_X1 port map( A1 => n4405, A2 => n11494, ZN => n12307);
   U3131 : NAND2_X1 port map( A1 => n11658, A2 => n11657, ZN => n12162);
   U2239 : NAND2_X1 port map( A1 => n6248, A2 => n10100, ZN => n3653);
   U10478 : NAND2_X1 port map( A1 => n10584, A2 => n3533, ZN => n12354);
   U8188 : OR2_X1 port map( A1 => n11279, A2 => n11278, ZN => n11795);
   U17369 : INV_X1 port map( A => n11801, ZN => n12286);
   U5650 : OR3_X1 port map( A1 => n4844, A2 => n12200, A3 => n12202, ZN => 
                           n5524);
   U1454 : CLKBUF_X1 port map( A => n12286, Z => n12401);
   U3089 : OAI22_X1 port map( A1 => n5079, A2 => n11673, B1 => n11848, B2 => 
                           n11672, ZN => n11846);
   U234 : NAND2_X1 port map( A1 => n11936, A2 => n11935, ZN => n13265);
   U3102 : OR2_X1 port map( A1 => n1493, A2 => n11550, ZN => n11160);
   U79 : OAI211_X1 port map( C1 => n11518, C2 => n11674, A => n11517, B => 
                           n11516, ZN => n12780);
   U1990 : AND2_X1 port map( A1 => n2355, A2 => n4711, ZN => n6645);
   U1410 : OAI21_X1 port map( B1 => n11846, B2 => n11679, A => n11678, ZN => 
                           n13553);
   U256 : AND2_X1 port map( A1 => n11504, A2 => n11503, ZN => n12722);
   U2081 : XNOR2_X1 port map( A => n13123, B => n13124, ZN => n14131);
   U1985 : XNOR2_X1 port map( A => n13135, B => n3097, ZN => n14325);
   U417 : XNOR2_X1 port map( A => n13399, B => n2875, ZN => n2974);
   U18094 : XNOR2_X1 port map( A => n12494, B => n12493, ZN => n14429);
   U18469 : NAND3_X1 port map( A1 => n28625, A2 => n14286, A3 => n14281, ZN => 
                           n12936);
   U18167 : XNOR2_X1 port map( A => n12565, B => n12564, ZN => n14318);
   U2980 : OR2_X1 port map( A1 => n14350, A2 => n13825, ZN => n1748);
   U1980 : OR2_X1 port map( A1 => n14240, A2 => n563, ZN => n14244);
   U10034 : OR2_X1 port map( A1 => n14244, A2 => n15199, ZN => n14245);
   U819 : OAI21_X1 port map( B1 => n4122, B2 => n4121, A => n13125, ZN => 
                           n15073);
   U372 : AOI21_X1 port map( B1 => n14067, B2 => n14328, A => n14066, ZN => 
                           n15285);
   U19343 : OAI211_X1 port map( C1 => n14386, C2 => n14385, A => n14384, B => 
                           n14383, ZN => n15275);
   U14236 : CLKBUF_X1 port map( A => n14806, Z => n28493);
   U420 : NAND3_X1 port map( A1 => n645, A2 => n643, A3 => n642, ZN => n15438);
   U6879 : OR2_X1 port map( A1 => n5635, A2 => n15456, ZN => n14797);
   U4646 : BUF_X1 port map( A => n13979, Z => n14740);
   U2921 : NAND2_X1 port map( A1 => n974, A2 => n973, ZN => n15185);
   U10271 : MUX2_X1 port map( A => n14988, B => n14987, S => n15155, Z => 
                           n16519);
   U1639 : OAI211_X1 port map( C1 => n14559, C2 => n14558, A => n14557, B => 
                           n14556, ZN => n16618);
   U686 : AND2_X1 port map( A1 => n6673, A2 => n6672, ZN => n16467);
   U2872 : OR2_X1 port map( A1 => n13984, A2 => n13983, ZN => n15788);
   U19692 : OAI21_X1 port map( B1 => n1809, B2 => n14958, A => n14957, ZN => 
                           n16296);
   U6796 : NAND3_X1 port map( A1 => n150, A2 => n14758, A3 => n14759, ZN => 
                           n16578);
   U2866 : INV_X1 port map( A => n15618, ZN => n16400);
   U214 : NAND3_X1 port map( A1 => n5, A2 => n14867, A3 => n2, ZN => n16456);
   U11559 : NOR2_X1 port map( A1 => n5596, A2 => n15172, ZN => n16264);
   U5849 : XNOR2_X1 port map( A => n15838, B => n15837, ZN => n17556);
   U4538 : XNOR2_X1 port map( A => n16158, B => n16157, ZN => n17464);
   U1053 : XNOR2_X1 port map( A => n4588, B => n16055, ZN => n17283);
   U20127 : BUF_X1 port map( A => n16943, Z => n17549);
   U2814 : INV_X1 port map( A => n17433, ZN => n17440);
   U965 : XNOR2_X1 port map( A => n15258, B => n15257, ZN => n6002);
   U2783 : BUF_X1 port map( A => n16883, Z => n17527);
   U328 : OR2_X1 port map( A1 => n17432, A2 => n17431, ZN => n31);
   U6976 : OR2_X1 port map( A1 => n17781, A2 => n17782, ZN => n4044);
   U1267 : AND2_X1 port map( A1 => n16966, A2 => n6224, ZN => n17858);
   U20249 : NOR2_X1 port map( A1 => n18063, A2 => n18064, ZN => n15939);
   U6428 : OR2_X1 port map( A1 => n18186, A2 => n527, ZN => n2135);
   U2685 : OR2_X1 port map( A1 => n757, A2 => n18343, ZN => n4077);
   U8519 : OAI211_X1 port map( C1 => n17676, C2 => n18487, A => n17675, B => 
                           n2459, ZN => n3444);
   U2680 : OAI211_X1 port map( C1 => n4943, C2 => n5223, A => n3349, B => n3350
                           , ZN => n16990);
   U731 : NOR2_X1 port map( A1 => n18714, A2 => n18713, ZN => n19075);
   U524 : AND2_X1 port map( A1 => n17723, A2 => n17722, ZN => n19656);
   U2659 : NAND3_X1 port map( A1 => n18436, A2 => n18435, A3 => n18434, ZN => 
                           n19207);
   U2629 : XNOR2_X1 port map( A => n5523, B => n5520, ZN => n20295);
   U2630 : XNOR2_X1 port map( A => n18775, B => n6667, ZN => n19761);
   U22372 : XNOR2_X1 port map( A => n19223, B => n19224, ZN => n20342);
   U21923 : XNOR2_X1 port map( A => n18673, B => n18674, ZN => n20374);
   U2614 : XNOR2_X1 port map( A => n5224, B => n17171, ZN => n20404);
   U691 : XNOR2_X1 port map( A => n18694, B => n18693, ZN => n20373);
   U6105 : OR2_X1 port map( A1 => n4245, A2 => n19928, ZN => n20645);
   U7077 : OR2_X1 port map( A1 => n20645, A2 => n5783, ZN => n5781);
   U2533 : NAND3_X1 port map( A1 => n20257, A2 => n20256, A3 => n1564, ZN => 
                           n21429);
   U2543 : INV_X1 port map( A => n20966, ZN => n21217);
   U22855 : OAI21_X1 port map( B1 => n19942, B2 => n19955, A => n19941, ZN => 
                           n21400);
   U23260 : INV_X1 port map( A => n21343, ZN => n21242);
   U2506 : BUF_X1 port map( A => n21014, Z => n22402);
   U1904 : NAND2_X1 port map( A1 => n20058, A2 => n20057, ZN => n21213);
   U2514 : OR2_X1 port map( A1 => n19893, A2 => n19894, ZN => n21567);
   U2481 : AND3_X1 port map( A1 => n6733, A2 => n20768, A3 => n6731, ZN => 
                           n22240);
   U24385 : XNOR2_X1 port map( A => n22327, B => n22328, ZN => n22651);
   U24216 : XNOR2_X1 port map( A => n22118, B => n22117, ZN => n22121);
   U2424 : BUF_X1 port map( A => n23102, Z => n23431);
   U227 : XNOR2_X1 port map( A => n22484, B => n22483, ZN => n28460);
   U5614 : XNOR2_X1 port map( A => n21873, B => n21874, ZN => n1914);
   U1895 : XNOR2_X1 port map( A => n21057, B => n21056, ZN => n23679);
   U161 : BUF_X1 port map( A => n23213, Z => n23403);
   U488 : XNOR2_X1 port map( A => n21928, B => n21927, ZN => n23799);
   U22929 : OAI21_X1 port map( B1 => n28390, B2 => n2138, A => n23313, ZN => 
                           n23565);
   U1678 : AND2_X1 port map( A1 => n23264, A2 => n23265, ZN => n25005);
   U24827 : MUX2_X1 port map( A => n23007, B => n23524, S => n23663, Z => 
                           n23009);
   U11924 : NAND2_X1 port map( A1 => n23264, A2 => n23265, ZN => n28415);
   U25233 : NOR2_X1 port map( A1 => n23782, A2 => n23781, ZN => n24801);
   U168 : OAI21_X1 port map( B1 => n23232, B2 => n1862, A => n23231, ZN => 
                           n24651);
   U1555 : OAI211_X1 port map( C1 => n23695, C2 => n5482, A => n5481, B => 
                           n5480, ZN => n24809);
   U4283 : NOR2_X1 port map( A1 => n22948, A2 => n22947, ZN => n24542);
   U174 : INV_X1 port map( A => n24378, ZN => n1828);
   U12517 : MUX2_X1 port map( A => n23133, B => n23132, S => n23678, Z => 
                           n24532);
   U12955 : AND2_X2 port map( A1 => n24544, A2 => n2054, ZN => n24547);
   U25549 : OAI211_X1 port map( C1 => n24237, C2 => n24236, A => n24235, B => 
                           n24234, ZN => n25745);
   U437 : MUX2_X1 port map( A => n24156, B => n24649, S => n3061, Z => n25261);
   U1544 : AOI21_X1 port map( B1 => n23027, B2 => n24310, A => n23026, ZN => 
                           n25910);
   U4492 : NAND2_X1 port map( A1 => n24080, A2 => n1128, ZN => n25251);
   U438 : BUF_X1 port map( A => n25844, Z => n363);
   U22309 : OAI21_X1 port map( B1 => n1777, B2 => n1828, A => n23094, ZN => 
                           n28628);
   U5081 : NAND3_X1 port map( A1 => n1495, A2 => n1653, A3 => n1652, ZN => 
                           n25262);
   U25089 : XNOR2_X1 port map( A => n23414, B => n23413, ZN => n26793);
   U2266 : XNOR2_X1 port map( A => n25078, B => n25077, ZN => n26920);
   U15484 : XNOR2_X1 port map( A => n25765, B => n25766, ZN => n26989);
   U7456 : INV_X1 port map( A => n26911, ZN => n5625);
   U6338 : AND2_X1 port map( A1 => n3589, A2 => n3590, ZN => n27819);
   U2193 : OR2_X1 port map( A1 => n27725, A2 => n27724, ZN => n26889);
   U2206 : AND2_X1 port map( A1 => n1944, A2 => n5373, ZN => n27382);
   U22972 : BUF_X1 port map( A => n27997, Z => n28636);
   U12488 : CLKBUF_X1 port map( A => n27913, Z => n1843);
   U2097 : CLKBUF_X1 port map( A => Key(30), Z => n3423);
   U1603 : CLKBUF_X1 port map( A => Key(144), Z => n28327);
   U11983 : NAND2_X1 port map( A1 => n10687, A2 => n10963, ZN => n10966);
   U3138 : OR2_X1 port map( A1 => n10168, A2 => n10167, ZN => n12125);
   U1558 : OR2_X1 port map( A1 => n11877, A2 => n10868, ZN => n1630);
   U1455 : NAND2_X1 port map( A1 => n6645, A2 => n11361, ZN => n6647);
   U13059 : CLKBUF_X1 port map( A => n17541, Z => n28454);
   U11129 : INV_X1 port map( A => n17478, ZN => n3883);
   U20340 : INV_X1 port map( A => n16904, ZN => n17710);
   U21390 : OAI21_X1 port map( B1 => n17736, B2 => n17735, A => n17734, ZN => 
                           n17965);
   U2608 : INV_X1 port map( A => n20324, ZN => n502);
   U2588 : OR2_X1 port map( A1 => n20020, A2 => n19795, ZN => n19796);
   U1508 : AOI21_X1 port map( B1 => n3973, B2 => n3974, A => n20586, ZN => 
                           n21134);
   U8285 : NAND2_X2 port map( A1 => n21611, A2 => n21610, ZN => n21326);
   U2353 : INV_X1 port map( A => n24367, ZN => n23897);
   U10287 : NOR2_X1 port map( A1 => n24650, A2 => n24155, ZN => n24524);
   U5925 : BUF_X1 port map( A => n26850, Z => n26849);
   U4002 : NOR2_X1 port map( A1 => n27898, A2 => n26510, ZN => n27904);
   U143 : NOR2_X1 port map( A1 => n28403, A2 => n27818, ZN => n27812);
   U26338 : NOR2_X1 port map( A1 => n27433, A2 => n27439, ZN => n27432);
   U870 : AND3_X2 port map( A1 => n2626, A2 => n2625, A3 => n2629, ZN => n8504)
                           ;
   U27190 : OR2_X2 port map( A1 => n5640, A2 => n5643, ZN => n16498);
   U453 : AND3_X2 port map( A1 => n782, A2 => n778, A3 => n781, ZN => n18242);
   U8286 : OR2_X2 port map( A1 => n7409, A2 => n2491, ZN => n9133);
   U8399 : NAND2_X2 port map( A1 => n2772, A2 => n7894, ZN => n8658);
   U1400 : BUF_X2 port map( A => n17474, Z => n16725);
   U21643 : AND2_X2 port map( A1 => n18207, A2 => n18208, ZN => n19491);
   U4311 : BUF_X1 port map( A => n19855, Z => n20552);
   U3012 : BUF_X2 port map( A => n13744, Z => n14254);
   U409 : OAI211_X2 port map( C1 => n13769, C2 => n15199, A => n13741, B => 
                           n13740, ZN => n15379);
   U11685 : AND2_X2 port map( A1 => n4390, A2 => n10744, ZN => n11671);
   U3282 : OAI21_X2 port map( B1 => n9002, B2 => n9200, A => n4302, ZN => 
                           n10426);
   U1160 : NAND4_X2 port map( A1 => n7735, A2 => n7031, A3 => n7032, A4 => 
                           n3115, ZN => n8874);
   U5074 : AND2_X2 port map( A1 => n1490, A2 => n1489, ZN => n13380);
   U9006 : OAI211_X2 port map( C1 => n21544, C2 => n21543, A => n2725, B => 
                           n2724, ZN => n21980);
   U45 : AND4_X2 port map( A1 => n2857, A2 => n2856, A3 => n17507, A4 => n2858,
                           ZN => n520);
   U1252 : AOI21_X2 port map( B1 => n8791, B2 => n8787, A => n8723, ZN => n9877
                           );
   U1084 : BUF_X2 port map( A => n23867, Z => n24716);
   U1520 : BUF_X2 port map( A => n11037, Z => n279);
   U1063 : OAI211_X2 port map( C1 => n12162, C2 => n10897, A => n10896, B => 
                           n11843, ZN => n13556);
   U25717 : OR2_X2 port map( A1 => n28689, A2 => n7757, ZN => n10022);
   U5069 : OR2_X2 port map( A1 => n19884, A2 => n19885, ZN => n4193);
   U466 : AND3_X2 port map( A1 => n1307, A2 => n1306, A3 => n2234, ZN => n18017
                           );
   U8411 : NAND3_X2 port map( A1 => n11342, A2 => n11343, A3 => n2580, ZN => 
                           n12281);
   U1615 : XNOR2_X2 port map( A => n18004, B => n18005, ZN => n20200);
   U24300 : AND2_X2 port map( A1 => n22217, A2 => n22216, ZN => n24735);
   U17451 : BUF_X2 port map( A => n13017, Z => n12894);
   U1125 : NAND2_X2 port map( A1 => n17874, A2 => n1034, ZN => n19643);
   U4436 : AND2_X2 port map( A1 => n1102, A2 => n1101, ZN => n13260);
   U3278 : OAI211_X2 port map( C1 => n9105, C2 => n9104, A => n4969, B => n9121
                           , ZN => n4714);
   U112 : NOR2_X1 port map( A1 => n3127, A2 => n3128, ZN => n9430);
   U10250 : AND2_X2 port map( A1 => n3392, A2 => n3391, ZN => n24383);
   U5852 : AND4_X2 port map( A1 => n17189, A2 => n4168, A3 => n4480, A4 => 
                           n4241, ZN => n18410);
   U9677 : XNOR2_X2 port map( A => n18363, B => n18362, ZN => n20546);
   U7358 : BUF_X2 port map( A => n7192, Z => n7985);
   U10892 : AND2_X2 port map( A1 => n6076, A2 => n6078, ZN => n19225);
   U3879 : NOR2_X2 port map( A1 => n5626, A2 => n5627, ZN => n2209);
   U1989 : XNOR2_X2 port map( A => n13409, B => n13408, ZN => n1368);
   U9136 : XNOR2_X2 port map( A => n13605, B => n13604, ZN => n17425);
   U14976 : OR2_X2 port map( A1 => n7392, A2 => n7391, ZN => n9132);
   U1278 : AND2_X2 port map( A1 => n2947, A2 => n10109, ZN => n11990);
   U912 : NAND3_X2 port map( A1 => n15442, A2 => n5681, A3 => n15443, ZN => 
                           n16303);
   U1301 : NOR2_X2 port map( A1 => n27900, A2 => n27899, ZN => n27919);
   U1043 : OAI21_X2 port map( B1 => n7961, B2 => n7960, A => n3368, ZN => n8666
                           );
   U9858 : OAI211_X2 port map( C1 => n8496, C2 => n8495, A => n8494, B => n8493
                           , ZN => n9771);
   U571 : BUF_X2 port map( A => n7040, Z => n7982);
   U4367 : NAND3_X2 port map( A1 => n1107, A2 => n11916, A3 => n11917, ZN => 
                           n13482);
   U14504 : AND2_X2 port map( A1 => n7014, A2 => n7013, ZN => n8881);
   U7409 : AOI21_X2 port map( B1 => n16754, B2 => n16753, A => n16752, ZN => 
                           n18179);
   U564 : AND3_X2 port map( A1 => n2162, A2 => n2073, A3 => n2160, ZN => n15780
                           );
   U3268 : NAND3_X2 port map( A1 => n8190, A2 => n8189, A3 => n8188, ZN => 
                           n9295);
   U3462 : XNOR2_X2 port map( A => Key(116), B => Plaintext(116), ZN => n7935);
   U897 : NAND3_X2 port map( A1 => n1020, A2 => n13304, A3 => n13303, ZN => 
                           n15690);
   U10092 : OAI21_X2 port map( B1 => n19746, B2 => n4362, A => n19745, ZN => 
                           n22141);
   U946 : AND2_X2 port map( A1 => n169, A2 => n168, ZN => n16579);
   U2662 : AND2_X2 port map( A1 => n17776, A2 => n17777, ZN => n19481);
   U1329 : AND2_X2 port map( A1 => n6743, A2 => n4733, ZN => n4298);
   U2891 : OAI21_X2 port map( B1 => n15180, B2 => n15181, A => n15179, ZN => 
                           n15850);
   U424 : XNOR2_X2 port map( A => n21206, B => n21205, ZN => n23131);
   U1716 : XNOR2_X2 port map( A => n15455, B => n15454, ZN => n17415);
   U21723 : OAI21_X2 port map( B1 => n18394, B2 => n18393, A => n18392, ZN => 
                           n18863);
   U14473 : XNOR2_X2 port map( A => n6997, B => Key(122), ZN => n7909);
   U1413 : NAND3_X1 port map( A1 => n4584, A2 => n7442, A3 => n7443, ZN => 
                           n9754);
   U12843 : NAND3_X1 port map( A1 => n9061, A2 => n9062, A3 => n9060, ZN => 
                           n5537);
   U16942 : OAI211_X1 port map( C1 => n11322, C2 => n11181, A => n10475, B => 
                           n10474, ZN => n12338);
   U3114 : AND2_X1 port map( A1 => n11428, A2 => n11426, ZN => n11487);
   U1072 : NAND3_X1 port map( A1 => n10885, A2 => n11028, A3 => n10886, ZN => 
                           n12164);
   U8134 : AND2_X1 port map( A1 => n2295, A2 => n2294, ZN => n15423);
   U5546 : OAI21_X1 port map( B1 => n15232, B2 => n15231, A => n15230, ZN => 
                           n16271);
   U19506 : NAND4_X1 port map( A1 => n14649, A2 => n14648, A3 => n14647, A4 => 
                           n14646, ZN => n15817);
   U109 : AND3_X1 port map( A1 => n16672, A2 => n16671, A3 => n16670, ZN => 
                           n17947);
   U3609 : OAI21_X1 port map( B1 => n19811, B2 => n20285, A => n19813, ZN => 
                           n20864);
   U13021 : NAND3_X1 port map( A1 => n24571, A2 => n24570, A3 => n24569, ZN => 
                           n25696);
   U1664 : OAI21_X2 port map( B1 => n26444, B2 => n26950, A => n26443, ZN => 
                           n27300);
   U10 : AOI21_X1 port map( B1 => n21225, B2 => n21224, A => n21223, ZN => 
                           n28517);
   U11 : AND2_X1 port map( A1 => n17060, A2 => n18337, ZN => n29204);
   U28 : BUF_X1 port map( A => n10816, Z => n28157);
   U151 : BUF_X1 port map( A => n10472, Z => n11183);
   U203 : AND4_X2 port map( A1 => n20731, A2 => n20732, A3 => n20730, A4 => 
                           n4776, ZN => n21990);
   U236 : INV_X2 port map( A => n15400, ZN => n28196);
   U238 : OAI211_X2 port map( C1 => n5956, C2 => n5285, A => n5284, B => n5283,
                           ZN => n15183);
   U240 : AND2_X2 port map( A1 => n16848, A2 => n16849, ZN => n18423);
   U265 : MUX2_X2 port map( A => n23869, B => n23868, S => n24720, Z => n26040)
                           ;
   U266 : AOI21_X2 port map( B1 => n14711, B2 => n14598, A => n14710, ZN => 
                           n16568);
   U283 : AND3_X2 port map( A1 => n3245, A2 => n23616, A3 => n23617, ZN => 
                           n24791);
   U330 : OAI211_X1 port map( C1 => n14006, C2 => n14007, A => n6106, B => 
                           n6105, ZN => n15431);
   U345 : XNOR2_X1 port map( A => n16449, B => n16305, ZN => n16154);
   U349 : BUF_X1 port map( A => n22953, Z => n23846);
   U356 : BUF_X1 port map( A => n20207, Z => n21674);
   U357 : OAI211_X1 port map( C1 => n17905, C2 => n18456, A => n3865, B => 
                           n3864, ZN => n19346);
   U358 : BUF_X1 port map( A => n26452, Z => n29105);
   U363 : NOR2_X1 port map( A1 => n15334, A2 => n15338, ZN => n28766);
   U376 : NOR2_X1 port map( A1 => n14569, A2 => n15071, ZN => n28767);
   U382 : XOR2_X1 port map( A => n15330, B => n15329, Z => n28768);
   U387 : OAI21_X2 port map( B1 => n19876, B2 => n19985, A => n19875, ZN => 
                           n21159);
   U389 : NOR2_X2 port map( A1 => n24774, A2 => n24773, ZN => n29046);
   U407 : XNOR2_X2 port map( A => n25524, B => n25523, ZN => n29058);
   U415 : OAI21_X2 port map( B1 => n5546, B2 => n26771, A => n6769, ZN => 
                           n27497);
   U416 : OAI21_X2 port map( B1 => n27116, B2 => n27115, A => n27114, ZN => 
                           n29049);
   U422 : OAI211_X2 port map( C1 => n17523, C2 => n18220, A => n17533, B => 
                           n1943, ZN => n19377);
   U427 : OAI211_X2 port map( C1 => n8771, C2 => n8770, A => n8769, B => n8768,
                           ZN => n9908);
   U434 : XNOR2_X2 port map( A => n13508, B => n13507, ZN => n14036);
   U441 : OAI211_X1 port map( C1 => n23072, C2 => n24712, A => n29249, B => 
                           n29248, ZN => n25908);
   U458 : NAND3_X2 port map( A1 => n3857, A2 => n3858, A3 => n21189, ZN => 
                           n22068);
   U465 : NOR2_X2 port map( A1 => n21238, A2 => n952, ZN => n22278);
   U481 : NAND3_X2 port map( A1 => n28274, A2 => n1654, A3 => n1424, ZN => 
                           n26070);
   U495 : XNOR2_X1 port map( A => Plaintext(137), B => Key(137), ZN => n8300);
   U508 : NAND2_X2 port map( A1 => n3647, A2 => n3646, ZN => n13338);
   U528 : BUF_X1 port map( A => n17175, Z => n28775);
   U530 : CLKBUF_X1 port map( A => n17175, Z => n28776);
   U531 : XNOR2_X1 port map( A => n16357, B => n16356, ZN => n17175);
   U573 : AND2_X1 port map( A1 => n572, A2 => n11754, ZN => n28878);
   U578 : AND2_X2 port map( A1 => n6084, A2 => n6082, ZN => n21448);
   U597 : OAI211_X2 port map( C1 => n9167, C2 => n9163, A => n8317, B => n8316,
                           ZN => n28488);
   U604 : NAND2_X2 port map( A1 => n828, A2 => n829, ZN => n15515);
   U620 : AND2_X1 port map( A1 => n25418, A2 => n26576, ZN => n26574);
   U622 : XNOR2_X1 port map( A => n9576, B => n9577, ZN => n9933);
   U628 : XNOR2_X2 port map( A => n18971, B => n18970, ZN => n20219);
   U637 : NAND2_X2 port map( A1 => n6557, A2 => n6558, ZN => n23126);
   U639 : XNOR2_X2 port map( A => n9483, B => n9482, ZN => n2690);
   U696 : NAND3_X2 port map( A1 => n2312, A2 => n1962, A3 => n3492, ZN => 
                           n22628);
   U719 : NOR2_X2 port map( A1 => n18352, A2 => n5920, ZN => n18900);
   U725 : XNOR2_X2 port map( A => n10400, B => n10399, ZN => n10431);
   U747 : INV_X2 port map( A => n852, ZN => n27357);
   U750 : XNOR2_X2 port map( A => n22367, B => n22366, ZN => n23621);
   U787 : XNOR2_X1 port map( A => n17684, B => n19336, ZN => n28140);
   U790 : XNOR2_X2 port map( A => n7007, B => Key(69), ZN => n7846);
   U811 : XNOR2_X1 port map( A => n9022, B => n9021, ZN => n5595);
   U820 : NOR2_X2 port map( A1 => n21434, A2 => n4311, ZN => n22333);
   U829 : AOI21_X2 port map( B1 => n10600, B2 => n10601, A => n10599, ZN => 
                           n11740);
   U891 : BUF_X2 port map( A => n24650, Z => n28785);
   U906 : OAI211_X1 port map( C1 => n23749, C2 => n23215, A => n5041, B => 
                           n3631, ZN => n24650);
   U929 : NAND3_X2 port map( A1 => n5609, A2 => n5610, A3 => n15646, ZN => 
                           n18489);
   U934 : XNOR2_X2 port map( A => n6968, B => Key(103), ZN => n7619);
   U950 : OAI211_X2 port map( C1 => n13128, C2 => n15082, A => n13127, B => 
                           n4169, ZN => n16476);
   U951 : NAND3_X2 port map( A1 => n28938, A2 => n8997, A3 => n3056, ZN => 
                           n9639);
   U963 : NOR2_X2 port map( A1 => n24495, A2 => n24494, ZN => n25849);
   U977 : XNOR2_X2 port map( A => n19581, B => n19580, ZN => n20323);
   U995 : XNOR2_X2 port map( A => n15570, B => n15569, ZN => n17336);
   U1018 : XNOR2_X2 port map( A => n9182, B => n9181, ZN => n11347);
   U1035 : OAI21_X2 port map( B1 => n19781, B2 => n19754, A => n19753, ZN => 
                           n22145);
   U1036 : NOR2_X2 port map( A1 => n21247, A2 => n21246, ZN => n22204);
   U1087 : XNOR2_X2 port map( A => n7043, B => Key(151), ZN => n7981);
   U1112 : OAI211_X2 port map( C1 => n8209, C2 => n7842, A => n1612, B => 
                           n28365, ZN => n8908);
   U1128 : INV_X1 port map( A => n24668, ZN => n4195);
   U1131 : NAND3_X1 port map( A1 => n21641, A2 => n21640, A3 => n3313, ZN => 
                           n22180);
   U1138 : INV_X1 port map( A => n22023, ZN => n28790);
   U1147 : INV_X1 port map( A => n21327, ZN => n28791);
   U1164 : OR2_X2 port map( A1 => n20741, A2 => n20736, ZN => n20858);
   U1168 : NAND3_X1 port map( A1 => n2135, A2 => n2136, A3 => n18191, ZN => 
                           n19486);
   U1170 : INV_X2 port map( A => n17798, ZN => n18456);
   U1175 : INV_X1 port map( A => n5891, ZN => n28792);
   U1177 : INV_X1 port map( A => n17354, ZN => n28793);
   U1192 : INV_X1 port map( A => n12354, ZN => n29209);
   U1201 : INV_X1 port map( A => n10875, ZN => n11220);
   U1211 : NAND2_X1 port map( A1 => n8562, A2 => n9144, ZN => n8937);
   U1217 : CLKBUF_X1 port map( A => Key(171), Z => n2986);
   U1219 : CLKBUF_X1 port map( A => Key(89), Z => n2477);
   U1229 : CLKBUF_X1 port map( A => Key(185), Z => n2465);
   U1234 : CLKBUF_X1 port map( A => Key(189), Z => n3554);
   U1236 : CLKBUF_X1 port map( A => Key(59), Z => n3223);
   U1263 : AND2_X1 port map( A1 => n4485, A2 => n27047, ZN => n27092);
   U1268 : AND2_X1 port map( A1 => n29029, A2 => n29030, ZN => n27944);
   U1279 : OAI21_X1 port map( B1 => n26253, B2 => n26735, A => n26252, ZN => 
                           n28066);
   U1315 : BUF_X1 port map( A => n25465, Z => n25782);
   U1316 : OAI21_X1 port map( B1 => n23144, B2 => n24229, A => n24895, ZN => 
                           n25134);
   U1339 : NAND3_X1 port map( A1 => n5293, A2 => n5292, A3 => n22499, ZN => 
                           n29109);
   U1340 : INV_X1 port map( A => n5763, ZN => n23284);
   U1344 : OR2_X1 port map( A1 => n22877, A2 => n23810, ZN => n5763);
   U1372 : INV_X1 port map( A => n23317, ZN => n28963);
   U1388 : BUF_X1 port map( A => n23250, Z => n28796);
   U1390 : AND2_X1 port map( A1 => n22174, A2 => n23587, ZN => n28824);
   U1398 : XNOR2_X1 port map( A => n21916, B => n21915, ZN => n23795);
   U1409 : OAI21_X1 port map( B1 => n21153, B2 => n21152, A => n21151, ZN => 
                           n22419);
   U1424 : OR2_X1 port map( A1 => n21462, A2 => n21457, ZN => n28941);
   U1426 : OAI21_X1 port map( B1 => n20998, B2 => n21217, A => n28979, ZN => 
                           n18788);
   U1427 : AND2_X1 port map( A1 => n4344, A2 => n28937, ZN => n21321);
   U1434 : NOR2_X1 port map( A1 => n22025, A2 => n22026, ZN => n22028);
   U1435 : NAND4_X1 port map( A1 => n21217, A2 => n21218, A3 => n19914, A4 => 
                           n28980, ZN => n28979);
   U1462 : AND2_X1 port map( A1 => n21135, A2 => n21134, ZN => n28937);
   U1463 : INV_X1 port map( A => n21394, ZN => n28797);
   U1466 : AND3_X1 port map( A1 => n28812, A2 => n29182, A3 => n29180, ZN => 
                           n21749);
   U1498 : OAI21_X1 port map( B1 => n28133, B2 => n20517, A => n28992, ZN => 
                           n19457);
   U1522 : XNOR2_X1 port map( A => n19121, B => n19120, ZN => n20498);
   U1527 : XNOR2_X1 port map( A => n19346, B => n19486, ZN => n19141);
   U1534 : AND2_X1 port map( A1 => n1708, A2 => n18177, ZN => n28981);
   U1537 : NAND3_X1 port map( A1 => n28827, A2 => n28826, A3 => n17999, ZN => 
                           n19428);
   U1541 : NAND2_X1 port map( A1 => n17785, A2 => n28978, ZN => n19378);
   U1567 : NAND3_X1 port map( A1 => n18080, A2 => n18079, A3 => n46, ZN => 
                           n19448);
   U1588 : OAI211_X1 port map( C1 => n15939, C2 => n15938, A => n15936, B => 
                           n29007, ZN => n19403);
   U1591 : AND2_X1 port map( A1 => n18423, A2 => n17802, ZN => n29274);
   U1600 : OR2_X1 port map( A1 => n16985, A2 => n18188, ZN => n29199);
   U1601 : OR2_X1 port map( A1 => n18170, A2 => n4044, ZN => n5203);
   U1605 : NAND2_X1 port map( A1 => n29203, A2 => n4583, ZN => n18338);
   U1616 : INV_X1 port map( A => n18135, ZN => n526);
   U1618 : NAND2_X1 port map( A1 => n16708, A2 => n1129, ZN => n18198);
   U1620 : AND2_X1 port map( A1 => n28831, A2 => n2600, ZN => n17132);
   U1630 : NAND2_X1 port map( A1 => n1088, A2 => n16818, ZN => n18172);
   U1631 : OR2_X1 port map( A1 => n2600, A2 => n17129, ZN => n5733);
   U1653 : INV_X1 port map( A => n17455, ZN => n28801);
   U1670 : NAND3_X1 port map( A1 => n28816, A2 => n1164, A3 => n28818, ZN => 
                           n16160);
   U1694 : AND3_X1 port map( A1 => n29012, A2 => n29011, A3 => n29010, ZN => 
                           n16395);
   U1696 : NAND2_X1 port map( A1 => n14951, A2 => n28896, ZN => n15999);
   U1720 : NOR2_X1 port map( A1 => n14682, A2 => n14681, ZN => n15802);
   U1721 : NOR2_X1 port map( A1 => n14952, A2 => n15082, ZN => n28897);
   U1735 : OR2_X1 port map( A1 => n14990, A2 => n14989, ZN => n3208);
   U1745 : AND3_X1 port map( A1 => n734, A2 => n735, A3 => n12936, ZN => n15082
                           );
   U1747 : INV_X1 port map( A => n15333, ZN => n28802);
   U1748 : BUF_X2 port map( A => n14981, Z => n28803);
   U1750 : OR2_X1 port map( A1 => n13699, A2 => n13306, ZN => n28950);
   U1762 : AND2_X1 port map( A1 => n13826, A2 => n14354, ZN => n28899);
   U1809 : INV_X1 port map( A => n14401, ZN => n28804);
   U1842 : INV_X1 port map( A => n14455, ZN => n28806);
   U1859 : NAND2_X1 port map( A1 => n2319, A2 => n11850, ZN => n12872);
   U1890 : NAND3_X1 port map( A1 => n29264, A2 => n11841, A3 => n4447, ZN => 
                           n12787);
   U1926 : OR2_X1 port map( A1 => n12030, A2 => n12031, ZN => n1192);
   U1939 : OAI22_X1 port map( A1 => n12299, A2 => n12300, B1 => n11769, B2 => 
                           n4197, ZN => n5020);
   U1956 : OR2_X1 port map( A1 => n11553, A2 => n11785, ZN => n29291);
   U1974 : AND3_X1 port map( A1 => n28811, A2 => n3449, A3 => n6361, ZN => 
                           n11751);
   U1983 : INV_X1 port map( A => n569, ZN => n28807);
   U2108 : NAND3_X1 port map( A1 => n2868, A2 => n2867, A3 => n6242, ZN => 
                           n11921);
   U2207 : AND2_X1 port map( A1 => n8109, A2 => n9245, ZN => n28911);
   U2216 : NAND2_X1 port map( A1 => n2310, A2 => n7346, ZN => n8185);
   U2219 : AND2_X1 port map( A1 => n2695, A2 => n28814, ZN => n8490);
   U2262 : INV_X1 port map( A => n8810, ZN => n28808);
   U2265 : NAND2_X1 port map( A1 => n29214, A2 => n7790, ZN => n8353);
   U2301 : NAND4_X1 port map( A1 => n7668, A2 => n901, A3 => n7667, A4 => n7666
                           , ZN => n8777);
   U2306 : MUX2_X1 port map( A => n7143, B => n7142, S => n7523, Z => n28913);
   U2329 : OR2_X1 port map( A1 => n7775, A2 => n7891, ZN => n5494);
   U2331 : XNOR2_X1 port map( A => n6971, B => Key(106), ZN => n7358);
   U2374 : INV_X1 port map( A => n9113, ZN => n28810);
   U2377 : OR2_X1 port map( A1 => n7017, A2 => n7690, ZN => n7502);
   U2435 : CLKBUF_X1 port map( A => n7851, Z => n371);
   U2445 : OR2_X1 port map( A1 => n8034, A2 => n7508, ZN => n8039);
   U2458 : AOI21_X1 port map( B1 => n9436, B2 => n8998, A => n9438, ZN => 
                           n28989);
   U2459 : OR2_X1 port map( A1 => n8868, A2 => n2006, ZN => n3788);
   U2463 : INV_X1 port map( A => n8490, ZN => n9099);
   U2477 : OAI211_X1 port map( C1 => n8036, C2 => n7514, A => n7513, B => n7512
                           , ZN => n8817);
   U2496 : OAI211_X1 port map( C1 => n8808, C2 => n28808, A => n29242, B => 
                           n29241, ZN => n2899);
   U2510 : AND2_X1 port map( A1 => n9213, A2 => n9212, ZN => n28858);
   U2540 : XNOR2_X1 port map( A => n10037, B => n9383, ZN => n10421);
   U2558 : AND2_X1 port map( A1 => n10808, A2 => n11149, ZN => n29263);
   U2578 : XNOR2_X1 port map( A => n10142, B => n10141, ZN => n11084);
   U2580 : INV_X1 port map( A => n12313, ZN => n12051);
   U2617 : NAND2_X1 port map( A1 => n10270, A2 => n28929, ZN => n28928);
   U2654 : OR2_X1 port map( A1 => n11486, A2 => n6482, ZN => n11793);
   U2669 : OR2_X1 port map( A1 => n12356, A2 => n11739, ZN => n919);
   U2693 : AND2_X1 port map( A1 => n11656, A2 => n28828, ZN => n11844);
   U2749 : MUX2_X1 port map( A => n10607, B => n10606, S => n10605, Z => n10608
                           );
   U2765 : OR2_X1 port map( A1 => n11853, A2 => n10905, ZN => n10906);
   U2766 : AND2_X1 port map( A1 => n11658, A2 => n11657, ZN => n28828);
   U2794 : OR2_X1 port map( A1 => n11911, A2 => n12363, ZN => n28961);
   U2800 : OAI21_X1 port map( B1 => n11639, B2 => n11672, A => n11671, ZN => 
                           n11518);
   U2806 : OR2_X1 port map( A1 => n11394, A2 => n11852, ZN => n28886);
   U2815 : OR2_X1 port map( A1 => n11686, A2 => n12000, ZN => n29175);
   U2817 : AND2_X1 port map( A1 => n11380, A2 => n11379, ZN => n28917);
   U2819 : INV_X1 port map( A => n29244, ZN => n29243);
   U2850 : NAND3_X1 port map( A1 => n11160, A2 => n11161, A3 => n1140, ZN => 
                           n13249);
   U2920 : BUF_X1 port map( A => n14171, Z => n29097);
   U2944 : AOI21_X1 port map( B1 => n6032, B2 => n13587, A => n58, ZN => n14041
                           );
   U2985 : OR2_X1 port map( A1 => n12744, A2 => n14465, ZN => n28936);
   U2987 : OR2_X1 port map( A1 => n14380, A2 => n14004, ZN => n14005);
   U3063 : OR2_X1 port map( A1 => n13824, A2 => n14126, ZN => n14357);
   U3070 : OR2_X1 port map( A1 => n14075, A2 => n14359, ZN => n28952);
   U3074 : OAI21_X1 port map( B1 => n14459, B2 => n13864, A => n13863, ZN => 
                           n15166);
   U3076 : NAND2_X1 port map( A1 => n14490, A2 => n14489, ZN => n15489);
   U3088 : INV_X1 port map( A => n15694, ZN => n29011);
   U3100 : OR2_X1 port map( A1 => n14837, A2 => n15290, ZN => n14521);
   U3121 : NOR2_X1 port map( A1 => n14601, A2 => n15284, ZN => n28842);
   U3134 : NOR2_X1 port map( A1 => n5596, A2 => n15172, ZN => n28406);
   U3151 : OAI21_X1 port map( B1 => n17160, B2 => n28497, A => n17162, ZN => 
                           n28852);
   U3175 : AND2_X1 port map( A1 => n17282, A2 => n17283, ZN => n29000);
   U3185 : INV_X1 port map( A => n17175, ZN => n16874);
   U3242 : OR2_X1 port map( A1 => n16614, A2 => n17496, ZN => n28993);
   U3255 : AND2_X1 port map( A1 => n4367, A2 => n4368, ZN => n17126);
   U3261 : AND2_X1 port map( A1 => n1880, A2 => n17249, ZN => n968);
   U3270 : INV_X1 port map( A => n16837, ZN => n17316);
   U3280 : OAI21_X1 port map( B1 => n1090, B2 => n29000, A => n29086, ZN => 
                           n28999);
   U3309 : OR2_X1 port map( A1 => n18710, A2 => n5023, ZN => n3766);
   U3334 : AND4_X2 port map( A1 => n16742, A2 => n16743, A3 => n16741, A4 => 
                           n16740, ZN => n18277);
   U3361 : BUF_X1 port map( A => n18057, Z => n1861);
   U3372 : OR2_X1 port map( A1 => n17403, A2 => n16904, ZN => n15934);
   U3408 : AOI22_X1 port map( A1 => n1963, A2 => n17996, B1 => n18382, B2 => 
                           n17997, ZN => n28826);
   U3449 : OR2_X1 port map( A1 => n18349, A2 => n18000, ZN => n28827);
   U3476 : NAND3_X1 port map( A1 => n4120, A2 => n4119, A3 => n5992, ZN => 
                           n18653);
   U3478 : XNOR2_X1 port map( A => n19603, B => n18767, ZN => n18768);
   U3548 : AND2_X1 port map( A1 => n20148, A2 => n20146, ZN => n28849);
   U3555 : OR2_X1 port map( A1 => n21090, A2 => n5817, ZN => n21931);
   U3558 : INV_X1 port map( A => n20286, ZN => n29166);
   U3566 : XNOR2_X1 port map( A => n18917, B => n18916, ZN => n29134);
   U3573 : XNOR2_X1 port map( A => n19169, B => n19168, ZN => n20495);
   U3596 : OAI21_X1 port map( B1 => n20307, B2 => n20305, A => n19948, ZN => 
                           n5194);
   U3600 : INV_X1 port map( A => n18919, ZN => n4877);
   U3617 : OR2_X1 port map( A1 => n29235, A2 => n20398, ZN => n20402);
   U3619 : INV_X1 port map( A => n1875, ZN => n28891);
   U3631 : OR2_X1 port map( A1 => n21539, A2 => n21503, ZN => n28991);
   U3637 : NAND2_X1 port map( A1 => n19930, A2 => n29183, ZN => n29182);
   U3638 : OR2_X1 port map( A1 => n20459, A2 => n20273, ZN => n29184);
   U3639 : CLKBUF_X1 port map( A => n28555, Z => n20117);
   U3646 : OR2_X1 port map( A1 => n20338, A2 => n29601, ZN => n28982);
   U3652 : NOR3_X1 port map( A1 => n20767, A2 => n29531, A3 => n20766, ZN => 
                           n21153);
   U3709 : INV_X1 port map( A => n21376, ZN => n29228);
   U3786 : OAI211_X1 port map( C1 => n21553, C2 => n21547, A => n1621, B => 
                           n28890, ZN => n21556);
   U3817 : INV_X1 port map( A => n21990, ZN => n22763);
   U3826 : AND2_X1 port map( A1 => n20712, A2 => n21269, ZN => n29256);
   U3847 : OR2_X1 port map( A1 => n23767, A2 => n23765, ZN => n23333);
   U3883 : INV_X1 port map( A => n22078, ZN => n28914);
   U3897 : OR2_X1 port map( A1 => n23267, A2 => n28581, ZN => n23217);
   U3898 : INV_X1 port map( A => n23353, ZN => n4232);
   U3909 : BUF_X1 port map( A => n22877, Z => n23808);
   U3910 : OR2_X1 port map( A1 => n23493, A2 => n23795, ZN => n23196);
   U3920 : MUX2_X1 port map( A => n23230, B => n23229, S => n22949, Z => n23231
                           );
   U3966 : INV_X1 port map( A => n24243, ZN => n24239);
   U3990 : OR2_X1 port map( A1 => n24246, A2 => n3061, ZN => n29002);
   U3993 : OR2_X1 port map( A1 => n24466, A2 => n24578, ZN => n29013);
   U4017 : OR2_X1 port map( A1 => n24612, A2 => n23922, ZN => n4639);
   U4049 : OR2_X1 port map( A1 => n462, A2 => n21303, ZN => n29015);
   U4086 : MUX2_X1 port map( A => n24048, B => n24047, S => n469, Z => n24049);
   U4136 : INV_X1 port map( A => n24532, ZN => n24894);
   U4137 : AND3_X1 port map( A1 => n24411, A2 => n24413, A3 => n24410, ZN => 
                           n2261);
   U4139 : OAI21_X1 port map( B1 => n4573, B2 => n4575, A => n4572, ZN => 
                           n24797);
   U4147 : AND2_X1 port map( A1 => n26868, A2 => n26865, ZN => n26870);
   U4152 : XNOR2_X1 port map( A => n25448, B => n25447, ZN => n26748);
   U4171 : BUF_X1 port map( A => n25365, Z => n26489);
   U4174 : INV_X1 port map( A => n27382, ZN => n29218);
   U4176 : OR2_X1 port map( A1 => n27591, A2 => n27594, ZN => n28967);
   U4204 : AND3_X1 port map( A1 => n25048, A2 => n25047, A3 => n25050, ZN => 
                           n28834);
   U4221 : CLKBUF_X1 port map( A => Key(71), Z => n3422);
   U4274 : XOR2_X1 port map( A => n10182, B => n10181, Z => n1851);
   U4285 : OR2_X1 port map( A1 => n10740, A2 => n10806, ZN => n28811);
   U4293 : OR2_X1 port map( A1 => n19931, A2 => n5783, ZN => n28812);
   U4307 : OR2_X1 port map( A1 => n20395, A2 => n20400, ZN => n28813);
   U4312 : AND2_X1 port map( A1 => n4834, A2 => n4833, ZN => n28814);
   U4330 : OR2_X1 port map( A1 => n24978, A2 => n24976, ZN => n28815);
   U4347 : OR2_X1 port map( A1 => n15395, A2 => n14633, ZN => n28816);
   U4357 : AND2_X1 port map( A1 => n15233, A2 => n15234, ZN => n28817);
   U4368 : INV_X1 port map( A => n7192, ZN => n7644);
   U4381 : INV_X1 port map( A => n2238, ZN => n29241);
   U4382 : NAND2_X1 port map( A1 => n7622, A2 => n7623, ZN => n9206);
   U4397 : INV_X1 port map( A => n14429, ZN => n28986);
   U4405 : OR2_X1 port map( A1 => n15391, A2 => n15390, ZN => n28818);
   U4406 : XNOR2_X1 port map( A => n16049, B => n16048, ZN => n16860);
   U4415 : OR2_X1 port map( A1 => n18170, A2 => n18168, ZN => n28819);
   U4419 : XOR2_X1 port map( A => n18748, B => n18747, Z => n28820);
   U4426 : XNOR2_X1 port map( A => n19531, B => n19530, ZN => n20265);
   U4427 : INV_X1 port map( A => n20702, ZN => n28980);
   U4446 : INV_X1 port map( A => n20619, ZN => n28894);
   U4451 : INV_X1 port map( A => n21932, ZN => n28916);
   U4455 : OR2_X1 port map( A1 => n23209, A2 => n22984, ZN => n28821);
   U4466 : OR2_X1 port map( A1 => n26374, A2 => n26440, ZN => n28822);
   U4476 : OR2_X1 port map( A1 => n29330, A2 => n26800, ZN => n28823);
   U4481 : NAND3_X1 port map( A1 => n21157, A2 => n21156, A3 => n20744, ZN => 
                           n19877);
   U4488 : NAND2_X1 port map( A1 => n23715, A2 => n28824, ZN => n23263);
   U4494 : NAND2_X1 port map( A1 => n9057, A2 => n9058, ZN => n9258);
   U4498 : NAND2_X1 port map( A1 => n1174, A2 => n28825, ZN => n11505);
   U4517 : OR2_X1 port map( A1 => n11320, A2 => n4650, ZN => n28825);
   U4518 : NAND2_X1 port map( A1 => n15222, A2 => n15223, ZN => n15351);
   U4525 : NAND3_X1 port map( A1 => n21597, A2 => n21598, A3 => n5720, ZN => 
                           n5719);
   U4548 : NAND3_X1 port map( A1 => n10959, A2 => n10958, A3 => n10778, ZN => 
                           n10603);
   U4567 : NAND3_X1 port map( A1 => n11820, A2 => n4028, A3 => n11816, ZN => 
                           n11823);
   U4569 : NAND2_X1 port map( A1 => n8234, A2 => n7358, ZN => n8239);
   U4578 : NAND2_X1 port map( A1 => n23969, A2 => n24479, ZN => n23553);
   U4585 : NAND2_X1 port map( A1 => n24046, A2 => n23968, ZN => n23969);
   U4618 : INV_X1 port map( A => n17070, ZN => n17072);
   U4661 : NAND2_X1 port map( A1 => n17829, A2 => n4270, ZN => n17070);
   U4678 : NOR2_X1 port map( A1 => n23311, A2 => n28829, ZN => n28358);
   U4688 : INV_X1 port map( A => n23556, ZN => n28829);
   U4701 : NAND2_X1 port map( A1 => n23628, A2 => n23309, ZN => n23556);
   U4720 : OAI21_X1 port map( B1 => n17616, B2 => n17615, A => n17613, ZN => 
                           n17306);
   U4754 : NAND3_X1 port map( A1 => n17305, A2 => n29152, A3 => n17421, ZN => 
                           n17613);
   U4759 : MUX2_X1 port map( A => n27425, B => n27429, S => n27424, Z => n27431
                           );
   U4774 : NAND2_X1 port map( A1 => n28491, A2 => n501, ZN => n20021);
   U4779 : OAI21_X2 port map( B1 => n20465, B2 => n21534, A => n20464, ZN => 
                           n22302);
   U4789 : OAI211_X1 port map( C1 => n20218, C2 => n20496, A => n6834, B => 
                           n20217, ZN => n2798);
   U4792 : NAND2_X1 port map( A1 => n20496, A2 => n20493, ZN => n20217);
   U4816 : XNOR2_X1 port map( A => n5809, B => n28830, ZN => n21353);
   U4841 : XNOR2_X1 port map( A => n19424, B => n19425, ZN => n28830);
   U4857 : NAND3_X1 port map( A1 => n459, A2 => n5168, A3 => n24017, ZN => 
                           n5218);
   U4865 : NAND2_X1 port map( A1 => n6423, A2 => n6424, ZN => n3459);
   U4881 : NAND2_X1 port map( A1 => n24142, A2 => n24144, ZN => n23931);
   U4902 : AND3_X2 port map( A1 => n3538, A2 => n17905, A3 => n3539, ZN => 
                           n19626);
   U4905 : NAND2_X1 port map( A1 => n1337, A2 => n4801, ZN => n10527);
   U4917 : NAND2_X1 port map( A1 => n28801, A2 => n16797, ZN => n2600);
   U4918 : NAND2_X1 port map( A1 => n17128, A2 => n17451, ZN => n28831);
   U4934 : NAND3_X2 port map( A1 => n28832, A2 => n7419, A3 => n7417, ZN => 
                           n9996);
   U4957 : NAND2_X1 port map( A1 => n7416, A2 => n714, ZN => n28832);
   U4964 : NAND3_X1 port map( A1 => n2464, A2 => n4907, A3 => n11205, ZN => 
                           n28875);
   U4984 : NAND2_X1 port map( A1 => n25052, A2 => n28833, ZN => Ciphertext(100)
                           );
   U5006 : NAND2_X1 port map( A1 => n25049, A2 => n28834, ZN => n28833);
   U5040 : NAND2_X1 port map( A1 => n9070, A2 => n8857, ZN => n9069);
   U5076 : NAND3_X1 port map( A1 => n5544, A2 => n21565, A3 => n20862, ZN => 
                           n2918);
   U5106 : NAND3_X1 port map( A1 => n18032, A2 => n18160, A3 => n18156, ZN => 
                           n28973);
   U5158 : NAND2_X1 port map( A1 => n17866, A2 => n28836, ZN => n17870);
   U5160 : NAND3_X1 port map( A1 => n511, A2 => n5690, A3 => n18216, ZN => 
                           n28836);
   U5171 : NAND2_X1 port map( A1 => n17485, A2 => n5737, ZN => n5736);
   U5172 : NAND2_X1 port map( A1 => n21198, A2 => n21509, ZN => n21535);
   U5174 : NAND2_X1 port map( A1 => n15237, A2 => n694, ZN => n28837);
   U5176 : NAND2_X1 port map( A1 => n5266, A2 => n10681, ZN => n28838);
   U5178 : NAND2_X1 port map( A1 => n5264, A2 => n10970, ZN => n28839);
   U5185 : OAI21_X1 port map( B1 => n8971, B2 => n8970, A => n28840, ZN => 
                           n9540);
   U5210 : NAND2_X1 port map( A1 => n8969, A2 => n8968, ZN => n28840);
   U5218 : NAND3_X2 port map( A1 => n15287, A2 => n5930, A3 => n28841, ZN => 
                           n16575);
   U5224 : NAND2_X1 port map( A1 => n14696, A2 => n28842, ZN => n28841);
   U5235 : NAND2_X1 port map( A1 => n7814, A2 => n2273, ZN => n8064);
   U5294 : NAND2_X1 port map( A1 => n136, A2 => n23514, ZN => n28844);
   U5307 : NOR2_X1 port map( A1 => n8540, A2 => n6901, ZN => n28845);
   U5327 : AND2_X2 port map( A1 => n28847, A2 => n6394, ZN => n22363);
   U5353 : NAND3_X1 port map( A1 => n6396, A2 => n21272, A3 => n6397, ZN => 
                           n28847);
   U5355 : NAND2_X1 port map( A1 => n830, A2 => n14273, ZN => n828);
   U5363 : NAND2_X1 port map( A1 => n827, A2 => n14361, ZN => n830);
   U5365 : NAND2_X1 port map( A1 => n7248, A2 => n8052, ZN => n1010);
   U5409 : OR2_X1 port map( A1 => n8381, A2 => n8735, ZN => n7575);
   U5460 : AND3_X2 port map( A1 => n9816, A2 => n9814, A3 => n9815, ZN => 
                           n11819);
   U5461 : AND2_X1 port map( A1 => n9438, A2 => n8995, ZN => n29221);
   U5526 : NAND2_X1 port map( A1 => n6894, A2 => n28848, ZN => n19012);
   U5529 : NAND2_X1 port map( A1 => n20145, A2 => n28849, ZN => n28848);
   U5535 : NAND2_X1 port map( A1 => n20985, A2 => n20913, ZN => n20921);
   U5536 : NAND2_X1 port map( A1 => n27480, A2 => n27492, ZN => n27475);
   U5545 : OAI21_X1 port map( B1 => n24977, B2 => n24258, A => n28815, ZN => 
                           n24981);
   U5554 : INV_X1 port map( A => n8794, ZN => n4839);
   U5580 : NAND2_X1 port map( A1 => n9037, A2 => n9034, ZN => n8794);
   U5583 : INV_X1 port map( A => n28852, ZN => n28851);
   U5602 : NAND2_X1 port map( A1 => n28853, A2 => n11261, ZN => n3326);
   U5633 : NAND2_X1 port map( A1 => n2754, A2 => n2755, ZN => n28853);
   U5634 : NAND2_X1 port map( A1 => n28855, A2 => n28854, ZN => n23133);
   U5668 : NAND2_X1 port map( A1 => n23366, A2 => n23364, ZN => n28854);
   U5675 : NAND2_X1 port map( A1 => n2921, A2 => n28604, ZN => n28855);
   U5700 : NAND2_X1 port map( A1 => n986, A2 => n988, ZN => n5445);
   U5710 : NOR2_X2 port map( A1 => n6198, A2 => n24298, ZN => n25760);
   U5718 : NAND2_X1 port map( A1 => n11274, A2 => n11034, ZN => n11035);
   U5726 : NAND2_X1 port map( A1 => n14569, A2 => n14570, ZN => n6320);
   U5742 : NAND2_X1 port map( A1 => n14967, A2 => n14964, ZN => n28856);
   U5747 : NAND2_X1 port map( A1 => n7658, A2 => n7659, ZN => n28857);
   U5763 : NAND2_X1 port map( A1 => n3325, A2 => n3326, ZN => n11887);
   U5897 : INV_X1 port map( A => n1096, ZN => n1356);
   U5914 : NAND3_X1 port map( A1 => n28950, A2 => n13309, A3 => n13697, ZN => 
                           n1096);
   U5941 : OR2_X1 port map( A1 => n14349, A2 => n14354, ZN => n6511);
   U5953 : NAND2_X1 port map( A1 => n3911, A2 => n20049, ZN => n20050);
   U5980 : OAI21_X2 port map( B1 => n9215, B2 => n9214, A => n28858, ZN => 
                           n10356);
   U5996 : NAND3_X1 port map( A1 => n22996, A2 => n23643, A3 => n23641, ZN => 
                           n22258);
   U6046 : NAND2_X1 port map( A1 => n9201, A2 => n9206, ZN => n28860);
   U6089 : INV_X1 port map( A => n9206, ZN => n28862);
   U6146 : NAND2_X1 port map( A1 => n16602, A2 => n17518, ZN => n3811);
   U6188 : NAND3_X1 port map( A1 => n5333, A2 => n6509, A3 => n6508, ZN => 
                           n21483);
   U6231 : NAND2_X1 port map( A1 => n18128, A2 => n18124, ZN => n18127);
   U6236 : OAI211_X2 port map( C1 => n12260, C2 => n12261, A => n12258, B => 
                           n28863, ZN => n12762);
   U6309 : OAI211_X1 port map( C1 => n13993, C2 => n14578, A => n15098, B => 
                           n28864, ZN => n12629);
   U6327 : NAND2_X1 port map( A1 => n14578, A2 => n15097, ZN => n28864);
   U6393 : NAND2_X1 port map( A1 => n13358, A2 => n13914, ZN => n28866);
   U6406 : NAND2_X1 port map( A1 => n24602, A2 => n24734, ZN => n5454);
   U6434 : NAND2_X1 port map( A1 => n1992, A2 => n6663, ZN => n3239);
   U6442 : NAND2_X1 port map( A1 => n4979, A2 => n17181, ZN => n16707);
   U6443 : AOI21_X1 port map( B1 => n2286, B2 => n23697, A => n28867, ZN => 
                           n6942);
   U6444 : NAND2_X1 port map( A1 => n23532, A2 => n6903, ZN => n28867);
   U6556 : NOR2_X2 port map( A1 => n13743, A2 => n4026, ZN => n15382);
   U6578 : XNOR2_X1 port map( A => n28869, B => n19210, ZN => n19213);
   U6611 : INV_X1 port map( A => n19212, ZN => n28869);
   U6683 : INV_X1 port map( A => n694, ZN => n28871);
   U6689 : NAND2_X1 port map( A1 => n28766, A2 => n694, ZN => n28872);
   U6737 : NAND2_X1 port map( A1 => n26984, A2 => n28019, ZN => n28005);
   U6773 : NAND2_X1 port map( A1 => n24228, A2 => n24532, ZN => n24895);
   U6808 : NAND2_X1 port map( A1 => n5030, A2 => n484, ZN => n5029);
   U6809 : AND2_X1 port map( A1 => n18107, A2 => n18106, ZN => n29156);
   U6849 : NAND3_X1 port map( A1 => n28874, A2 => n12299, A3 => n11767, ZN => 
                           n11366);
   U6856 : NAND2_X1 port map( A1 => n11769, A2 => n12302, ZN => n28874);
   U6864 : NAND3_X1 port map( A1 => n1657, A2 => n17258, A3 => n1574, ZN => 
                           n16670);
   U6865 : NAND2_X1 port map( A1 => n28875, A2 => n11208, ZN => n12053);
   U6895 : NAND3_X1 port map( A1 => n28627, A2 => n10806, A3 => n28876, ZN => 
                           n10543);
   U6899 : INV_X1 port map( A => n10808, ZN => n28876);
   U6919 : NAND2_X1 port map( A1 => n10726, A2 => n1879, ZN => n10727);
   U6942 : NAND2_X1 port map( A1 => n2194, A2 => n2748, ZN => n2193);
   U6944 : NAND2_X1 port map( A1 => n2649, A2 => n24390, ZN => n24691);
   U6959 : NAND3_X1 port map( A1 => n893, A2 => n14833, A3 => n15036, ZN => 
                           n14097);
   U7110 : NAND2_X1 port map( A1 => n3849, A2 => n28241, ZN => n28877);
   U7124 : NAND2_X1 port map( A1 => n11686, A2 => n28878, ZN => n11687);
   U7126 : AOI21_X1 port map( B1 => n28879, B2 => n15466, A => n15464, ZN => 
                           n15467);
   U7178 : NAND2_X1 port map( A1 => n4515, A2 => n15463, ZN => n28879);
   U7349 : NAND2_X1 port map( A1 => n11954, A2 => n4018, ZN => n4017);
   U7372 : OAI22_X1 port map( A1 => n2137, A2 => n58, B1 => n13999, B2 => n5918
                           , ZN => n6446);
   U7390 : NAND2_X1 port map( A1 => n14036, A2 => n29089, ZN => n2137);
   U7391 : NAND2_X1 port map( A1 => n20886, A2 => n21587, ZN => n21589);
   U7509 : NAND2_X1 port map( A1 => n2250, A2 => n8350, ZN => n28882);
   U7620 : OAI22_X2 port map( A1 => n17871, A2 => n18063, B1 => n18303, B2 => 
                           n18061, ZN => n19727);
   U7683 : OAI211_X2 port map( C1 => n8766, C2 => n8765, A => n9564, B => n2168
                           , ZN => n9710);
   U7695 : AOI22_X1 port map( A1 => n15074, A2 => n15073, B1 => n15076, B2 => 
                           n15075, ZN => n15080);
   U7709 : NAND2_X1 port map( A1 => n24653, A2 => n3061, ZN => n24245);
   U7722 : OR2_X2 port map( A1 => n23225, A2 => n23224, ZN => n3061);
   U7732 : NOR2_X2 port map( A1 => n26626, A2 => n5685, ZN => n27977);
   U7744 : NAND2_X1 port map( A1 => n5686, A2 => n5687, ZN => n5685);
   U7747 : INV_X1 port map( A => n15980, ZN => n539);
   U7748 : XNOR2_X1 port map( A => n15979, B => n6455, ZN => n15980);
   U7771 : NAND2_X1 port map( A1 => n13615, A2 => n3346, ZN => n15001);
   U7796 : OAI21_X1 port map( B1 => n16936, B2 => n16935, A => n17155, ZN => 
                           n28883);
   U7898 : NAND2_X1 port map( A1 => n21656, A2 => n20833, ZN => n2641);
   U7939 : NAND2_X1 port map( A1 => n28005, A2 => n28885, ZN => n26986);
   U7985 : NAND2_X1 port map( A1 => n28017, A2 => n445, ZN => n28885);
   U8008 : NOR2_X2 port map( A1 => n10967, A2 => n10968, ZN => n349);
   U8016 : NAND2_X1 port map( A1 => n11393, A2 => n28886, ZN => n13025);
   U8042 : NAND2_X1 port map( A1 => n3509, A2 => n29150, ZN => n28887);
   U8055 : NAND2_X1 port map( A1 => n28888, A2 => n4951, ZN => n22862);
   U8082 : NAND2_X1 port map( A1 => n29175, A2 => n11478, ZN => n12954);
   U8096 : OR2_X1 port map( A1 => n10913, A2 => n10735, ZN => n10607);
   U8149 : NAND3_X1 port map( A1 => n11215, A2 => n11216, A3 => n11214, ZN => 
                           n12313);
   U8193 : NAND2_X1 port map( A1 => n37, A2 => n39, ZN => n11326);
   U8198 : NAND2_X1 port map( A1 => n8177, A2 => n8173, ZN => n7290);
   U8203 : OAI21_X2 port map( B1 => n16840, B2 => n16839, A => n28889, ZN => 
                           n18190);
   U8229 : NAND2_X1 port map( A1 => n1405, A2 => n29550, ZN => n28889);
   U8239 : NAND2_X1 port map( A1 => n21547, A2 => n28891, ZN => n28890);
   U8262 : NAND2_X1 port map( A1 => n15207, A2 => n15202, ZN => n5515);
   U8269 : NAND2_X1 port map( A1 => n20346, A2 => n20347, ZN => n20348);
   U8289 : NAND2_X1 port map( A1 => n28489, A2 => n20511, ZN => n20347);
   U8350 : NAND3_X2 port map( A1 => n13634, A2 => n13635, A3 => n4689, ZN => 
                           n4688);
   U8353 : NAND3_X2 port map( A1 => n73, A2 => n20727, A3 => n3252, ZN => 
                           n22845);
   U8381 : OR2_X1 port map( A1 => n20430, A2 => n28894, ZN => n20622);
   U8404 : OR2_X1 port map( A1 => n4346, A2 => n1931, ZN => n10896);
   U8445 : INV_X1 port map( A => n12593, ZN => n5069);
   U8451 : NAND2_X1 port map( A1 => n29009, A2 => n2587, ZN => n12593);
   U8470 : NAND2_X1 port map( A1 => n28895, A2 => n5674, ZN => n5673);
   U8471 : OAI21_X1 port map( B1 => n6147, B2 => n9016, A => n5676, ZN => 
                           n28895);
   U8473 : INV_X1 port map( A => n12346, ZN => n10649);
   U8488 : NOR2_X1 port map( A1 => n21273, A2 => n6934, ZN => n21274);
   U8491 : AND2_X1 port map( A1 => n21373, A2 => n21372, ZN => n6934);
   U8497 : NAND2_X1 port map( A1 => n3776, A2 => n10722, ZN => n11486);
   U8498 : NOR2_X1 port map( A1 => n28767, A2 => n28897, ZN => n28896);
   U8501 : OAI21_X1 port map( B1 => n20359, B2 => n20238, A => n20243, ZN => 
                           n28898);
   U8529 : NAND3_X1 port map( A1 => n9039, A2 => n9243, A3 => n9248, ZN => 
                           n8694);
   U8578 : NAND2_X1 port map( A1 => n14355, A2 => n28899, ZN => n6873);
   U8587 : NAND2_X1 port map( A1 => n28902, A2 => n28900, ZN => n18084);
   U8613 : INV_X1 port map( A => n374, ZN => n28901);
   U8617 : NAND2_X1 port map( A1 => n18082, A2 => n374, ZN => n28902);
   U8626 : XNOR2_X1 port map( A => n28903, B => n3662, ZN => Ciphertext(18));
   U8628 : AOI22_X1 port map( A1 => n26961, A2 => n27410, B1 => n28607, B2 => 
                           n26962, ZN => n28903);
   U8643 : NAND2_X1 port map( A1 => n2518, A2 => n11085, ZN => n10165);
   U8648 : NAND2_X1 port map( A1 => n23929, A2 => n24588, ZN => n1283);
   U8649 : OR2_X2 port map( A1 => n28245, A2 => n14925, ZN => n16323);
   U8657 : NOR2_X2 port map( A1 => n23670, A2 => n23671, ZN => n24812);
   U8665 : NAND3_X1 port map( A1 => n13255, A2 => n13578, A3 => n13254, ZN => 
                           n6812);
   U8675 : NAND3_X2 port map( A1 => n3484, A2 => n29176, A3 => n28904, ZN => 
                           n18034);
   U8679 : NAND2_X1 port map( A1 => n28906, A2 => n28905, ZN => n28904);
   U8717 : INV_X1 port map( A => n17301, ZN => n28905);
   U8719 : INV_X1 port map( A => n17300, ZN => n28906);
   U8720 : NAND3_X1 port map( A1 => n29174, A2 => n980, A3 => n24076, ZN => 
                           n25398);
   U8732 : NAND2_X1 port map( A1 => n28909, A2 => n28907, ZN => n25243);
   U8742 : OR2_X1 port map( A1 => n27395, A2 => n28908, ZN => n28907);
   U8749 : INV_X1 port map( A => n26191, ZN => n28908);
   U8765 : NAND2_X1 port map( A1 => n27395, A2 => n27393, ZN => n28909);
   U8778 : NAND2_X1 port map( A1 => n28910, A2 => n10448, ZN => n2272);
   U8793 : NAND2_X1 port map( A1 => n6542, A2 => n10110, ZN => n28910);
   U8806 : XNOR2_X2 port map( A => n16599, B => n180, ZN => n17518);
   U8840 : NAND2_X1 port map( A1 => n9039, A2 => n28911, ZN => n8697);
   U8849 : NAND2_X1 port map( A1 => n29177, A2 => n17434, ZN => n28912);
   U8894 : XNOR2_X1 port map( A => n22079, B => n28914, ZN => n28622);
   U8928 : NAND3_X1 port map( A1 => n6586, A2 => n6585, A3 => n6584, ZN => 
                           n6741);
   U8934 : XNOR2_X1 port map( A => n10183, B => n10232, ZN => n9606);
   U8940 : NAND2_X1 port map( A1 => n28915, A2 => n20951, ZN => n20957);
   U8969 : NAND2_X1 port map( A1 => n21931, A2 => n28916, ZN => n28915);
   U8983 : OAI21_X2 port map( B1 => n11382, B2 => n11381, A => n28917, ZN => 
                           n13297);
   U9032 : NAND2_X1 port map( A1 => n24539, A2 => n24540, ZN => n24548);
   U9039 : OAI21_X1 port map( B1 => n26209, B2 => n283, A => n25665, ZN => 
                           n25632);
   U9101 : OAI211_X1 port map( C1 => n24162, C2 => n24802, A => n24503, B => 
                           n28918, ZN => n24165);
   U9169 : NAND2_X1 port map( A1 => n24162, A2 => n28919, ZN => n28918);
   U9216 : INV_X1 port map( A => n24806, ZN => n28919);
   U9218 : NAND2_X1 port map( A1 => n24681, A2 => n24391, ZN => n28262);
   U9261 : OAI211_X2 port map( C1 => n24381, C2 => n24380, A => n2905, B => 
                           n2906, ZN => n25352);
   U9265 : AOI21_X1 port map( B1 => n4826, B2 => n28920, A => n7641, ZN => 
                           n4825);
   U9279 : NAND2_X1 port map( A1 => n7985, A2 => n7642, ZN => n28920);
   U9294 : OR2_X2 port map( A1 => n1056, A2 => n8461, ZN => n9930);
   U9319 : AND2_X1 port map( A1 => n13653, A2 => n14327, ZN => n13799);
   U9324 : INV_X1 port map( A => n8767, ZN => n28921);
   U9327 : NAND2_X1 port map( A1 => n28921, A2 => n9425, ZN => n8769);
   U9329 : AND3_X2 port map( A1 => n28924, A2 => n28923, A3 => n28922, ZN => 
                           n24484);
   U9336 : NAND2_X1 port map( A1 => n6941, A2 => n23458, ZN => n28922);
   U9341 : NAND2_X1 port map( A1 => n23117, A2 => n23460, ZN => n28923);
   U9363 : INV_X1 port map( A => n11220, ZN => n28929);
   U9390 : NOR2_X1 port map( A1 => n10280, A2 => n28931, ZN => n28930);
   U9394 : AND2_X1 port map( A1 => n10269, A2 => n11220, ZN => n28931);
   U9398 : AND2_X2 port map( A1 => n1316, A2 => n1317, ZN => n12813);
   U9402 : OR2_X1 port map( A1 => n422, A2 => n16809, ZN => n29195);
   U9420 : NAND2_X1 port map( A1 => n2922, A2 => n28252, ZN => n20434);
   U9447 : NAND2_X1 port map( A1 => n17688, A2 => n1708, ZN => n853);
   U9467 : NAND2_X1 port map( A1 => n21579, A2 => n21578, ZN => n5139);
   U9557 : NAND2_X1 port map( A1 => n8049, A2 => n8131, ZN => n28933);
   U9586 : NAND2_X1 port map( A1 => n7556, A2 => n7127, ZN => n28934);
   U9592 : NAND3_X2 port map( A1 => n28935, A2 => n3885, A3 => n3884, ZN => 
                           n18215);
   U9618 : NAND2_X1 port map( A1 => n2559, A2 => n2560, ZN => n28935);
   U9629 : NAND2_X1 port map( A1 => n21392, A2 => n21632, ZN => n21634);
   U9652 : NAND3_X1 port map( A1 => n4754, A2 => n23119, A3 => n24479, ZN => 
                           n23120);
   U9682 : NAND3_X1 port map( A1 => n14281, A2 => n14082, A3 => n14081, ZN => 
                           n14088);
   U9685 : NAND3_X2 port map( A1 => n17245, A2 => n17244, A3 => n17243, ZN => 
                           n2855);
   U9687 : OAI22_X1 port map( A1 => n15337, A2 => n15338, B1 => n15339, B2 => 
                           n5777, ZN => n15340);
   U9688 : NAND2_X1 port map( A1 => n15233, A2 => n15333, ZN => n15337);
   U9731 : AND4_X2 port map( A1 => n6528, A2 => n21045, A3 => n21044, A4 => 
                           n21043, ZN => n22488);
   U9732 : NAND2_X1 port map( A1 => n1715, A2 => n1714, ZN => n1207);
   U9734 : NAND2_X1 port map( A1 => n4304, A2 => n9208, ZN => n28938);
   U9754 : NOR2_X1 port map( A1 => n24699, A2 => n28939, ZN => n711);
   U9756 : INV_X1 port map( A => n24771, ZN => n28939);
   U9793 : NAND2_X1 port map( A1 => n24768, A2 => n24697, ZN => n24771);
   U9828 : NAND3_X1 port map( A1 => n22255, A2 => n22256, A3 => n23645, ZN => 
                           n22257);
   U9851 : NAND2_X1 port map( A1 => n7640, A2 => n7980, ZN => n7647);
   U9857 : NAND2_X1 port map( A1 => n7644, A2 => n7981, ZN => n7640);
   U9878 : NAND2_X1 port map( A1 => n29005, A2 => n14338, ZN => n14339);
   U9912 : NAND2_X1 port map( A1 => n2948, A2 => n10730, ZN => n2947);
   U9943 : NAND2_X1 port map( A1 => n2929, A2 => n3033, ZN => n26462);
   U9944 : NAND3_X1 port map( A1 => n24655, A2 => n3061, A3 => n24651, ZN => 
                           n6223);
   U9947 : NAND3_X2 port map( A1 => n28940, A2 => n28941, A3 => n6213, ZN => 
                           n21728);
   U9953 : NAND3_X1 port map( A1 => n21571, A2 => n20754, A3 => n21457, ZN => 
                           n28940);
   U9954 : XNOR2_X2 port map( A => n7049, B => Key(159), ZN => n1938);
   U9984 : OAI211_X1 port map( C1 => n5234, C2 => n18391, A => n18390, B => 
                           n18389, ZN => n18392);
   U10004 : NAND2_X1 port map( A1 => n17732, A2 => n5234, ZN => n18390);
   U10008 : NAND2_X1 port map( A1 => n3844, A2 => n3846, ZN => n16192);
   U10009 : NAND2_X1 port map( A1 => n3845, A2 => n13865, ZN => n3844);
   U10061 : AOI21_X2 port map( B1 => n711, B2 => n28942, A => n24701, ZN => 
                           n25927);
   U10090 : NAND2_X1 port map( A1 => n3054, A2 => n24700, ZN => n28942);
   U10120 : NAND2_X1 port map( A1 => n20867, A2 => n21497, ZN => n28943);
   U10132 : AOI21_X1 port map( B1 => n3442, B2 => n3441, A => n28944, ZN => 
                           n11247);
   U10164 : OAI211_X1 port map( C1 => n16337, C2 => n2158, A => n2157, B => 
                           n28945, ZN => n2155);
   U10178 : NAND2_X1 port map( A1 => n16337, A2 => n538, ZN => n28945);
   U10201 : NAND2_X1 port map( A1 => n28947, A2 => n28946, ZN => n17011);
   U10213 : NAND3_X1 port map( A1 => n29088, A2 => n5891, A3 => n17428, ZN => 
                           n28946);
   U10246 : NAND2_X1 port map( A1 => n17006, A2 => n28792, ZN => n28947);
   U10247 : NOR2_X1 port map( A1 => n17942, A2 => n17762, ZN => n1442);
   U10294 : NAND2_X1 port map( A1 => n23518, A2 => n23519, ZN => n23520);
   U10331 : NAND2_X1 port map( A1 => n26801, A2 => n28823, ZN => n28948);
   U10342 : NAND3_X1 port map( A1 => n10408, A2 => n2891, A3 => n2892, ZN => 
                           n29273);
   U10407 : OR2_X1 port map( A1 => n23360, A2 => n23676, ZN => n2888);
   U10418 : NAND2_X1 port map( A1 => n2909, A2 => n21672, ZN => n3903);
   U10474 : XNOR2_X1 port map( A => n26073, B => n2350, ZN => n25367);
   U10489 : NOR2_X1 port map( A1 => n7534, A2 => n8014, ZN => n3031);
   U10490 : NAND2_X1 port map( A1 => n8013, A2 => n7743, ZN => n7534);
   U10518 : INV_X1 port map( A => n27101, ZN => n3542);
   U10519 : AND2_X1 port map( A1 => n28949, A2 => n27101, ZN => n3236);
   U10521 : NOR2_X2 port map( A1 => n26854, A2 => n27839, ZN => n27101);
   U10533 : INV_X1 port map( A => n27100, ZN => n28949);
   U10541 : NAND2_X1 port map( A1 => n14295, A2 => n13306, ZN => n13309);
   U10542 : OAI211_X1 port map( C1 => n23431, C2 => n408, A => n23430, B => 
                           n28951, ZN => n1073);
   U10552 : NAND2_X1 port map( A1 => n4178, A2 => n23431, ZN => n28951);
   U10560 : NAND3_X1 port map( A1 => n13618, A2 => n13617, A3 => n13616, ZN => 
                           n28953);
   U10568 : NAND2_X1 port map( A1 => n10990, A2 => n10995, ZN => n10693);
   U10591 : NAND2_X1 port map( A1 => n24634, A2 => n24635, ZN => n24243);
   U10637 : NOR2_X1 port map( A1 => n23792, A2 => n23790, ZN => n28954);
   U10646 : INV_X1 port map( A => n23495, ZN => n28955);
   U10662 : NAND2_X1 port map( A1 => n1121, A2 => n17027, ZN => n1120);
   U10670 : NAND2_X1 port map( A1 => n5219, A2 => n884, ZN => n24612);
   U10677 : NAND2_X1 port map( A1 => n17930, A2 => n1863, ZN => n19508);
   U10685 : OR3_X1 port map( A1 => n1910, A2 => n8077, A3 => n8058, ZN => n7807
                           );
   U10700 : XNOR2_X1 port map( A => n28956, B => n22619, ZN => n6017);
   U10702 : NAND3_X1 port map( A1 => n2665, A2 => n6015, A3 => n2667, ZN => 
                           n28956);
   U10703 : OAI211_X2 port map( C1 => n23299, C2 => n23300, A => n5712, B => 
                           n5713, ZN => n24404);
   U10732 : NOR2_X1 port map( A1 => n5181, A2 => n20149, ZN => n20741);
   U10768 : NAND3_X1 port map( A1 => n21561, A2 => n21465, A3 => n21464, ZN => 
                           n28958);
   U10797 : INV_X1 port map( A => n10345, ZN => n9612);
   U10800 : NAND2_X1 port map( A1 => n203, A2 => n6688, ZN => n10345);
   U10876 : NAND2_X1 port map( A1 => n28960, A2 => n16906, ZN => n1721);
   U10882 : NAND2_X1 port map( A1 => n17228, A2 => n1723, ZN => n28960);
   U10909 : OAI211_X1 port map( C1 => n11907, C2 => n12359, A => n919, B => 
                           n12363, ZN => n28962);
   U10954 : NAND3_X1 port map( A1 => n28963, A2 => n23640, A3 => n22996, ZN => 
                           n2622);
   U10966 : OAI211_X1 port map( C1 => n11262, C2 => n29122, A => n11265, B => 
                           n6631, ZN => n12293);
   U10967 : XNOR2_X1 port map( A => n19254, B => n28964, ZN => n4307);
   U10979 : XNOR2_X1 port map( A => n19383, B => n28965, ZN => n28964);
   U10982 : INV_X1 port map( A => n18737, ZN => n28965);
   U11027 : NOR2_X1 port map( A1 => n28966, A2 => n29026, ZN => n23965);
   U11042 : INV_X1 port map( A => n24583, ZN => n28966);
   U11043 : OAI21_X2 port map( B1 => n21978, B2 => n23607, A => n21977, ZN => 
                           n24583);
   U11054 : OAI22_X1 port map( A1 => n27266, A2 => n27596, B1 => n26346, B2 => 
                           n28967, ZN => n27269);
   U11084 : NAND2_X1 port map( A1 => n26372, A2 => n28970, ZN => n28969);
   U11107 : INV_X1 port map( A => n26266, ZN => n28970);
   U11121 : INV_X1 port map( A => n463, ZN => n28971);
   U11161 : NAND3_X1 port map( A1 => n28971, A2 => n24775, A3 => n24779, ZN => 
                           n3836);
   U11204 : NAND2_X1 port map( A1 => n3564, A2 => n4778, ZN => n15184);
   U11214 : NAND3_X1 port map( A1 => n3432, A2 => n3502, A3 => n23734, ZN => 
                           n2481);
   U11232 : AOI22_X2 port map( A1 => n17521, A2 => n17520, B1 => n17519, B2 => 
                           n796, ZN => n18227);
   U11253 : XNOR2_X2 port map( A => n2257, B => n19690, ZN => n20440);
   U11262 : OAI21_X2 port map( B1 => n4586, B2 => n13464, A => n28972, ZN => 
                           n13789);
   U11268 : NAND2_X1 port map( A1 => n14148, A2 => n14376, ZN => n28972);
   U11286 : OAI21_X1 port map( B1 => n4854, B2 => n18033, A => n28973, ZN => 
                           n17827);
   U11300 : NAND2_X1 port map( A1 => n4959, A2 => n28974, ZN => n20861);
   U11376 : NAND3_X1 port map( A1 => n20858, A2 => n21157, A3 => n21156, ZN => 
                           n28974);
   U11454 : NAND3_X1 port map( A1 => n27664, A2 => n28347, A3 => n27661, ZN => 
                           n28373);
   U11462 : OAI21_X1 port map( B1 => n20572, B2 => n20571, A => n20570, ZN => 
                           n20715);
   U11474 : NAND3_X1 port map( A1 => n29557, A2 => n28975, A3 => n27225, ZN => 
                           n4526);
   U11477 : INV_X1 port map( A => n4528, ZN => n28975);
   U11516 : NAND2_X1 port map( A1 => n11168, A2 => n10820, ZN => n4107);
   U11517 : XNOR2_X1 port map( A => n28977, B => n25322, ZN => n24608);
   U11560 : NAND2_X1 port map( A1 => n947, A2 => n946, ZN => n28977);
   U11561 : OR2_X1 port map( A1 => n21092, A2 => n18919, ZN => n19870);
   U11579 : NAND3_X1 port map( A1 => n14, A2 => n21158, A3 => n21157, ZN => n13
                           );
   U11583 : NAND3_X1 port map( A1 => n29238, A2 => n2330, A3 => n28819, ZN => 
                           n28978);
   U11601 : NOR2_X2 port map( A1 => n18176, A2 => n28981, ZN => n18880);
   U11634 : AOI21_X1 port map( B1 => n7650, B2 => n7651, A => n7649, ZN => 
                           n7654);
   U11656 : NAND2_X1 port map( A1 => n437, A2 => n29082, ZN => n7650);
   U11767 : NAND3_X1 port map( A1 => n8299, A2 => n8298, A3 => n8297, ZN => 
                           n2405);
   U11783 : NAND2_X1 port map( A1 => n1018, A2 => n1017, ZN => n4005);
   U11820 : NAND2_X1 port map( A1 => n14254, A2 => n29312, ZN => n4376);
   U11876 : NAND3_X1 port map( A1 => n2450, A2 => n17358, A3 => n2449, ZN => 
                           n1752);
   U11963 : NAND3_X1 port map( A1 => n23546, A2 => n4773, A3 => n4772, ZN => 
                           n28983);
   U11966 : NAND2_X1 port map( A1 => n28985, A2 => n28984, ZN => n14610);
   U12008 : NAND2_X1 port map( A1 => n14306, A2 => n14429, ZN => n28984);
   U12037 : NAND2_X1 port map( A1 => n28987, A2 => n28986, ZN => n28985);
   U12053 : NAND2_X1 port map( A1 => n14305, A2 => n4837, ZN => n28987);
   U12060 : NAND2_X1 port map( A1 => n9437, A2 => n28988, ZN => n10045);
   U12111 : NAND2_X1 port map( A1 => n28990, A2 => n28989, ZN => n28988);
   U12113 : NAND2_X1 port map( A1 => n9435, A2 => n9434, ZN => n28990);
   U12121 : NAND2_X1 port map( A1 => n28185, A2 => n28991, ZN => n21193);
   U12123 : NAND2_X1 port map( A1 => n21356, A2 => n28126, ZN => n28992);
   U12151 : XNOR2_X1 port map( A => n29519, B => n3462, ZN => n22412);
   U12201 : NAND3_X1 port map( A1 => n28994, A2 => n3629, A3 => n28993, ZN => 
                           n18312);
   U12213 : NAND2_X1 port map( A1 => n5587, A2 => n29373, ZN => n28994);
   U12220 : NAND2_X1 port map( A1 => n28198, A2 => n28995, ZN => n4181);
   U12221 : NOR2_X1 port map( A1 => n14845, A2 => n28996, ZN => n28995);
   U12227 : INV_X1 port map( A => n15285, ZN => n28996);
   U12231 : OAI21_X1 port map( B1 => n7709, B2 => n7737, A => n28998, ZN => 
                           n7713);
   U12309 : NAND2_X1 port map( A1 => n16859, A2 => n28999, ZN => n17802);
   U12319 : NAND2_X1 port map( A1 => n569, A2 => n12305, ZN => n1238);
   U12349 : MUX2_X1 port map( A => n9095, B => n8665, S => n8490, Z => n8668);
   U12366 : AOI21_X1 port map( B1 => n10920, B2 => n10718, A => n29001, ZN => 
                           n10050);
   U12390 : NAND2_X1 port map( A1 => n10031, A2 => n3862, ZN => n29001);
   U12426 : NAND2_X1 port map( A1 => n24248, A2 => n24155, ZN => n24246);
   U12436 : NAND2_X1 port map( A1 => n24524, A2 => n3061, ZN => n29003);
   U12439 : NAND3_X1 port map( A1 => n29004, A2 => n23921, A3 => n4783, ZN => 
                           n24858);
   U12441 : NAND2_X1 port map( A1 => n3295, A2 => n24582, ZN => n29004);
   U12465 : NAND3_X1 port map( A1 => n5190, A2 => n5189, A3 => n15311, ZN => 
                           n29005);
   U12471 : OAI211_X2 port map( C1 => n21381, C2 => n21380, A => n4265, B => 
                           n29006, ZN => n22625);
   U12474 : NAND2_X1 port map( A1 => n21380, A2 => n21253, ZN => n29006);
   U12484 : NAND2_X1 port map( A1 => n15939, A2 => n18061, ZN => n29007);
   U12504 : NAND2_X1 port map( A1 => n29008, A2 => n16874, ZN => n4291);
   U12510 : NAND2_X1 port map( A1 => n1262, A2 => n29512, ZN => n21726);
   U12512 : AND2_X2 port map( A1 => n2396, A2 => n3619, ZN => n22387);
   U12514 : AOI22_X1 port map( A1 => n12429, A2 => n12428, B1 => n10586, B2 => 
                           n10587, ZN => n29009);
   U12524 : NAND2_X1 port map( A1 => n1886, A2 => n15084, ZN => n29010);
   U12546 : NAND2_X1 port map( A1 => n15693, A2 => n15692, ZN => n29012);
   U12599 : NAND2_X1 port map( A1 => n21019, A2 => n22023, ZN => n22025);
   U12618 : OAI21_X1 port map( B1 => n24055, B2 => n24054, A => n29013, ZN => 
                           n24056);
   U12665 : OAI21_X1 port map( B1 => n29015, B2 => n29545, A => n29014, ZN => 
                           n24026);
   U12705 : NAND2_X1 port map( A1 => n24022, A2 => n462, ZN => n29014);
   U12762 : BUF_X1 port map( A => n26459, Z => n28476);
   U12793 : AOI22_X2 port map( A1 => n23191, A2 => n23757, B1 => n5741, B2 => 
                           n23190, ZN => n24635);
   U12866 : XNOR2_X1 port map( A => n19326, B => n19325, ZN => n20625);
   U12902 : XNOR2_X1 port map( A => n25841, B => n25842, ZN => n27120);
   U12921 : INV_X1 port map( A => n27092, ZN => n27920);
   U12938 : OAI211_X1 port map( C1 => n28550, C2 => n24747, A => n24267, B => 
                           n24266, ZN => n29017);
   U12949 : NOR2_X2 port map( A1 => n20657, A2 => n20656, ZN => n28550);
   U12960 : BUF_X1 port map( A => n23432, Z => n29018);
   U12982 : XNOR2_X1 port map( A => n3983, B => n22660, ZN => n23432);
   U12998 : AND2_X1 port map( A1 => n21415, A2 => n29019, ZN => n21050);
   U13011 : NAND2_X1 port map( A1 => n21413, A2 => n20663, ZN => n29019);
   U13013 : MUX2_X1 port map( A => n23914, B => n23913, S => n24667, Z => 
                           n23915);
   U13046 : XNOR2_X1 port map( A => n22530, B => n22529, ZN => n23297);
   U13069 : AND3_X1 port map( A1 => n3177, A2 => n26618, A3 => n26619, ZN => 
                           n29021);
   U13086 : NAND3_X1 port map( A1 => n3177, A2 => n26618, A3 => n26619, ZN => 
                           n27979);
   U13125 : OR2_X1 port map( A1 => n29104, A2 => n20041, ZN => n20089);
   U13232 : NAND2_X1 port map( A1 => n6492, A2 => n6026, ZN => n29022);
   U13233 : OR2_X1 port map( A1 => n24496, A2 => n5004, ZN => n24207);
   U13237 : OAI22_X1 port map( A1 => n6857, A2 => n5221, B1 => n27054, B2 => 
                           n1971, ZN => n28025);
   U13252 : INV_X1 port map( A => n5234, ZN => n29023);
   U13288 : INV_X1 port map( A => n5234, ZN => n29024);
   U13296 : BUF_X1 port map( A => n26746, Z => n28563);
   U13317 : XNOR2_X2 port map( A => n26027, B => n26026, ZN => n26865);
   U13322 : OAI21_X1 port map( B1 => n22129, B2 => n28474, A => n22128, ZN => 
                           n29025);
   U13395 : OR2_X1 port map( A1 => n26308, A2 => n26307, ZN => n29027);
   U13396 : OAI21_X1 port map( B1 => n22129, B2 => n28474, A => n22128, ZN => 
                           n24577);
   U13409 : XOR2_X1 port map( A => n24276, B => n24275, Z => n29028);
   U13491 : OR2_X1 port map( A1 => n29075, A2 => n29500, ZN => n27066);
   U13507 : AND2_X1 port map( A1 => n5114, A2 => n5112, ZN => n29029);
   U13516 : OR3_X1 port map( A1 => n27074, A2 => n26992, A3 => n27076, ZN => 
                           n29030);
   U13538 : AND2_X1 port map( A1 => n3254, A2 => n25556, ZN => n29031);
   U13543 : MUX2_X1 port map( A => n25462, B => n25461, S => n5760, Z => n25472
                           );
   U13545 : AND3_X1 port map( A1 => n26669, A2 => n26531, A3 => n27417, ZN => 
                           n26535);
   U13546 : MUX2_X1 port map( A => n29560, B => n28548, S => n26210, Z => 
                           n26719);
   U13577 : AND2_X1 port map( A1 => n25600, A2 => n25599, ZN => n29032);
   U13582 : AND2_X1 port map( A1 => n25600, A2 => n25599, ZN => n28038);
   U13583 : BUF_X1 port map( A => n26028, Z => n28534);
   U13599 : OAI211_X1 port map( C1 => n24894, C2 => n23984, A => n29269, B => 
                           n29268, ZN => n26028);
   U13678 : OAI21_X2 port map( B1 => n26219, B2 => n26716, A => n26218, ZN => 
                           n28063);
   U13708 : AOI21_X2 port map( B1 => n26269, B2 => n26775, A => n26268, ZN => 
                           n27594);
   U13709 : BUF_X1 port map( A => n27052, Z => n28446);
   U13712 : NAND2_X1 port map( A1 => n23813, A2 => n1239, ZN => n29033);
   U13740 : OR2_X1 port map( A1 => n17257, A2 => n17256, ZN => n29034);
   U13748 : AND2_X1 port map( A1 => n17972, A2 => n17973, ZN => n29035);
   U13753 : NOR2_X1 port map( A1 => n18034, A2 => n18033, ZN => n18164);
   U13756 : OR2_X1 port map( A1 => n17743, A2 => n18034, ZN => n29289);
   U13764 : XOR2_X1 port map( A => n21979, B => n22880, Z => n21986);
   U13766 : OAI211_X2 port map( C1 => n20846, C2 => n20841, A => n20845, B => 
                           n3555, ZN => n22703);
   U13781 : OAI211_X1 port map( C1 => n220, C2 => n24464, A => n24462, B => 
                           n24463, ZN => n29053);
   U13796 : OAI211_X1 port map( C1 => n220, C2 => n24464, A => n24462, B => 
                           n24463, ZN => n25889);
   U13810 : XNOR2_X1 port map( A => n12767, B => n12766, ZN => n29036);
   U13876 : XNOR2_X1 port map( A => n12767, B => n12766, ZN => n29037);
   U13881 : OAI211_X1 port map( C1 => n18240, C2 => n17290, A => n17289, B => 
                           n17288, ZN => n29038);
   U13882 : OAI211_X1 port map( C1 => n18240, C2 => n17290, A => n17289, B => 
                           n17288, ZN => n18935);
   U13923 : AOI22_X1 port map( A1 => n24407, A2 => n3797, B1 => n24086, B2 => 
                           n24085, ZN => n25913);
   U13965 : XNOR2_X1 port map( A => n19039, B => n19381, ZN => n6569);
   U13976 : INV_X1 port map( A => n500, ZN => n29040);
   U14001 : XNOR2_X1 port map( A => n18637, B => n18636, ZN => n29041);
   U14040 : XOR2_X1 port map( A => n22907, B => n22906, Z => n29042);
   U14063 : OR2_X1 port map( A1 => n20862, A2 => n29236, ZN => n4543);
   U14090 : XNOR2_X1 port map( A => n21986, B => n21985, ZN => n23735);
   U14100 : OAI211_X1 port map( C1 => n23035, C2 => n23034, A => n4935, B => 
                           n4934, ZN => n24704);
   U14111 : BUF_X1 port map( A => n26466, Z => n280);
   U14113 : NAND2_X1 port map( A1 => n2484, A2 => n16832, ZN => n29044);
   U14120 : NAND2_X1 port map( A1 => n2484, A2 => n16832, ZN => n19561);
   U14124 : XOR2_X1 port map( A => n18991, B => n18992, Z => n18997);
   U14125 : XOR2_X1 port map( A => n19245, B => n19669, Z => n17597);
   U14135 : XNOR2_X1 port map( A => n15598, B => n15599, ZN => n29045);
   U14151 : INV_X1 port map( A => n22053, ZN => n22731);
   U14181 : NOR2_X2 port map( A1 => n1008, A2 => n26324, ZN => n27795);
   U14262 : NOR2_X1 port map( A1 => n24774, A2 => n24773, ZN => n29047);
   U14285 : AND2_X1 port map( A1 => n446, A2 => n27377, ZN => n29219);
   U14361 : XNOR2_X1 port map( A => n26064, B => n26063, ZN => n29048);
   U14391 : NOR2_X1 port map( A1 => n27902, A2 => n26848, ZN => n26852);
   U14417 : BUF_X1 port map( A => n26579, Z => n28477);
   U14496 : AND2_X1 port map( A1 => n26926, A2 => n26579, ZN => n26929);
   U14502 : XOR2_X1 port map( A => n10368, B => n9703, Z => n9708);
   U14503 : AND2_X1 port map( A1 => n24095, A2 => n4532, ZN => n29051);
   U14522 : AND2_X1 port map( A1 => n4532, A2 => n24095, ZN => n23874);
   U14544 : AND2_X1 port map( A1 => n28669, A2 => n5422, ZN => n29052);
   U14581 : AND2_X1 port map( A1 => n28669, A2 => n5422, ZN => n27352);
   U14721 : XNOR2_X1 port map( A => n24787, B => n24786, ZN => n29054);
   U14741 : OR2_X1 port map( A1 => n26200, A2 => n26235, ZN => n29055);
   U14788 : BUF_X1 port map( A => n29052, Z => n27351);
   U14810 : AND4_X1 port map( A1 => n679, A2 => n16893, A3 => n16892, A4 => 
                           n16894, ZN => n29057);
   U14862 : OR2_X1 port map( A1 => n17113, A2 => n29539, ZN => n3099);
   U14870 : XNOR2_X1 port map( A => n28311, B => n1987, ZN => n29059);
   U14881 : XNOR2_X1 port map( A => n28311, B => n1987, ZN => n14008);
   U14935 : XNOR2_X1 port map( A => n26037, B => n26036, ZN => n29060);
   U15010 : XNOR2_X1 port map( A => n22565, B => n22564, ZN => n22566);
   U15060 : AOI22_X1 port map( A1 => n26611, A2 => n28394, B1 => n295, B2 => 
                           n26610, ZN => n5651);
   U15074 : XNOR2_X1 port map( A => n25483, B => n25482, ZN => n29062);
   U15084 : OR2_X1 port map( A1 => n26626, A2 => n5685, ZN => n29063);
   U15100 : XNOR2_X1 port map( A => n25483, B => n25482, ZN => n27050);
   U15101 : OAI21_X1 port map( B1 => n11359, B2 => n12401, A => n11358, ZN => 
                           n29064);
   U15114 : INV_X1 port map( A => n2656, ZN => n29065);
   U15150 : OAI21_X1 port map( B1 => n11359, B2 => n12401, A => n11358, ZN => 
                           n12746);
   U15157 : AOI21_X1 port map( B1 => n16968, B2 => n6130, A => n6126, ZN => 
                           n17889);
   U15167 : XNOR2_X1 port map( A => n18866, B => n18865, ZN => n29066);
   U15169 : OAI21_X1 port map( B1 => n24414, B2 => n4136, A => n2261, ZN => 
                           n29067);
   U15174 : XNOR2_X1 port map( A => n18866, B => n18865, ZN => n20161);
   U15175 : OAI21_X1 port map( B1 => n24414, B2 => n4136, A => n2261, ZN => 
                           n25550);
   U15191 : NOR2_X1 port map( A1 => n25797, A2 => n25800, ZN => n29069);
   U15216 : NOR2_X1 port map( A1 => n25797, A2 => n25800, ZN => n25729);
   U15227 : XNOR2_X1 port map( A => n25163, B => n25164, ZN => n29071);
   U15380 : XNOR2_X1 port map( A => n25163, B => n25164, ZN => n26952);
   U15381 : BUF_X1 port map( A => n17296, Z => n29072);
   U15447 : AOI21_X1 port map( B1 => n24034, B2 => n24033, A => n24032, ZN => 
                           n29073);
   U15458 : AOI21_X1 port map( B1 => n24034, B2 => n24033, A => n24032, ZN => 
                           n25886);
   U15520 : OAI21_X1 port map( B1 => n3671, B2 => n24513, A => n3618, ZN => 
                           n29193);
   U15553 : XNOR2_X1 port map( A => n22237, B => n22236, ZN => n29074);
   U15554 : XNOR2_X1 port map( A => n22237, B => n22236, ZN => n23642);
   U15693 : XOR2_X1 port map( A => n25700, B => n25699, Z => n29075);
   U15844 : XOR2_X1 port map( A => n25700, B => n25699, Z => n29076);
   U15907 : CLKBUF_X1 port map( A => n25344, Z => n26737);
   U15930 : XNOR2_X1 port map( A => n9346, B => n9347, ZN => n29077);
   U15938 : XNOR2_X1 port map( A => n9346, B => n9347, ZN => n29078);
   U16008 : BUF_X1 port map( A => n22783, Z => n29079);
   U16039 : XNOR2_X1 port map( A => n7058, B => Key(167), ZN => n29081);
   U16071 : XNOR2_X1 port map( A => n7058, B => Key(167), ZN => n29082);
   U16216 : XNOR2_X1 port map( A => n1257, B => n1258, ZN => n29083);
   U16217 : XNOR2_X1 port map( A => n7058, B => Key(167), ZN => n7876);
   U16250 : XNOR2_X1 port map( A => n1257, B => n1258, ZN => n16811);
   U16251 : NAND3_X1 port map( A1 => n15034, A2 => n15035, A3 => n15033, ZN => 
                           n29084);
   U16340 : NAND3_X1 port map( A1 => n15034, A2 => n15035, A3 => n15033, ZN => 
                           n15966);
   U16360 : NAND2_X1 port map( A1 => n26395, A2 => n56, ZN => n29085);
   U16375 : NAND2_X1 port map( A1 => n26395, A2 => n56, ZN => n27572);
   U16437 : XOR2_X1 port map( A => n16049, B => n16048, Z => n29086);
   U16444 : XOR2_X1 port map( A => n22053, B => n22052, Z => n29087);
   U16445 : INV_X1 port map( A => n6013, ZN => n29088);
   U16688 : XOR2_X1 port map( A => n13477, B => n13476, Z => n29089);
   U16689 : NAND3_X2 port map( A1 => n2051, A2 => n26233, A3 => n26232, ZN => 
                           n28067);
   U16785 : NAND2_X1 port map( A1 => n27164, A2 => n5993, ZN => n29090);
   U16824 : NAND2_X1 port map( A1 => n27164, A2 => n5993, ZN => n29091);
   U16832 : NAND2_X1 port map( A1 => n27164, A2 => n5993, ZN => n27673);
   U16883 : OR2_X1 port map( A1 => n26635, A2 => n26634, ZN => n29092);
   U16901 : NOR2_X2 port map( A1 => n26578, A2 => n26577, ZN => n29093);
   U16957 : NOR2_X1 port map( A1 => n26578, A2 => n26577, ZN => n27494);
   U16960 : MUX2_X1 port map( A => n21027, B => n21026, S => n23016, Z => 
                           n21060);
   U17016 : NOR2_X1 port map( A1 => n146, A2 => n23904, ZN => n29094);
   U17032 : NOR2_X1 port map( A1 => n146, A2 => n23904, ZN => n25246);
   U17036 : OAI21_X1 port map( B1 => n28617, B2 => n8262, A => n8261, ZN => 
                           n29096);
   U17070 : OAI21_X1 port map( B1 => n28617, B2 => n8262, A => n8261, ZN => 
                           n8954);
   U17072 : XNOR2_X1 port map( A => n11546, B => n11545, ZN => n14171);
   U17114 : XNOR2_X1 port map( A => n15883, B => n15882, ZN => n29098);
   U17127 : XNOR2_X1 port map( A => n25439, B => n25438, ZN => n29099);
   U17150 : XNOR2_X1 port map( A => n25439, B => n25438, ZN => n29100);
   U17222 : BUF_X1 port map( A => n21696, Z => n29101);
   U17265 : XNOR2_X1 port map( A => n22622, B => n22623, ZN => n29102);
   U17270 : XNOR2_X1 port map( A => n22622, B => n22623, ZN => n23806);
   U17318 : NOR2_X1 port map( A1 => n24733, A2 => n3725, ZN => n29103);
   U17376 : NOR2_X1 port map( A1 => n24733, A2 => n3725, ZN => n25531);
   U17383 : XNOR2_X1 port map( A => n18747, B => n18748, ZN => n29104);
   U17384 : XNOR2_X1 port map( A => n13182, B => n13183, ZN => n29107);
   U17393 : XNOR2_X1 port map( A => n7008, B => Key(71), ZN => n7011);
   U17406 : XNOR2_X1 port map( A => n13182, B => n13183, ZN => n13920);
   U17457 : XNOR2_X1 port map( A => n24937, B => n25560, ZN => n27703);
   U17472 : XNOR2_X1 port map( A => n21456, B => n21455, ZN => n23427);
   U17479 : NAND2_X1 port map( A1 => n20035, A2 => n29186, ZN => n22643);
   U17498 : NAND3_X1 port map( A1 => n5293, A2 => n5292, A3 => n22499, ZN => 
                           n24613);
   U17598 : BUF_X1 port map( A => n8237, Z => n29110);
   U17604 : XNOR2_X1 port map( A => n6969, B => Key(104), ZN => n8237);
   U17606 : BUF_X1 port map( A => n26089, Z => n29111);
   U17618 : OAI22_X1 port map( A1 => n23951, A2 => n23950, B1 => n5004, B2 => 
                           n24810, ZN => n26089);
   U17715 : XNOR2_X1 port map( A => n22361, B => n22360, ZN => n960);
   U17716 : XNOR2_X1 port map( A => n7085, B => Key(4), ZN => n29112);
   U17802 : XNOR2_X1 port map( A => n7085, B => Key(4), ZN => n7891);
   U17959 : BUF_X1 port map( A => n23733, Z => n1862);
   U18090 : BUF_X1 port map( A => n23562, Z => n29115);
   U18120 : XNOR2_X1 port map( A => n18742, B => n18741, ZN => n20090);
   U18139 : BUF_X2 port map( A => n11288, Z => n29116);
   U18354 : XNOR2_X1 port map( A => n10326, B => n10325, ZN => n11288);
   U18470 : NOR2_X1 port map( A1 => n26293, A2 => n26294, ZN => n29117);
   U18476 : NOR2_X1 port map( A1 => n26293, A2 => n26294, ZN => n29118);
   U18735 : NOR2_X1 port map( A1 => n26293, A2 => n26294, ZN => n27768);
   U18820 : XNOR2_X1 port map( A => Key(44), B => Plaintext(44), ZN => n29119);
   U18974 : OR2_X1 port map( A1 => n23782, A2 => n23781, ZN => n29120);
   U18981 : XNOR2_X1 port map( A => Key(44), B => Plaintext(44), ZN => n8136);
   U18999 : MUX2_X2 port map( A => n21102, B => n21101, S => n28916, Z => 
                           n22768);
   U19073 : INV_X1 port map( A => n28091, ZN => n29121);
   U19094 : AOI22_X1 port map( A1 => n26732, A2 => n1623, B1 => n26730, B2 => 
                           n29579, ZN => n28091);
   U19113 : INV_X1 port map( A => n20333, ZN => n28186);
   U19118 : XNOR2_X1 port map( A => n1141, B => n9628, ZN => n29122);
   U19127 : XNOR2_X1 port map( A => n1141, B => n9628, ZN => n11260);
   U19235 : XOR2_X1 port map( A => n18863, B => n18395, Z => n29124);
   U19317 : BUF_X1 port map( A => n19562, Z => n29125);
   U19338 : XOR2_X1 port map( A => n22385, B => n22384, Z => n29126);
   U19351 : OAI211_X1 port map( C1 => n17224, C2 => n16908, A => n16917, B => 
                           n16835, ZN => n19562);
   U19389 : XOR2_X1 port map( A => n16209, B => n16210, Z => n29127);
   U19398 : AOI22_X1 port map( A1 => n22989, A2 => n22990, B1 => n23624, B2 => 
                           n22988, ZN => n29128);
   U19440 : AOI22_X1 port map( A1 => n22989, A2 => n22990, B1 => n23624, B2 => 
                           n22988, ZN => n24436);
   U19475 : NAND3_X1 port map( A1 => n28362, A2 => n3359, A3 => n28361, ZN => 
                           n29129);
   U19517 : NAND3_X1 port map( A1 => n28362, A2 => n3359, A3 => n28361, ZN => 
                           n26073);
   U19543 : XNOR2_X1 port map( A => Key(68), B => Plaintext(68), ZN => n29130);
   U19548 : XNOR2_X1 port map( A => Key(68), B => Plaintext(68), ZN => n8023);
   U19687 : AND2_X1 port map( A1 => n10884, A2 => n11282, ZN => n29212);
   U19695 : XOR2_X1 port map( A => n22335, B => n22336, Z => n29131);
   U19732 : AOI22_X1 port map( A1 => n1362, A2 => n17314, B1 => n1361, B2 => 
                           n29550, ZN => n17826);
   U19733 : XNOR2_X1 port map( A => n24866, B => n24865, ZN => n29132);
   U19734 : XNOR2_X1 port map( A => n12412, B => n12411, ZN => n29133);
   U19835 : XNOR2_X1 port map( A => n18916, B => n18917, ZN => n21092);
   U19840 : NOR2_X2 port map( A1 => n28103, A2 => n5037, ZN => n28089);
   U19856 : XOR2_X1 port map( A => n10149, B => n9619, Z => n9906);
   U19911 : XNOR2_X1 port map( A => n21999, B => n22812, ZN => n29136);
   U19912 : XNOR2_X1 port map( A => Key(119), B => Plaintext(119), ZN => n9113)
                           ;
   U20079 : OAI21_X1 port map( B1 => n11143, B2 => n11142, A => n1452, ZN => 
                           n29137);
   U20140 : BUF_X1 port map( A => n17565, Z => n29138);
   U20284 : XNOR2_X1 port map( A => n2790, B => n16267, ZN => n17565);
   U20316 : OR2_X1 port map( A1 => n29330, A2 => n26280, ZN => n26801);
   U20341 : OAI21_X1 port map( B1 => n11644, B2 => n11643, A => n11642, ZN => 
                           n29140);
   U20444 : NOR2_X1 port map( A1 => n11636, A2 => n11633, ZN => n11673);
   U20544 : OAI21_X1 port map( B1 => n11644, B2 => n11643, A => n11642, ZN => 
                           n13012);
   U20743 : CLKBUF_X3 port map( A => n27378, Z => n295);
   U20822 : XNOR2_X1 port map( A => n15827, B => n15826, ZN => n29142);
   U20831 : INV_X1 port map( A => n19838, ZN => n29143);
   U20839 : XNOR2_X1 port map( A => n15827, B => n15826, ZN => n17557);
   U20843 : XNOR2_X1 port map( A => n17813, B => n17812, ZN => n29144);
   U20879 : XNOR2_X1 port map( A => n18563, B => n18564, ZN => n29145);
   U20950 : XNOR2_X1 port map( A => n18564, B => n18563, ZN => n29146);
   U20959 : XNOR2_X1 port map( A => n9599, B => n9600, ZN => n29149);
   U20984 : AND2_X1 port map( A1 => n11126, A2 => n10114, ZN => n11403);
   U21031 : AND2_X1 port map( A1 => n29618, A2 => n22452, ZN => n29169);
   U21051 : OAI21_X1 port map( B1 => n15298, B2 => n15297, A => n15296, ZN => 
                           n29151);
   U21079 : XNOR2_X1 port map( A => n15330, B => n15329, ZN => n29152);
   U21099 : OAI21_X1 port map( B1 => n15298, B2 => n15297, A => n15296, ZN => 
                           n16580);
   U21116 : OAI211_X1 port map( C1 => n13888, C2 => n14313, A => n13887, B => 
                           n3602, ZN => n29153);
   U21117 : AOI21_X1 port map( B1 => n3634, B2 => n24459, A => n24458, ZN => 
                           n29154);
   U21174 : AOI21_X1 port map( B1 => n3634, B2 => n24459, A => n24458, ZN => 
                           n29155);
   U21177 : OAI211_X1 port map( C1 => n13888, C2 => n14313, A => n13887, B => 
                           n3602, ZN => n15160);
   U21179 : AOI21_X1 port map( B1 => n3634, B2 => n24459, A => n24458, ZN => 
                           n25759);
   U21180 : NAND2_X1 port map( A1 => n18456, A2 => n29156, ZN => n3865);
   U21242 : OR3_X1 port map( A1 => n27492, A2 => n27494, A3 => n27497, ZN => 
                           n27500);
   U21251 : XOR2_X1 port map( A => n22115, B => n22114, Z => n29157);
   U21272 : INV_X1 port map( A => n2433, ZN => n29158);
   U21348 : XNOR2_X1 port map( A => n25452, B => n25451, ZN => n29159);
   U21367 : NOR2_X1 port map( A1 => n25472, A2 => n28670, ZN => n29160);
   U21384 : NOR2_X1 port map( A1 => n25472, A2 => n28670, ZN => n29161);
   U21386 : NOR2_X1 port map( A1 => n25472, A2 => n28670, ZN => n28024);
   U21422 : NAND2_X1 port map( A1 => n4305, A2 => n9211, ZN => n9207);
   U21423 : XNOR2_X1 port map( A => n29163, B => n22761, ZN => n22767);
   U21447 : XNOR2_X1 port map( A => n22758, B => n22757, ZN => n29163);
   U21487 : NAND2_X1 port map( A1 => n29165, A2 => n29164, ZN => n20767);
   U21565 : NAND2_X1 port map( A1 => n20287, A2 => n20286, ZN => n29164);
   U21591 : NAND2_X1 port map( A1 => n20288, A2 => n29166, ZN => n29165);
   U21621 : NOR3_X1 port map( A1 => n29168, A2 => n26536, A3 => n26535, ZN => 
                           Ciphertext(25));
   U21632 : NAND2_X1 port map( A1 => n28605, A2 => n8200, ZN => n28246);
   U21722 : NAND2_X1 port map( A1 => n7423, A2 => n3112, ZN => n7370);
   U21826 : NAND3_X1 port map( A1 => n3161, A2 => n11349, A3 => n11355, ZN => 
                           n11354);
   U21889 : NAND2_X1 port map( A1 => n10765, A2 => n10764, ZN => n13109);
   U22216 : NAND2_X1 port map( A1 => n13889, A2 => n29153, ZN => n29171);
   U22218 : NAND2_X1 port map( A1 => n13890, A2 => n545, ZN => n29172);
   U22347 : NAND2_X1 port map( A1 => n4835, A2 => n15464, ZN => n29173);
   U22363 : NAND2_X1 port map( A1 => n24073, A2 => n24072, ZN => n29174);
   U22390 : NAND2_X1 port map( A1 => n5856, A2 => n23418, ZN => n23097);
   U22437 : NAND2_X1 port map( A1 => n4274, A2 => n4275, ZN => n10545);
   U22474 : NAND3_X1 port map( A1 => n386, A2 => n4306, A3 => n28408, ZN => 
                           n5358);
   U22506 : NAND2_X1 port map( A1 => n17873, A2 => n17938, ZN => n17874);
   U22514 : NAND3_X1 port map( A1 => n17416, A2 => n5430, A3 => n17413, ZN => 
                           n29176);
   U22573 : NAND3_X1 port map( A1 => n21661, A2 => n21654, A3 => n21655, ZN => 
                           n20835);
   U22692 : NAND2_X1 port map( A1 => n529, A2 => n17439, ZN => n29177);
   U22799 : NAND2_X1 port map( A1 => n17846, A2 => n18137, ZN => n17848);
   U22807 : NAND2_X1 port map( A1 => n8590, A2 => n8973, ZN => n8597);
   U22818 : NAND2_X1 port map( A1 => n21449, A2 => n21448, ZN => n29178);
   U22819 : NAND2_X1 port map( A1 => n29179, A2 => n11873, ZN => n12849);
   U22829 : NAND2_X1 port map( A1 => n6305, A2 => n6304, ZN => n29179);
   U22837 : NAND2_X1 port map( A1 => n29181, A2 => n20265, ZN => n29180);
   U22840 : NAND2_X1 port map( A1 => n6202, A2 => n6204, ZN => n29181);
   U22848 : INV_X1 port map( A => n20265, ZN => n29183);
   U22904 : NAND3_X1 port map( A1 => n28745, A2 => n18486, A3 => n18493, ZN => 
                           n1997);
   U22910 : NAND2_X1 port map( A1 => n20478, A2 => n20477, ZN => n20232);
   U22915 : XNOR2_X2 port map( A => n15560, B => n15559, ZN => n17338);
   U22987 : NAND3_X1 port map( A1 => n412, A2 => n21678, A3 => n21448, ZN => 
                           n2909);
   U22988 : NAND2_X1 port map( A1 => n29185, A2 => n585, ZN => n2954);
   U22996 : NAND2_X1 port map( A1 => n11026, A2 => n11027, ZN => n29185);
   U23024 : OAI211_X1 port map( C1 => n21633, C2 => n21631, A => n21036, B => 
                           n28797, ZN => n29186);
   U23054 : NAND2_X1 port map( A1 => n24155, A2 => n28785, ZN => n24249);
   U23086 : NAND4_X1 port map( A1 => n25671, A2 => n25672, A3 => n29188, A4 => 
                           n29187, ZN => n25675);
   U23087 : NAND2_X1 port map( A1 => n25658, A2 => n27350, ZN => n29187);
   U23120 : NAND2_X1 port map( A1 => n27351, A2 => n25657, ZN => n29188);
   U23288 : NAND2_X1 port map( A1 => n23535, A2 => n23531, ZN => n5481);
   U23311 : OR2_X1 port map( A1 => n24237, A2 => n29642, ZN => n6238);
   U23384 : NAND2_X1 port map( A1 => n29189, A2 => n28821, ZN => n24155);
   U23385 : NAND2_X1 port map( A1 => n23608, A2 => n23211, ZN => n29189);
   U23434 : NAND2_X1 port map( A1 => n3549, A2 => n17364, ZN => n16760);
   U23435 : NAND2_X1 port map( A1 => n17234, A2 => n17368, ZN => n17364);
   U23506 : NAND2_X1 port map( A1 => n1576, A2 => n512, ZN => n29191);
   U23535 : NAND2_X1 port map( A1 => n1577, A2 => n16862, ZN => n29192);
   U23543 : NAND2_X2 port map( A1 => n29193, A2 => n24519, ZN => n25909);
   U23563 : NAND2_X1 port map( A1 => n28284, A2 => n28285, ZN => n26578);
   U23587 : NOR2_X2 port map( A1 => n5194, A2 => n19962, ZN => n21472);
   U23683 : NAND2_X1 port map( A1 => n4914, A2 => n1574, ZN => n29194);
   U23684 : AND3_X2 port map( A1 => n19185, A2 => n29197, A3 => n29196, ZN => 
                           n21372);
   U23723 : NAND2_X1 port map( A1 => n19179, A2 => n19863, ZN => n29196);
   U23724 : NAND2_X1 port map( A1 => n1041, A2 => n19867, ZN => n29197);
   U23756 : OAI211_X2 port map( C1 => n1750, C2 => n9410, A => n29198, B => 
                           n6505, ZN => n10271);
   U23806 : NAND2_X1 port map( A1 => n9040, A2 => n9410, ZN => n29198);
   U23938 : NAND3_X1 port map( A1 => n2422, A2 => n10699, A3 => n2423, ZN => 
                           n11491);
   U23965 : NAND3_X1 port map( A1 => n16830, A2 => n2485, A3 => n16829, ZN => 
                           n2484);
   U24032 : NAND3_X1 port map( A1 => n10754, A2 => n11152, A3 => n10804, ZN => 
                           n10755);
   U24033 : NAND3_X1 port map( A1 => n12022, A2 => n29209, A3 => n12428, ZN => 
                           n1369);
   U24079 : NAND3_X1 port map( A1 => n6434, A2 => n6307, A3 => n14310, ZN => 
                           n6433);
   U24098 : NAND2_X1 port map( A1 => n5981, A2 => n14393, ZN => n29201);
   U24135 : NOR2_X1 port map( A1 => n29202, A2 => n11831, ZN => n11832);
   U24137 : NOR3_X1 port map( A1 => n6281, A2 => n12207, A3 => n12206, ZN => 
                           n29202);
   U24228 : NAND2_X1 port map( A1 => n465, A2 => n24633, ZN => n24560);
   U24268 : NAND3_X1 port map( A1 => n15322, A2 => n15327, A3 => n15013, ZN => 
                           n1106);
   U24326 : NAND2_X1 port map( A1 => n1068, A2 => n27955, ZN => n29277);
   U24334 : NAND3_X1 port map( A1 => n18158, A2 => n18160, A3 => n18159, ZN => 
                           n18161);
   U24392 : NOR2_X1 port map( A1 => n4214, A2 => n29204, ZN => n17061);
   U24431 : NAND2_X1 port map( A1 => n7750, A2 => n8161, ZN => n7157);
   U24623 : NAND2_X1 port map( A1 => n29206, A2 => n29205, ZN => n16840);
   U24624 : NAND2_X1 port map( A1 => n17312, A2 => n29550, ZN => n29205);
   U24713 : NAND2_X1 port map( A1 => n16836, A2 => n17560, ZN => n29206);
   U24747 : NAND2_X1 port map( A1 => n15514, A2 => n15515, ZN => n15277);
   U24807 : NAND2_X1 port map( A1 => n14886, A2 => n29207, ZN => n6668);
   U24811 : OR2_X1 port map( A1 => n14972, A2 => n14969, ZN => n29207);
   U24813 : INV_X1 port map( A => n10816, ZN => n28207);
   U24890 : XNOR2_X1 port map( A => n8479, B => n8480, ZN => n10816);
   U24909 : NAND3_X1 port map( A1 => n512, A2 => n17802, A3 => n29507, ZN => 
                           n227);
   U24928 : NAND3_X1 port map( A1 => n28820, A2 => n20039, A3 => n20090, ZN => 
                           n6410);
   U24964 : OR2_X1 port map( A1 => n22991, A2 => n23563, ZN => n22993);
   U24972 : NAND2_X1 port map( A1 => n15436, A2 => n15300, ZN => n14664);
   U24976 : NAND2_X1 port map( A1 => n17508, A2 => n17829, ZN => n28323);
   U24977 : OAI21_X1 port map( B1 => n10568, B2 => n10623, A => n11896, ZN => 
                           n29208);
   U24987 : NAND2_X1 port map( A1 => n29210, A2 => n29209, ZN => n26);
   U24994 : NAND2_X1 port map( A1 => n11467, A2 => n12428, ZN => n29210);
   U25003 : OAI211_X2 port map( C1 => n15268, C2 => n15494, A => n14619, B => 
                           n29211, ZN => n16399);
   U25023 : NAND2_X1 port map( A1 => n11283, A2 => n29212, ZN => n10380);
   U25047 : NAND2_X1 port map( A1 => n10779, A2 => n10966, ZN => n10782);
   U25127 : NAND2_X1 port map( A1 => n6556, A2 => n24538, ZN => n24539);
   U25140 : NAND3_X1 port map( A1 => n6692, A2 => n6691, A3 => n8979, ZN => 
                           n203);
   U25141 : OAI21_X1 port map( B1 => n7784, B2 => n2670, A => n7783, ZN => 
                           n29214);
   U25193 : NAND2_X1 port map( A1 => n454, A2 => n4820, ZN => n6435);
   U25216 : NAND2_X1 port map( A1 => n27908, A2 => n27092, ZN => n27883);
   U25242 : NAND3_X1 port map( A1 => n11930, A2 => n568, A3 => n12267, ZN => 
                           n1491);
   U25243 : MUX2_X1 port map( A => n17767, B => n18387, S => n18388, Z => 
                           n17736);
   U25269 : NAND2_X1 port map( A1 => n29215, A2 => n10488, ZN => n10648);
   U25294 : NAND2_X1 port map( A1 => n10485, A2 => n11057, ZN => n29215);
   U25305 : OAI21_X1 port map( B1 => n2425, B2 => n2029, A => n8958, ZN => 
                           n8624);
   U25345 : OR2_X1 port map( A1 => n18414, A2 => n18121, ZN => n3915);
   U25360 : NAND2_X1 port map( A1 => n27381, A2 => n29217, ZN => n27385);
   U25400 : OAI21_X1 port map( B1 => n27376, B2 => n29219, A => n29218, ZN => 
                           n29217);
   U25401 : NAND2_X1 port map( A1 => n29220, A2 => n22878, ZN => n24278);
   U25408 : NAND4_X1 port map( A1 => n1151, A2 => n1284, A3 => n2202, A4 => 
                           n1150, ZN => n29220);
   U25495 : NAND2_X1 port map( A1 => n28332, A2 => n28334, ZN => n11180);
   U25496 : NAND2_X1 port map( A1 => n9435, A2 => n29221, ZN => n7683);
   U25541 : NAND3_X1 port map( A1 => n15029, A2 => n15430, A3 => n15028, ZN => 
                           n15035);
   U25551 : AOI22_X2 port map( A1 => n9693, A2 => n28405, B1 => n9694, B2 => 
                           n592, ZN => n12186);
   U25589 : NAND2_X1 port map( A1 => n29222, A2 => n9060, ZN => n8107);
   U25607 : OAI21_X1 port map( B1 => n9059, B2 => n9064, A => n8397, ZN => 
                           n29222);
   U25704 : NAND2_X1 port map( A1 => n29223, A2 => n17434, ZN => n4428);
   U25723 : NAND2_X1 port map( A1 => n17308, A2 => n16962, ZN => n29223);
   U25765 : NAND2_X1 port map( A1 => n21375, A2 => n21702, ZN => n29224);
   U25766 : NAND2_X1 port map( A1 => n29226, A2 => n29227, ZN => n29225);
   U25801 : INV_X1 port map( A => n21378, ZN => n29226);
   U25920 : INV_X2 port map( A => n21709, ZN => n29227);
   U25998 : OAI21_X1 port map( B1 => n7795, B2 => n7796, A => n29229, ZN => 
                           n7544);
   U25999 : NAND2_X1 port map( A1 => n7796, A2 => n7542, ZN => n29229);
   U26068 : NAND3_X1 port map( A1 => n29230, A2 => n7685, A3 => n7520, ZN => 
                           n7013);
   U26069 : NAND2_X1 port map( A1 => n7684, A2 => n7517, ZN => n29230);
   U26110 : AND3_X2 port map( A1 => n2270, A2 => n26335, A3 => n2269, ZN => 
                           n27818);
   U26172 : XNOR2_X2 port map( A => n6467, B => n19163, ZN => n5225);
   U26240 : OAI21_X1 port map( B1 => n27819, B2 => n29232, A => n29231, ZN => 
                           n26679);
   U26255 : NAND2_X1 port map( A1 => n27819, A2 => n27818, ZN => n29231);
   U26339 : INV_X1 port map( A => n27795, ZN => n29232);
   U26385 : NAND3_X1 port map( A1 => n20056, A2 => n6114, A3 => n20171, ZN => 
                           n29233);
   U26397 : NAND2_X1 port map( A1 => n11242, A2 => n11069, ZN => n10198);
   U26523 : NAND2_X1 port map( A1 => n7980, A2 => n7985, ZN => n7459);
   U26555 : OAI21_X1 port map( B1 => n20400, B2 => n20401, A => n20562, ZN => 
                           n29235);
   U26582 : INV_X1 port map( A => n28580, ZN => n29236);
   U26596 : NAND2_X1 port map( A1 => n21560, A2 => n5953, ZN => n20862);
   U26618 : NAND3_X1 port map( A1 => n5126, A2 => n28658, A3 => n29315, ZN => 
                           n4472);
   U26649 : NAND2_X1 port map( A1 => n28542, A2 => n26948, ZN => n6469);
   U26716 : NAND2_X1 port map( A1 => n1333, A2 => n1332, ZN => n29237);
   U26769 : NAND2_X1 port map( A1 => n2329, A2 => n1708, ZN => n29238);
   U26783 : AND3_X2 port map( A1 => n29239, A2 => n11766, A3 => n6725, ZN => 
                           n15108);
   U26910 : NAND2_X1 port map( A1 => n11765, A2 => n293, ZN => n29239);
   U27074 : NAND3_X1 port map( A1 => n7074, A2 => n7884, A3 => n7882, ZN => 
                           n7076);
   U27089 : NAND2_X1 port map( A1 => n9083, A2 => n9082, ZN => n7490);
   U27141 : NAND2_X1 port map( A1 => n2099, A2 => n8270, ZN => n9083);
   U27142 : XNOR2_X2 port map( A => n20471, B => n20472, ZN => n23531);
   U27143 : AOI21_X2 port map( B1 => n17231, B2 => n871, A => n17230, ZN => 
                           n18148);
   U27253 : NAND2_X1 port map( A1 => n2357, A2 => n12162, ZN => n12171);
   U27269 : OR2_X1 port map( A1 => n17383, A2 => n17384, ZN => n29240);
   U27271 : NAND2_X1 port map( A1 => n8808, A2 => n8809, ZN => n29242);
   U27272 : NAND2_X1 port map( A1 => n4195, A2 => n24669, ZN => n4194);
   U27304 : OR3_X1 port map( A1 => n18042, A2 => n18421, A3 => n29507, ZN => 
                           n18425);
   U27339 : NAND2_X1 port map( A1 => n29245, A2 => n29243, ZN => n13191);
   U27344 : OAI21_X1 port map( B1 => n12004, B2 => n11760, A => n11758, ZN => 
                           n29244);
   U27354 : OAI21_X1 port map( B1 => n11757, B2 => n11756, A => n12004, ZN => 
                           n29245);
   U27425 : NAND2_X1 port map( A1 => n14424, A2 => n14425, ZN => n4523);
   U27487 : NAND2_X1 port map( A1 => n29246, A2 => n28813, ZN => n21676);
   U27513 : NAND2_X1 port map( A1 => n20211, A2 => n20210, ZN => n29246);
   U27519 : NAND2_X1 port map( A1 => n24351, A2 => n24712, ZN => n29248);
   U27547 : NAND2_X1 port map( A1 => n23070, A2 => n28416, ZN => n29249);
   U27582 : NAND3_X1 port map( A1 => n2281, A2 => n23816, A3 => n28609, ZN => 
                           n3990);
   U27600 : NOR2_X1 port map( A1 => n29251, A2 => n23819, ZN => n23822);
   U27611 : NAND2_X1 port map( A1 => n407, A2 => n23290, ZN => n29251);
   U27727 : NAND2_X1 port map( A1 => n21669, A2 => n22401, ZN => n2072);
   U27729 : XNOR2_X2 port map( A => Key(80), B => Plaintext(80), ZN => n7690);
   U27751 : NAND2_X1 port map( A1 => n29253, A2 => n23100, ZN => n23101);
   U27776 : OAI21_X1 port map( B1 => n23098, B2 => n23097, A => n23096, ZN => 
                           n29253);
   U27790 : INV_X1 port map( A => n24813, ZN => n220);
   U27934 : NAND3_X1 port map( A1 => n29255, A2 => n5707, A3 => n5710, ZN => 
                           n5704);
   U28001 : NAND2_X1 port map( A1 => n5709, A2 => n11237, ZN => n29255);
   U28033 : NOR2_X2 port map( A1 => n29256, A2 => n1312, ZN => n22913);
   U28036 : NAND2_X1 port map( A1 => n7744, A2 => n7743, ZN => n7524);
   U28110 : NAND2_X1 port map( A1 => n29257, A2 => n11538, ZN => n6146);
   U28124 : NAND2_X1 port map( A1 => n11685, A2 => n11540, ZN => n29257);
   U28125 : OAI21_X1 port map( B1 => n6906, B2 => n2107, A => n24195, ZN => 
                           n24197);
   U28153 : NAND2_X1 port map( A1 => n24644, A2 => n24642, ZN => n24195);
   U28154 : NAND2_X1 port map( A1 => n14613, A2 => n14612, ZN => n14614);
   U28160 : NAND2_X1 port map( A1 => n7685, A2 => n7844, ZN => n7686);
   U28164 : OAI211_X2 port map( C1 => n21321, C2 => n21137, A => n21589, B => 
                           n4962, ZN => n22418);
   U28166 : NOR2_X1 port map( A1 => n29258, A2 => n27432, ZN => n25426);
   U28176 : OAI21_X1 port map( B1 => n26829, B2 => n27434, A => n26708, ZN => 
                           n29258);
   U28197 : AOI21_X1 port map( B1 => n6194, B2 => n6197, A => n6196, ZN => 
                           n29259);
   U28199 : XNOR2_X1 port map( A => n29261, B => n29260, ZN => Ciphertext(153))
                           ;
   U28205 : INV_X1 port map( A => n27894, ZN => n29260);
   U28213 : OAI211_X1 port map( C1 => n27892, C2 => n27893, A => n27891, B => 
                           n27890, ZN => n29261);
   U28216 : NOR2_X2 port map( A1 => n29262, A2 => n20442, ZN => n21513);
   U28217 : AOI22_X1 port map( A1 => n20439, A2 => n20438, B1 => n20436, B2 => 
                           n29508, ZN => n29262);
   U28218 : NAND2_X1 port map( A1 => n6864, A2 => n6865, ZN => n4238);
   U28219 : NAND2_X1 port map( A1 => n10742, A2 => n29263, ZN => n4274);
   U28220 : NAND2_X1 port map( A1 => n223, A2 => n14894, ZN => n3360);
   U28221 : NOR2_X2 port map( A1 => n21517, A2 => n21518, ZN => n22615);
   U28222 : NAND2_X1 port map( A1 => n71, A2 => n4448, ZN => n29264);
   U28223 : NAND3_X1 port map( A1 => n20189, A2 => n6261, A3 => n19959, ZN => 
                           n6260);
   U28224 : XNOR2_X1 port map( A => n15849, B => n2465, ZN => n15851);
   U28225 : NAND2_X1 port map( A1 => n3777, A2 => n14875, ZN => n15849);
   U28226 : NAND2_X1 port map( A1 => n27156, A2 => n28180, ZN => n27158);
   U28227 : NAND2_X1 port map( A1 => n17687, A2 => n20417, ZN => n20418);
   U28229 : NAND2_X1 port map( A1 => n21623, A2 => n22141, ZN => n29265);
   U28230 : NAND2_X1 port map( A1 => n27663, A2 => n27661, ZN => n27652);
   U28231 : NOR2_X2 port map( A1 => n23278, A2 => n23279, ZN => n24083);
   U28234 : NAND2_X1 port map( A1 => n21708, A2 => n496, ZN => n6104);
   U28235 : NAND2_X1 port map( A1 => n21703, A2 => n21277, ZN => n21708);
   U28236 : NAND2_X1 port map( A1 => n6086, A2 => n20406, ZN => n6085);
   U28237 : AND2_X2 port map( A1 => n3308, A2 => n7335, ZN => n8562);
   U28240 : NAND2_X1 port map( A1 => n5054, A2 => n5055, ZN => n3648);
   U28242 : NAND2_X1 port map( A1 => n14417, A2 => n14418, ZN => n14449);
   U28243 : NAND2_X1 port map( A1 => n19052, A2 => n29584, ZN => n19057);
   U28244 : NAND2_X1 port map( A1 => n24894, A2 => n23982, ZN => n29268);
   U28245 : NAND2_X1 port map( A1 => n24295, A2 => n24294, ZN => n29269);
   U28246 : NAND3_X1 port map( A1 => n1268, A2 => n1267, A3 => n1269, ZN => 
                           n1266);
   U28247 : NAND4_X2 port map( A1 => n6216, A2 => n6217, A3 => n29271, A4 => 
                           n29270, ZN => n16185);
   U28248 : NAND2_X1 port map( A1 => n15502, A2 => n14923, ZN => n29270);
   U28249 : NAND2_X1 port map( A1 => n14707, A2 => n15506, ZN => n29271);
   U28250 : NAND2_X1 port map( A1 => n1739, A2 => n25656, ZN => n28669);
   U28251 : NOR2_X1 port map( A1 => n26738, A2 => n26737, ZN => n1739);
   U28252 : INV_X1 port map( A => n7847, ZN => n7260);
   U28253 : NAND2_X1 port map( A1 => n7846, A2 => n8024, ZN => n7847);
   U28254 : NAND2_X1 port map( A1 => n26686, A2 => n395, ZN => n29288);
   U28255 : NAND2_X1 port map( A1 => n27300, A2 => n26879, ZN => n26686);
   U28256 : NAND2_X1 port map( A1 => n29272, A2 => n18334, ZN => n18336);
   U28257 : NAND2_X1 port map( A1 => n18333, A2 => n817, ZN => n29272);
   U28258 : XNOR2_X1 port map( A => n29273, B => n10409, ZN => n10414);
   U28259 : NAND3_X1 port map( A1 => n3877, A2 => n18423, A3 => n1942, ZN => 
                           n3876);
   U28260 : NAND2_X1 port map( A1 => n29274, A2 => n16862, ZN => n5495);
   U28261 : NAND3_X1 port map( A1 => n2789, A2 => n7511, A3 => n2788, ZN => 
                           n3683);
   U28262 : XNOR2_X1 port map( A => n29275, B => n28097, ZN => Ciphertext(189))
                           ;
   U28263 : NAND3_X1 port map( A1 => n28095, A2 => n3470, A3 => n3469, ZN => 
                           n29275);
   U28264 : NAND2_X1 port map( A1 => n29276, A2 => n11140, ZN => n1452);
   U28265 : NAND2_X1 port map( A1 => n11138, A2 => n11139, ZN => n29276);
   U28266 : OR2_X1 port map( A1 => n11473, A2 => n10648, ZN => n12345);
   U28267 : INV_X1 port map( A => n14570, ZN => n15076);
   U28268 : NAND2_X1 port map( A1 => n14874, A2 => n15071, ZN => n14570);
   U28269 : NAND2_X1 port map( A1 => n142, A2 => n602, ZN => n8130);
   U28270 : XNOR2_X1 port map( A => n29277, B => n27957, ZN => Ciphertext(162))
                           ;
   U28272 : AOI22_X1 port map( A1 => n1684, A2 => n27364, B1 => n26496, B2 => 
                           n27370, ZN => n29278);
   U28273 : NAND2_X1 port map( A1 => n7919, A2 => n7619, ZN => n7430);
   U28274 : AOI21_X1 port map( B1 => n19898, B2 => n3009, A => n19897, ZN => 
                           n21124);
   U28275 : AND3_X2 port map( A1 => n26154, A2 => n26153, A3 => n29279, ZN => 
                           n27465);
   U28276 : NAND3_X1 port map( A1 => n28286, A2 => n25418, A3 => n6826, ZN => 
                           n29279);
   U28277 : NAND2_X1 port map( A1 => n29281, A2 => n29280, ZN => n26744);
   U28278 : NAND2_X1 port map( A1 => n26739, A2 => n26235, ZN => n29280);
   U28279 : NAND2_X1 port map( A1 => n26738, A2 => n26737, ZN => n29281);
   U28280 : OAI211_X2 port map( C1 => n20846, C2 => n6247, A => n5175, B => 
                           n29282, ZN => n22279);
   U28281 : NAND3_X1 port map( A1 => n19904, A2 => n21125, A3 => n21461, ZN => 
                           n29282);
   U28282 : OAI211_X1 port map( C1 => n26608, C2 => n27458, A => n29284, B => 
                           n29283, ZN => n26609);
   U28283 : NAND2_X1 port map( A1 => n26605, A2 => n27447, ZN => n29283);
   U28284 : NAND2_X1 port map( A1 => n27458, A2 => n26606, ZN => n29284);
   U28285 : NAND2_X1 port map( A1 => n29286, A2 => n29285, ZN => n26630);
   U28286 : OR3_X1 port map( A1 => n29481, A2 => n26733, A3 => n26995, ZN => 
                           n29285);
   U28287 : NAND2_X1 port map( A1 => n26628, A2 => n26995, ZN => n29286);
   U28289 : AOI22_X1 port map( A1 => n26887, A2 => n5425, B1 => n29288, B2 => 
                           n29287, ZN => n26446);
   U28290 : INV_X1 port map( A => n444, ZN => n29287);
   U28291 : OAI21_X1 port map( B1 => n18157, B2 => n17744, A => n29289, ZN => 
                           n2501);
   U28292 : NOR2_X1 port map( A1 => n17614, A2 => n17616, ZN => n17307);
   U28293 : NAND2_X1 port map( A1 => n6001, A2 => n17303, ZN => n17614);
   U28294 : NAND2_X1 port map( A1 => n29290, A2 => n15399, ZN => n6262);
   U28296 : NAND2_X1 port map( A1 => n3900, A2 => n29291, ZN => n3166);
   U28297 : NOR2_X2 port map( A1 => n2534, A2 => n29292, ZN => n21268);
   U28298 : NAND2_X1 port map( A1 => n28383, A2 => n28384, ZN => n29292);
   U28299 : NAND2_X1 port map( A1 => n1109, A2 => n1110, ZN => n21013);
   U28302 : NAND3_X1 port map( A1 => n29121, A2 => n29056, A3 => n28089, ZN => 
                           n28080);
   U28303 : OAI22_X1 port map( A1 => n27204, A2 => n27547, B1 => n27205, B2 => 
                           n28422, ZN => n27206);
   U28305 : XNOR2_X1 port map( A => n15721, B => n15722, ZN => n17362);
   U28307 : INV_X1 port map( A => n20351, ZN => n21553);
   U28308 : XOR2_X1 port map( A => n24868, B => n24869, Z => n29293);
   U2951 : AOI21_X2 port map( B1 => n12673, B2 => n190, A => n12672, ZN => 
                           n15103);
   U1024 : OAI21_X2 port map( B1 => n22975, B2 => n22974, A => n22973, ZN => 
                           n24434);
   U827 : OR2_X2 port map( A1 => n15479, A2 => n15478, ZN => n16319);
   U9166 : OAI211_X2 port map( C1 => n8130, C2 => n8129, A => n8128, B => n8127
                           , ZN => n2845);
   U18281 : BUF_X2 port map( A => n12711, Z => n14204);
   U3585 : NAND2_X2 port map( A1 => n4111, A2 => n6874, ZN => n8642);
   U1493 : NAND3_X2 port map( A1 => n28982, A2 => n5865, A3 => n1132, ZN => 
                           n21549);
   U270 : BUF_X2 port map( A => n26841, Z => n27088);
   U1724 : INV_X2 port map( A => n20425, ZN => n21823);
   U28187 : NAND2_X2 port map( A1 => n28756, A2 => n15210, ZN => n16404);
   U1359 : AND2_X2 port map( A1 => n5462, A2 => n12243, ZN => n13054);
   U3064 : AND3_X2 port map( A1 => n2682, A2 => n6280, A3 => n2685, ZN => 
                           n13523);
   U2375 : BUF_X1 port map( A => n7838, Z => n7700);
   U1126 : NOR2_X2 port map( A1 => n23597, A2 => n23467, ZN => n24975);
   U730 : NAND3_X2 port map( A1 => n20126, A2 => n20127, A3 => n20128, ZN => 
                           n5827);
   U426 : BUF_X1 port map( A => n10318, Z => n11076);
   U2606 : BUF_X1 port map( A => n19787, Z => n20632);
   U1531 : XNOR2_X2 port map( A => n19177, B => n19178, ZN => n20496);
   U1343 : XNOR2_X2 port map( A => n13023, B => n13022, ZN => n14362);
   U5227 : XNOR2_X2 port map( A => n1619, B => n18641, ZN => n20209);
   U10374 : NAND3_X2 port map( A1 => n28372, A2 => n8010, A3 => n8011, ZN => 
                           n9504);
   U9320 : AOI22_X2 port map( A1 => n5022, A2 => n18406, B1 => n18709, B2 => 
                           n18407, ZN => n18948);
   U619 : AND2_X2 port map( A1 => n10841, A2 => n10840, ZN => n12244);
   U2538 : AND2_X2 port map( A1 => n3855, A2 => n21435, ZN => n21442);
   U9076 : OAI21_X2 port map( B1 => n17180, B2 => n1801, A => n17178, ZN => 
                           n18411);
   U659 : OAI21_X2 port map( B1 => n23219, B2 => n23610, A => n23218, ZN => 
                           n24248);
   U312 : BUF_X2 port map( A => n8608, Z => n9532);
   U678 : BUF_X2 port map( A => n17679, Z => n18478);
   U1274 : BUF_X1 port map( A => n21729, Z => n1929);
   U2913 : AND3_X2 port map( A1 => n4519, A2 => n4521, A3 => n14430, ZN => 
                           n15506);
   U789 : NOR2_X2 port map( A1 => n2201, A2 => n22744, ZN => n24551);
   U10018 : AOI21_X2 port map( B1 => n18347, B2 => n18346, A => n18345, ZN => 
                           n18680);
   U1500 : NAND3_X2 port map( A1 => n17510, A2 => n5807, A3 => n17511, ZN => 
                           n17592);
   U7022 : AND3_X2 port map( A1 => n4795, A2 => n5399, A3 => n16763, ZN => 
                           n18441);
   U2528 : AND2_X2 port map( A1 => n19987, A2 => n19988, ZN => n20663);
   U3572 : BUF_X1 port map( A => n19795, Z => n20261);
   U3562 : OR2_X2 port map( A1 => n674, A2 => n23274, ZN => n25008);
   U1648 : NAND2_X2 port map( A1 => n689, A2 => n23944, ZN => n25708);
   U16940 : OR2_X2 port map( A1 => n10471, A2 => n10470, ZN => n12339);
   U5184 : XNOR2_X2 port map( A => n15367, B => n15368, ZN => n17298);
   U1222 : NAND2_X2 port map( A1 => n5550, A2 => n3719, ZN => n19617);
   U618 : BUF_X2 port map( A => n11385, Z => n12991);
   U1569 : INV_X2 port map( A => n18408, ZN => n28798);
   U82 : NAND2_X1 port map( A1 => n20739, A2 => n20737, ZN => n21156);
   U11124 : XNOR2_X2 port map( A => n4989, B => n5566, ZN => n3880);
   U10641 : INV_X1 port map( A => n3829, ZN => n11137);
   U5413 : INV_X2 port map( A => n5023, ZN => n18709);
   U2539 : NOR2_X2 port map( A1 => n18890, A2 => n18889, ZN => n20988);
   U19671 : INV_X1 port map( A => n14921, ZN => n16038);
   U1224 : BUF_X2 port map( A => n20013, Z => n20510);
   U1622 : BUF_X2 port map( A => n27408, Z => n28177);
   U1416 : OAI211_X2 port map( C1 => n29228, C2 => n29227, A => n29225, B => 
                           n29224, ZN => n22464);
   U4094 : BUF_X1 port map( A => n26682, Z => n27434);
   U809 : BUF_X1 port map( A => n12955, Z => n13218);
   U1744 : NAND2_X2 port map( A1 => n28953, A2 => n28952, ZN => n15127);
   U18138 : NAND2_X2 port map( A1 => n14907, A2 => n14905, ZN => n15098);
   U3141 : NAND3_X2 port map( A1 => n9055, A2 => n9054, A3 => n9056, ZN => 
                           n12200);
   U1672 : AND3_X2 port map( A1 => n5445, A2 => n5444, A3 => n14515, ZN => 
                           n15828);
   U340 : MUX2_X2 port map( A => n20297, B => n20296, S => n20295, Z => n21308)
                           ;
   U7244 : OAI21_X2 port map( B1 => n22277, B2 => n23636, A => n5457, ZN => 
                           n22356);
   U1002 : NOR2_X2 port map( A1 => n1339, A2 => n22014, ZN => n22923);
   U15066 : BUF_X1 port map( A => n23633, Z => n29061);
   U1519 : OR2_X2 port map( A1 => n21275, A2 => n21283, ZN => n21709);
   U26 : OAI211_X2 port map( C1 => n6933, C2 => n4633, A => n4632, B => n4631, 
                           ZN => n22882);
   U1480 : NAND2_X2 port map( A1 => n20715, A2 => n20713, ZN => n21591);
   U11677 : BUF_X1 port map( A => n26350, Z => n28410);
   U2352 : BUF_X1 port map( A => n10008, Z => n28616);
   U2163 : NAND2_X2 port map( A1 => n11792, A2 => n28701, ZN => n13020);
   U2641 : INV_X2 port map( A => n2571, ZN => n19198);
   U2361 : NAND4_X1 port map( A1 => n8986, A2 => n8985, A3 => n8988, A4 => 
                           n8987, ZN => n10258);
   U3354 : NAND2_X2 port map( A1 => n4695, A2 => n4698, ZN => n9531);
   U1647 : AND2_X2 port map( A1 => n28256, A2 => n28255, ZN => n25509);
   U1114 : NOR2_X2 port map( A1 => n27062, A2 => n27061, ZN => n27905);
   U9848 : NAND3_X2 port map( A1 => n15424, A2 => n15418, A3 => n15419, ZN => 
                           n16569);
   U956 : NAND2_X2 port map( A1 => n10899, A2 => n172, ZN => n13101);
   U3649 : INV_X2 port map( A => n21657, ZN => n6275);
   U11637 : NAND2_X2 port map( A1 => n25359, A2 => n25357, ZN => n27366);
   U13179 : MUX2_X2 port map( A => n26760, B => n25276, S => n26755, Z => 
                           n25359);
   U796 : XNOR2_X2 port map( A => n22834, B => n22833, ZN => n23290);
   U1322 : AND2_X2 port map( A1 => n5885, A2 => n5884, ZN => n24631);
   U1560 : OAI21_X2 port map( B1 => n15736, B2 => n15737, A => n15735, ZN => 
                           n19103);
   U866 : OAI21_X1 port map( B1 => n14412, B2 => n14411, A => n4001, ZN => 
                           n14922);
   U6631 : OR2_X1 port map( A1 => n2382, A2 => n7084, ZN => n4675);
   U2938 : OAI21_X2 port map( B1 => n13259, B2 => n14312, A => n2331, ZN => 
                           n14563);
   U3830 : NAND3_X2 port map( A1 => n908, A2 => n4473, A3 => n907, ZN => n24388
                           );
   U25124 : OAI211_X2 port map( C1 => n23510, C2 => n24081, A => n23509, B => 
                           n23508, ZN => n25324);
   U1638 : MUX2_X2 port map( A => n8332, B => n8331, S => n8763, Z => n10137);
   U1540 : XNOR2_X2 port map( A => n9945, B => n9944, ZN => n10461);
   U1907 : NAND3_X2 port map( A1 => n15080, A2 => n15079, A3 => n28221, ZN => 
                           n15865);
   U617 : BUF_X1 port map( A => n10657, Z => n10872);
   U1083 : BUF_X2 port map( A => n23422, Z => n23344);
   U9543 : NAND3_X2 port map( A1 => n3051, A2 => n8750, A3 => n3050, ZN => 
                           n10149);
   U3594 : XNOR2_X2 port map( A => n18742, B => n18741, ZN => n29114);
   U13051 : AND3_X2 port map( A1 => n5749, A2 => n5750, A3 => n5748, ZN => 
                           n25819);
   U3000 : XNOR2_X2 port map( A => n10772, B => n10773, ZN => n14107);
   U2879 : NAND2_X2 port map( A1 => n11425, A2 => n11424, ZN => n12420);
   U14814 : XNOR2_X2 port map( A => n7203, B => Key(134), ZN => n7400);
   U102 : AND3_X2 port map( A1 => n1597, A2 => n15130, A3 => n15129, ZN => 
                           n3661);
   U1491 : AOI21_X1 port map( B1 => n14183, B2 => n14470, A => n5598, ZN => 
                           n15165);
   U13203 : XNOR2_X2 port map( A => n6707, B => n13927, ZN => n5891);
   U5292 : OAI21_X1 port map( B1 => n12452, B2 => n12451, A => n1671, ZN => 
                           n15097);
   U931 : NAND2_X2 port map( A1 => n11987, A2 => n163, ZN => n13543);
   U11329 : NAND2_X2 port map( A1 => n10521, A2 => n4068, ZN => n11449);
   U3465 : INV_X1 port map( A => n2984, ZN => n624);
   U4478 : XNOR2_X1 port map( A => n26099, B => n26098, ZN => n27137);
   U4475 : NOR3_X1 port map( A1 => n27147, A2 => n27142, A3 => n26858, ZN => 
                           n27687);
   U2885 : OAI211_X2 port map( C1 => n14690, C2 => n14689, A => n14688, B => 
                           n14687, ZN => n16238);
   U24 : MUX2_X2 port map( A => n20111, B => n20110, S => n20323, Z => n20898);
   U4355 : CLKBUF_X3 port map( A => n9313, Z => n9997);
   U362 : BUF_X1 port map( A => n18492, Z => n28632);
   U1732 : BUF_X2 port map( A => n25059, Z => n365);
   U1984 : BUF_X1 port map( A => n13595, Z => n14372);
   U26381 : AOI22_X2 port map( A1 => n26178, A2 => n26455, B1 => n25416, B2 => 
                           n25415, ZN => n26830);
   U22103 : XNOR2_X2 port map( A => n18873, B => n18872, ZN => n20157);
   U27041 : NAND2_X2 port map( A1 => n28712, A2 => n4242, ZN => n22888);
   U22730 : INV_X1 port map( A => n19787, ZN => n20635);
   U1124 : BUF_X1 port map( A => n24739, Z => n29050);
   U3086 : MUX2_X2 port map( A => n12040, B => n12039, S => n375, Z => n13171);
   U9491 : AOI21_X2 port map( B1 => n23079, B2 => n23080, A => n6580, ZN => 
                           n23994);
   U11723 : NAND2_X2 port map( A1 => n2314, A2 => n17122, ZN => n17846);
   U1142 : OAI21_X2 port map( B1 => n18844, B2 => n18843, A => n18842, ZN => 
                           n20816);
   U2816 : BUF_X1 port map( A => n17098, Z => n17101);
   U1407 : AND2_X2 port map( A1 => n23719, A2 => n23718, ZN => n24517);
   U10604 : XNOR2_X2 port map( A => n7572, B => n7573, ZN => n11146);
   U22633 : INV_X1 port map( A => n19938, ZN => n20281);
   U12822 : NAND3_X2 port map( A1 => n13676, A2 => n13675, A3 => n5519, ZN => 
                           n15388);
   U943 : OAI211_X2 port map( C1 => n6785, C2 => n7618, A => n3490, B => n3489,
                           ZN => n329);
   U1869 : INV_X1 port map( A => n6309, ZN => n24729);
   U10708 : OR2_X1 port map( A1 => n7707, A2 => n371, ZN => n4160);
   U1456 : BUF_X2 port map( A => n26507, Z => n27084);
   U12305 : BUF_X1 port map( A => n23700, Z => n28428);
   U182 : AND3_X2 port map( A1 => n2072, A2 => n3474, A3 => n3475, ZN => n22542
                           );
   U7564 : NAND2_X2 port map( A1 => n2552, A2 => n26844, ZN => n27827);
   U14609 : INV_X1 port map( A => n7072, ZN => n7886);
   U4305 : AOI21_X1 port map( B1 => n20707, B2 => n20706, A => n20705, ZN => 
                           n22798);
   U6191 : NAND3_X2 port map( A1 => n23895, A2 => n2265, A3 => n2266, ZN => 
                           n25532);
   U14436 : NOR2_X1 port map( A1 => n4466, A2 => n4465, ZN => n22661);
   U5145 : AND3_X2 port map( A1 => n1553, A2 => n1554, A3 => n5428, ZN => 
                           n18263);
   U2566 : AND4_X2 port map( A1 => n2177, A2 => n2179, A3 => n2082, A4 => n2182
                           , ZN => n21311);
   U2871 : AOI22_X2 port map( A1 => n14820, A2 => n14819, B1 => n15444, B2 => 
                           n14818, ZN => n16605);
   U676 : NAND2_X2 port map( A1 => n20037, A2 => n3136, ZN => n22023);
   U6988 : INV_X2 port map( A => n20225, ZN => n20500);
   U21720 : XNOR2_X2 port map( A => n18385, B => n18386, ZN => n20290);
   U1715 : BUF_X2 port map( A => n20375, Z => n351);
   U5161 : NAND3_X2 port map( A1 => n8783, A2 => n9006, A3 => n1566, ZN => 
                           n9716);
   U6164 : MUX2_X1 port map( A => n23548, B => n23547, S => n24772, Z => n23549
                           );
   U1833 : CLKBUF_X1 port map( A => Key(5), Z => n3219);
   U1226 : CLKBUF_X1 port map( A => Key(100), Z => n29247);
   U1814 : CLKBUF_X1 port map( A => Key(143), Z => n3049);
   U51 : CLKBUF_X1 port map( A => Key(183), Z => n3722);
   U2113 : CLKBUF_X1 port map( A => Key(102), Z => n26665);
   U1832 : CLKBUF_X1 port map( A => Key(6), Z => n3087);
   U14531 : XNOR2_X1 port map( A => Key(55), B => Plaintext(55), ZN => n7507);
   U1230 : CLKBUF_X1 port map( A => Key(0), Z => n1215);
   U5760 : XNOR2_X1 port map( A => Key(54), B => Plaintext(54), ZN => n7514);
   U1235 : CLKBUF_X1 port map( A => Key(175), Z => n3062);
   U3446 : XNOR2_X1 port map( A => Key(174), B => Plaintext(174), ZN => n7071);
   U14670 : XNOR2_X1 port map( A => Key(9), B => Plaintext(9), ZN => n7320);
   U14450 : XNOR2_X1 port map( A => Key(98), B => Plaintext(98), ZN => n7363);
   U14418 : XNOR2_X1 port map( A => Key(112), B => Plaintext(112), ZN => n8213)
                           ;
   U933 : XNOR2_X1 port map( A => Key(182), B => Plaintext(182), ZN => n7092);
   U675 : XNOR2_X1 port map( A => n7098, B => Key(17), ZN => n7759);
   U16341 : INV_X1 port map( A => n1196, ZN => n24906);
   U247 : XNOR2_X1 port map( A => n6972, B => Key(102), ZN => n8232);
   U14590 : XNOR2_X1 port map( A => n7057, B => Key(166), ZN => n7999);
   U14568 : XNOR2_X1 port map( A => n7045, B => Key(157), ZN => n7965);
   U14598 : XNOR2_X1 port map( A => n7062, B => Key(162), ZN => n7992);
   U14699 : XNOR2_X1 port map( A => n7128, B => Key(46), ZN => n8131);
   U14469 : XNOR2_X1 port map( A => n6995, B => Key(120), ZN => n7628);
   U132 : BUF_X1 port map( A => n7110, Z => n7898);
   U14542 : XNOR2_X1 port map( A => n7028, B => Key(64), ZN => n7521);
   U3414 : BUF_X1 port map( A => n8290, Z => n7915);
   U2413 : XNOR2_X1 port map( A => n7016, B => Key(88), ZN => n7837);
   U3403 : BUF_X1 port map( A => n7404, Z => n7976);
   U781 : OR2_X1 port map( A1 => n7324, A2 => n7325, ZN => n8579);
   U694 : NAND3_X1 port map( A1 => n7951, A2 => n7950, A3 => n117, ZN => n9107)
                           ;
   U4546 : OR2_X1 port map( A1 => n8026, A2 => n8025, ZN => n8899);
   U2453 : MUX2_X1 port map( A => n7762, B => n7761, S => n7760, Z => n7765);
   U1377 : OR2_X1 port map( A1 => n7944, A2 => n7945, ZN => n8914);
   U4183 : NAND2_X1 port map( A1 => n7772, A2 => n3183, ZN => n8351);
   U680 : OAI21_X1 port map( B1 => n7152, B2 => n8148, A => n7151, ZN => n9247)
                           ;
   U3388 : OR2_X1 port map( A1 => n7429, A2 => n7428, ZN => n9075);
   U14453 : OAI21_X1 port map( B1 => n6983, B2 => n6982, A => n6981, ZN => 
                           n9229);
   U665 : NAND3_X1 port map( A1 => n3185, A2 => n2221, A3 => n2222, ZN => n8502
                           );
   U4505 : NAND3_X1 port map( A1 => n6802, A2 => n6801, A3 => n7593, ZN => 
                           n8414);
   U15204 : OAI211_X1 port map( C1 => n7732, C2 => n7733, A => n7731, B => 
                           n7730, ZN => n9186);
   U3348 : NAND2_X1 port map( A1 => n8152, A2 => n1512, ZN => n8983);
   U1167 : OR2_X1 port map( A1 => n7599, A2 => n7598, ZN => n8788);
   U1065 : OR2_X1 port map( A1 => n7713, A2 => n7712, ZN => n9029);
   U1442 : OAI211_X1 port map( C1 => n7673, C2 => n8275, A => n7672, B => n7671
                           , ZN => n8996);
   U1349 : OR2_X1 port map( A1 => n2506, A2 => n7131, ZN => n9041);
   U1586 : NOR2_X1 port map( A1 => n3445, A2 => n155, ZN => n28606);
   U1549 : BUF_X1 port map( A => n7726, Z => n9188);
   U861 : OR2_X1 port map( A1 => n732, A2 => n7739, ZN => n8782);
   U410 : AND2_X1 port map( A1 => n7904, A2 => n7903, ZN => n8635);
   U3343 : NAND2_X1 port map( A1 => n7972, A2 => n7973, ZN => n8665);
   U159 : MUX2_X1 port map( A => n7217, B => n7214, S => n29673, Z => n9228);
   U8448 : NAND2_X1 port map( A1 => n2424, A2 => n2059, ZN => n8719);
   U654 : NAND2_X1 port map( A1 => n6199, A2 => n7242, ZN => n8608);
   U1098 : BUF_X1 port map( A => n7175, Z => n8537);
   U3333 : AND2_X1 port map( A1 => n1042, A2 => n7195, ZN => n8685);
   U3366 : AND2_X1 port map( A1 => n7558, A2 => n7559, ZN => n8872);
   U8480 : OR2_X1 port map( A1 => n8785, A2 => n8414, ZN => n8438);
   U6238 : OR2_X1 port map( A1 => n9063, A2 => n9062, ZN => n5536);
   U86 : OR2_X1 port map( A1 => n8943, A2 => n8944, ZN => n2168);
   U910 : NAND3_X1 port map( A1 => n8489, A2 => n6318, A3 => n6317, ZN => 
                           n10386);
   U8663 : MUX2_X1 port map( A => n8437, B => n8436, S => n9210, Z => n9735);
   U15739 : OR2_X1 port map( A1 => n8646, A2 => n8762, ZN => n10406);
   U834 : OR2_X1 port map( A1 => n9011, A2 => n9010, ZN => n9512);
   U533 : OR2_X1 port map( A1 => n9341, A2 => n2229, ZN => n9979);
   U868 : OR2_X1 port map( A1 => n8895, A2 => n8894, ZN => n9824);
   U136 : AND3_X1 port map( A1 => n2247, A2 => n3755, A3 => n28882, ZN => n9648
                           );
   U5888 : OR2_X1 port map( A1 => n127, A2 => n8713, ZN => n9575);
   U556 : NAND2_X1 port map( A1 => n9415, A2 => n9414, ZN => n10392);
   U5623 : MUX2_X1 port map( A => n8442, B => n8441, S => n8440, Z => n1920);
   U15283 : OR2_X1 port map( A1 => n7956, A2 => n7955, ZN => n10357);
   U3276 : NAND3_X1 port map( A1 => n3182, A2 => n8841, A3 => n3181, ZN => 
                           n10272);
   U9258 : NAND2_X1 port map( A1 => n8618, A2 => n2907, ZN => n10043);
   U3291 : OR2_X1 port map( A1 => n5308, A2 => n8645, ZN => n10184);
   U2564 : OAI21_X1 port map( B1 => n8662, B2 => n5677, A => n5673, ZN => 
                           n10134);
   U740 : OAI211_X1 port map( C1 => n9227, C2 => n9228, A => n9225, B => n9226,
                           ZN => n10335);
   U15807 : XNOR2_X1 port map( A => n9295, B => n26656, ZN => n8772);
   U4121 : OAI21_X1 port map( B1 => n8356, B2 => n8431, A => n971, ZN => n10282
                           );
   U5645 : XNOR2_X1 port map( A => n10321, B => n2845, ZN => n9770);
   U3267 : NAND2_X1 port map( A1 => n2334, A2 => n2336, ZN => n10294);
   U3274 : NAND3_X1 port map( A1 => n8387, A2 => n8386, A3 => n8385, ZN => 
                           n10074);
   U10996 : NAND2_X1 port map( A1 => n3781, A2 => n3780, ZN => n10208);
   U1448 : OAI21_X1 port map( B1 => n29147, B2 => n8198, A => n8197, ZN => 
                           n10060);
   U2143 : XNOR2_X1 port map( A => n9908, B => n10021, ZN => n10319);
   U516 : XNOR2_X1 port map( A => n9916, B => n9698, ZN => n10342);
   U16058 : XNOR2_X1 port map( A => n9280, B => n9279, ZN => n10705);
   U2333 : XNOR2_X1 port map( A => n5401, B => n5400, ZN => n11135);
   U16011 : XNOR2_X1 port map( A => n9217, B => n9216, ZN => n11349);
   U1667 : XNOR2_X1 port map( A => n9651, B => n9652, ZN => n11267);
   U3220 : XNOR2_X1 port map( A => n9159, B => n9158, ZN => n10847);
   U451 : XNOR2_X1 port map( A => n9898, B => n9897, ZN => n11120);
   U3217 : XNOR2_X1 port map( A => n10378, B => n10377, ZN => n11281);
   U269 : BUF_X1 port map( A => n10096, Z => n29150);
   U3189 : XNOR2_X1 port map( A => n3437, B => n5860, ZN => n10958);
   U217 : XNOR2_X1 port map( A => n9792, B => n9791, ZN => n10995);
   U1338 : XNOR2_X1 port map( A => n5562, B => n10286, ZN => n11290);
   U9884 : OR2_X1 port map( A1 => n11237, A2 => n11010, ZN => n11234);
   U669 : XNOR2_X1 port map( A => n4590, B => n4589, ZN => n11165);
   U3200 : XNOR2_X1 port map( A => n9361, B => n9360, ZN => n10962);
   U1000 : BUF_X2 port map( A => n11064, Z => n11069);
   U198 : XNOR2_X1 port map( A => n9328, B => n9327, ZN => n10913);
   U7569 : BUF_X1 port map( A => n10097, Z => n11114);
   U2665 : NOR2_X1 port map( A1 => n11199, A2 => n28207, ZN => n10749);
   U3201 : BUF_X1 port map( A => n10855, Z => n11308);
   U17250 : OAI211_X1 port map( C1 => n10989, C2 => n10988, A => n10987, B => 
                           n10986, ZN => n12249);
   U3164 : MUX2_X1 port map( A => n10631, B => n9848, S => n10783, Z => n9865);
   U17119 : OR2_X1 port map( A1 => n10737, A2 => n10736, ZN => n11426);
   U860 : NAND2_X1 port map( A1 => n3165, A2 => n10092, ZN => n10905);
   U6206 : NAND3_X1 port map( A1 => n1080, A2 => n10633, A3 => n10634, ZN => 
                           n12218);
   U3158 : AOI22_X1 port map( A1 => n11224, A2 => n11223, B1 => n11222, B2 => 
                           n11221, ZN => n12320);
   U2006 : OAI211_X1 port map( C1 => n10822, C2 => n28208, A => n10824, B => 
                           n6885, ZN => n12146);
   U4145 : NAND2_X1 port map( A1 => n1214, A2 => n3018, ZN => n12058);
   U1587 : AND3_X1 port map( A1 => n10217, A2 => n10216, A3 => n10215, ZN => 
                           n11824);
   U4024 : AND2_X1 port map( A1 => n898, A2 => n1146, ZN => n12271);
   U2140 : OR2_X1 port map( A1 => n10762, A2 => n6918, ZN => n11405);
   U838 : OR2_X1 port map( A1 => n10654, A2 => n10653, ZN => n1986);
   U2875 : NOR2_X1 port map( A1 => n11636, A2 => n11633, ZN => n29139);
   U4349 : OAI21_X1 port map( B1 => n4815, B2 => n4325, A => n4328, ZN => 
                           n12156);
   U1487 : AND3_X1 port map( A1 => n3815, A2 => n4800, A3 => n3814, ZN => 
                           n12111);
   U745 : OR2_X1 port map( A1 => n11660, A2 => n10895, ZN => n11377);
   U717 : NAND3_X1 port map( A1 => n4710, A2 => n10511, A3 => n6271, ZN => 
                           n11500);
   U229 : NAND2_X1 port map( A1 => n28282, A2 => n28283, ZN => n6482);
   U7444 : NAND3_X1 port map( A1 => n3373, A2 => n8623, A3 => n8622, ZN => 
                           n12203);
   U13632 : INV_X1 port map( A => n11794, ZN => n10717);
   U1797 : AND3_X1 port map( A1 => n2943, A2 => n11102, A3 => n1945, ZN => 
                           n12516);
   U3112 : BUF_X1 port map( A => n11390, Z => n11851);
   U5451 : NAND2_X1 port map( A1 => n1786, A2 => n1787, ZN => n12251);
   U187 : AND2_X1 port map( A1 => n11495, A2 => n11493, ZN => n569);
   U55 : BUF_X1 port map( A => n11878, Z => n287);
   U17867 : NAND2_X1 port map( A1 => n12198, A2 => n12189, ZN => n12131);
   U5971 : BUF_X1 port map( A => n11859, Z => n11943);
   U7578 : BUF_X1 port map( A => n12307, Z => n4197);
   U4540 : NAND2_X1 port map( A1 => n10604, A2 => n3322, ZN => n12356);
   U6298 : INV_X1 port map( A => n12307, ZN => n12300);
   U11157 : OR2_X1 port map( A1 => n3910, A2 => n3908, ZN => n4341);
   U7445 : INV_X1 port map( A => n12203, ZN => n4844);
   U3125 : INV_X1 port map( A => n11058, ZN => n12267);
   U652 : BUF_X1 port map( A => n11505, Z => n12400);
   U3127 : BUF_X1 port map( A => n11419, Z => n11785);
   U16436 : BUF_X1 port map( A => n9692, Z => n12109);
   U5761 : NAND2_X1 port map( A1 => n11887, A2 => n11886, ZN => n12327);
   U6287 : OR2_X1 port map( A1 => n11622, A2 => n11194, ZN => n11580);
   U10185 : MUX2_X1 port map( A => n10118, B => n10117, S => n12507, Z => 
                           n13167);
   U10906 : NAND3_X1 port map( A1 => n11909, A2 => n28962, A3 => n28961, ZN => 
                           n13413);
   U1095 : NAND3_X1 port map( A1 => n11573, A2 => n11572, A3 => n3745, ZN => 
                           n13291);
   U1169 : AND2_X1 port map( A1 => n3795, A2 => n3794, ZN => n13493);
   U5628 : OAI211_X1 port map( C1 => n11485, C2 => n11484, A => n11483, B => 
                           n11612, ZN => n13244);
   U20964 : NOR2_X1 port map( A1 => n12185, A2 => n12184, ZN => n13261);
   U1190 : OAI211_X1 port map( C1 => n11711, C2 => n5169, A => n3688, B => 
                           n11414, ZN => n12723);
   U590 : OAI21_X1 port map( B1 => n12225, B2 => n12224, A => n12223, ZN => 
                           n13285);
   U12374 : AND2_X1 port map( A1 => n5096, A2 => n5095, ZN => n13236);
   U2954 : NAND2_X1 port map( A1 => n11475, A2 => n3592, ZN => n13018);
   U13713 : OAI21_X1 port map( B1 => n6481, B2 => n6478, A => n11721, ZN => 
                           n13067);
   U1265 : NAND2_X1 port map( A1 => n3566, A2 => n233, ZN => n13159);
   U3056 : XNOR2_X1 port map( A => n13166, B => n13219, ZN => n13522);
   U1307 : BUF_X1 port map( A => n12752, Z => n12783);
   U1100 : OAI21_X1 port map( B1 => n1401, B2 => n12431, A => n12430, ZN => 
                           n13369);
   U8956 : XNOR2_X1 port map( A => n13523, B => n1885, ZN => n12454);
   U1846 : NAND2_X1 port map( A1 => n10651, A2 => n10650, ZN => n12560);
   U759 : XNOR2_X1 port map( A => n12719, B => n12720, ZN => n13933);
   U3031 : XNOR2_X1 port map( A => n12970, B => n12969, ZN => n14091);
   U817 : XNOR2_X1 port map( A => n12476, B => n12477, ZN => n12480);
   U1288 : XNOR2_X1 port map( A => n12540, B => n12539, ZN => n14426);
   U18060 : XNOR2_X1 port map( A => n12463, B => n12464, ZN => n14217);
   U3034 : BUF_X1 port map( A => n13755, Z => n14475);
   U3036 : XNOR2_X1 port map( A => n12139, B => n12138, ZN => n14166);
   U3001 : XNOR2_X1 port map( A => n2962, B => n3110, ZN => n14435);
   U91 : BUF_X1 port map( A => n13749, Z => n14261);
   U3009 : XNOR2_X1 port map( A => n13065, B => n13064, ZN => n14351);
   U994 : XNOR2_X1 port map( A => n12984, B => n12983, ZN => n14358);
   U1308 : BUF_X1 port map( A => n13686, Z => n14415);
   U758 : XNOR2_X1 port map( A => n2173, B => n2171, ZN => n14376);
   U2978 : OAI21_X1 port map( B1 => n13696, B2 => n13656, A => n13655, ZN => 
                           n14743);
   U972 : OR2_X1 port map( A1 => n14042, A2 => n14041, ZN => n14600);
   U18988 : OAI21_X1 port map( B1 => n13696, B2 => n14325, A => n13695, ZN => 
                           n14115);
   U10527 : MUX2_X1 port map( A => n13165, B => n13164, S => n14328, Z => 
                           n15692);
   U23940 : NAND3_X1 port map( A1 => n1345, A2 => n14329, A3 => n1344, ZN => 
                           n15306);
   U751 : NOR2_X1 port map( A1 => n13665, A2 => n2373, ZN => n14514);
   U2961 : INV_X1 port map( A => n14115, ZN => n15138);
   U1361 : AND2_X1 port map( A1 => n13905, A2 => n13904, ZN => n14807);
   U28161 : NAND3_X1 port map( A1 => n28754, A2 => n1016, A3 => n28753, ZN => 
                           n14773);
   U3187 : INV_X1 port map( A => n14600, ZN => n14601);
   U2955 : AND2_X1 port map( A1 => n4163, A2 => n14277, ZN => n14763);
   U2973 : OR2_X1 port map( A1 => n14378, A2 => n14377, ZN => n15511);
   U1743 : AND3_X1 port map( A1 => n12758, A2 => n14471, A3 => n28936, ZN => 
                           n15101);
   U225 : OR2_X1 port map( A1 => n6446, A2 => n13590, ZN => n15400);
   U2969 : AOI22_X1 port map( A1 => n13746, A2 => n13745, B1 => n14076, B2 => 
                           n4376, ZN => n15383);
   U1642 : OAI211_X1 port map( C1 => n14009, C2 => n5404, A => n6614, B => 
                           n6613, ZN => n14826);
   U226 : AND2_X1 port map( A1 => n14830, A2 => n14834, ZN => n15292);
   U5803 : NAND2_X1 port map( A1 => n13705, A2 => n3435, ZN => n15250);
   U9541 : NAND2_X1 port map( A1 => n1627, A2 => n14472, ZN => n15491);
   U11705 : OR2_X1 port map( A1 => n13979, A2 => n14743, ZN => n14744);
   U18975 : NOR2_X1 port map( A1 => n14990, A2 => n14989, ZN => n15395);
   U1162 : AOI21_X1 port map( B1 => n5823, B2 => n293, A => n5820, ZN => n14986
                           );
   U6391 : OAI21_X1 port map( B1 => n5834, B2 => n13336, A => n28866, ZN => 
                           n14882);
   U3081 : NOR2_X1 port map( A1 => n13596, A2 => n13597, ZN => n13638);
   U876 : NAND2_X1 port map( A1 => n2562, A2 => n2561, ZN => n15174);
   U6901 : INV_X2 port map( A => n15311, ZN => n14851);
   U2915 : BUF_X1 port map( A => n14518, Z => n15036);
   U895 : INV_X1 port map( A => n14518, ZN => n3827);
   U4766 : INV_X1 port map( A => n14575, ZN => n15105);
   U3120 : NOR2_X1 port map( A1 => n3208, A2 => n15387, ZN => n14994);
   U15633 : OAI211_X1 port map( C1 => n14968, C2 => n14961, A => n13787, B => 
                           n13786, ZN => n16284);
   U1492 : OR2_X1 port map( A1 => n15495, A2 => n15491, ZN => n264);
   U1710 : AND3_X1 port map( A1 => n29173, A2 => n29172, A3 => n29171, ZN => 
                           n16634);
   U537 : NAND2_X1 port map( A1 => n88, A2 => n14794, ZN => n16509);
   U892 : AND4_X1 port map( A1 => n5052, A2 => n5051, A3 => n14919, A4 => n5050
                           , ZN => n15977);
   U2881 : NOR2_X1 port map( A1 => n14828, A2 => n14829, ZN => n16526);
   U621 : NAND2_X1 port map( A1 => n3682, A2 => n15364, ZN => n16230);
   U9696 : NAND2_X1 port map( A1 => n15220, A2 => n15221, ZN => n15642);
   U4770 : NAND2_X1 port map( A1 => n15270, A2 => n1243, ZN => n16242);
   U3900 : AOI21_X1 port map( B1 => n13978, B2 => n15014, A => n13977, ZN => 
                           n16146);
   U2877 : OR2_X1 port map( A1 => n4720, A2 => n4718, ZN => n15618);
   U1688 : AND2_X1 port map( A1 => n14626, A2 => n14627, ZN => n16043);
   U1264 : OR2_X1 port map( A1 => n15149, A2 => n15148, ZN => n16051);
   U1690 : NAND3_X1 port map( A1 => n28837, A2 => n15240, A3 => n2885, ZN => 
                           n16105);
   U10506 : NAND3_X1 port map( A1 => n4417, A2 => n3550, A3 => n14599, ZN => 
                           n16233);
   U509 : NAND2_X1 port map( A1 => n82, A2 => n1964, ZN => n16589);
   U1683 : XNOR2_X1 port map( A => n15846, B => n15845, ZN => n16908);
   U1960 : XNOR2_X1 port map( A => n14720, B => n14721, ZN => n17393);
   U2823 : XNOR2_X1 port map( A => n16573, B => n16572, ZN => n17516);
   U67 : BUF_X1 port map( A => n15551, Z => n17348);
   U1243 : XNOR2_X1 port map( A => n15684, B => n15683, ZN => n17548);
   U19897 : XNOR2_X1 port map( A => n15429, B => n15428, ZN => n17411);
   U2839 : XNOR2_X1 port map( A => n15913, B => n15912, ZN => n17572);
   U10567 : XNOR2_X1 port map( A => n16515, B => n16516, ZN => n17450);
   U595 : XNOR2_X1 port map( A => n15776, B => n15775, ZN => n17543);
   U713 : XNOR2_X1 port map( A => n16195, B => n16194, ZN => n16888);
   U1650 : BUF_X1 port map( A => n17466, Z => n28800);
   U10409 : XNOR2_X1 port map( A => n6502, B => n16380, ZN => n17375);
   U2810 : INV_X1 port map( A => n4316, ZN => n17229);
   U1273 : BUF_X1 port map( A => n16137, Z => n17262);
   U3149 : BUF_X1 port map( A => n16837, Z => n17562);
   U10593 : MUX2_X1 port map( A => n16905, B => n17706, S => n4156, Z => n18268
                           );
   U3287 : OAI21_X1 port map( B1 => n17194, B2 => n5260, A => n17193, ZN => 
                           n18121);
   U26675 : AOI22_X1 port map( A1 => n3169, A2 => n3172, B1 => n16725, B2 => 
                           n16660, ZN => n16663);
   U616 : MUX2_X1 port map( A => n16886, B => n16885, S => n17158, Z => n18516)
                           ;
   U2769 : INV_X1 port map( A => n19562, ZN => n527);
   U4223 : OR2_X1 port map( A1 => n16688, A2 => n16689, ZN => n18342);
   U1844 : NAND2_X1 port map( A1 => n14507, A2 => n17009, ZN => n18306);
   U2731 : AND3_X1 port map( A1 => n16979, A2 => n6538, A3 => n16978, ZN => 
                           n18081);
   U1614 : OAI21_X1 port map( B1 => n17161, B2 => n17386, A => n28851, ZN => 
                           n18376);
   U473 : NAND3_X1 port map( A1 => n4702, A2 => n4700, A3 => n4699, ZN => 
                           n18276);
   U6121 : AND3_X1 port map( A1 => n3811, A2 => n3812, A3 => n5620, ZN => 
                           n18356);
   U1943 : OR2_X1 port map( A1 => n17144, A2 => n17145, ZN => n5383);
   U4793 : NAND2_X1 port map( A1 => n1264, A2 => n16692, ZN => n18344);
   U457 : NAND2_X1 port map( A1 => n5250, A2 => n783, ZN => n17969);
   U56 : OR2_X1 port map( A1 => n17306, A2 => n17307, ZN => n17620);
   U1242 : BUF_X1 port map( A => n17826, Z => n18160);
   U27347 : NAND2_X1 port map( A1 => n6175, A2 => n6176, ZN => n18527);
   U27746 : NAND2_X1 port map( A1 => n28728, A2 => n1367, ZN => n16985);
   U2719 : AND2_X1 port map( A1 => n2702, A2 => n4280, ZN => n18260);
   U1619 : AND2_X1 port map( A1 => n29240, A2 => n4040, ZN => n18248);
   U1753 : BUF_X1 port map( A => n18522, Z => n373);
   U9048 : AND2_X1 port map( A1 => n5326, A2 => n5327, ZN => n18286);
   U6979 : NOR2_X1 port map( A1 => n18298, A2 => n18063, ZN => n2791);
   U78 : INV_X1 port map( A => n17207, ZN => n17835);
   U100 : OR2_X1 port map( A1 => n18304, A2 => n17679, ZN => n18012);
   U21364 : AOI21_X1 port map( B1 => n16898, B2 => n18276, A => n18279, ZN => 
                           n18206);
   U2677 : NAND2_X1 port map( A1 => n16901, A2 => n16900, ZN => n19111);
   U884 : OAI211_X1 port map( C1 => n18163, C2 => n18164, A => n18162, B => 
                           n18161, ZN => n19678);
   U2681 : OAI21_X1 port map( B1 => n6326, B2 => n18454, A => n18453, ZN => 
                           n19220);
   U351 : NAND2_X1 port map( A1 => n40, A2 => n18287, ZN => n19695);
   U1220 : NAND2_X1 port map( A1 => n2214, A2 => n2212, ZN => n18638);
   U2643 : NAND2_X1 port map( A1 => n2566, A2 => n17841, ZN => n19704);
   U1760 : NAND2_X1 port map( A1 => n28733, A2 => n17648, ZN => n19108);
   U1713 : OAI21_X1 port map( B1 => n18359, B2 => n18360, A => n18358, ZN => 
                           n18798);
   U1051 : AND2_X1 port map( A1 => n1784, A2 => n17981, ZN => n18959);
   U21921 : XNOR2_X1 port map( A => n19111, B => n2889, ZN => n18671);
   U21441 : XNOR2_X1 port map( A => n28447, B => n19706, ZN => n19285);
   U6079 : INV_X1 port map( A => n18867, ZN => n19087);
   U4051 : NAND2_X1 port map( A1 => n916, A2 => n913, ZN => n19697);
   U22429 : XNOR2_X1 port map( A => n19312, B => n19311, ZN => n20626);
   U9673 : XNOR2_X1 port map( A => n19264, B => n3111, ZN => n20601);
   U1341 : XNOR2_X1 port map( A => n19684, B => n19683, ZN => n20607);
   U468 : XNOR2_X1 port map( A => n19722, B => n19721, ZN => n20614);
   U303 : XNOR2_X1 port map( A => n19494, B => n19493, ZN => n20444);
   U9769 : XNOR2_X1 port map( A => n18771, B => n19455, ZN => n20063);
   U1922 : BUF_X1 port map( A => n19995, Z => n20478);
   U773 : BUF_X1 port map( A => n28140, Z => n28779);
   U273 : BUF_X1 port map( A => n20224, Z => n297);
   U8041 : BUF_X1 port map( A => n17954, Z => n20311);
   U4723 : BUF_X1 port map( A => n19928, Z => n20449);
   U3608 : NOR3_X1 port map( A1 => n20545, A2 => n20546, A3 => n20547, ZN => 
                           n21585);
   U690 : MUX2_X1 port map( A => n20543, B => n20542, S => n20541, Z => n21586)
                           ;
   U3516 : AND2_X1 port map( A1 => n5302, A2 => n5305, ZN => n21047);
   U534 : OAI21_X1 port map( B1 => n20411, B2 => n20410, A => n20409, ZN => 
                           n21503);
   U25346 : OAI21_X1 port map( B1 => n18833, B2 => n20097, A => n28326, ZN => 
                           n20878);
   U7131 : BUF_X1 port map( A => n20722, Z => n21598);
   U23326 : BUF_X2 port map( A => n20782, Z => n21551);
   U252 : OR2_X1 port map( A1 => n20254, A2 => n28295, ZN => n21014);
   U2553 : AND2_X1 port map( A1 => n2747, A2 => n5376, ZN => n21534);
   U593 : AND3_X1 port map( A1 => n20566, A2 => n20564, A3 => n20565, ZN => 
                           n5684);
   U1916 : MUX2_X1 port map( A => n19742, B => n19741, S => n19740, Z => n22140
                           );
   U4621 : NAND3_X1 port map( A1 => n19853, A2 => n19854, A3 => n19852, ZN => 
                           n21574);
   U1910 : OR2_X1 port map( A1 => n19998, A2 => n6028, ZN => n21171);
   U419 : NOR2_X1 port map( A1 => n1099, A2 => n1335, ZN => n20783);
   U19739 : OR2_X1 port map( A1 => n28662, A2 => n28661, ZN => n28584);
   U1913 : NAND3_X1 port map( A1 => n20004, A2 => n6137, A3 => n20003, ZN => 
                           n21408);
   U2484 : OR2_X1 port map( A1 => n1327, A2 => n21749, ZN => n5975);
   U22532 : NOR2_X1 port map( A1 => n19459, A2 => n19458, ZN => n21717);
   U1773 : OR2_X1 port map( A1 => n21645, A2 => n497, ZN => n21237);
   U2483 : OAI21_X1 port map( B1 => n21685, B2 => n21684, A => n21683, ZN => 
                           n22221);
   U10007 : AOI21_X1 port map( B1 => n21405, B2 => n21404, A => n21403, ZN => 
                           n22411);
   U7087 : MUX2_X1 port map( A => n18549, B => n18548, S => n28440, Z => n21825
                           );
   U588 : OAI21_X1 port map( B1 => n20364, B2 => n20365, A => n20363, ZN => 
                           n22472);
   U10079 : NAND2_X1 port map( A1 => n21201, A2 => n3288, ZN => n22854);
   U2474 : AND2_X1 port map( A1 => n1084, A2 => n1083, ZN => n22414);
   U2475 : AND3_X1 port map( A1 => n6694, A2 => n6695, A3 => n6696, ZN => 
                           n22437);
   U761 : AND4_X1 port map( A1 => n21486, A2 => n21488, A3 => n6369, A4 => 
                           n21487, ZN => n22337);
   U927 : NAND3_X1 port map( A1 => n6350, A2 => n21444, A3 => n6349, ZN => 
                           n22479);
   U1423 : AOI21_X1 port map( B1 => n21214, B2 => n21213, A => n872, ZN => 
                           n22783);
   U218 : NOR2_X1 port map( A1 => n18788, A2 => n18787, ZN => n2805);
   U1585 : NAND2_X1 port map( A1 => n21285, A2 => n21284, ZN => n22501);
   U1538 : AND3_X1 port map( A1 => n6041, A2 => n6040, A3 => n6039, ZN => 
                           n22710);
   U5415 : OAI211_X1 port map( C1 => n20530, C2 => n20531, A => n20529, B => 
                           n20528, ZN => n22750);
   U1901 : NAND2_X1 port map( A1 => n2991, A2 => n2988, ZN => n22525);
   U145 : XNOR2_X1 port map( A => n21948, B => n274, ZN => n23606);
   U1178 : XNOR2_X1 port map( A => n4760, B => n21803, ZN => n23769);
   U3913 : XNOR2_X1 port map( A => n22385, B => n22384, ZN => n23566);
   U908 : XNOR2_X1 port map( A => n21968, B => n21969, ZN => n23607);
   U1706 : XNOR2_X1 port map( A => n22005, B => n22004, ZN => n2141);
   U13805 : XNOR2_X1 port map( A => n22795, B => n22794, ZN => n23416);
   U13034 : BUF_X1 port map( A => n23297, Z => n29020);
   U1513 : BUF_X1 port map( A => n22946, Z => n23741);
   U2400 : BUF_X1 port map( A => n23233, Z => n23714);
   U224 : BUF_X1 port map( A => n23280, Z => n28418);
   U1677 : OR2_X1 port map( A1 => n23088, A2 => n23087, ZN => n24378);
   U901 : NAND2_X1 port map( A1 => n22176, A2 => n22175, ZN => n24582);
   U777 : OR2_X1 port map( A1 => n5346, A2 => n23208, ZN => n138);
   U13361 : OAI21_X1 port map( B1 => n22129, B2 => n28474, A => n22128, ZN => 
                           n29026);
   U9865 : NAND3_X1 port map( A1 => n6764, A2 => n6763, A3 => n1965, ZN => 
                           n24391);
   U2351 : OR2_X1 port map( A1 => n2835, A2 => n2076, ZN => n24800);
   U271 : NAND2_X1 port map( A1 => n1446, A2 => n28695, ZN => n24081);
   U1334 : OAI211_X1 port map( C1 => n23035, C2 => n23034, A => n4935, B => 
                           n4934, ZN => n29043);
   U1662 : NAND2_X1 port map( A1 => n5456, A2 => n28224, ZN => n24602);
   U9787 : AND2_X1 port map( A1 => n2818, A2 => n2817, ZN => n24420);
   U26111 : AND2_X1 port map( A1 => n23730, A2 => n23731, ZN => n24520);
   U14362 : BUF_X1 port map( A => n23932, Z => n24597);
   U435 : BUF_X1 port map( A => n25908, Z => n28769);
   U14356 : AOI21_X1 port map( B1 => n23975, B2 => n23974, A => n23973, ZN => 
                           n25187);
   U1389 : AND2_X1 port map( A1 => n964, A2 => n967, ZN => n26100);
   U207 : OAI211_X1 port map( C1 => n4749, C2 => n4748, A => n24147, B => 
                           n24148, ZN => n26093);
   U1473 : XNOR2_X1 port map( A => n25111, B => n25110, ZN => n26800);
   U2260 : XNOR2_X1 port map( A => n25707, B => n25706, ZN => n27069);
   U6580 : AND2_X1 port map( A1 => n26865, A2 => n27110, ZN => n27152);
   U27064 : MUX2_X1 port map( A => n26351, B => n26350, S => n27701, Z => 
                           n26355);
   U26887 : AND2_X1 port map( A1 => n26128, A2 => n27161, ZN => n27707);
   U10327 : OAI21_X1 port map( B1 => n26365, B2 => n28948, A => n26363, ZN => 
                           n27632);
   U1221 : NAND2_X1 port map( A1 => n2966, A2 => n26564, ZN => n27496);
   U16604 : NAND2_X1 port map( A1 => n26243, A2 => n26244, ZN => n28543);
   U1238 : CLKBUF_X1 port map( A => Key(153), Z => n3537);
   U14692 : XNOR2_X1 port map( A => Key(43), B => Plaintext(43), ZN => n8048);
   U4207 : BUF_X1 port map( A => Key(161), Z => n3787);
   U2473 : BUF_X1 port map( A => Key(134), Z => n28693);
   U3497 : BUF_X1 port map( A => Key(70), Z => n3036);
   U2063 : BUF_X1 port map( A => Key(79), Z => n26214);
   U1829 : BUF_X1 port map( A => Key(131), Z => n3491);
   U1604 : BUF_X2 port map( A => Key(186), Z => n3015);
   U4208 : CLKBUF_X1 port map( A => Key(162), Z => n3196);
   U8405 : OR2_X1 port map( A1 => n2406, A2 => n6999, ZN => n9045);
   U1205 : OR2_X1 port map( A1 => n7339, A2 => n7338, ZN => n9144);
   U2227 : NOR2_X1 port map( A1 => n7661, A2 => n28857, ZN => n8995);
   U3387 : INV_X1 port map( A => n29303, ZN => n610);
   U11936 : OR2_X1 port map( A1 => n4671, A2 => n7319, ZN => n8327);
   U157 : NAND2_X1 port map( A1 => n3179, A2 => n7617, ZN => n9196);
   U124 : BUF_X1 port map( A => n9363, Z => n284);
   U3325 : INV_X1 port map( A => n8384, ZN => n8739);
   U2379 : NAND2_X1 port map( A1 => n28751, A2 => n2480, ZN => n8741);
   U14462 : NAND2_X1 port map( A1 => n7482, A2 => n7483, ZN => n28500);
   U5458 : OAI211_X1 port map( C1 => n1792, C2 => n1794, A => n1789, B => n2844
                           , ZN => n9696);
   U1367 : OAI211_X1 port map( C1 => n9169, C2 => n8250, A => n8249, B => n8248
                           , ZN => n10178);
   U517 : OAI21_X1 port map( B1 => n2713, B2 => n8339, A => n2712, ZN => n9698)
                           ;
   U643 : NAND2_X1 port map( A1 => n5867, A2 => n3678, ZN => n9991);
   U3254 : NAND2_X1 port map( A1 => n8255, A2 => n8254, ZN => n10059);
   U3192 : XNOR2_X1 port map( A => n9912, B => n9911, ZN => n11124);
   U1800 : INV_X1 port map( A => n10993, ZN => n3454);
   U1660 : BUF_X1 port map( A => n11226, Z => n333);
   U2018 : INV_X1 port map( A => n11086, ZN => n433);
   U2013 : BUF_X1 port map( A => n10528, Z => n11261);
   U1565 : INV_X2 port map( A => n11140, ZN => n3862);
   U688 : BUF_X1 port map( A => n9344, Z => n10916);
   U8343 : OAI22_X1 port map( A1 => n10881, A2 => n10880, B1 => n5063, B2 => 
                           n10641, ZN => n12166);
   U16995 : MUX2_X1 port map( A => n10565, B => n10564, S => n11196, Z => 
                           n10567);
   U3545 : NAND2_X1 port map( A1 => n2351, A2 => n3807, ZN => n11782);
   U9362 : AND2_X1 port map( A1 => n28930, A2 => n28928, ZN => n11730);
   U1194 : INV_X2 port map( A => n11500, ZN => n390);
   U1256 : NOR2_X1 port map( A1 => n11673, A2 => n11671, ZN => n11677);
   U3775 : INV_X1 port map( A => n12233, ZN => n776);
   U3084 : NAND3_X1 port map( A1 => n6550, A2 => n6551, A3 => n6549, ZN => 
                           n13461);
   U2183 : AND3_X1 port map( A1 => n3200, A2 => n3202, A3 => n2074, ZN => 
                           n12854);
   U8733 : NAND3_X1 port map( A1 => n6561, A2 => n10770, A3 => n2538, ZN => 
                           n13547);
   U5788 : BUF_X2 port map( A => n12954, Z => n12763);
   U1993 : NAND4_X1 port map( A1 => n12171, A2 => n12170, A3 => n12168, A4 => 
                           n12169, ZN => n13113);
   U1254 : NAND2_X1 port map( A1 => n2979, A2 => n12323, ZN => n13272);
   U18116 : XNOR2_X1 port map( A => n12521, B => n12919, ZN => n13434);
   U5993 : XNOR2_X1 port map( A => n12975, B => n12974, ZN => n14365);
   U1546 : INV_X1 port map( A => n15194, ZN => n28172);
   U1810 : INV_X1 port map( A => n13953, ZN => n28805);
   U1982 : AOI22_X1 port map( A1 => n14065, A2 => n14324, B1 => n14328, B2 => 
                           n14327, ZN => n13696);
   U1987 : INV_X2 port map( A => n14200, ZN => n427);
   U5809 : AOI21_X1 port map( B1 => n5796, B2 => n308, A => n14371, ZN => 
                           n14697);
   U19252 : AOI22_X1 port map( A1 => n14124, A2 => n14123, B1 => n308, B2 => 
                           n14121, ZN => n14153);
   U202 : AOI21_X1 port map( B1 => n13768, B2 => n13769, A => n15193, ZN => 
                           n14961);
   U949 : MUX2_X1 port map( A => n14595, B => n14594, S => n14593, Z => n14762)
                           ;
   U59 : AND2_X1 port map( A1 => n912, A2 => n14096, ZN => n14518);
   U25597 : NAND2_X1 port map( A1 => n14203, A2 => n28684, ZN => n15338);
   U350 : NAND2_X1 port map( A1 => n15346, A2 => n15344, ZN => n15222);
   U14278 : OR2_X1 port map( A1 => n14903, A2 => n14902, ZN => n15100);
   U2825 : BUF_X1 port map( A => n16691, Z => n17476);
   U2788 : INV_X1 port map( A => n16944, ZN => n5398);
   U10024 : AND2_X1 port map( A1 => n6013, A2 => n17424, ZN => n16846);
   U1951 : NAND3_X1 port map( A1 => n16277, A2 => n4653, A3 => n4654, ZN => 
                           n1384);
   U11426 : NAND2_X1 port map( A1 => n4155, A2 => n4154, ZN => n17771);
   U2734 : NAND2_X1 port map( A1 => n5518, A2 => n5517, ZN => n17977);
   U2757 : OR2_X1 port map( A1 => n17042, A2 => n17041, ZN => n18334);
   U3485 : INV_X1 port map( A => n15810, ZN => n18298);
   U1839 : NAND3_X1 port map( A1 => n2375, A2 => n6554, A3 => n6553, ZN => 
                           n18020);
   U939 : BUF_X1 port map( A => n17695, Z => n18279);
   U386 : INV_X1 port map( A => n18017, ZN => n524);
   U569 : CLKBUF_X1 port map( A => n17207, Z => n18126);
   U9098 : OAI21_X1 port map( B1 => n2791, B2 => n18303, A => n18302, ZN => 
                           n19631);
   U8367 : NAND3_X1 port map( A1 => n2457, A2 => n16189, A3 => n5417, ZN => 
                           n5416);
   U1345 : AND2_X1 port map( A1 => n6655, A2 => n6654, ZN => n18735);
   U5162 : NAND2_X1 port map( A1 => n16821, A2 => n28254, ZN => n18395);
   U21575 : OAI211_X1 port map( C1 => n18147, C2 => n18049, A => n18048, B => 
                           n18047, ZN => n19421);
   U1737 : XNOR2_X1 port map( A => n19051, B => n19050, ZN => n20475);
   U22712 : NOR2_X1 port map( A1 => n19985, A2 => n29066, ZN => n20163);
   U1027 : INV_X2 port map( A => n20133, ZN => n415);
   U10214 : NAND2_X1 port map( A1 => n18847, A2 => n835, ZN => n20875);
   U3960 : NAND3_X1 port map( A1 => n2872, A2 => n3411, A3 => n5469, ZN => 
                           n21221);
   U1132 : INV_X1 port map( A => n20864, ZN => n28789);
   U7106 : INV_X1 port map( A => n21581, ZN => n5142);
   U22817 : OAI211_X1 port map( C1 => n21452, C2 => n21451, A => n1445, B => 
                           n29178, ZN => n22334);
   U27 : MUX2_X1 port map( A => n20856, B => n20855, S => n21143, Z => n22526);
   U1033 : OAI21_X1 port map( B1 => n18851, B2 => n29553, A => n18850, ZN => 
                           n6520);
   U8276 : AND3_X1 port map( A1 => n5634, A2 => n21107, A3 => n21108, ZN => 
                           n22052);
   U9514 : NAND2_X1 port map( A1 => n21050, A2 => n3039, ZN => n22820);
   U12935 : NAND3_X1 port map( A1 => n2299, A2 => n19803, A3 => n4225, ZN => 
                           n28450);
   U24256 : INV_X1 port map( A => n23262, ZN => n23716);
   U2427 : CLKBUF_X1 port map( A => n22954, Z => n23845);
   U2404 : INV_X1 port map( A => n6227, ZN => n4231);
   U1468 : BUF_X1 port map( A => n23745, Z => n24516);
   U20339 : MUX2_X1 port map( A => n23866, B => n23865, S => n28531, Z => 
                           n25790);
   U13900 : CLKBUF_X1 port map( A => n25913, Z => n29039);
   U1060 : NAND2_X2 port map( A1 => n6055, A2 => n24587, ZN => n945);
   U25579 : NOR2_X1 port map( A1 => n24286, A2 => n24285, ZN => n25341);
   U1209 : AND4_X1 port map( A1 => n5118, A2 => n5117, A3 => n5115, A4 => n2997
                           , ZN => n25820);
   U26202 : INV_X1 port map( A => n26440, ZN => n26775);
   U5111 : OR2_X1 port map( A1 => n26502, A2 => n3632, ZN => n27852);
   U1612 : AND3_X1 port map( A1 => n6627, A2 => n26759, A3 => n6626, ZN => 
                           n28107);
   U2186 : CLKBUF_X1 port map( A => n27582, Z => n27586);
   U1001 : AOI21_X2 port map( B1 => n11738, B2 => n11737, A => n11736, ZN => 
                           n13511);
   U9975 : AND3_X2 port map( A1 => n2547, A2 => n7929, A3 => n8214, ZN => n8669
                           );
   U14673 : XNOR2_X2 port map( A => Key(10), B => Plaintext(10), ZN => n7342);
   U5636 : MUX2_X2 port map( A => n17559, B => n17558, S => n29142, Z => n18251
                           );
   U1299 : AND3_X2 port map( A1 => n5081, A2 => n16778, A3 => n16777, ZN => 
                           n18106);
   U10548 : OAI21_X2 port map( B1 => n4000, B2 => n11753, A => n11752, ZN => 
                           n12699);
   U1202 : AND2_X2 port map( A1 => n4904, A2 => n4903, ZN => n11622);
   U9516 : OAI211_X2 port map( C1 => n3082, C2 => n6573, A => n11579, B => 
                           n6572, ZN => n15415);
   U885 : NAND2_X2 port map( A1 => n722, A2 => n11464, ZN => n12817);
   U1189 : BUF_X2 port map( A => n6988, Z => n7821);
   U10359 : OR2_X2 port map( A1 => n5073, A2 => n14397, ZN => n15265);
   U9835 : NAND2_X2 port map( A1 => n18119, A2 => n268, ZN => n21692);
   U8364 : XNOR2_X2 port map( A => n2387, B => Key(164), ZN => n7997);
   U5117 : NAND3_X2 port map( A1 => n6412, A2 => n14782, A3 => n2047, ZN => 
                           n16321);
   U313 : OR2_X2 port map( A1 => n17237, A2 => n17238, ZN => n18433);
   U542 : BUF_X2 port map( A => n7285, Z => n7796);
   U2160 : AND2_X2 port map( A1 => n28720, A2 => n28719, ZN => n12696);
   U1275 : NOR2_X2 port map( A1 => n1929, A2 => n21736, ZN => n21388);
   U183 : XNOR2_X2 port map( A => n7205, B => Key(136), ZN => n7655);
   U1804 : AND2_X2 port map( A1 => n8240, A2 => n8241, ZN => n8963);
   U852 : AND3_X2 port map( A1 => n3525, A2 => n3524, A3 => n3523, ZN => n19615
                           );
   U483 : NOR2_X2 port map( A1 => n9730, A2 => n28269, ZN => n12198);
   U3921 : NAND2_X2 port map( A1 => n7005, A2 => n7006, ZN => n8699);
   U61 : AND3_X2 port map( A1 => n4614, A2 => n4612, A3 => n4613, ZN => n17942)
                           ;
   U655 : NOR2_X2 port map( A1 => n23130, A2 => n23129, ZN => n25738);
   U9015 : NAND3_X2 port map( A1 => n3979, A2 => n2730, A3 => n3977, ZN => 
                           n16305);
   U565 : NAND2_X2 port map( A1 => n13764, A2 => n2408, ZN => n15202);
   U687 : BUF_X2 port map( A => n14407, Z => n14332);
   U200 : OR2_X2 port map( A1 => n23032, A2 => n23151, ZN => n24706);
   U133 : INV_X2 port map( A => n6958, ZN => n7925);
   U15740 : NAND2_X2 port map( A1 => n10407, A2 => n10406, ZN => n10283);
   U3126 : AND2_X2 port map( A1 => n2749, A2 => n11783, ZN => n11550);
   U1928 : AND2_X2 port map( A1 => n12368, A2 => n12369, ZN => n14937);
   U23 : BUF_X2 port map( A => n21775, Z => n23788);
   U2343 : NOR2_X2 port map( A1 => n9239, A2 => n9240, ZN => n9352);
   U2830 : BUF_X2 port map( A => n16730, Z => n17497);
   U832 : OAI21_X2 port map( B1 => n1237, B2 => n7287, A => n7286, ZN => n8891)
                           ;
   U526 : XNOR2_X2 port map( A => n16220, B => n16219, ZN => n17139);
   U31 : NAND2_X2 port map( A1 => n4813, A2 => n20073, ZN => n22013);
   U10898 : MUX2_X2 port map( A => n24385, B => n24384, S => n4195, Z => n26071
                           );
   U1402 : BUF_X2 port map( A => n15018, Z => n15022);
   U21435 : OAI211_X2 port map( C1 => n17810, C2 => n18195, A => n17809, B => 
                           n17808, ZN => n19679);
   U842 : AND4_X2 port map( A1 => n4203, A2 => n4206, A3 => n4202, A4 => n4201,
                           ZN => n22245);
   U12983 : AND4_X2 port map( A1 => n15267, A2 => n5721, A3 => n5722, A4 => 
                           n5723, ZN => n16084);
   U3205 : XNOR2_X2 port map( A => n10084, B => n10083, ZN => n11152);
   U24938 : XNOR2_X2 port map( A => n18728, B => n5586, ZN => n20039);
   U2937 : OR2_X2 port map( A1 => n13975, A2 => n13974, ZN => n15321);
   U3240 : XNOR2_X2 port map( A => n9812, B => n9510, ZN => n11038);
   U1807 : AND3_X2 port map( A1 => n5919, A2 => n5921, A3 => n2048, ZN => 
                           n18383);
   U1405 : NAND2_X2 port map( A1 => n9556, A2 => n9557, ZN => n12206);
   U633 : OR2_X2 port map( A1 => n8949, A2 => n8948, ZN => n10371);
   U19217 : MUX2_X2 port map( A => n14035, B => n14034, S => n14033, Z => 
                           n15284);
   U28241 : OAI211_X2 port map( C1 => n14423, C2 => n14422, A => n14449, B => 
                           n14448, ZN => n15503);
   U733 : XNOR2_X2 port map( A => n7009, B => Key(66), ZN => n8024);
   U1200 : OR2_X2 port map( A1 => n3280, A2 => n21936, ZN => n22811);
   U15590 : MUX2_X2 port map( A => n8447, B => n8446, S => n9187, Z => n10298);
   U635 : BUF_X2 port map( A => n10853, Z => n1933);
   U13431 : OAI21_X2 port map( B1 => n6143, B2 => n14170, A => n6142, ZN => 
                           n14666);
   U1610 : NAND2_X2 port map( A1 => n29237, A2 => n4564, ZN => n18173);
   U430 : NAND3_X2 port map( A1 => n3076, A2 => n3077, A3 => n5668, ZN => 
                           n21090);
   U10767 : NAND2_X2 port map( A1 => n24670, A2 => n4603, ZN => n25869);
   U18966 : BUF_X2 port map( A => n13674, Z => n14498);
   U8804 : NAND2_X2 port map( A1 => n4970, A2 => n10557, ZN => n12000);
   U14887 : AND3_X2 port map( A1 => n7264, A2 => n7263, A3 => n7262, ZN => 
                           n8944);
   U3346 : AND2_X2 port map( A1 => n1007, A2 => n7213, ZN => n9221);
   U114 : OAI21_X2 port map( B1 => n984, B2 => n23038, A => n23037, ZN => 
                           n24707);
   U2888 : NAND2_X2 port map( A1 => n6456, A2 => n15317, ZN => n16625);
   U20139 : OAI21_X2 port map( B1 => n24038, B2 => n24039, A => n24037, ZN => 
                           n28592);
   U3124 : INV_X2 port map( A => n11195, ZN => n6706);
   U262 : BUF_X2 port map( A => n12607, Z => n13699);
   U63 : NAND3_X2 port map( A1 => n18073, A2 => n4846, A3 => n4845, ZN => 
                           n18508);
   U16244 : XNOR2_X2 port map( A => n9463, B => n9464, ZN => n10929);
   U2294 : NAND3_X2 port map( A1 => n818, A2 => n23912, A3 => n812, ZN => 
                           n25372);
   U1108 : AND3_X2 port map( A1 => n6256, A2 => n18514, A3 => n6255, ZN => 
                           n18652);
   U990 : AND3_X2 port map( A1 => n17461, A2 => n17462, A3 => n17460, ZN => 
                           n18213);
   U3075 : AND2_X2 port map( A1 => n4276, A2 => n12074, ZN => n12377);
   U1392 : BUF_X2 port map( A => n23049, Z => n23193);
   U1712 : XNOR2_X2 port map( A => n20279, B => n20280, ZN => n23067);
   U18588 : XNOR2_X2 port map( A => n13100, B => n6922, ZN => n14346);
   U1892 : XNOR2_X2 port map( A => n21747, B => n21746, ZN => n23787);
   U703 : NAND2_X2 port map( A1 => n3733, A2 => n13991, ZN => n16295);
   U14667 : OR2_X2 port map( A1 => n7113, A2 => n7112, ZN => n8826);
   U392 : NAND2_X2 port map( A1 => n21139, A2 => n3534, ZN => n22822);
   U23141 : OAI211_X2 port map( C1 => n29521, C2 => n20514, A => n20513, B => 
                           n20512, ZN => n21612);
   U869 : NAND2_X2 port map( A1 => n2227, A2 => n1163, ZN => n12332);
   U1180 : OR2_X2 port map( A1 => n7190, A2 => n7189, ZN => n8687);
   U574 : XNOR2_X2 port map( A => n21846, B => n21845, ZN => n23776);
   U139 : NAND2_X2 port map( A1 => n24418, A2 => n24419, ZN => n25737);
   U11087 : XNOR2_X2 port map( A => n21169, B => n21170, ZN => n23672);
   U18174 : XNOR2_X2 port map( A => n12571, B => n6923, ZN => n14314);
   U3397 : BUF_X2 port map( A => n7106, Z => n7895);
   U5534 : BUF_X2 port map( A => n12712, Z => n14460);
   U560 : MUX2_X2 port map( A => n16751, B => n16750, S => n28454, Z => n18096)
                           ;
   U3186 : AND2_X2 port map( A1 => n17143, A2 => n17138, ZN => n17088);
   U8731 : AND3_X2 port map( A1 => n2087, A2 => n4087, A3 => n2847, ZN => 
                           n12042);
   U1104 : OR2_X2 port map( A1 => n7505, A2 => n7504, ZN => n8819);
   U1073 : AND3_X2 port map( A1 => n5385, A2 => n20507, A3 => n20508, ZN => 
                           n21327);
   U370 : AND2_X2 port map( A1 => n1294, A2 => n8789, ZN => n9934);
   U28134 : XNOR2_X2 port map( A => n15842, B => n15841, ZN => n17554);
   U11101 : XNOR2_X2 port map( A => n6051, B => n13431, ZN => n3860);
   U8862 : MUX2_X2 port map( A => n9077, B => n9076, S => n9075, Z => n9695);
   U4700 : BUF_X2 port map( A => n16724, Z => n17477);
   U11029 : XNOR2_X2 port map( A => n9835, B => n9834, ZN => n10989);
   U3272 : INV_X2 port map( A => n9785, ZN => n9677);
   U2292 : INV_X2 port map( A => n24272, ZN => n26095);
   U1470 : XNOR2_X2 port map( A => n25070, B => n4810, ZN => n26919);
   U2408 : AND2_X2 port map( A1 => n23651, A2 => n23472, ZN => n1740);
   U3136 : AND3_X2 port map( A1 => n6778, A2 => n6780, A3 => n6777, ZN => 
                           n12304);
   U2744 : OAI21_X2 port map( B1 => n17085, B2 => n2609, A => n17084, ZN => 
                           n18595);
   U12795 : XNOR2_X2 port map( A => n21584, B => n21583, ZN => n23666);
   U2618 : XNOR2_X2 port map( A => n19091, B => n19090, ZN => n20483);
   U1543 : AND2_X2 port map( A1 => n6313, A2 => n6312, ZN => n22248);
   U178 : MUX2_X2 port map( A => n24154, B => n24153, S => n23597, Z => n25366)
                           ;
   U23404 : OAI21_X2 port map( B1 => n20905, B2 => n20904, A => n20903, ZN => 
                           n22459);
   U1535 : NAND2_X2 port map( A1 => n28727, A2 => n14946, ZN => n15949);
   U3933 : NAND3_X2 port map( A1 => n860, A2 => n4016, A3 => n11957, ZN => 
                           n13488);
   U11168 : AND2_X2 port map( A1 => n15349, A2 => n15345, ZN => n15046);
   U1231 : AND3_X2 port map( A1 => n24478, A2 => n24477, A3 => n24476, ZN => 
                           n5146);
   U980 : XNOR2_X2 port map( A => n13492, B => n13491, ZN => n5918);
   U2878 : OR2_X2 port map( A1 => n3925, A2 => n3923, ZN => n1967);
   U2024 : AND3_X2 port map( A1 => n8822, A2 => n1813, A3 => n8821, ZN => n9505
                           );
   U7787 : NAND2_X2 port map( A1 => n28883, A2 => n16938, ZN => n18529);
   U16435 : XNOR2_X2 port map( A => n9690, B => n9691, ZN => n11053);
   U4855 : NAND4_X2 port map( A1 => n8640, A2 => n8641, A3 => n8842, A4 => 
                           n1311, ZN => n9746);
   U1163 : OAI211_X2 port map( C1 => n6640, C2 => n6639, A => n13466, B => 
                           n3613, ZN => n14972);
   U5890 : XNOR2_X2 port map( A => n9299, B => n9300, ZN => n10976);
   U3216 : XNOR2_X2 port map( A => n16317, B => n16316, ZN => n17062);
   U677 : NOR2_X2 port map( A1 => n8374, A2 => n8373, ZN => n10330);
   U23881 : INV_X2 port map( A => n22618, ZN => n22724);
   U1708 : AND3_X2 port map( A1 => n28259, A2 => n20246, A3 => n28258, ZN => 
                           n22618);
   U6509 : INV_X2 port map( A => n21649, ZN => n22610);
   U3154 : OAI211_X2 port map( C1 => n6021, C2 => n11130, A => n11129, B => 
                           n11128, ZN => n11778);
   U2943 : AND2_X2 port map( A1 => n1321, A2 => n14548, ZN => n15171);
   U28304 : BUF_X2 port map( A => n13824, Z => n13826);
   U2718 : AND2_X2 port map( A1 => n17096, A2 => n17095, ZN => n18144);
   U4429 : XNOR2_X2 port map( A => n19366, B => n19365, ZN => n20619);
   U1292 : BUF_X2 port map( A => n16289, Z => n321);
   U2005 : OR2_X2 port map( A1 => n10812, A2 => n10813, ZN => n11715);
   U297 : AOI21_X2 port map( B1 => n18036, B2 => n17745, A => n17622, ZN => 
                           n18738);
   U12120 : NAND2_X2 port map( A1 => n26803, A2 => n3075, ZN => n27277);
   U9761 : NOR2_X2 port map( A1 => n20337, A2 => n3144, ZN => n21177);
   U148 : AND2_X2 port map( A1 => n15194, A2 => n14241, ZN => n14172);
   U815 : XNOR2_X2 port map( A => n11481, B => n11480, ZN => n14241);
   U2373 : XNOR2_X2 port map( A => Key(119), B => Plaintext(119), ZN => n29135)
                           ;
   U577 : XNOR2_X2 port map( A => n16490, B => n16489, ZN => n17484);
   U985 : OAI21_X2 port map( B1 => n7908, B2 => n8651, A => n7907, ZN => n4479)
                           ;
   U384 : OR2_X2 port map( A1 => n839, A2 => n8344, ZN => n10138);
   U272 : AND3_X2 port map( A1 => n28292, A2 => n18227, A3 => n28672, ZN => 
                           n5439);
   U3402 : BUF_X2 port map( A => n7072, Z => n7580);
   U13726 : AND3_X2 port map( A1 => n15277, A2 => n15278, A3 => n6493, ZN => 
                           n15545);
   U442 : AOI21_X2 port map( B1 => n19817, B2 => n19816, A => n1970, ZN => 
                           n21493);
   U9471 : MUX2_X2 port map( A => n23328, B => n23327, S => n23474, Z => n24677
                           );
   U1934 : NAND3_X2 port map( A1 => n5843, A2 => n5842, A3 => n16664, ZN => 
                           n1741);
   U2293 : NAND2_X2 port map( A1 => n3206, A2 => n2473, ZN => n26118);
   U27119 : NOR2_X2 port map( A1 => n26417, A2 => n26416, ZN => n27255);
   U208 : OAI21_X2 port map( B1 => n23479, B2 => n23478, A => n23477, ZN => 
                           n24779);
   U3477 : XNOR2_X2 port map( A => Key(2), B => Plaintext(2), ZN => n7089);
   U11002 : XNOR2_X2 port map( A => n15610, B => n15609, ZN => n17385);
   U14687 : XNOR2_X2 port map( A => n7123, B => Key(40), ZN => n8143);
   U19888 : OAI21_X2 port map( B1 => n15416, B2 => n223, A => n15414, ZN => 
                           n16649);
   U1655 : OAI211_X2 port map( C1 => n11062, C2 => n11061, A => n11060, B => 
                           n11059, ZN => n12827);
   U3245 : XNOR2_X2 port map( A => n9497, B => n9496, ZN => n11315);
   U1239 : NAND2_X2 port map( A1 => n1298, A2 => n1297, ZN => n8760);
   U3654 : NOR2_X1 port map( A1 => n3760, A2 => n3759, ZN => n3758);
   U553 : XNOR2_X2 port map( A => n19068, B => n19067, ZN => n20481);
   U8225 : AND2_X2 port map( A1 => n6093, A2 => n6094, ZN => n9028);
   U22984 : INV_X1 port map( A => n20207, ZN => n21678);
   U255 : AND2_X2 port map( A1 => n17789, A2 => n17788, ZN => n18181);
   U447 : XNOR2_X2 port map( A => n18631, B => n18632, ZN => n20401);
   U2667 : AND2_X2 port map( A1 => n2775, A2 => n2774, ZN => n19370);
   U322 : NOR2_X2 port map( A1 => n10168, A2 => n10167, ZN => n1890);
   U640 : INV_X2 port map( A => n18782, ZN => n19592);
   U641 : OR2_X2 port map( A1 => n18427, A2 => n18428, ZN => n18782);
   U657 : NAND4_X2 port map( A1 => n1791, A2 => n5957, A3 => n8333, A4 => n1790
                           , ZN => n10171);
   U184 : OAI211_X2 port map( C1 => n11558, C2 => n3946, A => n3944, B => 
                           n11557, ZN => n13364);
   U10840 : MUX2_X2 port map( A => n17311, B => n17310, S => n17440, Z => 
                           n18156);
   U2740 : AND2_X2 port map( A1 => n5107, A2 => n2030, ZN => n17989);
   U1656 : AND2_X2 port map( A1 => n2106, A2 => n2105, ZN => n26004);
   U5736 : OAI211_X2 port map( C1 => n14967, C2 => n14968, A => n14966, B => 
                           n28856, ZN => n16534);
   U1061 : NAND2_X2 port map( A1 => n195, A2 => n3578, ZN => n22791);
   U1210 : INV_X2 port map( A => n11247, ZN => n12049);
   U2365 : OR2_X2 port map( A1 => n5626, A2 => n5627, ZN => n24643);
   U287 : NAND2_X2 port map( A1 => n12126, A2 => n13203, ZN => n13406);
   U1383 : BUF_X2 port map( A => n19678, Z => n19464);
   U1970 : NOR2_X2 port map( A1 => n14733, A2 => n14115, ZN => n14512);
   U5930 : BUF_X2 port map( A => n6958, Z => n7625);
   U27246 : OR3_X2 port map( A1 => n26596, A2 => n27875, A3 => n27865, ZN => 
                           n26597);
   U2403 : BUF_X2 port map( A => n23245, Z => n23577);
   U3379 : OR2_X2 port map( A1 => n7833, A2 => n7834, ZN => n8910);
   U3050 : BUF_X1 port map( A => n12388, Z => n12684);
   U2298 : MUX2_X2 port map( A => n24399, B => n24398, S => n24676, Z => n25900
                           );
   U16703 : AOI21_X2 port map( B1 => n10054, B2 => n10053, A => n10052, ZN => 
                           n11853);
   U3266 : OAI211_X2 port map( C1 => n8761, C2 => n8569, A => n7387, B => n7386
                           , ZN => n10364);
   U13669 : NAND2_X2 port map( A1 => n10533, A2 => n6430, ZN => n6432);
   U19744 : NAND2_X2 port map( A1 => n15064, A2 => n15063, ZN => n16619);
   U14444 : XNOR2_X2 port map( A => n6978, B => Key(97), ZN => n7634);
   U296 : BUF_X2 port map( A => n27081, Z => n27085);
   U4545 : NAND3_X2 port map( A1 => n1805, A2 => n23044, A3 => n23043, ZN => 
                           n1808);
   U13124 : OAI21_X2 port map( B1 => n20912, B2 => n21607, A => n20911, ZN => 
                           n22123);
   U3384 : OR2_X1 port map( A1 => n8315, A2 => n8314, ZN => n8802);
   U367 : AND4_X1 port map( A1 => n7270, A2 => n7272, A3 => n7269, A4 => n7271,
                           ZN => n8762);
   U1590 : BUF_X1 port map( A => Key(167), Z => n27225);
   U501 : BUF_X1 port map( A => n9913, Z => n11121);
   U580 : BUF_X1 port map( A => n13837, Z => n14150);
   U2929 : NAND3_X1 port map( A1 => n5641, A2 => n2969, A3 => n5642, ZN => 
                           n14916);
   U1972 : OAI21_X1 port map( B1 => n13736, B2 => n557, A => n13735, ZN => 
                           n15371);
   U1497 : BUF_X2 port map( A => n15085, Z => n323);
   U8561 : AND2_X1 port map( A1 => n14501, A2 => n6797, ZN => n15494);
   U6023 : INV_X1 port map( A => n15108, ZN => n15406);
   U2940 : BUF_X1 port map( A => n14621, Z => n15502);
   U12513 : OAI21_X1 port map( B1 => n13950, B2 => n14667, A => n13949, ZN => 
                           n16564);
   U1965 : MUX2_X1 port map( A => n14525, B => n14524, S => n550, Z => n16405);
   U20056 : BUF_X1 port map( A => n15617, Z => n16636);
   U1193 : AND2_X1 port map( A1 => n3917, A2 => n3919, ZN => n16556);
   U46 : OAI21_X1 port map( B1 => n16705, B2 => n28574, A => n16704, ZN => 
                           n18449);
   U2721 : AND2_X1 port map( A1 => n16441, A2 => n16440, ZN => n18467);
   U12232 : AOI21_X2 port map( B1 => n17503, B2 => n17504, A => n4963, ZN => 
                           n18393);
   U1503 : BUF_X2 port map( A => n17534, Z => n17842);
   U3841 : AND2_X1 port map( A1 => n16663, A2 => n824, ZN => n18311);
   U755 : BUF_X1 port map( A => n19556, Z => n28144);
   U189 : AND2_X1 port map( A1 => n28898, A2 => n4793, ZN => n21656);
   U1181 : BUF_X1 port map( A => n22765, Z => n28162);
   U7245 : INV_X1 port map( A => n22356, ZN => n24744);
   U4 : BUF_X1 port map( A => n25182, Z => n25441);
   U5 : NAND3_X1 port map( A1 => n29352, A2 => n153, A3 => n24126, ZN => n26110
                           );
   U13 : NOR2_X1 port map( A1 => n1330, A2 => n1329, ZN => n20814);
   U15 : INV_X1 port map( A => n17881, ZN => n17883);
   U17 : AND3_X1 port map( A1 => n5894, A2 => n5893, A3 => n13925, ZN => n16090
                           );
   U19 : XNOR2_X1 port map( A => n12703, B => n12702, ZN => n14459);
   U20 : BUF_X1 port map( A => n5595, Z => n29316);
   U36 : BUF_X2 port map( A => n18613, Z => n20383);
   U37 : OR2_X2 port map( A1 => n26744, A2 => n26743, ZN => n29056);
   U38 : NOR2_X2 port map( A1 => n23346, A2 => n23345, ZN => n24074);
   U71 : OR2_X2 port map( A1 => n6181, A2 => n11869, ZN => n11457);
   U80 : AND3_X2 port map( A1 => n6260, A2 => n28215, A3 => n6259, ZN => n21675
                           );
   U101 : NOR2_X1 port map( A1 => n20860, A2 => n20861, ZN => n22670);
   U104 : BUF_X2 port map( A => n25267, Z => n26757);
   U107 : MUX2_X2 port map( A => n12533, B => n12532, S => n13872, Z => n14907)
                           ;
   U110 : NAND2_X2 port map( A1 => n15273, A2 => n15954, ZN => n16387);
   U116 : NAND2_X2 port map( A1 => n8467, A2 => n29439, ZN => n9964);
   U117 : AOI211_X2 port map( C1 => n11232, C2 => n9709, A => n10621, B => 
                           n28568, ZN => n10626);
   U125 : NAND2_X2 port map( A1 => n10608, A2 => n29710, ZN => n12362);
   U131 : NAND2_X2 port map( A1 => n3563, A2 => n3562, ZN => n22891);
   U134 : OAI22_X2 port map( A1 => n20697, A2 => n20983, B1 => n20698, B2 => 
                           n20699, ZN => n22796);
   U138 : XNOR2_X2 port map( A => n13544, B => n29798, ZN => n13572);
   U141 : BUF_X2 port map( A => n16993, Z => n29299);
   U144 : NOR2_X2 port map( A1 => n19750, A2 => n20383, ZN => n20571);
   U152 : AOI21_X2 port map( B1 => n24004, B2 => n24547, A => n24003, ZN => 
                           n26109);
   U156 : NAND4_X2 port map( A1 => n13680, A2 => n13681, A3 => n14187, A4 => 
                           n13679, ZN => n15144);
   U162 : OAI21_X2 port map( B1 => n3529, B2 => n29718, A => n6335, ZN => 
                           n17818);
   U163 : OR2_X2 port map( A1 => n29794, A2 => n7526, ZN => n8593);
   U169 : OAI21_X2 port map( B1 => n15191, B2 => n15190, A => n15189, ZN => 
                           n16407);
   U170 : XNOR2_X2 port map( A => n15876, B => n15875, ZN => n17568);
   U180 : AND2_X2 port map( A1 => n26431, A2 => n26382, ZN => n26380);
   U230 : BUF_X2 port map( A => n12053, Z => n285);
   U251 : OAI211_X2 port map( C1 => n14804, C2 => n14803, A => n14805, B => 
                           n785, ZN => n4504);
   U259 : XNOR2_X2 port map( A => n25023, B => n25022, ZN => n27181);
   U260 : AND2_X2 port map( A1 => n20617, A2 => n20618, ZN => n19890);
   U261 : BUF_X2 port map( A => n26728, Z => n29501);
   U263 : AND2_X2 port map( A1 => n4597, A2 => n4594, ZN => n24758);
   U264 : XNOR2_X2 port map( A => n7073, B => Key(179), ZN => n7887);
   U274 : BUF_X2 port map( A => n25998, Z => n27368);
   U281 : AOI21_X2 port map( B1 => n12090, B2 => n12089, A => n430, ZN => 
                           n12995);
   U286 : INV_X2 port map( A => n2155, ZN => n18465);
   U288 : AND3_X2 port map( A1 => n28983, A2 => n4768, A3 => n4770, ZN => 
                           n24745);
   U289 : INV_X2 port map( A => n19843, ZN => n29315);
   U290 : AND2_X2 port map( A1 => n1832, A2 => n20864, ZN => n21183);
   U294 : AOI21_X2 port map( B1 => n21469, B2 => n28155, A => n29435, ZN => 
                           n22677);
   U298 : NOR2_X2 port map( A1 => n12995, A2 => n12101, ZN => n13331);
   U304 : OAI211_X2 port map( C1 => n8882, C2 => n8881, A => n8880, B => n8879,
                           ZN => n1852);
   U309 : AND2_X1 port map( A1 => n26434, A2 => n26433, ZN => n29493);
   U321 : AND3_X1 port map( A1 => n26453, A2 => n6736, A3 => n2043, ZN => 
                           n29542);
   U360 : INV_X1 port map( A => n25633, ZN => n27386);
   U379 : AND2_X1 port map( A1 => n21655, A2 => n21656, ZN => n29334);
   U385 : OR2_X1 port map( A1 => n14702, A2 => n14916, ZN => n15268);
   U390 : AND2_X1 port map( A1 => n18471, A2 => n18467, ZN => n18315);
   U401 : BUF_X1 port map( A => n26575, Z => n29576);
   U412 : OR2_X1 port map( A1 => n6578, A2 => n20219, ZN => n2096);
   U413 : BUF_X1 port map( A => n24214, Z => n29307);
   U431 : BUF_X1 port map( A => n24214, Z => n29309);
   U432 : OAI211_X1 port map( C1 => n8430, C2 => n7809, A => n7808, B => n7807,
                           ZN => n9550);
   U436 : CLKBUF_X1 port map( A => n11646, Z => n11712);
   U454 : CLKBUF_X1 port map( A => n15167, Z => n15474);
   U456 : XOR2_X1 port map( A => n16372, B => n16371, Z => n29294);
   U472 : NOR2_X2 port map( A1 => n17870, A2 => n17869, ZN => n18760);
   U485 : OAI211_X2 port map( C1 => n19764, C2 => n29491, A => n19763, B => 
                           n1699, ZN => n21118);
   U487 : AOI22_X1 port map( A1 => n21480, A2 => n29314, B1 => n21478, B2 => 
                           n21479, ZN => n21649);
   U489 : NOR2_X2 port map( A1 => n22930, A2 => n22929, ZN => n24593);
   U494 : AOI21_X2 port map( B1 => n22454, B2 => n22453, A => n29169, ZN => 
                           n24614);
   U496 : XNOR2_X2 port map( A => n25073, B => n26104, ZN => n26782);
   U498 : OAI21_X2 port map( B1 => n19063, B2 => n19062, A => n19061, ZN => 
                           n21703);
   U499 : XNOR2_X2 port map( A => n7202, B => Key(133), ZN => n7657);
   U502 : OAI21_X2 port map( B1 => n23105, B2 => n23301, A => n23104, ZN => 
                           n24209);
   U523 : AOI21_X2 port map( B1 => n11292, B2 => n10663, A => n10327, ZN => 
                           n12177);
   U529 : XNOR2_X2 port map( A => n13326, B => n13327, ZN => n13730);
   U546 : BUF_X1 port map( A => n23450, Z => n29295);
   U554 : BUF_X1 port map( A => n23450, Z => n29296);
   U558 : XNOR2_X1 port map( A => n22695, B => n22696, ZN => n23450);
   U570 : NOR2_X2 port map( A1 => n7044, A2 => n4825, ZN => n8808);
   U579 : AND3_X2 port map( A1 => n19911, A2 => n5938, A3 => n29265, ZN => 
                           n22330);
   U581 : AOI22_X2 port map( A1 => n7224, A2 => n7465, B1 => n7223, B2 => n7222
                           , ZN => n9220);
   U596 : CLKBUF_X1 port map( A => n16993, Z => n29297);
   U600 : CLKBUF_X1 port map( A => n16993, Z => n29298);
   U615 : XNOR2_X1 port map( A => n14592, B => n14591, ZN => n16993);
   U629 : MUX2_X2 port map( A => n14880, B => n14879, S => n15691, Z => n15982)
                           ;
   U630 : XNOR2_X2 port map( A => n19908, B => n19909, ZN => n23529);
   U631 : NAND3_X2 port map( A1 => n5975, A2 => n19943, A3 => n5976, ZN => 
                           n22265);
   U638 : XNOR2_X2 port map( A => n7029, B => Key(61), ZN => n8032);
   U644 : XNOR2_X2 port map( A => n12845, B => n12844, ZN => n14193);
   U646 : OR2_X2 port map( A1 => n7435, A2 => n7434, ZN => n9070);
   U647 : CLKBUF_X1 port map( A => n359, Z => n29300);
   U664 : BUF_X1 port map( A => n359, Z => n29301);
   U666 : BUF_X1 port map( A => n359, Z => n29302);
   U673 : XNOR2_X1 port map( A => Plaintext(158), B => Key(158), ZN => n359);
   U692 : XNOR2_X2 port map( A => n29451, B => Key(169), ZN => n441);
   U693 : XNOR2_X2 port map( A => n10182, B => n10181, ZN => n11242);
   U707 : INV_X1 port map( A => n11192, ZN => n11355);
   U711 : CLKBUF_X1 port map( A => n9123, Z => n29303);
   U712 : BUF_X2 port map( A => n9123, Z => n29304);
   U714 : XNOR2_X2 port map( A => n22505, B => n22504, ZN => n22531);
   U716 : NAND3_X2 port map( A1 => n7848, A2 => n7847, A3 => n29771, ZN => 
                           n9014);
   U724 : CLKBUF_X1 port map( A => n13946, Z => n29305);
   U727 : BUF_X2 port map( A => n13946, Z => n29306);
   U728 : XNOR2_X1 port map( A => n12048, B => n12047, ZN => n13946);
   U729 : XNOR2_X2 port map( A => n12825, B => n6343, ZN => n14194);
   U742 : NOR2_X2 port map( A1 => n14839, A2 => n14840, ZN => n15887);
   U748 : BUF_X1 port map( A => n24214, Z => n29308);
   U762 : AOI22_X1 port map( A1 => n23473, A2 => n23654, B1 => n28391, B2 => 
                           n23471, ZN => n24214);
   U764 : CLKBUF_X1 port map( A => n28606, Z => n29310);
   U770 : BUF_X1 port map( A => n28606, Z => n29311);
   U774 : XNOR2_X2 port map( A => n6208, B => Key(168), ZN => n7591);
   U788 : BUF_X2 port map( A => n22494, Z => n23839);
   U791 : OAI21_X2 port map( B1 => n8601, B2 => n9062, A => n8600, ZN => n9601)
                           ;
   U792 : NAND2_X2 port map( A1 => n5243, A2 => n5239, ZN => n8828);
   U795 : NAND2_X2 port map( A1 => n2895, A2 => n12372, ZN => n16310);
   U797 : OAI21_X2 port map( B1 => n11490, B2 => n11489, A => n11488, ZN => 
                           n13263);
   U805 : NOR2_X2 port map( A1 => n5320, A2 => n23255, ZN => n24368);
   U813 : XNOR2_X2 port map( A => n7026, B => Key(62), ZN => n7265);
   U816 : OAI211_X2 port map( C1 => n17664, C2 => n17665, A => n5700, B => 
                           n5701, ZN => n19465);
   U818 : XNOR2_X2 port map( A => n12175, B => n12174, ZN => n14260);
   U823 : XNOR2_X2 port map( A => n10049, B => n6107, ZN => n10919);
   U824 : AOI21_X2 port map( B1 => n13996, B2 => n13995, A => n13994, ZN => 
                           n16062);
   U825 : BUF_X2 port map( A => n28588, Z => n29312);
   U826 : XNOR2_X2 port map( A => n7052, B => Key(171), ZN => n7231);
   U828 : XNOR2_X2 port map( A => Key(118), B => Plaintext(118), ZN => n7933);
   U830 : XNOR2_X2 port map( A => n13344, B => n13345, ZN => n13912);
   U835 : OAI21_X2 port map( B1 => n4022, B2 => n8274, A => n8273, ZN => n8958)
                           ;
   U840 : XNOR2_X2 port map( A => Key(70), B => Plaintext(70), ZN => n7844);
   U841 : XNOR2_X2 port map( A => n6989, B => Key(91), ZN => n7822);
   U844 : NAND2_X2 port map( A1 => n938, A2 => n1171, ZN => n10183);
   U862 : NAND4_X2 port map( A1 => n14537, A2 => n14538, A3 => n14536, A4 => 
                           n14535, ZN => n15927);
   U872 : XNOR2_X2 port map( A => n7061, B => Key(163), ZN => n7995);
   U874 : AOI21_X2 port map( B1 => n7344, B2 => n4051, A => n7343, ZN => n8563)
                           ;
   U879 : OAI22_X2 port map( A1 => n6811, A2 => n6429, B1 => n18254, B2 => 
                           n28370, ZN => n28516);
   U880 : XNOR2_X2 port map( A => n21952, B => n21953, ZN => n23247);
   U886 : OAI21_X2 port map( B1 => n6346, B2 => n20803, A => n6345, ZN => 
                           n22903);
   U888 : BUF_X2 port map( A => n21359, Z => n28586);
   U917 : XNOR2_X2 port map( A => Key(142), B => Plaintext(142), ZN => n8280);
   U919 : XNOR2_X2 port map( A => n12656, B => n12655, ZN => n14452);
   U928 : XNOR2_X2 port map( A => n12552, B => n12553, ZN => n14317);
   U935 : XNOR2_X2 port map( A => Key(117), B => Plaintext(117), ZN => n7614);
   U944 : OAI211_X2 port map( C1 => n6716, C2 => n6019, A => n6243, B => n2935,
                           ZN => n19632);
   U945 : NAND2_X2 port map( A1 => n4192, A2 => n4905, ZN => n6314);
   U952 : OAI22_X2 port map( A1 => n8538, A2 => n28845, B1 => n8542, B2 => 
                           n8731, ZN => n9626);
   U957 : XNOR2_X2 port map( A => n18257, B => n18258, ZN => n20547);
   U962 : XNOR2_X2 port map( A => n16474, B => n16475, ZN => n17505);
   U966 : XNOR2_X2 port map( A => n8125, B => n8126, ZN => n11330);
   U967 : OAI21_X2 port map( B1 => n9192, B2 => n9191, A => n9190, ZN => n10072
                           );
   U971 : XNOR2_X2 port map( A => n16413, B => n16412, ZN => n17181);
   U974 : XNOR2_X2 port map( A => n16098, B => n15521, ZN => n17414);
   U975 : XNOR2_X2 port map( A => Key(183), B => Plaintext(183), ZN => n7172);
   U976 : OAI21_X2 port map( B1 => n21181, B2 => n21180, A => n879, ZN => 
                           n22514);
   U981 : XNOR2_X2 port map( A => n7046, B => Key(156), ZN => n7675);
   U982 : NOR2_X2 port map( A1 => n26462, A2 => n6221, ZN => n27426);
   U984 : MUX2_X2 port map( A => n10095, B => n10094, S => n10905, Z => n13219)
                           ;
   U996 : OAI211_X2 port map( C1 => n5040, C2 => n12134, A => n5039, B => n5038
                           , ZN => n13459);
   U997 : NOR2_X2 port map( A1 => n29351, A2 => n21830, ZN => n24726);
   U1017 : XNOR2_X2 port map( A => Key(127), B => Plaintext(127), ZN => n7618);
   U1019 : OAI211_X2 port map( C1 => n8609, C2 => n7419, A => n6405, B => n6404
                           , ZN => n4713);
   U1025 : OAI211_X2 port map( C1 => n8463, C2 => n7120, A => n7119, B => n2410
                           , ZN => n9799);
   U1034 : OAI211_X2 port map( C1 => n4895, C2 => n4896, A => n6873, B => n4894
                           , ZN => n15456);
   U1037 : AND3_X2 port map( A1 => n1676, A2 => n2451, A3 => n1675, ZN => 
                           n24373);
   U1044 : AOI21_X2 port map( B1 => n21529, B2 => n21528, A => n1263, ZN => 
                           n24751);
   U1046 : XNOR2_X2 port map( A => n19259, B => n4307, ZN => n4569);
   U1047 : XNOR2_X2 port map( A => n7008, B => Key(71), ZN => n29106);
   U1054 : XNOR2_X2 port map( A => n9459, B => n9458, ZN => n10932);
   U1069 : XNOR2_X2 port map( A => n12446, B => n12445, ZN => n14402);
   U1070 : OAI22_X2 port map( A1 => n3201, A2 => n11854, B1 => n3307, B2 => 
                           n3306, ZN => n12978);
   U1081 : XNOR2_X2 port map( A => n14954, B => n14955, ZN => n17437);
   U1088 : XNOR2_X2 port map( A => Plaintext(32), B => Key(32), ZN => n7349);
   U1109 : NOR2_X2 port map( A1 => n4343, A2 => n21324, ZN => n22386);
   U1111 : OR2_X1 port map( A1 => n442, A2 => n27625, ZN => n29463);
   U1115 : INV_X1 port map( A => n4823, ZN => n27458);
   U1116 : OAI211_X1 port map( C1 => n2140, C2 => n1950, A => n2139, B => n2038
                           , ZN => n27628);
   U1130 : INV_X1 port map( A => n24433, ZN => n29726);
   U1150 : INV_X1 port map( A => n23525, ZN => n23663);
   U1156 : INV_X1 port map( A => n21291, ZN => n29313);
   U1159 : INV_X1 port map( A => n21387, ZN => n29314);
   U1165 : NAND2_X1 port map( A1 => n29425, A2 => n18446, ZN => n19219);
   U1212 : NAND2_X1 port map( A1 => n3597, A2 => n17764, ZN => n2759);
   U1213 : INV_X2 port map( A => n14894, ZN => n3362);
   U1225 : AND3_X1 port map( A1 => n13723, A2 => n13722, A3 => n2144, ZN => 
                           n15372);
   U1248 : INV_X2 port map( A => n14317, ZN => n14313);
   U1255 : NAND3_X1 port map( A1 => n29466, A2 => n11966, A3 => n2976, ZN => 
                           n13209);
   U1271 : NAND2_X1 port map( A1 => n12154, A2 => n29705, ZN => n13433);
   U1276 : INV_X2 port map( A => n12428, ZN => n29735);
   U1284 : BUF_X1 port map( A => n12577, Z => n28202);
   U1286 : OR2_X1 port map( A1 => n7035, A2 => n7034, ZN => n10297);
   U1290 : BUF_X1 port map( A => n7114, Z => n8824);
   U1291 : OAI21_X1 port map( B1 => n7999, B2 => n7881, A => n5363, ZN => n8500
                           );
   U1298 : AND2_X1 port map( A1 => n7844, A2 => n29321, ZN => n29772);
   U1306 : BUF_X1 port map( A => Key(39), Z => n3083);
   U1309 : CLKBUF_X1 port map( A => Key(62), Z => n2350);
   U1310 : BUF_X1 port map( A => Key(53), Z => n27422);
   U1312 : BUF_X1 port map( A => Key(165), Z => n3565);
   U1313 : BUF_X1 port map( A => Key(45), Z => n3643);
   U1314 : BUF_X2 port map( A => n8300, Z => n29317);
   U1320 : OR2_X1 port map( A1 => n307, A2 => n26817, ZN => n29389);
   U1328 : NAND2_X1 port map( A1 => n26137, A2 => n26136, ZN => n27711);
   U1330 : BUF_X2 port map( A => n28091, Z => n28794);
   U1331 : NAND4_X1 port map( A1 => n6302, A2 => n6300, A3 => n26327, A4 => 
                           n6301, ZN => n27807);
   U1336 : AND3_X1 port map( A1 => n768, A2 => n28100, A3 => n767, ZN => n28111
                           );
   U1337 : AND3_X1 port map( A1 => n29454, A2 => n28822, A3 => n28969, ZN => 
                           n27571);
   U1346 : OAI21_X1 port map( B1 => n4739, B2 => n28410, A => n28398, ZN => 
                           n27650);
   U1354 : INV_X1 port map( A => n27551, ZN => n29445);
   U1366 : AND2_X1 port map( A1 => n29778, A2 => n5300, ZN => n27859);
   U1375 : OAI21_X1 port map( B1 => n6823, B2 => n26574, A => n6825, ZN => 
                           n6824);
   U1378 : BUF_X1 port map( A => n27120, Z => n29016);
   U1397 : BUF_X1 port map( A => n27044, Z => n28130);
   U1399 : XNOR2_X1 port map( A => n25539, B => n25538, ZN => n28783);
   U1411 : INV_X1 port map( A => n26079, ZN => n29410);
   U1419 : AND2_X1 port map( A1 => n5101, A2 => n5104, ZN => n25921);
   U1420 : OR2_X1 port map( A1 => n24128, A2 => n5752, ZN => n29352);
   U1431 : INV_X1 port map( A => n28223, ZN => n29677);
   U1432 : AND2_X1 port map( A1 => n5647, A2 => n5646, ZN => n24544);
   U1438 : AND3_X1 port map( A1 => n6764, A2 => n6763, A3 => n1965, ZN => 
                           n29471);
   U1452 : AND3_X1 port map( A1 => n23653, A2 => n5555, A3 => n23652, ZN => 
                           n24794);
   U1483 : AND3_X1 port map( A1 => n23359, A2 => n23358, A3 => n6628, ZN => 
                           n24666);
   U1490 : AOI22_X1 port map( A1 => n23316, A2 => n28390, B1 => n23317, B2 => 
                           n23565, ZN => n28635);
   U1499 : BUF_X1 port map( A => n22566, Z => n29564);
   U1505 : OR2_X1 port map( A1 => n22458, A2 => n28183, ZN => n29729);
   U1510 : XNOR2_X1 port map( A => n22254, B => n22253, ZN => n23640);
   U1516 : BUF_X1 port map( A => n23773, Z => n29641);
   U1518 : INV_X1 port map( A => n28582, ZN => n29402);
   U1525 : XNOR2_X1 port map( A => n6520, B => n22670, ZN => n22828);
   U1526 : AOI22_X1 port map( A1 => n21115, A2 => n1897, B1 => n21114, B2 => 
                           n21463, ZN => n29519);
   U1536 : INV_X1 port map( A => n20857, ZN => n21157);
   U1547 : INV_X1 port map( A => n20756, ZN => n21463);
   U1554 : INV_X1 port map( A => n20786, ZN => n29586);
   U1556 : NAND3_X1 port map( A1 => n3972, A2 => n21134, A3 => n3971, ZN => 
                           n20886);
   U1562 : NAND2_X1 port map( A1 => n19866, A2 => n29348, ZN => n21155);
   U1571 : OAI211_X1 port map( C1 => n19972, C2 => n19973, A => n29347, B => 
                           n29346, ZN => n21387);
   U1577 : AND2_X1 port map( A1 => n20334, A2 => n20626, ZN => n20006);
   U1581 : BUF_X2 port map( A => n19766, Z => n21091);
   U1583 : BUF_X1 port map( A => n21353, Z => n28491);
   U1592 : XNOR2_X1 port map( A => n5005, B => n5006, ZN => n20441);
   U1633 : AND3_X1 port map( A1 => n29386, A2 => n6483, A3 => n29385, ZN => 
                           n18778);
   U1643 : INV_X1 port map( A => n3444, ZN => n29318);
   U1668 : OAI21_X1 port map( B1 => n18297, B2 => n18296, A => n18295, ZN => 
                           n19482);
   U1693 : NAND2_X1 port map( A1 => n2501, A2 => n2498, ZN => n19332);
   U1704 : OR2_X1 port map( A1 => n17014, A2 => n18600, ZN => n4419);
   U1707 : OR2_X1 port map( A1 => n1436, A2 => n17765, ZN => n3597);
   U1714 : OR2_X1 port map( A1 => n17976, A2 => n521, ZN => n29715);
   U1722 : AND2_X1 port map( A1 => n29191, A2 => n29192, ZN => n16868);
   U1726 : OR2_X1 port map( A1 => n17746, A2 => n29663, ZN => n17809);
   U1728 : BUF_X2 port map( A => n18601, Z => n28142);
   U1741 : OAI21_X1 port map( B1 => n5287, B2 => n5288, A => n29674, ZN => 
                           n18304);
   U1749 : OR2_X1 port map( A1 => n18507, A2 => n18508, ZN => n29350);
   U1756 : NAND2_X1 port map( A1 => n17499, A2 => n18226, ZN => n18388);
   U1757 : INV_X1 port map( A => n18195, ZN => n29663);
   U1763 : INV_X1 port map( A => n18530, ZN => n29336);
   U1778 : OAI21_X1 port map( B1 => n16748, B2 => n17350, A => n17349, ZN => 
                           n18090);
   U1782 : NOR2_X1 port map( A1 => n16806, A2 => n16668, ZN => n16850);
   U1783 : BUF_X1 port map( A => n17250, Z => n29503);
   U1791 : XNOR2_X1 port map( A => n15832, B => n15831, ZN => n17553);
   U1806 : XNOR2_X1 port map( A => n14603, B => n14602, ZN => n14629);
   U1840 : XNOR2_X1 port map( A => n15995, B => n15996, ZN => n17248);
   U1847 : XNOR2_X1 port map( A => n16480, B => n1967, ZN => n15973);
   U1849 : AND3_X1 port map( A1 => n29326, A2 => n1000, A3 => n1006, ZN => 
                           n15971);
   U1866 : INV_X1 port map( A => n16322, ZN => n29319);
   U1871 : NOR2_X1 port map( A1 => n15022, A2 => n15303, ZN => n14657);
   U1883 : OR2_X1 port map( A1 => n15223, A2 => n15224, ZN => n29355);
   U1888 : AND2_X1 port map( A1 => n1111, A2 => n13584, ZN => n14944);
   U1903 : AND3_X1 port map( A1 => n3357, A2 => n3356, A3 => n29325, ZN => 
                           n15132);
   U1906 : OR2_X1 port map( A1 => n1660, A2 => n13900, ZN => n29682);
   U1908 : AND2_X1 port map( A1 => n14415, A2 => n14215, ZN => n29760);
   U1935 : OR2_X1 port map( A1 => n4893, A2 => n13826, ZN => n14125);
   U1962 : OR2_X1 port map( A1 => n14484, A2 => n29305, ZN => n14167);
   U1967 : INV_X1 port map( A => n14480, ZN => n29320);
   U1976 : NAND2_X1 port map( A1 => n12029, A2 => n1192, ZN => n12913);
   U1996 : OAI21_X1 port map( B1 => n11588, B2 => n11589, A => n29354, ZN => 
                           n13061);
   U2029 : AND2_X1 port map( A1 => n4997, A2 => n4996, ZN => n12632);
   U2045 : OAI211_X1 port map( C1 => n11521, C2 => n11836, A => n11520, B => 
                           n29670, ZN => n13270);
   U2053 : AND2_X1 port map( A1 => n11990, A2 => n12508, ZN => n29671);
   U2091 : OR2_X1 port map( A1 => n29462, A2 => n29460, ZN => n12315);
   U2096 : NAND3_X1 port map( A1 => n10583, A2 => n10581, A3 => n10582, ZN => 
                           n12022);
   U2099 : AND2_X1 port map( A1 => n5704, A2 => n5705, ZN => n12150);
   U2102 : INV_X1 port map( A => n11896, ZN => n29461);
   U2138 : NAND2_X1 port map( A1 => n8577, A2 => n4440, ZN => n9763);
   U2152 : NAND3_X1 port map( A1 => n29393, A2 => n749, A3 => n8613, ZN => n748
                           );
   U2157 : NAND2_X1 port map( A1 => n8854, A2 => n8853, ZN => n9619);
   U2211 : AND3_X1 port map( A1 => n9537, A2 => n29660, A3 => n29661, ZN => 
                           n10033);
   U2212 : BUF_X2 port map( A => n10222, Z => n301);
   U2214 : NAND2_X1 port map( A1 => n6172, A2 => n29650, ZN => n9794);
   U2230 : INV_X1 port map( A => n8500, ZN => n29416);
   U2242 : AND3_X1 port map( A1 => n8017, A2 => n6807, A3 => n8020, ZN => n9122
                           );
   U2243 : NAND2_X1 port map( A1 => n7469, A2 => n29756, ZN => n8726);
   U2246 : INV_X1 port map( A => n24166, ZN => n5490);
   U2248 : XNOR2_X1 port map( A => n7153, B => Key(31), ZN => n8165);
   U2257 : XNOR2_X1 port map( A => n7218, B => Key(130), ZN => n6782);
   U2268 : OR2_X1 port map( A1 => n7162, A2 => n7320, ZN => n7769);
   U2275 : XNOR2_X1 port map( A => Key(59), B => Plaintext(59), ZN => n29629);
   U2277 : INV_X1 port map( A => n7850, ZN => n29321);
   U2290 : AND2_X1 port map( A1 => n7468, A2 => n7467, ZN => n29756);
   U2291 : XNOR2_X1 port map( A => Key(50), B => Plaintext(50), ZN => n7141);
   U2299 : OR2_X1 port map( A1 => n9196, A2 => n9206, ZN => n28861);
   U2346 : INV_X1 port map( A => n8891, ZN => n8887);
   U2402 : AOI22_X1 port map( A1 => n6689, A2 => n8591, B1 => n8975, B2 => n607
                           , ZN => n6688);
   U2420 : OR2_X1 port map( A1 => n9126, A2 => n284, ZN => n29650);
   U2428 : OR2_X1 port map( A1 => n8956, A2 => n8955, ZN => n8625);
   U2438 : OAI21_X1 port map( B1 => n604, B2 => n8770, A => n8579, ZN => n9582)
                           ;
   U2444 : CLKBUF_X1 port map( A => n8586, Z => n29147);
   U2469 : OAI21_X1 port map( B1 => n9137, B2 => n8552, A => n8551, ZN => n9851
                           );
   U2512 : OR2_X1 port map( A1 => n11045, A2 => n11267, ZN => n2754);
   U2513 : XNOR2_X1 port map( A => n10022, B => n9550, ZN => n10179);
   U2515 : XNOR2_X1 port map( A => n10043, B => n27422, ZN => n9750);
   U2522 : BUF_X1 port map( A => n9863, Z => n10957);
   U2523 : XNOR2_X1 port map( A => n9960, B => n9959, ZN => n10497);
   U2536 : XNOR2_X1 port map( A => n9600, B => n9599, ZN => n29148);
   U2547 : AND3_X1 port map( A1 => n3801, A2 => n3800, A3 => n3805, ZN => 
                           n12097);
   U2554 : XNOR2_X1 port map( A => n9813, B => n9812, ZN => n10991);
   U2567 : BUF_X1 port map( A => n10747, Z => n10563);
   U2571 : OR2_X1 port map( A1 => n10696, A2 => n10980, ZN => n2422);
   U2658 : OR2_X1 port map( A1 => n11782, A2 => n11419, ZN => n1493);
   U2675 : INV_X1 port map( A => n12111, ZN => n6281);
   U2679 : BUF_X1 port map( A => n11730, Z => n13206);
   U2690 : NAND3_X1 port map( A1 => n29208, A2 => n3103, A3 => n11899, ZN => 
                           n12352);
   U2703 : AND2_X1 port map( A1 => n11947, A2 => n11945, ZN => n11861);
   U2732 : OAI21_X1 port map( B1 => n11008, B2 => n11009, A => n3013, ZN => 
                           n12070);
   U2750 : NOR2_X1 port map( A1 => n11869, A2 => n11867, ZN => n11501);
   U2775 : AND2_X1 port map( A1 => n12207, A2 => n12211, ZN => n12115);
   U2778 : AND2_X1 port map( A1 => n11587, A2 => n11586, ZN => n29354);
   U2824 : CLKBUF_X1 port map( A => n11058, Z => n11435);
   U2845 : INV_X1 port map( A => n11878, ZN => n567);
   U2848 : NAND2_X1 port map( A1 => n2272, A2 => n2271, ZN => n10453);
   U2853 : OAI21_X1 port map( B1 => n12516, B2 => n11567, A => n11566, ZN => 
                           n3871);
   U2856 : NAND2_X1 port map( A1 => n12293, A2 => n12290, ZN => n12289);
   U2898 : XNOR2_X1 port map( A => n13413, B => n11912, ZN => n13274);
   U2908 : OAI21_X1 port map( B1 => n14213, B2 => n14402, A => n14212, ZN => 
                           n15239);
   U2911 : XNOR2_X1 port map( A => n12897, B => n12898, ZN => n14082);
   U2965 : BUF_X1 port map( A => n14479, Z => n293);
   U2974 : MUX2_X1 port map( A => n14154, B => n14155, S => n29037, Z => n15346
                           );
   U3010 : OAI211_X1 port map( C1 => n14480, C2 => n293, A => n14478, B => 
                           n14477, ZN => n15485);
   U3048 : OR2_X1 port map( A1 => n15250, A2 => n15135, ZN => n14729);
   U3062 : OR2_X1 port map( A1 => n14639, A2 => n14874, ZN => n15081);
   U3069 : BUF_X1 port map( A => n15001, Z => n14998);
   U3072 : NAND2_X1 port map( A1 => n3012, A2 => n3010, ZN => n15224);
   U3080 : AOI21_X1 port map( B1 => n15091, B2 => n15690, A => n15694, ZN => 
                           n15089);
   U3083 : OR2_X1 port map( A1 => n15041, A2 => n15040, ZN => n28306);
   U3140 : OR2_X1 port map( A1 => n15245, A2 => n15244, ZN => n29675);
   U3143 : OAI211_X1 port map( C1 => n15168, C2 => n15473, A => n14801, B => 
                           n15472, ZN => n3856);
   U3184 : AND4_X2 port map( A1 => n6332, A2 => n6333, A3 => n15016, A4 => 
                           n15017, ZN => n16283);
   U3226 : XNOR2_X1 port map( A => n16509, B => n16585, ZN => n16119);
   U3230 : XNOR2_X1 port map( A => n15865, B => n15092, ZN => n16598);
   U3248 : OR2_X1 port map( A1 => n17293, A2 => n17401, ZN => n5487);
   U3289 : OR2_X1 port map( A1 => n17120, A2 => n16811, ZN => n17116);
   U3304 : XNOR2_X1 port map( A => n16336, B => n16335, ZN => n17491);
   U3389 : INV_X1 port map( A => n17498, ZN => n538);
   U3440 : XNOR2_X1 port map( A => n16021, B => n16020, ZN => n17018);
   U3451 : INV_X1 port map( A => n17275, ZN => n29421);
   U3466 : XOR2_X1 port map( A => n15604, B => n15603, Z => n28497);
   U3486 : OR2_X1 port map( A1 => n29373, A2 => n17491, ZN => n17493);
   U3488 : INV_X1 port map( A => n17720, ZN => n17431);
   U3512 : XNOR2_X1 port map( A => n15748, B => n15749, ZN => n29550);
   U3552 : BUF_X1 port map( A => n17433, Z => n29566);
   U3569 : OR2_X1 port map( A1 => n6927, A2 => n2656, ZN => n2216);
   U3571 : OR2_X1 port map( A1 => n16986, A2 => n18087, ZN => n18186);
   U3581 : INV_X1 port map( A => n16611, ZN => n518);
   U3589 : OR2_X1 port map( A1 => n17842, A2 => n18241, ZN => n17757);
   U3590 : OR2_X1 port map( A1 => n18448, A2 => n18447, ZN => n29425);
   U3601 : OR2_X1 port map( A1 => n18143, A2 => n18144, ZN => n2635);
   U3673 : OR2_X1 port map( A1 => n5589, A2 => n6484, ZN => n29385);
   U3681 : AOI22_X1 port map( A1 => n18381, A2 => n18382, B1 => n5670, B2 => 
                           n17883, ZN => n3207);
   U3685 : BUF_X1 port map( A => n17793, Z => n18445);
   U3687 : NAND2_X1 port map( A1 => n3874, A2 => n3876, ZN => n19278);
   U3699 : BUF_X1 port map( A => n20017, Z => n28489);
   U3734 : INV_X1 port map( A => n20568, ZN => n97);
   U3744 : OR2_X1 port map( A1 => n97, A2 => n19833, ZN => n20570);
   U3754 : OAI21_X1 port map( B1 => n19867, B2 => n499, A => n20491, ZN => 
                           n29349);
   U3780 : INV_X1 port map( A => n20227, ZN => n29426);
   U3796 : BUF_X1 port map( A => n20484, Z => n29527);
   U3802 : AND2_X1 port map( A1 => n29315, A2 => n18838, ZN => n19779);
   U3844 : BUF_X1 port map( A => n21355, Z => n28126);
   U3848 : INV_X1 port map( A => n506, ZN => n29707);
   U3878 : AND2_X1 port map( A1 => n20488, A2 => n19093, ZN => n20359);
   U3888 : AND2_X1 port map( A1 => n28236, A2 => n28235, ZN => n29659);
   U3895 : NAND2_X1 port map( A1 => n3551, A2 => n20301, ZN => n29531);
   U3896 : NOR2_X1 port map( A1 => n21410, A2 => n20663, ZN => n21230);
   U3925 : OAI211_X1 port map( C1 => n20460, C2 => n28408, A => n4568, B => 
                           n29184, ZN => n21509);
   U3939 : OR2_X1 port map( A1 => n20728, A2 => n21292, ZN => n3252);
   U3959 : OR2_X1 port map( A1 => n21481, A2 => n21483, ZN => n21579);
   U3968 : OR2_X1 port map( A1 => n20979, A2 => n20978, ZN => n29591);
   U3981 : NAND3_X1 port map( A1 => n5139, A2 => n5141, A3 => n5140, ZN => 
                           n21987);
   U4007 : XNOR2_X1 port map( A => n29763, B => n22884, ZN => n5862);
   U4016 : INV_X1 port map( A => n21798, ZN => n29417);
   U4020 : XNOR2_X1 port map( A => n22121, B => n22120, ZN => n28484);
   U4033 : OR2_X1 port map( A1 => n5883, A2 => n23517, ZN => n29358);
   U4037 : BUF_X1 port map( A => n23156, Z => n23779);
   U4056 : CLKBUF_X1 port map( A => n23525, Z => n29123);
   U4163 : INV_X1 port map( A => n23386, ZN => n22084);
   U4173 : XNOR2_X1 port map( A => n21799, B => n29417, ZN => n28554);
   U4213 : BUF_X1 port map( A => n23629, Z => n23636);
   U4214 : CLKBUF_X1 port map( A => n22174, Z => n23260);
   U4233 : BUF_X1 port map( A => n24409, Z => n28524);
   U4238 : OR2_X1 port map( A1 => n23803, A2 => n23541, ZN => n6763);
   U4255 : OAI22_X1 port map( A1 => n4686, A2 => n23660, B1 => n405, B2 => 
                           n23659, ZN => n24813);
   U4257 : NAND2_X1 port map( A1 => n29259, A2 => n6195, ZN => n24629);
   U4259 : AOI21_X1 port map( B1 => n23846, B2 => n22455, A => n23843, ZN => 
                           n22129);
   U4260 : INV_X1 port map( A => n22931, ZN => n23819);
   U4272 : OR2_X1 port map( A1 => n29128, A2 => n24347, ZN => n29727);
   U4289 : BUF_X1 port map( A => n24813, Z => n24810);
   U4300 : OAI211_X1 port map( C1 => n23500, C2 => n5355, A => n5353, B => 
                           n5354, ZN => n23945);
   U4314 : CLKBUF_X1 port map( A => Key(126), Z => n4029);
   U4359 : MUX2_X1 port map( A => n3671, B => n23752, S => n24420, Z => n23753)
                           ;
   U4363 : OR2_X1 port map( A1 => n29028, A2 => n26466, ZN => n25617);
   U4378 : XNOR2_X1 port map( A => n26043, B => n26042, ZN => n26050);
   U4390 : XNOR2_X1 port map( A => n26071, B => n1459, ZN => n25541);
   U4404 : OR2_X1 port map( A1 => n29479, A2 => n26240, ZN => n29388);
   U4418 : NOR2_X1 port map( A1 => n1874, A2 => n26740, ZN => n29459);
   U4457 : XNOR2_X1 port map( A => n23919, B => n23920, ZN => n26449);
   U4461 : OR2_X1 port map( A1 => n26791, A2 => n23862, ZN => n28709);
   U4467 : XOR2_X1 port map( A => n24989, B => n24988, Z => n28535);
   U4504 : CLKBUF_X1 port map( A => n1907, Z => n29487);
   U4543 : INV_X1 port map( A => n27663, ZN => n29449);
   U4555 : XNOR2_X1 port map( A => n26078, B => n29410, ZN => n29633);
   U4556 : OR2_X1 port map( A1 => n29480, A2 => n29121, ZN => n29681);
   U4566 : AND2_X1 port map( A1 => n6492, A2 => n6026, ZN => n29070);
   U4568 : OR3_X1 port map( A1 => n27442, A2 => n27433, A3 => n26682, ZN => 
                           n25423);
   U4581 : MUX2_X1 port map( A => n27180, B => n27179, S => n27178, Z => n27661
                           );
   U4598 : OAI211_X1 port map( C1 => n5299, C2 => n26511, A => n5297, B => 
                           n29615, ZN => n29778);
   U4610 : NAND2_X1 port map( A1 => n26337, A2 => n5485, ZN => n27817);
   U4628 : CLKBUF_X1 port map( A => Key(133), Z => n2389);
   U4669 : INV_X1 port map( A => n1193, ZN => n26713);
   U4677 : CLKBUF_X1 port map( A => Key(84), Z => n1225);
   U4683 : CLKBUF_X1 port map( A => Key(31), Z => n3414);
   U4684 : CLKBUF_X1 port map( A => Key(7), Z => n1079);
   U4690 : CLKBUF_X1 port map( A => Key(36), Z => n3256);
   U4691 : CLKBUF_X1 port map( A => Key(124), Z => n2960);
   U4725 : AND3_X1 port map( A1 => n17898, A2 => n18356, A3 => n18355, ZN => 
                           n29322);
   U4732 : AND2_X1 port map( A1 => n673, A2 => n28481, ZN => n29323);
   U4744 : INV_X1 port map( A => n9530, ZN => n29662);
   U4753 : INV_X1 port map( A => n8749, ZN => n29395);
   U4757 : NAND2_X1 port map( A1 => n28674, A2 => n28913, ZN => n8693);
   U4761 : AND2_X1 port map( A1 => n4095, A2 => n5717, ZN => n29324);
   U4772 : OR2_X1 port map( A1 => n14080, A2 => n561, ZN => n29325);
   U4776 : INV_X1 port map( A => n14278, ZN => n29691);
   U4788 : NAND2_X1 port map( A1 => n15120, A2 => n1904, ZN => n29326);
   U4798 : INV_X1 port map( A => n15144, ZN => n29380);
   U4830 : INV_X1 port map( A => n17470, ZN => n29406);
   U4861 : XNOR2_X1 port map( A => n16181, B => n16180, ZN => n17280);
   U4869 : INV_X1 port map( A => n17280, ZN => n29737);
   U4874 : CLKBUF_X1 port map( A => n19054, Z => n20177);
   U4878 : AND2_X1 port map( A1 => n18529, A2 => n29335, ZN => n29327);
   U4882 : AND2_X1 port map( A1 => n3551, A2 => n20301, ZN => n29328);
   U4886 : OR3_X1 port map( A1 => n21709, A2 => n21372, A3 => n21277, ZN => 
                           n29329);
   U4895 : INV_X1 port map( A => n21211, ZN => n29364);
   U4896 : NOR2_X1 port map( A1 => n1330, A2 => n1329, ZN => n29488);
   U4898 : INV_X1 port map( A => n24373, ZN => n29340);
   U4987 : INV_X1 port map( A => n24258, ZN => n24976);
   U4991 : OAI211_X1 port map( C1 => n23466, C2 => n23465, A => n23464, B => 
                           n23463, ZN => n24258);
   U5031 : INV_X1 port map( A => n27364, ZN => n29387);
   U5042 : XOR2_X1 port map( A => n25093, B => n25092, Z => n29330);
   U5055 : BUF_X1 port map( A => n27028, Z => n306);
   U5061 : OR3_X1 port map( A1 => n27417, A2 => n26531, A3 => n26530, ZN => 
                           n29331);
   U5070 : NAND2_X1 port map( A1 => n26195, A2 => n27393, ZN => n29332);
   U5073 : NAND2_X1 port map( A1 => n3967, A2 => n19798, ZN => n20756);
   U5114 : NOR2_X2 port map( A1 => n11581, A2 => n6848, ZN => n12881);
   U5148 : NAND3_X2 port map( A1 => n20836, A2 => n20835, A3 => n29333, ZN => 
                           n6458);
   U5175 : NAND2_X1 port map( A1 => n6275, A2 => n29334, ZN => n29333);
   U5177 : NAND3_X1 port map( A1 => n29336, A2 => n4280, A3 => n4281, ZN => 
                           n29335);
   U5193 : NAND2_X1 port map( A1 => n29337, A2 => n23399, ZN => n751);
   U5211 : NAND2_X1 port map( A1 => n754, A2 => n755, ZN => n29337);
   U5234 : OR2_X1 port map( A1 => n17030, A2 => n17357, ZN => n4279);
   U5239 : OAI21_X1 port map( B1 => n27025, B2 => n24364, A => n29338, ZN => 
                           n27033);
   U5247 : NAND2_X1 port map( A1 => n27029, A2 => n27025, ZN => n29338);
   U5252 : OAI21_X2 port map( B1 => n2726, B2 => n14114, A => n14113, ZN => 
                           n16329);
   U5304 : OAI21_X1 port map( B1 => n23995, B2 => n29340, A => n29339, ZN => 
                           n23905);
   U5305 : NAND2_X1 port map( A1 => n23995, A2 => n24380, ZN => n29339);
   U5319 : NAND2_X1 port map( A1 => n29341, A2 => n23235, ZN => n23236);
   U5324 : NAND2_X1 port map( A1 => n23584, A2 => n23260, ZN => n29341);
   U5326 : NAND3_X1 port map( A1 => n1836, A2 => n11874, A3 => n11360, ZN => 
                           n2355);
   U5335 : OR2_X1 port map( A1 => n24577, A2 => n6741, ZN => n1204);
   U5369 : OAI21_X1 port map( B1 => n18429, B2 => n420, A => n29342, ZN => 
                           n29797);
   U5403 : NAND3_X1 port map( A1 => n2853, A2 => n2855, A3 => n18431, ZN => 
                           n29342);
   U5489 : NAND4_X2 port map( A1 => n6547, A2 => n2816, A3 => n6548, A4 => 
                           n24424, ZN => n25864);
   U5490 : OAI22_X1 port map( A1 => n15146, A2 => n3208, B1 => n1326, B2 => 
                           n15145, ZN => n15149);
   U5495 : NAND2_X1 port map( A1 => n17557, A2 => n17553, ZN => n17224);
   U5530 : NAND2_X2 port map( A1 => n29343, A2 => n26144, ZN => n27725);
   U5532 : NOR2_X1 port map( A1 => n26141, A2 => n26142, ZN => n29343);
   U5542 : NAND2_X1 port map( A1 => n14833, A2 => n893, ZN => n15291);
   U5543 : NAND2_X1 port map( A1 => n14095, A2 => n6000, ZN => n14833);
   U5548 : NAND2_X1 port map( A1 => n17123, A2 => n29344, ZN => n17125);
   U5561 : NAND3_X1 port map( A1 => n17477, A2 => n1816, A3 => n3883, ZN => 
                           n29344);
   U5606 : NAND2_X1 port map( A1 => n7159, A2 => n29345, ZN => n10346);
   U5714 : OR2_X1 port map( A1 => n7160, A2 => n7161, ZN => n29345);
   U5716 : MUX2_X1 port map( A => n24726, B => n24596, S => n24725, Z => n21944
                           );
   U5729 : NAND2_X1 port map( A1 => n29733, A2 => n21864, ZN => n24725);
   U5798 : NAND2_X1 port map( A1 => n19973, A2 => n20295, ZN => n29346);
   U5826 : NAND2_X1 port map( A1 => n19970, A2 => n20290, ZN => n29347);
   U5883 : NAND2_X1 port map( A1 => n20857, A2 => n21155, ZN => n3762);
   U5901 : INV_X1 port map( A => n29349, ZN => n29348);
   U5995 : NAND2_X1 port map( A1 => n27188, A2 => n26401, ZN => n26360);
   U6011 : NAND3_X1 port map( A1 => n3360, A2 => n15108, A3 => n3361, ZN => 
                           n3919);
   U6018 : NAND2_X1 port map( A1 => n16868, A2 => n16867, ZN => n18761);
   U6030 : OAI211_X1 port map( C1 => n18512, C2 => n418, A => n29350, B => 
                           n18516, ZN => n6256);
   U6038 : NAND2_X1 port map( A1 => n28353, A2 => n6461, ZN => n29351);
   U6053 : NAND3_X2 port map( A1 => n16786, A2 => n1226, A3 => n16785, ZN => 
                           n18107);
   U6058 : XNOR2_X1 port map( A => n25891, B => n5146, ZN => n24487);
   U6063 : NOR2_X2 port map( A1 => n6420, A2 => n6422, ZN => n25891);
   U6091 : XNOR2_X2 port map( A => n29353, B => n22850, ZN => n28182);
   U6125 : INV_X1 port map( A => n22849, ZN => n29353);
   U6133 : NAND3_X1 port map( A1 => n24578, A2 => n24468, A3 => n24582, ZN => 
                           n6421);
   U6181 : NAND2_X1 port map( A1 => n1631, A2 => n24617, ZN => n24024);
   U6204 : AND2_X2 port map( A1 => n29658, A2 => n29659, ZN => n21192);
   U6225 : OR2_X2 port map( A1 => n28337, A2 => n1210, ZN => n6095);
   U6228 : NAND3_X1 port map( A1 => n5669, A2 => n273, A3 => n4235, ZN => n5817
                           );
   U6261 : INV_X1 port map( A => n25659, ZN => n25660);
   U6263 : XNOR2_X1 port map( A => n25296, B => n25297, ZN => n25659);
   U6290 : NAND2_X1 port map( A1 => n15226, A2 => n29355, ZN => n15231);
   U6313 : XNOR2_X1 port map( A => n19687, B => n19688, ZN => n29769);
   U6352 : NAND4_X2 port map( A1 => n5235, A2 => n5232, A3 => n5231, A4 => 
                           n17768, ZN => n19687);
   U6387 : NAND2_X1 port map( A1 => n18511, A2 => n18512, ZN => n18513);
   U6395 : NAND2_X1 port map( A1 => n24236, A2 => n24568, ZN => n23176);
   U6403 : NAND2_X1 port map( A1 => n24643, A2 => n24638, ZN => n24236);
   U6469 : NAND2_X1 port map( A1 => n29356, A2 => n6600, ZN => n6597);
   U6477 : OAI21_X1 port map( B1 => n24162, B2 => n28522, A => n24802, ZN => 
                           n29356);
   U6501 : OAI21_X1 port map( B1 => n23211, B2 => n22985, A => n29357, ZN => 
                           n2621);
   U6516 : NAND3_X1 port map( A1 => n23604, A2 => n23583, A3 => n23578, ZN => 
                           n29357);
   U6550 : NAND2_X1 port map( A1 => n21159, A2 => n20744, ZN => n20746);
   U6568 : NAND2_X1 port map( A1 => n5881, A2 => n29358, ZN => n5885);
   U6596 : NAND3_X1 port map( A1 => n29359, A2 => n19802, A3 => n20631, ZN => 
                           n21464);
   U6613 : NAND2_X1 port map( A1 => n6059, A2 => n20012, ZN => n29359);
   U6615 : NAND2_X1 port map( A1 => n14426, A2 => n4522, ZN => n13704);
   U6643 : NOR2_X2 port map( A1 => n23907, A2 => n3028, ZN => n26055);
   U6644 : NAND3_X2 port map( A1 => n29361, A2 => n3059, A3 => n29360, ZN => 
                           n25577);
   U6666 : NAND2_X1 port map( A1 => n29323, A2 => n24653, ZN => n29360);
   U6676 : OR2_X1 port map( A1 => n24006, A2 => n24653, ZN => n29361);
   U6704 : AND2_X2 port map( A1 => n3231, A2 => n3230, ZN => n28456);
   U6722 : NAND2_X1 port map( A1 => n14413, A2 => n14414, ZN => n14446);
   U6780 : NAND2_X1 port map( A1 => n12481, A2 => n14444, ZN => n14413);
   U6946 : NAND2_X1 port map( A1 => n14754, A2 => n29362, ZN => n16495);
   U6954 : OAI21_X1 port map( B1 => n14750, B2 => n14751, A => n15243, ZN => 
                           n29362);
   U7025 : NAND3_X1 port map( A1 => n5927, A2 => n20141, A3 => n21088, ZN => 
                           n1245);
   U7058 : OAI211_X2 port map( C1 => n23542, C2 => n23541, A => n2326, B => 
                           n712, ZN => n24768);
   U7073 : NAND2_X1 port map( A1 => n29477, A2 => n2070, ZN => n5618);
   U7095 : OR2_X1 port map( A1 => n5023, A2 => n18708, ZN => n863);
   U7100 : NAND2_X1 port map( A1 => n15095, A2 => n15096, ZN => n2497);
   U7184 : NOR2_X1 port map( A1 => n17992, A2 => n17994, ZN => n17881);
   U7195 : OAI22_X1 port map( A1 => n241, A2 => n17339, B1 => n5226, B2 => 
                           n17342, ZN => n17992);
   U7201 : NAND3_X2 port map( A1 => n3648, A2 => n4409, A3 => n4410, ZN => 
                           n22286);
   U7224 : INV_X1 port map( A => n22294, ZN => n22027);
   U7280 : NAND2_X1 port map( A1 => n29364, A2 => n29363, ZN => n22294);
   U7346 : INV_X1 port map( A => n21208, ZN => n29363);
   U7398 : NAND3_X1 port map( A1 => n15293, A2 => n3827, A3 => n15291, ZN => 
                           n14520);
   U7405 : NAND2_X1 port map( A1 => n29366, A2 => n29365, ZN => n26349);
   U7423 : NAND2_X1 port map( A1 => n26347, A2 => n27585, ZN => n29365);
   U7424 : NAND2_X1 port map( A1 => n26348, A2 => n27591, ZN => n29366);
   U7472 : AND2_X2 port map( A1 => n3713, A2 => n29367, ZN => n25826);
   U7491 : INV_X1 port map( A => n29368, ZN => n29367);
   U7492 : OAI21_X1 port map( B1 => n3715, B2 => n464, A => n3714, ZN => n29368
                           );
   U7518 : OAI21_X1 port map( B1 => n23628, B2 => n23632, A => n23040, ZN => 
                           n22277);
   U7528 : NAND3_X1 port map( A1 => n122, A2 => n18087, A3 => n123, ZN => 
                           n28892);
   U7593 : NOR2_X1 port map( A1 => n20616, A2 => n19920, ZN => n20430);
   U7604 : XNOR2_X2 port map( A => n19358, B => n19357, ZN => n20616);
   U7631 : NAND2_X1 port map( A1 => n19825, A2 => n19826, ZN => n1832);
   U7679 : NAND2_X1 port map( A1 => n26567, A2 => n26912, ZN => n4455);
   U7686 : AND3_X2 port map( A1 => n3130, A2 => n3129, A3 => n2431, ZN => 
                           n11640);
   U7745 : NAND2_X1 port map( A1 => n18197, A2 => n18193, ZN => n18194);
   U7772 : NAND2_X1 port map( A1 => n29369, A2 => n6494, ZN => n20749);
   U7789 : NAND2_X1 port map( A1 => n4472, A2 => n19848, ZN => n29369);
   U7809 : NAND3_X1 port map( A1 => n16729, A2 => n2578, A3 => n2579, ZN => 
                           n4705);
   U7815 : OAI22_X2 port map( A1 => n21165, A2 => n21166, B1 => n21326, B2 => 
                           n159, ZN => n22506);
   U7828 : MUX2_X1 port map( A => n29139, B => n11671, S => n11640, Z => n11402
                           );
   U7878 : NAND2_X1 port map( A1 => n5868, A2 => n8523, ZN => n5867);
   U7896 : OAI21_X1 port map( B1 => n24579, B2 => n24578, A => n24469, ZN => 
                           n6422);
   U7963 : XNOR2_X1 port map( A => n29370, B => n2389, ZN => Ciphertext(8));
   U7982 : NAND2_X1 port map( A1 => n1681, A2 => n29278, ZN => n29370);
   U7983 : NAND2_X1 port map( A1 => n11239, A2 => n29371, ZN => n28944);
   U8005 : NAND3_X1 port map( A1 => n11235, A2 => n11237, A3 => n11236, ZN => 
                           n29371);
   U8021 : AND2_X2 port map( A1 => n29372, A2 => n7311, ZN => n9425);
   U8029 : NAND3_X1 port map( A1 => n7307, A2 => n4438, A3 => n4439, ZN => 
                           n29372);
   U8034 : INV_X1 port map( A => n16612, ZN => n29373);
   U8047 : OAI211_X2 port map( C1 => n4539, C2 => n10693, A => n4537, B => 
                           n10692, ZN => n12303);
   U8048 : NAND2_X1 port map( A1 => n8163, A2 => n8164, ZN => n8172);
   U8064 : NAND3_X1 port map( A1 => n747, A2 => n746, A3 => n7895, ZN => n997);
   U8066 : NAND3_X1 port map( A1 => n28839, A2 => n29374, A3 => n28838, ZN => 
                           n11739);
   U8085 : AOI22_X1 port map( A1 => n10612, A2 => n10972, B1 => n10969, B2 => 
                           n5267, ZN => n29374);
   U8104 : NAND2_X1 port map( A1 => n29375, A2 => n196, ZN => n27634);
   U8141 : NAND2_X1 port map( A1 => n2414, A2 => n2415, ZN => n29375);
   U8144 : NAND2_X1 port map( A1 => n16739, A2 => n16738, ZN => n18204);
   U8151 : NAND2_X1 port map( A1 => n8167, A2 => n7298, ZN => n8169);
   U8177 : NAND2_X1 port map( A1 => n29376, A2 => n21463, ZN => n2299);
   U8180 : NAND2_X1 port map( A1 => n4224, A2 => n4223, ZN => n29376);
   U8196 : NAND2_X1 port map( A1 => n29377, A2 => n18260, ZN => n2705);
   U8204 : OAI21_X1 port map( B1 => n17699, B2 => n18535, A => n18259, ZN => 
                           n29377);
   U8264 : OAI21_X1 port map( B1 => n16824, B2 => n17291, A => n28729, ZN => 
                           n28728);
   U8284 : NOR2_X1 port map( A1 => n17395, A2 => n17397, ZN => n17291);
   U8290 : AND2_X2 port map( A1 => n1373, A2 => n1656, ZN => n18241);
   U8291 : NAND2_X1 port map( A1 => n29433, A2 => n6464, ZN => n29432);
   U8293 : OR2_X2 port map( A1 => n17608, A2 => n3847, ZN => n18799);
   U8295 : NAND3_X1 port map( A1 => n6020, A2 => n11702, A3 => n4844, ZN => 
                           n11705);
   U8314 : NAND3_X1 port map( A1 => n11952, A2 => n11944, A3 => n11943, ZN => 
                           n2440);
   U8323 : NAND2_X1 port map( A1 => n4455, A2 => n29378, ZN => n1021);
   U8371 : NAND2_X1 port map( A1 => n26786, A2 => n26565, ZN => n29378);
   U8375 : INV_X1 port map( A => n14633, ZN => n14722);
   U8383 : NAND2_X1 port map( A1 => n29379, A2 => n15389, ZN => n14634);
   U8446 : NAND2_X1 port map( A1 => n14633, A2 => n29380, ZN => n29379);
   U8459 : NAND2_X1 port map( A1 => n14992, A2 => n15387, ZN => n14633);
   U8479 : NAND2_X1 port map( A1 => n28871, A2 => n28817, ZN => n29787);
   U8482 : NOR2_X2 port map( A1 => n29382, A2 => n29381, ZN => n25386);
   U8487 : OAI22_X1 port map( A1 => n24311, A2 => n24390, B1 => n24312, B2 => 
                           n2649, ZN => n29381);
   U8513 : AND2_X1 port map( A1 => n24314, A2 => n24682, ZN => n29382);
   U8528 : NAND2_X1 port map( A1 => n28901, A2 => n18083, ZN => n28900);
   U8541 : OR2_X1 port map( A1 => n19938, A2 => n19810, ZN => n29706);
   U8544 : OAI211_X1 port map( C1 => n4232, C2 => n23140, A => n23012, B => 
                           n29383, ZN => n23014);
   U8550 : NAND3_X1 port map( A1 => n23011, A2 => n4232, A3 => n23351, ZN => 
                           n29383);
   U8575 : NOR2_X2 port map( A1 => n3732, A2 => n5972, ZN => n13262);
   U8597 : OR2_X1 port map( A1 => n17155, A2 => n17336, ZN => n6336);
   U8603 : OAI21_X1 port map( B1 => n27443, B2 => n26833, A => n26832, ZN => 
                           n26834);
   U8605 : NAND3_X1 port map( A1 => n20982, A2 => n21008, A3 => n21809, ZN => 
                           n2259);
   U8606 : NAND2_X1 port map( A1 => n3637, A2 => n29384, ZN => n7693);
   U8619 : NAND3_X1 port map( A1 => n7691, A2 => n7818, A3 => n7690, ZN => 
                           n29384);
   U8631 : NOR2_X1 port map( A1 => n17900, A2 => n29322, ZN => n29386);
   U8632 : NAND3_X1 port map( A1 => n29541, A2 => n28562, A3 => n29387, ZN => 
                           n5359);
   U8637 : NAND4_X2 port map( A1 => n6882, A2 => n6881, A3 => n20260, A4 => 
                           n6883, ZN => n5151);
   U8640 : XNOR2_X1 port map( A => n16255, B => n16126, ZN => n16499);
   U8642 : NAND3_X2 port map( A1 => n15325, A2 => n3626, A3 => n3627, ZN => 
                           n16255);
   U8647 : NAND2_X1 port map( A1 => n25649, A2 => n29388, ZN => n25975);
   U8661 : OAI211_X2 port map( C1 => n6341, C2 => n6113, A => n29233, B => 
                           n29739, ZN => n20786);
   U8668 : NAND3_X1 port map( A1 => n5084, A2 => n5083, A3 => n6484, ZN => 
                           n5082);
   U8669 : NAND2_X1 port map( A1 => n23426, A2 => n23339, ZN => n6197);
   U8697 : NAND3_X1 port map( A1 => n4133, A2 => n26816, A3 => n29389, ZN => 
                           n4925);
   U8726 : NAND3_X1 port map( A1 => n3440, A2 => n623, A3 => n3439, ZN => n1729
                           );
   U8740 : NAND2_X1 port map( A1 => n4545, A2 => n521, ZN => n3440);
   U8741 : NAND2_X1 port map( A1 => n29390, A2 => n1202, ZN => n23967);
   U8762 : NAND2_X1 port map( A1 => n23965, A2 => n24582, ZN => n29390);
   U8772 : NAND2_X1 port map( A1 => n28133, A2 => n28610, ZN => n20328);
   U8773 : NAND2_X1 port map( A1 => n29391, A2 => n21163, ZN => n20731);
   U8784 : INV_X1 port map( A => n21162, ZN => n29391);
   U8826 : NAND2_X1 port map( A1 => n21334, A2 => n21612, ZN => n21162);
   U8833 : AND3_X2 port map( A1 => n29392, A2 => n26383, A3 => n1029, ZN => 
                           n27551);
   U8851 : NAND2_X1 port map( A1 => n26379, A2 => n26425, ZN => n29392);
   U8856 : NAND2_X1 port map( A1 => n28860, A2 => n28861, ZN => n7639);
   U8858 : NAND2_X1 port map( A1 => n8611, A2 => n29394, ZN => n29393);
   U8885 : NAND2_X1 port map( A1 => n9532, A2 => n29395, ZN => n29394);
   U8905 : OR2_X1 port map( A1 => n9037, A2 => n8792, ZN => n3353);
   U8906 : XNOR2_X1 port map( A => n19462, B => n19299, ZN => n19077);
   U8916 : NAND2_X2 port map( A1 => n6036, A2 => n28877, ZN => n19462);
   U8920 : NOR2_X2 port map( A1 => n16988, A2 => n29396, ZN => n19408);
   U8932 : NAND2_X1 port map( A1 => n28892, A2 => n2444, ZN => n29396);
   U8938 : AND3_X2 port map( A1 => n1299, A2 => n6597, A3 => n6595, ZN => 
                           n25928);
   U8944 : AND2_X2 port map( A1 => n1462, A2 => n1460, ZN => n21410);
   U8955 : NAND2_X1 port map( A1 => n12990, A2 => n12150, ZN => n12994);
   U8984 : INV_X1 port map( A => n10793, ZN => n12990);
   U8986 : NAND3_X2 port map( A1 => n29397, A2 => n23451, A3 => n23452, ZN => 
                           n24972);
   U8987 : OAI21_X1 port map( B1 => n23444, B2 => n23443, A => n4794, ZN => 
                           n29397);
   U9007 : NAND2_X1 port map( A1 => n1249, A2 => n1250, ZN => n24153);
   U9035 : NAND3_X1 port map( A1 => n29398, A2 => n26210, A3 => n26209, ZN => 
                           n29657);
   U9049 : NAND2_X1 port map( A1 => n26723, A2 => n26208, ZN => n29398);
   U9085 : OAI21_X1 port map( B1 => n24248, B2 => n24523, A => n24030, ZN => 
                           n24006);
   U9088 : NAND2_X1 port map( A1 => n28785, A2 => n24248, ZN => n24030);
   U9147 : NAND2_X1 port map( A1 => n3145, A2 => n1078, ZN => n22681);
   U9180 : NAND2_X1 port map( A1 => n3701, A2 => n18505, ZN => n18517);
   U9194 : OAI21_X1 port map( B1 => n26772, B2 => n26771, A => n29399, ZN => 
                           n26773);
   U9202 : NAND3_X1 port map( A1 => n28421, A2 => n26768, A3 => n26935, ZN => 
                           n29399);
   U9227 : NAND2_X1 port map( A1 => n26940, A2 => n26941, ZN => n26772);
   U9244 : XNOR2_X1 port map( A => n25134, B => n25133, ZN => n25136);
   U9247 : AND2_X2 port map( A1 => n29401, A2 => n29400, ZN => n25133);
   U9255 : NAND2_X1 port map( A1 => n24149, A2 => n29050, ZN => n29400);
   U9274 : NAND2_X1 port map( A1 => n23935, A2 => n24744, ZN => n29401);
   U9291 : NAND3_X1 port map( A1 => n29403, A2 => n760, A3 => n29402, ZN => 
                           n23616);
   U9307 : INV_X1 port map( A => n476, ZN => n29403);
   U9321 : NAND2_X1 port map( A1 => n29404, A2 => n19931, ZN => n4268);
   U9322 : NAND2_X1 port map( A1 => n19573, A2 => n6205, ZN => n29404);
   U9323 : NAND2_X1 port map( A1 => n23363, A2 => n23673, ZN => n23361);
   U9328 : NAND2_X1 port map( A1 => n29407, A2 => n29405, ZN => n16602);
   U9345 : NAND2_X1 port map( A1 => n17106, A2 => n29406, ZN => n29405);
   U9356 : NAND2_X1 port map( A1 => n17083, A2 => n17470, ZN => n29407);
   U9357 : NAND3_X1 port map( A1 => n29408, A2 => n28208, A3 => n4107, ZN => 
                           n248);
   U9359 : NAND2_X1 port map( A1 => n11331, A2 => n11169, ZN => n29408);
   U9367 : XNOR2_X1 port map( A => n29409, B => Key(13), ZN => Ciphertext(128))
                           ;
   U9378 : NAND2_X1 port map( A1 => n96, A2 => n26341, ZN => n29409);
   U9384 : NAND2_X1 port map( A1 => n29411, A2 => n8500, ZN => n8115);
   U9482 : INV_X1 port map( A => n8116, ZN => n29411);
   U9490 : OAI211_X2 port map( C1 => n11894, C2 => n10794, A => n10798, B => 
                           n29412, ZN => n12088);
   U9492 : NAND2_X1 port map( A1 => n10796, A2 => n11893, ZN => n29412);
   U9497 : XNOR2_X1 port map( A => n29413, B => n27534, ZN => Ciphertext(58));
   U9499 : NAND2_X1 port map( A1 => n27532, A2 => n27533, ZN => n29413);
   U9504 : NAND2_X1 port map( A1 => n29415, A2 => n29414, ZN => n7908);
   U9528 : NAND2_X1 port map( A1 => n8652, A2 => n8500, ZN => n29414);
   U9533 : NAND2_X1 port map( A1 => n8655, A2 => n29416, ZN => n29415);
   U9535 : NAND3_X1 port map( A1 => n28912, A2 => n16926, A3 => n15069, ZN => 
                           n29674);
   U9542 : NAND3_X1 port map( A1 => n23584, A2 => n23710, A3 => n380, ZN => 
                           n6154);
   U9549 : NAND2_X1 port map( A1 => n29418, A2 => n29332, ZN => n27387);
   U9585 : NOR2_X1 port map( A1 => n27392, A2 => n29419, ZN => n29418);
   U9632 : NOR2_X1 port map( A1 => n25621, A2 => n6685, ZN => n29419);
   U9638 : OAI211_X1 port map( C1 => n4681, C2 => n6465, A => n29421, B => 
                           n29420, ZN => n5107);
   U9644 : NAND2_X1 port map( A1 => n4681, A2 => n17277, ZN => n29420);
   U9678 : XNOR2_X2 port map( A => n5433, B => n5434, ZN => n26935);
   U9719 : NAND3_X1 port map( A1 => n11705, A2 => n6073, A3 => n29422, ZN => 
                           n3438);
   U9729 : NAND2_X1 port map( A1 => n12205, A2 => n11703, ZN => n29422);
   U9737 : NAND2_X1 port map( A1 => n16791, A2 => n16792, ZN => n17798);
   U9774 : NAND2_X1 port map( A1 => n20025, A2 => n20026, ZN => n21632);
   U9781 : OR2_X1 port map( A1 => n10544, A2 => n11149, ZN => n1064);
   U9794 : NAND2_X1 port map( A1 => n24113, A2 => n24111, ZN => n23870);
   U9840 : NOR2_X1 port map( A1 => n19656, A2 => n19659, ZN => n19606);
   U9842 : NAND3_X1 port map( A1 => n7580, A2 => n7887, A3 => n7581, ZN => 
                           n7083);
   U9874 : OAI21_X1 port map( B1 => n9211, B2 => n8995, A => n8994, ZN => n8436
                           );
   U9883 : NAND2_X1 port map( A1 => n9211, A2 => n8996, ZN => n8994);
   U9888 : NAND3_X1 port map( A1 => n29424, A2 => n29423, A3 => n11112, ZN => 
                           n2351);
   U9907 : NAND2_X1 port map( A1 => n5109, A2 => n11111, ZN => n29423);
   U9909 : NAND2_X1 port map( A1 => n243, A2 => n242, ZN => n29424);
   U9917 : NAND2_X1 port map( A1 => n16715, A2 => n16716, ZN => n18197);
   U9961 : OAI211_X1 port map( C1 => n17196, C2 => n29546, A => n16714, B => 
                           n4283, ZN => n16715);
   U10012 : AOI21_X1 port map( B1 => n29427, B2 => n29426, A => n20008, ZN => 
                           n20010);
   U10030 : NAND2_X1 port map( A1 => n4991, A2 => n6156, ZN => n29427);
   U10032 : AND2_X1 port map( A1 => n6309, A2 => n24726, ZN => n4749);
   U10059 : NAND3_X1 port map( A1 => n17339, A2 => n17340, A3 => n17338, ZN => 
                           n17341);
   U10063 : OAI21_X1 port map( B1 => n26532, B2 => n26528, A => n29331, ZN => 
                           n29168);
   U10068 : NAND2_X1 port map( A1 => n29429, A2 => n29428, ZN => n19801);
   U10070 : NAND2_X1 port map( A1 => n19800, A2 => n29601, ZN => n29428);
   U10077 : NAND2_X1 port map( A1 => n19799, A2 => n1624, ZN => n29429);
   U10110 : NAND2_X1 port map( A1 => n29431, A2 => n29430, ZN => n15767);
   U10121 : NAND2_X1 port map( A1 => n532, A2 => n17316, ZN => n29430);
   U10139 : NAND2_X1 port map( A1 => n790, A2 => n17562, ZN => n29431);
   U10157 : NOR2_X2 port map( A1 => n6635, A2 => n19801, ZN => n21465);
   U10159 : XNOR2_X1 port map( A => n29432, B => n26287, ZN => Ciphertext(84));
   U10187 : OR2_X1 port map( A1 => n26286, A2 => n26346, ZN => n29433);
   U10195 : OAI21_X1 port map( B1 => n325, B2 => n27711, A => n29434, ZN => 
                           n27713);
   U10200 : NAND2_X1 port map( A1 => n325, A2 => n27716, ZN => n29434);
   U10207 : NAND2_X1 port map( A1 => n28958, A2 => n21467, ZN => n29435);
   U10208 : OAI21_X1 port map( B1 => n29437, B2 => n1931, A => n29436, ZN => 
                           n12106);
   U10212 : NAND2_X1 port map( A1 => n12104, A2 => n1931, ZN => n29436);
   U10225 : NOR2_X1 port map( A1 => n11656, A2 => n12162, ZN => n29437);
   U10263 : NAND3_X1 port map( A1 => n23296, A2 => n29020, A3 => n22864, ZN => 
                           n5712);
   U10283 : NAND2_X1 port map( A1 => n23837, A2 => n23391, ZN => n23281);
   U10291 : NAND3_X1 port map( A1 => n8027, A2 => n8029, A3 => n8028, ZN => 
                           n29464);
   U10325 : NAND2_X1 port map( A1 => n29438, A2 => n724, ZN => n22393);
   U10385 : NAND2_X1 port map( A1 => n726, A2 => n22392, ZN => n29438);
   U10452 : NOR2_X1 port map( A1 => n27286, A2 => n27287, ZN => n26811);
   U10455 : NOR2_X2 port map( A1 => n26795, A2 => n26796, ZN => n27287);
   U10472 : NAND3_X1 port map( A1 => n8465, A2 => n8464, A3 => n8826, ZN => 
                           n29439);
   U10477 : MUX2_X1 port map( A => n18398, B => n18231, S => n18233, Z => 
                           n18235);
   U10540 : NAND4_X2 port map( A1 => n4987, A2 => n4988, A3 => n5459, A4 => 
                           n5458, ZN => n18233);
   U10546 : OR2_X2 port map( A1 => n29440, A2 => n17922, ZN => n19413);
   U10580 : AOI21_X1 port map( B1 => n17919, B2 => n17920, A => n18357, ZN => 
                           n29440);
   U10616 : NAND3_X2 port map( A1 => n29441, A2 => n5979, A3 => n5977, ZN => 
                           n15447);
   U10623 : NAND3_X1 port map( A1 => n29201, A2 => n28805, A3 => n5980, ZN => 
                           n29441);
   U10632 : NAND2_X1 port map( A1 => n26404, A2 => n29442, ZN => n26406);
   U10633 : NAND3_X1 port map( A1 => n2433, A2 => n29444, A3 => n29443, ZN => 
                           n29442);
   U10645 : NAND2_X1 port map( A1 => n27553, A2 => n27551, ZN => n29443);
   U10649 : NAND2_X1 port map( A1 => n27552, A2 => n29445, ZN => n29444);
   U10650 : NAND2_X1 port map( A1 => n1120, A2 => n1122, ZN => n29203);
   U10653 : NAND2_X1 port map( A1 => n29446, A2 => n7235, ZN => n6382);
   U10661 : OAI21_X1 port map( B1 => n7232, B2 => n6384, A => n2833, ZN => 
                           n29446);
   U10664 : INV_X1 port map( A => n25617, ZN => n27394);
   U10688 : OAI211_X2 port map( C1 => n19982, C2 => n18886, A => n18884, B => 
                           n18885, ZN => n21288);
   U10697 : NAND2_X1 port map( A1 => n29448, A2 => n29447, ZN => n27666);
   U10705 : NAND2_X1 port map( A1 => n27664, A2 => n27663, ZN => n29447);
   U10718 : NAND2_X1 port map( A1 => n29450, A2 => n29449, ZN => n29448);
   U10751 : NAND2_X1 port map( A1 => n27674, A2 => n28655, ZN => n29450);
   U10753 : INV_X1 port map( A => Plaintext(169), ZN => n29451);
   U10761 : INV_X1 port map( A => n21971, ZN => n22555);
   U10763 : XNOR2_X1 port map( A => n21801, B => n20798, ZN => n21971);
   U10764 : AND2_X2 port map( A1 => n29453, A2 => n29452, ZN => n21364);
   U10773 : NAND2_X1 port map( A1 => n19240, A2 => n28489, ZN => n29452);
   U10785 : NAND2_X1 port map( A1 => n19241, A2 => n20511, ZN => n29453);
   U10789 : NAND2_X1 port map( A1 => n26373, A2 => n26266, ZN => n29454);
   U10818 : NAND2_X1 port map( A1 => n14101, A2 => n14105, ZN => n6563);
   U10821 : NAND2_X1 port map( A1 => n29455, A2 => n113, ZN => n4803);
   U10864 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => n29455);
   U10885 : NAND2_X1 port map( A1 => n21184, A2 => n21497, ZN => n21186);
   U10888 : XNOR2_X2 port map( A => n21891, B => n21892, ZN => n23800);
   U10893 : NAND2_X1 port map( A1 => n27386, A2 => n27410, ZN => n27388);
   U10927 : NOR2_X2 port map( A1 => n25626, A2 => n4013, ZN => n27410);
   U10933 : OAI21_X1 port map( B1 => n23342, B2 => n23428, A => n29456, ZN => 
                           n23346);
   U10938 : NAND3_X1 port map( A1 => n23341, A2 => n23340, A3 => n28570, ZN => 
                           n29456);
   U10959 : OAI21_X1 port map( B1 => n530, B2 => n29636, A => n29457, ZN => 
                           n17164);
   U10997 : NAND2_X1 port map( A1 => n17374, A2 => n29635, ZN => n29457);
   U11012 : AND2_X1 port map( A1 => n20158, A2 => n20157, ZN => n19769);
   U11013 : NAND2_X1 port map( A1 => n4433, A2 => n4434, ZN => n4432);
   U11038 : NAND2_X1 port map( A1 => n2777, A2 => n739, ZN => n2774);
   U11052 : NAND2_X1 port map( A1 => n19772, A2 => n19771, ZN => n21144);
   U11060 : NAND2_X1 port map( A1 => n22963, A2 => n22964, ZN => n4672);
   U11070 : NAND3_X1 port map( A1 => n23696, A2 => n23693, A3 => n4086, ZN => 
                           n5480);
   U11083 : INV_X1 port map( A => n20814, ZN => n21266);
   U11114 : MUX2_X1 port map( A => n20878, B => n21269, S => n20814, Z => 
                           n18851);
   U11176 : NAND2_X1 port map( A1 => n29459, A2 => n29458, ZN => n798);
   U11215 : NAND2_X1 port map( A1 => n26204, A2 => n26235, ZN => n29458);
   U11224 : OR3_X1 port map( A1 => n17439, A2 => n17437, A3 => n17433, ZN => 
                           n1387);
   U11238 : OAI22_X1 port map( A1 => n11228, A2 => n29461, B1 => n11232, B2 => 
                           n11231, ZN => n29460);
   U11248 : NOR2_X1 port map( A1 => n11229, A2 => n11896, ZN => n29462);
   U11296 : NAND3_X1 port map( A1 => n3367, A2 => n3366, A3 => n29463, ZN => 
                           n196);
   U11301 : NAND3_X1 port map( A1 => n3153, A2 => n18063, A3 => n17672, ZN => 
                           n4347);
   U11334 : XNOR2_X1 port map( A => n26102, B => n3256, ZN => n26103);
   U11352 : AOI22_X2 port map( A1 => n24197, A2 => n6238, B1 => n24196, B2 => 
                           n6239, ZN => n26102);
   U11361 : NAND3_X2 port map( A1 => n29464, A2 => n8031, A3 => n4061, ZN => 
                           n9124);
   U11436 : OAI211_X2 port map( C1 => n5382, C2 => n15105, A => n5379, B => 
                           n29465, ZN => n16229);
   U11506 : NAND2_X1 port map( A1 => n5381, A2 => n15105, ZN => n29465);
   U11566 : NAND2_X1 port map( A1 => n28725, A2 => n11964, ZN => n29466);
   U11595 : NAND2_X1 port map( A1 => n11998, A2 => n11536, ZN => n11685);
   U11602 : AOI22_X2 port map( A1 => n10552, A2 => n10551, B1 => n10550, B2 => 
                           n10461, ZN => n11998);
   U11691 : AOI22_X2 port map( A1 => n18973, A2 => n2096, B1 => n18974, B2 => 
                           n19060, ZN => n21290);
   U11726 : BUF_X1 port map( A => n14416, Z => n29638);
   U11728 : XOR2_X1 port map( A => n23919, B => n23920, Z => n29467);
   U11731 : NAND2_X1 port map( A1 => n29696, A2 => n26164, ZN => n29468);
   U11736 : OR2_X1 port map( A1 => n26519, A2 => n29633, ZN => n27690);
   U11749 : NOR2_X1 port map( A1 => n26312, A2 => n6669, ZN => n27777);
   U11766 : NAND2_X1 port map( A1 => n29696, A2 => n26164, ZN => n27463);
   U11768 : INV_X1 port map( A => n26177, ZN => n29697);
   U11797 : XNOR2_X1 port map( A => n9856, B => n9855, ZN => n10983);
   U11811 : AND2_X1 port map( A1 => n26337, A2 => n5485, ZN => n29469);
   U11838 : BUF_X2 port map( A => n24078, Z => n29470);
   U11900 : MUX2_X1 port map( A => n23900, B => n23899, S => n24688, Z => 
                           n23904);
   U11975 : OAI21_X1 port map( B1 => n26160, B2 => n26161, A => n29697, ZN => 
                           n29696);
   U12001 : XNOR2_X1 port map( A => n24910, B => n24909, ZN => n27191);
   U12042 : AND2_X1 port map( A1 => n2263, A2 => n29472, ZN => n28590);
   U12043 : AND2_X1 port map( A1 => n2262, A2 => n29473, ZN => n29472);
   U12083 : INV_X1 port map( A => n26724, ZN => n29473);
   U12148 : XNOR2_X1 port map( A => n26049, B => n26050, ZN => n29474);
   U12155 : OR2_X1 port map( A1 => n27780, A2 => n29070, ZN => n29475);
   U12163 : XNOR2_X1 port map( A => n26049, B => n26050, ZN => n27110);
   U12164 : OR2_X1 port map( A1 => n29649, A2 => n14278, ZN => n4163);
   U12182 : OR2_X1 port map( A1 => n15420, A2 => n15103, ZN => n15419);
   U12228 : AND2_X1 port map( A1 => n16952, A2 => n17354, ZN => n29476);
   U12258 : XNOR2_X1 port map( A => n15638, B => n15637, ZN => n17354);
   U12260 : AOI22_X1 port map( A1 => n6610, A2 => n23390, B1 => n6279, B2 => 
                           n23837, ZN => n29477);
   U12296 : OR2_X1 port map( A1 => n27310, A2 => n29478, ZN => n29701);
   U12303 : OR2_X1 port map( A1 => n29493, A2 => n27308, ZN => n29478);
   U12327 : NAND2_X1 port map( A1 => n29748, A2 => n10865, ZN => n13552);
   U12363 : XOR2_X1 port map( A => n25258, B => n25259, Z => n29479);
   U12389 : NAND3_X1 port map( A1 => n6627, A2 => n26759, A3 => n6626, ZN => 
                           n29480);
   U12417 : XNOR2_X1 port map( A => n25594, B => n25593, ZN => n29481);
   U12419 : XOR2_X1 port map( A => n25594, B => n25593, Z => n29482);
   U12427 : AND2_X1 port map( A1 => n23097, A2 => n2452, ZN => n3612);
   U12429 : BUF_X2 port map( A => n27128, Z => n397);
   U12435 : XOR2_X1 port map( A => n15665, B => n15664, Z => n29483);
   U12437 : AND4_X1 port map( A1 => n17578, A2 => n3086, A3 => n3085, A4 => 
                           n3084, ZN => n29484);
   U12449 : INV_X1 port map( A => n17534, ZN => n18243);
   U12463 : OAI21_X1 port map( B1 => n24607, B2 => n24606, A => n24605, ZN => 
                           n29485);
   U12479 : OAI21_X1 port map( B1 => n24607, B2 => n24606, A => n24605, ZN => 
                           n25754);
   U12501 : INV_X1 port map( A => n11955, ZN => n571);
   U12505 : OR2_X1 port map( A1 => n26997, A2 => n26998, ZN => n29486);
   U12506 : XNOR2_X2 port map( A => n25568, B => n25567, ZN => n26998);
   U12562 : XNOR2_X1 port map( A => n24971, B => n24970, ZN => n1907);
   U12568 : AND2_X1 port map( A1 => n2263, A2 => n29472, ZN => n28115);
   U12580 : BUF_X1 port map( A => n25597, Z => n26229);
   U12585 : XNOR2_X1 port map( A => n24915, B => n24914, ZN => n27124);
   U12625 : INV_X1 port map( A => n24666, ZN => n29754);
   U12656 : OAI21_X1 port map( B1 => n1391, B2 => n1642, A => n1390, ZN => 
                           n24237);
   U12673 : OAI211_X1 port map( C1 => n20641, C2 => n1908, A => n19790, B => 
                           n19789, ZN => n21113);
   U12675 : AOI21_X1 port map( B1 => n21197, B2 => n21196, A => n21195, ZN => 
                           n29489);
   U12678 : AOI21_X1 port map( B1 => n21197, B2 => n21196, A => n21195, ZN => 
                           n29490);
   U12697 : AOI21_X1 port map( B1 => n21197, B2 => n21196, A => n21195, ZN => 
                           n22428);
   U12726 : INV_X1 port map( A => n3911, ZN => n29491);
   U12737 : BUF_X1 port map( A => n18845, Z => n19765);
   U12782 : OR2_X1 port map( A1 => n22286, A2 => n21213, ZN => n20666);
   U12849 : MUX2_X1 port map( A => n19989, B => n20165, S => n19993, Z => 
                           n19862);
   U12890 : BUF_X1 port map( A => n26717, Z => n283);
   U12892 : NAND3_X1 port map( A1 => n4516, A2 => n28, A3 => n27, ZN => n29492)
                           ;
   U12893 : NAND3_X1 port map( A1 => n4516, A2 => n28, A3 => n27, ZN => n18756)
                           ;
   U12905 : OR2_X1 port map( A1 => n4118, A2 => n17569, ZN => n17228);
   U12929 : OAI211_X1 port map( C1 => n11375, C2 => n11831, A => n3685, B => 
                           n3684, ZN => n29494);
   U12947 : OAI211_X1 port map( C1 => n11375, C2 => n11831, A => n3685, B => 
                           n3684, ZN => n29495);
   U12964 : OAI211_X1 port map( C1 => n11375, C2 => n11831, A => n3685, B => 
                           n3684, ZN => n13401);
   U12993 : NAND2_X1 port map( A1 => n18071, A2 => n18070, ZN => n29496);
   U13016 : XNOR2_X1 port map( A => n25907, B => n25906, ZN => n29497);
   U13017 : NAND2_X1 port map( A1 => n4095, A2 => n5717, ZN => n29498);
   U13033 : NAND2_X1 port map( A1 => n4095, A2 => n5717, ZN => n29499);
   U13039 : XNOR2_X1 port map( A => n3168, B => n25712, ZN => n29500);
   U13057 : XNOR2_X1 port map( A => n25236, B => n25235, ZN => n26728);
   U13068 : AND2_X1 port map( A1 => n16716, A2 => n16715, ZN => n29502);
   U13089 : XNOR2_X1 port map( A => n25681, B => n25396, ZN => n25807);
   U13094 : CLKBUF_X1 port map( A => n27871, Z => n29504);
   U13112 : BUF_X1 port map( A => n23874, Z => n24470);
   U13116 : OAI21_X1 port map( B1 => n29227, B2 => n21378, A => n29329, ZN => 
                           n29652);
   U13130 : XOR2_X1 port map( A => n16171, B => n15920, Z => n15924);
   U13153 : NAND4_X1 port map( A1 => n4076, A2 => n4077, A3 => n4075, A4 => 
                           n16694, ZN => n29505);
   U13174 : NAND4_X1 port map( A1 => n4076, A2 => n4077, A3 => n4075, A4 => 
                           n16694, ZN => n29506);
   U13175 : NAND4_X1 port map( A1 => n4076, A2 => n4077, A3 => n4075, A4 => 
                           n16694, ZN => n19707);
   U13180 : OAI211_X1 port map( C1 => n4865, C2 => n4866, A => n4864, B => 
                           n29738, ZN => n29507);
   U13196 : XNOR2_X1 port map( A => n6804, B => n19730, ZN => n29508);
   U13259 : OAI211_X1 port map( C1 => n4865, C2 => n4866, A => n4864, B => 
                           n29738, ZN => n18422);
   U13378 : XNOR2_X1 port map( A => n6804, B => n19730, ZN => n20437);
   U13379 : INV_X1 port map( A => n10383, ZN => n29509);
   U13386 : CLKBUF_X1 port map( A => n28174, Z => n29510);
   U13392 : AND2_X1 port map( A1 => n1907, A2 => n26387, ZN => n27167);
   U13397 : CLKBUF_X1 port map( A => n16449, Z => n29511);
   U13419 : OR2_X1 port map( A1 => n21303, A2 => n24745, ZN => n29512);
   U13421 : CLKBUF_X1 port map( A => n17571, Z => n29513);
   U13441 : OAI21_X1 port map( B1 => n21336, B2 => n21337, A => n21335, ZN => 
                           n29514);
   U13453 : OAI21_X1 port map( B1 => n21336, B2 => n21337, A => n21335, ZN => 
                           n22668);
   U13486 : CLKBUF_X1 port map( A => n27418, Z => n29515);
   U13513 : XOR2_X1 port map( A => n26972, B => n24166, Z => Ciphertext(27));
   U13524 : NAND2_X1 port map( A1 => n856, A2 => n18274, ZN => n19320);
   U13539 : OR2_X1 port map( A1 => n5540, A2 => n6268, ZN => n25203);
   U13584 : OAI21_X1 port map( B1 => n4955, B2 => n4957, A => n14110, ZN => 
                           n29516);
   U13601 : MUX2_X2 port map( A => n26226, B => n26225, S => n25453, Z => 
                           n28069);
   U13649 : CLKBUF_X1 port map( A => n27629, Z => n27626);
   U13663 : AOI21_X1 port map( B1 => n25241, B2 => n25240, A => n26464, ZN => 
                           n25242);
   U13664 : INV_X1 port map( A => n25065, ZN => n26114);
   U13667 : BUF_X1 port map( A => n23261, Z => n23715);
   U13668 : AND2_X2 port map( A1 => n5365, A2 => n16923, ZN => n18324);
   U13695 : XNOR2_X1 port map( A => n10430, B => n10429, ZN => n29517);
   U13699 : XNOR2_X1 port map( A => n10430, B => n10429, ZN => n11206);
   U13700 : OAI211_X2 port map( C1 => n23143, C2 => n4772, A => n3886, B => 
                           n2058, ZN => n24891);
   U13780 : OAI211_X1 port map( C1 => n20615, C2 => n20614, A => n20613, B => 
                           n20612, ZN => n21600);
   U13789 : XNOR2_X1 port map( A => n29485, B => n25714, ZN => n29518);
   U13819 : INV_X1 port map( A => n26614, ZN => n29520);
   U13840 : AOI22_X1 port map( A1 => n21115, A2 => n1897, B1 => n21114, B2 => 
                           n21463, ZN => n22410);
   U13871 : CLKBUF_X1 port map( A => n19785, Z => n29521);
   U13888 : NAND2_X1 port map( A1 => n26571, A2 => n26570, ZN => n29522);
   U13931 : NAND2_X1 port map( A1 => n26571, A2 => n26570, ZN => n29523);
   U13952 : NAND2_X1 port map( A1 => n26571, A2 => n26570, ZN => n27498);
   U13971 : XNOR2_X1 port map( A => n10282, B => n9648, ZN => n9748);
   U13981 : XOR2_X1 port map( A => n25518, B => n25519, Z => n29524);
   U13990 : AND2_X1 port map( A1 => n26227, A2 => n28063, ZN => n28055);
   U13992 : AOI21_X1 port map( B1 => n20298, B2 => n19903, A => n19902, ZN => 
                           n21459);
   U14000 : OAI211_X1 port map( C1 => n1809, C2 => n15170, A => n14553, B => 
                           n14552, ZN => n29525);
   U14073 : OAI211_X1 port map( C1 => n19058, C2 => n20056, A => n19056, B => 
                           n19057, ZN => n29526);
   U14123 : OAI211_X1 port map( C1 => n19058, C2 => n20056, A => n19056, B => 
                           n19057, ZN => n21277);
   U14129 : XNOR2_X1 port map( A => n19100, B => n19099, ZN => n20484);
   U14131 : XNOR2_X1 port map( A => n24130, B => n24131, ZN => n29528);
   U14147 : OR2_X1 port map( A1 => n26479, A2 => n26478, ZN => n29529);
   U14169 : XNOR2_X1 port map( A => n21456, B => n21455, ZN => n29108);
   U14257 : NAND2_X1 port map( A1 => n3551, A2 => n20301, ZN => n29530);
   U14276 : OAI21_X2 port map( B1 => n24993, B2 => n29487, A => n24992, ZN => 
                           n29532);
   U14294 : OAI21_X1 port map( B1 => n24993, B2 => n29487, A => n24992, ZN => 
                           n26671);
   U14370 : AOI21_X1 port map( B1 => n23204, B2 => n28596, A => n23203, ZN => 
                           n29533);
   U14381 : AOI21_X1 port map( B1 => n23204, B2 => n28596, A => n23203, ZN => 
                           n29534);
   U14406 : OR2_X1 port map( A1 => n28403, A2 => n27818, ZN => n29535);
   U14412 : XNOR2_X2 port map( A => n18797, B => n18796, ZN => n20155);
   U14499 : BUF_X1 port map( A => n26299, Z => n29536);
   U14529 : OAI22_X1 port map( A1 => n26300, A2 => n29497, B1 => n26301, B2 => 
                           n27060, ZN => n29537);
   U14594 : OAI22_X1 port map( A1 => n26300, A2 => n29497, B1 => n26301, B2 => 
                           n27060, ZN => n27773);
   U14652 : OR2_X1 port map( A1 => n25238, A2 => n25237, ZN => n29538);
   U14684 : OR2_X1 port map( A1 => n25238, A2 => n25237, ZN => n25998);
   U14689 : XNOR2_X1 port map( A => n16074, B => n16073, ZN => n29539);
   U14734 : OAI211_X1 port map( C1 => n19751, C2 => n28637, A => n4361, B => 
                           n3443, ZN => n29540);
   U14798 : XNOR2_X1 port map( A => n16074, B => n16073, ZN => n16541);
   U14835 : OAI211_X1 port map( C1 => n19751, C2 => n28637, A => n4361, B => 
                           n3443, ZN => n21625);
   U14864 : NAND2_X2 port map( A1 => n28680, A2 => n28217, ZN => n28015);
   U14882 : NOR2_X2 port map( A1 => n25243, A2 => n25242, ZN => n29541);
   U14902 : NOR2_X1 port map( A1 => n25243, A2 => n25242, ZN => n27371);
   U14919 : AND3_X1 port map( A1 => n26453, A2 => n6736, A3 => n2043, ZN => 
                           n27424);
   U14953 : BUF_X1 port map( A => n26119, Z => n29543);
   U14954 : AOI22_X1 port map( A1 => n23924, A2 => n24017, B1 => n459, B2 => 
                           n23923, ZN => n26119);
   U15041 : OR2_X1 port map( A1 => n20017, A2 => n20349, ZN => n20513);
   U15049 : XNOR2_X1 port map( A => n20960, B => n20959, ZN => n29544);
   U15051 : OR2_X1 port map( A1 => n21060, A2 => n21059, ZN => n29545);
   U15080 : XNOR2_X1 port map( A => n20960, B => n20959, ZN => n23683);
   U15085 : INV_X1 port map( A => n7404, ZN => n742);
   U15176 : XNOR2_X1 port map( A => n2567, B => n15641, ZN => n29546);
   U15220 : AND2_X1 port map( A1 => n3914, A2 => n17197, ZN => n29547);
   U15228 : AND3_X1 port map( A1 => n24, A2 => n5565, A3 => n5564, ZN => n29548
                           );
   U15323 : AND3_X1 port map( A1 => n24, A2 => n5565, A3 => n5564, ZN => n29549
                           );
   U15401 : AND3_X1 port map( A1 => n24, A2 => n5565, A3 => n5564, ZN => n22705
                           );
   U15417 : XNOR2_X1 port map( A => n15748, B => n15749, ZN => n17313);
   U15419 : XNOR2_X1 port map( A => n18572, B => n19649, ZN => n29551);
   U15440 : INV_X1 port map( A => n25421, ZN => n29552);
   U15468 : XNOR2_X1 port map( A => n18572, B => n19649, ZN => n28526);
   U15470 : XNOR2_X1 port map( A => n22943, B => n22942, ZN => n26576);
   U15471 : OR2_X1 port map( A1 => n2534, A2 => n29292, ZN => n29553);
   U15487 : NAND3_X1 port map( A1 => n17325, A2 => n3248, A3 => n17326, ZN => 
                           n29554);
   U15490 : NAND3_X1 port map( A1 => n17325, A2 => n3248, A3 => n17326, ZN => 
                           n19670);
   U15585 : OR2_X1 port map( A1 => n17234, A2 => n17361, ZN => n17044);
   U15658 : XNOR2_X2 port map( A => n18559, B => n18560, ZN => n20081);
   U15708 : OR3_X1 port map( A1 => n11195, A2 => n4341, A3 => n12257, ZN => 
                           n5661);
   U15717 : NOR2_X1 port map( A1 => n28358, A2 => n878, ZN => n29555);
   U15811 : NOR2_X1 port map( A1 => n28358, A2 => n878, ZN => n24395);
   U15812 : INV_X1 port map( A => n4809, ZN => n29556);
   U15813 : OR2_X1 port map( A1 => n27502, A2 => n4808, ZN => n29557);
   U15845 : CLKBUF_X1 port map( A => n13874, Z => n29558);
   U15878 : XNOR2_X1 port map( A => n16030, B => n16029, ZN => n29559);
   U15926 : XNOR2_X1 port map( A => n16030, B => n16029, ZN => n17102);
   U16094 : XNOR2_X1 port map( A => n25314, B => n25313, ZN => n29560);
   U16368 : XNOR2_X1 port map( A => n25314, B => n25313, ZN => n26721);
   U16414 : NOR2_X1 port map( A1 => n15848, A2 => n1241, ZN => n29561);
   U16415 : NOR2_X1 port map( A1 => n20820, A2 => n20819, ZN => n29562);
   U16480 : NOR2_X1 port map( A1 => n15848, A2 => n1241, ZN => n18060);
   U16534 : NOR2_X1 port map( A1 => n20820, A2 => n20819, ZN => n22426);
   U16646 : OAI211_X1 port map( C1 => n24743, C2 => n24744, A => n24742, B => 
                           n24741, ZN => n29563);
   U16912 : XNOR2_X1 port map( A => n12119, B => n12118, ZN => n29565);
   U16945 : XNOR2_X1 port map( A => n12119, B => n12118, ZN => n14165);
   U16959 : XNOR2_X1 port map( A => n14932, B => n1233, ZN => n17433);
   U17012 : OR3_X1 port map( A1 => n20589, A2 => n20314, A3 => n20585, ZN => 
                           n6931);
   U17018 : INV_X1 port map( A => n19827, ZN => n20589);
   U17035 : NOR2_X1 port map( A1 => n23009, A2 => n23008, ZN => n29567);
   U17047 : NOR2_X1 port map( A1 => n23009, A2 => n23008, ZN => n24390);
   U17068 : XNOR2_X2 port map( A => n12502, B => n12501, ZN => n12534);
   U17100 : XNOR2_X1 port map( A => n6998, B => Key(123), ZN => n29568);
   U17152 : INV_X1 port map( A => n28584, ZN => n29569);
   U17153 : NOR2_X1 port map( A1 => n28662, A2 => n28661, ZN => n21587);
   U17202 : AND2_X1 port map( A1 => n18060, A2 => n17671, ZN => n18301);
   U17329 : INV_X1 port map( A => n28009, ZN => n26984);
   U17330 : XNOR2_X1 port map( A => n25529, B => n25530, ZN => n29570);
   U17339 : OAI211_X1 port map( C1 => n15247, C2 => n14733, A => n14732, B => 
                           n14731, ZN => n29571);
   U17340 : XNOR2_X1 port map( A => n14749, B => n14748, ZN => n29572);
   U17341 : OAI211_X1 port map( C1 => n15247, C2 => n14733, A => n14732, B => 
                           n14731, ZN => n16172);
   U17379 : XNOR2_X1 port map( A => n14749, B => n14748, ZN => n17401);
   U17380 : XNOR2_X1 port map( A => n25093, B => n25092, ZN => n29573);
   U17428 : XNOR2_X1 port map( A => n3677, B => n5828, ZN => n29574);
   U17465 : XOR2_X1 port map( A => n25926, B => n25925, Z => n29575);
   U17542 : XNOR2_X1 port map( A => n9317, B => n9316, ZN => n29577);
   U17558 : BUF_X1 port map( A => n27573, Z => n29578);
   U17671 : XNOR2_X1 port map( A => n9317, B => n9316, ZN => n10971);
   U17739 : NOR2_X1 port map( A1 => n26377, A2 => n6723, ZN => n27573);
   U17747 : XNOR2_X1 port map( A => n25502, B => n25208, ZN => n29579);
   U17750 : XNOR2_X1 port map( A => n25502, B => n25208, ZN => n26731);
   U17751 : NAND3_X2 port map( A1 => n4587, A2 => n19936, A3 => n19937, ZN => 
                           n21645);
   U17790 : OAI21_X1 port map( B1 => n4954, B2 => n671, A => n4785, ZN => 
                           n29580);
   U17846 : AND2_X1 port map( A1 => n19771, A2 => n19772, ZN => n29581);
   U17853 : OAI21_X1 port map( B1 => n4954, B2 => n671, A => n4785, ZN => 
                           n19463);
   U18127 : INV_X1 port map( A => n29315, ZN => n29582);
   U18347 : XNOR2_X1 port map( A => n20839, B => n20838, ZN => n29583);
   U18717 : XNOR2_X2 port map( A => n25468, B => n25469, ZN => n26747);
   U18749 : BUF_X1 port map( A => n20053, Z => n29584);
   U18761 : XNOR2_X1 port map( A => n6122, B => n24900, ZN => n29585);
   U18918 : XNOR2_X1 port map( A => n6122, B => n24900, ZN => n2108);
   U18919 : XOR2_X1 port map( A => n18941, B => n18940, Z => n29587);
   U18976 : BUF_X1 port map( A => n27026, Z => n29588);
   U18980 : XNOR2_X1 port map( A => n13376, B => n13377, ZN => n29589);
   U18997 : XNOR2_X1 port map( A => n13376, B => n13377, ZN => n14016);
   U19128 : XOR2_X1 port map( A => n7218, B => Key(130), Z => n29590);
   U19148 : OR2_X1 port map( A1 => n2719, A2 => n18144, ZN => n2720);
   U19157 : BUF_X1 port map( A => n24215, Z => n29592);
   U19189 : AOI22_X1 port map( A1 => n23646, A2 => n6378, B1 => n23565, B2 => 
                           n23564, ZN => n24215);
   U19214 : BUF_X1 port map( A => n10875, Z => n29593);
   U19254 : OAI211_X1 port map( C1 => n4005, C2 => n17001, A => n4004, B => 
                           n6638, ZN => n29594);
   U19291 : OAI211_X1 port map( C1 => n4005, C2 => n17001, A => n4004, B => 
                           n6638, ZN => n29595);
   U19312 : OAI211_X1 port map( C1 => n4005, C2 => n17001, A => n4004, B => 
                           n6638, ZN => n18040);
   U19353 : OR2_X1 port map( A1 => n26186, A2 => n26182, ZN => n29596);
   U19372 : INV_X1 port map( A => n469, ZN => n29597);
   U19444 : XOR2_X1 port map( A => n16108, B => n16109, Z => n29598);
   U19458 : OAI21_X1 port map( B1 => n24623, B2 => n28223, A => n24621, ZN => 
                           n29599);
   U19465 : XNOR2_X1 port map( A => n14629, B => n14628, ZN => n29600);
   U19489 : BUF_X1 port map( A => n20506, Z => n29601);
   U19490 : XNOR2_X1 port map( A => n14629, B => n14628, ZN => n16992);
   U19572 : XNOR2_X2 port map( A => n22540, B => n22539, ZN => n29602);
   U19574 : XNOR2_X1 port map( A => n22540, B => n22539, ZN => n23831);
   U19735 : AOI21_X1 port map( B1 => n16928, B2 => n29566, A => n16927, ZN => 
                           n29603);
   U19755 : AOI21_X1 port map( B1 => n16928, B2 => n29566, A => n16927, ZN => 
                           n18325);
   U19765 : XNOR2_X1 port map( A => n12811, B => n12812, ZN => n29604);
   U19792 : XNOR2_X1 port map( A => n12811, B => n12812, ZN => n2728);
   U19800 : XNOR2_X1 port map( A => n15924, B => n15923, ZN => n29605);
   U19812 : OAI22_X1 port map( A1 => n24548, A2 => n24547, B1 => n24545, B2 => 
                           n24546, ZN => n29606);
   U19913 : OAI22_X1 port map( A1 => n24548, A2 => n24547, B1 => n24545, B2 => 
                           n24546, ZN => n25534);
   U19983 : XNOR2_X1 port map( A => n12381, B => n12382, ZN => n29607);
   U20011 : AND2_X2 port map( A1 => n29608, A2 => n29609, ZN => n19215);
   U20051 : AND2_X1 port map( A1 => n2901, A2 => n2031, ZN => n29608);
   U20055 : OR2_X1 port map( A1 => n17632, A2 => n17834, ZN => n29609);
   U20063 : XNOR2_X1 port map( A => n12381, B => n12382, ZN => n14331);
   U20114 : XNOR2_X1 port map( A => n19456, B => n19455, ZN => n21359);
   U20209 : XNOR2_X2 port map( A => n3649, B => n25371, ZN => n29610);
   U20261 : XNOR2_X1 port map( A => n3649, B => n25371, ZN => n26912);
   U20297 : XNOR2_X1 port map( A => n13289, B => n13288, ZN => n29611);
   U20342 : NOR2_X1 port map( A1 => n23753, A2 => n23754, ZN => n29612);
   U20344 : NOR2_X1 port map( A1 => n23753, A2 => n23754, ZN => n29613);
   U20429 : XNOR2_X1 port map( A => n13289, B => n13288, ZN => n14301);
   U20643 : NOR2_X1 port map( A1 => n23753, A2 => n23754, ZN => n26056);
   U20744 : BUF_X1 port map( A => n25913, Z => n29614);
   U20766 : OR2_X1 port map( A1 => n27898, A2 => n26510, ZN => n29615);
   U20855 : XNOR2_X1 port map( A => n19158, B => n19157, ZN => n29616);
   U20856 : CLKBUF_X1 port map( A => n26194, Z => n29617);
   U20857 : XNOR2_X1 port map( A => n19158, B => n19157, ZN => n20493);
   U20867 : XNOR2_X1 port map( A => n22083, B => n22082, ZN => n29618);
   U20886 : INV_X1 port map( A => n6150, ZN => n29619);
   U20936 : XNOR2_X1 port map( A => n22316, B => n22317, ZN => n29620);
   U20958 : XNOR2_X1 port map( A => n26124, B => n26123, ZN => n29621);
   U20968 : XNOR2_X1 port map( A => n26124, B => n26123, ZN => n27140);
   U21035 : XNOR2_X1 port map( A => n25726, B => n25725, ZN => n29622);
   U21194 : AOI21_X1 port map( B1 => n26991, B2 => n25770, A => n25769, ZN => 
                           n29623);
   U21198 : AND2_X1 port map( A1 => n7291, A2 => n7292, ZN => n7784);
   U21257 : OAI21_X1 port map( B1 => n23535, B2 => n23534, A => n6942, ZN => 
                           n29624);
   U21288 : XOR2_X1 port map( A => n19684, B => n19683, Z => n29625);
   U21307 : XOR2_X1 port map( A => n13135, B => n3097, Z => n29626);
   U21308 : XNOR2_X1 port map( A => n9952, B => n9951, ZN => n29627);
   U21322 : CLKBUF_X1 port map( A => n14401, Z => n29628);
   U21394 : XNOR2_X1 port map( A => Key(59), B => Plaintext(59), ZN => n8034);
   U21431 : XOR2_X1 port map( A => n16495, B => n14760, Z => n29630);
   U21462 : XOR2_X1 port map( A => n25171, B => n25170, Z => n29631);
   U21478 : BUF_X1 port map( A => n24111, Z => n24422);
   U21497 : XNOR2_X1 port map( A => n15556, B => n15555, ZN => n29632);
   U21610 : XNOR2_X1 port map( A => n15556, B => n15555, ZN => n17344);
   U21630 : OAI22_X1 port map( A1 => n23951, A2 => n23950, B1 => n5004, B2 => 
                           n24810, ZN => n29634);
   U21634 : XNOR2_X1 port map( A => n16372, B => n16371, ZN => n29635);
   U21651 : XNOR2_X1 port map( A => n16372, B => n16371, ZN => n29636);
   U21689 : BUF_X1 port map( A => n11056, Z => n29637);
   U21700 : XNOR2_X1 port map( A => n4592, B => n9659, ZN => n11056);
   U21769 : MUX2_X2 port map( A => n27126, B => n27127, S => n4109, Z => n27759
                           );
   U21770 : MUX2_X1 port map( A => n7800, B => n7898, S => n7801, Z => n7314);
   U21777 : XNOR2_X1 port map( A => n7103, B => Key(187), ZN => n7801);
   U21778 : XNOR2_X1 port map( A => n10363, B => n9401, ZN => n10425);
   U21797 : XNOR2_X2 port map( A => n14985, B => n14984, ZN => n17439);
   U21845 : XNOR2_X2 port map( A => n21942, B => n21941, ZN => n23789);
   U21994 : NAND4_X2 port map( A1 => n17377, A2 => n16875, A3 => n16877, A4 => 
                           n16876, ZN => n18507);
   U22057 : XOR2_X1 port map( A => Key(148), B => Plaintext(148), Z => n29639);
   U22060 : CLKBUF_X1 port map( A => n12554, Z => n29640);
   U22078 : OAI211_X1 port map( C1 => n23161, C2 => n23489, A => n28844, B => 
                           n3026, ZN => n29642);
   U22080 : OAI211_X1 port map( C1 => n23161, C2 => n23489, A => n28844, B => 
                           n3026, ZN => n29643);
   U22093 : OAI211_X1 port map( C1 => n23161, C2 => n23489, A => n28844, B => 
                           n3026, ZN => n24645);
   U22175 : XOR2_X1 port map( A => n18166, B => n18167, Z => n29644);
   U22188 : CLKBUF_X1 port map( A => n24644, Z => n29645);
   U22227 : OAI21_X1 port map( B1 => n23175, B2 => n23174, A => n23173, ZN => 
                           n24644);
   U22228 : XNOR2_X1 port map( A => n2638, B => Key(47), ZN => n29646);
   U22349 : NAND2_X1 port map( A1 => n29774, A2 => n29741, ZN => n29647);
   U22350 : XNOR2_X1 port map( A => n2638, B => Key(47), ZN => n7129);
   U22364 : XOR2_X1 port map( A => n9753, B => n9752, Z => n29648);
   U22382 : AOI21_X1 port map( B1 => n14358, B2 => n14273, A => n14271, ZN => 
                           n29649);
   U22457 : NAND2_X1 port map( A1 => n24686, A2 => n24687, ZN => n2649);
   U22530 : NAND3_X1 port map( A1 => n9031, A2 => n9029, A3 => n9030, ZN => 
                           n9032);
   U22657 : NAND2_X1 port map( A1 => n149, A2 => n23901, ZN => n148);
   U22714 : NOR2_X2 port map( A1 => n29652, A2 => n29651, ZN => n22698);
   U22721 : INV_X1 port map( A => n19188, ZN => n29651);
   U22733 : NAND3_X1 port map( A1 => n7709, A2 => n8032, A3 => n7734, ZN => 
                           n28998);
   U22743 : NAND2_X1 port map( A1 => n29653, A2 => n15372, ZN => n15378);
   U22788 : NAND2_X1 port map( A1 => n683, A2 => n15369, ZN => n29653);
   U22791 : OR2_X1 port map( A1 => n14147, A2 => n14148, ZN => n6254);
   U22822 : NAND2_X1 port map( A1 => n2302, A2 => n2303, ZN => n13179);
   U22876 : OAI21_X1 port map( B1 => n17980, B2 => n18709, A => n29654, ZN => 
                           n18249);
   U22892 : NAND2_X1 port map( A1 => n18709, A2 => n18248, ZN => n29654);
   U22894 : NOR2_X2 port map( A1 => n13033, A2 => n29655, ZN => n14948);
   U22911 : NAND2_X1 port map( A1 => n5351, A2 => n13024, ZN => n29655);
   U22918 : NOR2_X1 port map( A1 => n1725, A2 => n14657, ZN => n14669);
   U23006 : NAND3_X1 port map( A1 => n21484, A2 => n21575, A3 => n21485, ZN => 
                           n21486);
   U23047 : NAND3_X1 port map( A1 => n3454, A2 => n10991, A3 => n10992, ZN => 
                           n9814);
   U23049 : NAND3_X2 port map( A1 => n17049, A2 => n29709, A3 => n29708, ZN => 
                           n18333);
   U23083 : NAND2_X1 port map( A1 => n17263, A2 => n16995, ZN => n17266);
   U23152 : XNOR2_X2 port map( A => n14656, B => n14655, ZN => n17263);
   U23176 : NAND2_X1 port map( A1 => n10702, A2 => n28310, ZN => n10710);
   U23177 : NAND3_X1 port map( A1 => n21481, A2 => n21483, A3 => n21574, ZN => 
                           n21488);
   U23208 : NAND2_X1 port map( A1 => n29316, A2 => n11321, ZN => n11188);
   U23209 : XNOR2_X2 port map( A => n9053, B => n9052, ZN => n11321);
   U23216 : NAND3_X1 port map( A1 => n6706, A2 => n4341, A3 => n6687, ZN => 
                           n28863);
   U23217 : NAND3_X1 port map( A1 => n14901, A2 => n14906, A3 => n14904, ZN => 
                           n14679);
   U23219 : NAND2_X1 port map( A1 => n5733, A2 => n5734, ZN => n5732);
   U23284 : XNOR2_X1 port map( A => n29656, B => n21946, ZN => n21104);
   U23285 : XNOR2_X1 port map( A => n21083, B => n6520, ZN => n29656);
   U23286 : XNOR2_X2 port map( A => n22329, B => n1772, ZN => n23474);
   U23369 : OR2_X1 port map( A1 => n10484, A2 => n11258, ZN => n29722);
   U23370 : AND3_X2 port map( A1 => n29657, A2 => n26213, A3 => n26212, ZN => 
                           n27213);
   U23439 : NOR2_X1 port map( A1 => n21501, A2 => n21192, ZN => n21504);
   U23440 : NAND2_X1 port map( A1 => n20380, A2 => n20379, ZN => n29658);
   U23453 : NAND3_X1 port map( A1 => n20023, A2 => n28126, A3 => n19795, ZN => 
                           n3969);
   U23489 : NAND3_X2 port map( A1 => n29194, A2 => n16807, A3 => n29195, ZN => 
                           n18170);
   U23504 : OR2_X1 port map( A1 => n5200, A2 => n5222, ZN => n4943);
   U23514 : NAND2_X1 port map( A1 => n8321, A2 => n9530, ZN => n29660);
   U23583 : NAND2_X1 port map( A1 => n8322, A2 => n29662, ZN => n29661);
   U23590 : NAND2_X1 port map( A1 => n18449, A2 => n18198, ZN => n17746);
   U23638 : NAND3_X1 port map( A1 => n13935, A2 => n293, A3 => n29320, ZN => 
                           n642);
   U23731 : NAND2_X1 port map( A1 => n14614, A2 => n14615, ZN => n1310);
   U23732 : NAND2_X1 port map( A1 => n4799, A2 => n4837, ZN => n13705);
   U23733 : NAND2_X1 port map( A1 => n4627, A2 => n13704, ZN => n4799);
   U23738 : NAND2_X1 port map( A1 => n29664, A2 => n2554, ZN => n10591);
   U23741 : NAND2_X1 port map( A1 => n11005, A2 => n5573, ZN => n29664);
   U23966 : XNOR2_X1 port map( A => n29665, B => n2960, ZN => Ciphertext(137));
   U24053 : AOI22_X1 port map( A1 => n27250, A2 => n27828, B1 => n27826, B2 => 
                           n27249, ZN => n29665);
   U24062 : NAND2_X1 port map( A1 => n29667, A2 => n29666, ZN => n29749);
   U24080 : INV_X1 port map( A => n3817, ZN => n29666);
   U24134 : NAND2_X1 port map( A1 => n29669, A2 => n29668, ZN => n29667);
   U24145 : NAND2_X1 port map( A1 => n3820, A2 => n10833, ZN => n29668);
   U24184 : NAND2_X1 port map( A1 => n29148, A2 => n1338, ZN => n29669);
   U24207 : NAND2_X1 port map( A1 => n28349, A2 => n29671, ZN => n29670);
   U24303 : NAND2_X1 port map( A1 => n26728, A2 => n26481, ZN => n26726);
   U24331 : NAND2_X1 port map( A1 => n189, A2 => n192, ZN => n15349);
   U24351 : NAND2_X1 port map( A1 => n7478, A2 => n29672, ZN => n7483);
   U24399 : NAND2_X1 port map( A1 => n29673, A2 => n7477, ZN => n29672);
   U24481 : NAND2_X1 port map( A1 => n7975, A2 => n8275, ZN => n7477);
   U24495 : INV_X1 port map( A => n7976, ZN => n29673);
   U24620 : NAND3_X1 port map( A1 => n6003, A2 => n6004, A3 => n29675, ZN => 
                           n16360);
   U24679 : NAND2_X2 port map( A1 => n29676, A2 => n23927, ZN => n25328);
   U24751 : NAND2_X1 port map( A1 => n29678, A2 => n29677, ZN => n29676);
   U24764 : NAND2_X1 port map( A1 => n29512, A2 => n24751, ZN => n29678);
   U24828 : NAND2_X2 port map( A1 => n29679, A2 => n1304, ZN => n19702);
   U24829 : OAI21_X1 port map( B1 => n18448, B2 => n18097, A => n668, ZN => 
                           n29679);
   U24907 : OAI21_X1 port map( B1 => n28086, B2 => n28087, A => n29680, ZN => 
                           n3517);
   U24960 : NAND3_X1 port map( A1 => n91, A2 => n2021, A3 => n29681, ZN => 
                           n29680);
   U24961 : NAND2_X1 port map( A1 => n1659, A2 => n29682, ZN => n15009);
   U24978 : XNOR2_X1 port map( A => n14921, B => n15575, ZN => n16320);
   U25001 : AND2_X2 port map( A1 => n29684, A2 => n29683, ZN => n15575);
   U25002 : NAND2_X1 port map( A1 => n6320, A2 => n14574, ZN => n29683);
   U25013 : NAND2_X1 port map( A1 => n14573, A2 => n14572, ZN => n29684);
   U25017 : NOR2_X1 port map( A1 => n20173, A2 => n20178, ZN => n19002);
   U25018 : NAND3_X2 port map( A1 => n3282, A2 => n7294, A3 => n28696, ZN => 
                           n8336);
   U25037 : NAND2_X1 port map( A1 => n29685, A2 => n715, ZN => n19086);
   U25040 : NAND2_X1 port map( A1 => n17861, A2 => n2292, ZN => n29685);
   U25051 : NAND2_X1 port map( A1 => n29687, A2 => n29686, ZN => n8860);
   U25058 : NAND2_X1 port map( A1 => n9075, A2 => n9069, ZN => n29686);
   U25068 : NAND2_X1 port map( A1 => n8859, A2 => n28212, ZN => n29687);
   U25104 : NAND3_X1 port map( A1 => n15460, A2 => n15457, A3 => n15459, ZN => 
                           n2745);
   U25129 : NAND3_X1 port map( A1 => n13831, A2 => n13830, A3 => n29688, ZN => 
                           n14534);
   U25134 : NAND2_X1 port map( A1 => n29690, A2 => n29689, ZN => n29688);
   U25137 : AOI21_X1 port map( B1 => n14359, B2 => n14278, A => n13832, ZN => 
                           n29689);
   U25225 : NAND2_X1 port map( A1 => n28507, A2 => n29691, ZN => n29690);
   U25235 : NAND3_X1 port map( A1 => n2684, A2 => n2683, A3 => n6281, ZN => 
                           n2682);
   U25264 : OAI21_X1 port map( B1 => n29693, B2 => n22290, A => n29692, ZN => 
                           n20668);
   U25268 : NAND2_X1 port map( A1 => n22290, A2 => n20666, ZN => n29692);
   U25312 : INV_X1 port map( A => n20667, ZN => n29693);
   U25323 : NAND3_X1 port map( A1 => n7711, A2 => n8029, A3 => n618, ZN => 
                           n1032);
   U25336 : NAND2_X1 port map( A1 => n7734, A2 => n7265, ZN => n7711);
   U25354 : NOR2_X1 port map( A1 => n1019, A2 => n29694, ZN => n1389);
   U25382 : NOR2_X1 port map( A1 => n28257, A2 => n60, ZN => n29694);
   U25383 : NAND2_X1 port map( A1 => n29695, A2 => n24725, ZN => n24148);
   U25430 : INV_X1 port map( A => n6309, ZN => n29695);
   U25494 : NAND3_X2 port map( A1 => n29698, A2 => n12994, A3 => n3008, ZN => 
                           n13386);
   U25584 : NAND2_X1 port map( A1 => n10801, A2 => n12149, ZN => n29698);
   U25594 : NAND3_X1 port map( A1 => n28076, A2 => n29700, A3 => n29699, ZN => 
                           n28079);
   U25618 : INV_X1 port map( A => n28110, ZN => n29699);
   U25619 : NAND2_X1 port map( A1 => n28109, A2 => n28794, ZN => n29700);
   U25626 : NAND2_X1 port map( A1 => n1626, A2 => n1624, ZN => n21435);
   U25634 : NAND3_X1 port map( A1 => n17105, A2 => n17104, A3 => n17103, ZN => 
                           n18135);
   U25638 : NAND4_X1 port map( A1 => n29701, A2 => n1411, A3 => n1407, A4 => 
                           n27307, ZN => n1410);
   U25706 : NAND2_X1 port map( A1 => n2782, A2 => n14428, ZN => n13875);
   U25724 : AND2_X2 port map( A1 => n16022, A2 => n3729, ZN => n17762);
   U25727 : NAND2_X1 port map( A1 => n4871, A2 => n29702, ZN => n24533);
   U25866 : NAND3_X1 port map( A1 => n4892, A2 => n23146, A3 => n23457, ZN => 
                           n29702);
   U25913 : NAND3_X1 port map( A1 => n29703, A2 => n1949, A3 => n4096, ZN => 
                           n21642);
   U25959 : NAND2_X1 port map( A1 => n2487, A2 => n4278, ZN => n29703);
   U26011 : NAND2_X1 port map( A1 => n29704, A2 => n20221, ZN => n1413);
   U26039 : NAND2_X1 port map( A1 => n296, A2 => n20219, ZN => n29704);
   U26104 : NAND3_X1 port map( A1 => n15087, A2 => n13989, A3 => n15083, ZN => 
                           n13990);
   U26105 : NAND3_X1 port map( A1 => n14617, A2 => n14916, A3 => n14618, ZN => 
                           n29211);
   U26142 : OAI211_X2 port map( C1 => n12010, C2 => n14250, A => n12009, B => 
                           n5790, ZN => n14894);
   U26177 : NOR3_X1 port map( A1 => n15691, A2 => n15690, A3 => n14563, ZN => 
                           n15694);
   U26242 : NAND3_X1 port map( A1 => n28677, A2 => n28676, A3 => n12990, ZN => 
                           n29705);
   U26243 : OAI21_X1 port map( B1 => n20281, B2 => n29707, A => n29706, ZN => 
                           n19898);
   U26287 : OR2_X1 port map( A1 => n17236, A2 => n15731, ZN => n29708);
   U26324 : NAND2_X1 port map( A1 => n7410, A2 => n8925, ZN => n8926);
   U26328 : NAND2_X1 port map( A1 => n17047, A2 => n17365, ZN => n29709);
   U26337 : NAND2_X1 port map( A1 => n29712, A2 => n29711, ZN => n29710);
   U26373 : AOI21_X1 port map( B1 => n10912, B2 => n9348, A => n10609, ZN => 
                           n29711);
   U26374 : NAND2_X1 port map( A1 => n10915, A2 => n29078, ZN => n29712);
   U26414 : NAND2_X1 port map( A1 => n10898, A2 => n12361, ZN => n870);
   U26432 : NAND3_X1 port map( A1 => n3519, A2 => n4950, A3 => n28609, ZN => 
                           n28888);
   U26475 : OR2_X1 port map( A1 => n17428, A2 => n6013, ZN => n14226);
   U26487 : NAND3_X1 port map( A1 => n6097, A2 => n6098, A3 => n24489, ZN => 
                           n24102);
   U26496 : OAI21_X1 port map( B1 => n2018, B2 => n4586, A => n29713, ZN => 
                           n13596);
   U26544 : NAND3_X1 port map( A1 => n4586, A2 => n14376, A3 => n2849, ZN => 
                           n29713);
   U26546 : NAND2_X1 port map( A1 => n29714, A2 => n2594, ZN => n20675);
   U26547 : NAND2_X1 port map( A1 => n20007, A2 => n20623, ZN => n29714);
   U26572 : NAND2_X1 port map( A1 => n11580, A2 => n11954, ZN => n12260);
   U26583 : NAND4_X2 port map( A1 => n29715, A2 => n17443, A3 => n17445, A4 => 
                           n17444, ZN => n19468);
   U26840 : NAND2_X1 port map( A1 => n15466, A2 => n15463, ZN => n4734);
   U26853 : NAND4_X2 port map( A1 => n3228, A2 => n4500, A3 => n13870, A4 => 
                           n13869, ZN => n15466);
   U26854 : NAND3_X1 port map( A1 => n3934, A2 => n11162, A3 => n3935, ZN => 
                           n4037);
   U26855 : NOR2_X2 port map( A1 => n20675, A2 => n20670, ZN => n21394);
   U26873 : NAND3_X1 port map( A1 => n10523, A2 => n11269, A3 => n11275, ZN => 
                           n11270);
   U26884 : NAND2_X1 port map( A1 => n29717, A2 => n29716, ZN => n15590);
   U26903 : NAND2_X1 port map( A1 => n15581, A2 => n17339, ZN => n29716);
   U26904 : NAND2_X1 port map( A1 => n15582, A2 => n29718, ZN => n29717);
   U26905 : INV_X1 port map( A => n17339, ZN => n29718);
   U26908 : OR2_X2 port map( A1 => n4887, A2 => n19869, ZN => n20857);
   U26909 : NAND2_X1 port map( A1 => n9000, A2 => n9001, ZN => n4303);
   U26918 : NAND2_X1 port map( A1 => n9200, A2 => n329, ZN => n9001);
   U26935 : NAND2_X1 port map( A1 => n29719, A2 => n2232, ZN => n12019);
   U26958 : NAND2_X1 port map( A1 => n12018, A2 => n12017, ZN => n29719);
   U27024 : NAND2_X1 port map( A1 => n15, A2 => n1416, ZN => n9786);
   U27030 : NAND2_X1 port map( A1 => n8044, A2 => n8139, ZN => n8045);
   U27040 : NAND3_X1 port map( A1 => n16915, A2 => n186, A3 => n16914, ZN => 
                           n18326);
   U27050 : BUF_X2 port map( A => n25908, Z => n28771);
   U27062 : NAND2_X1 port map( A1 => n29721, A2 => n29720, ZN => n8801);
   U27068 : NAND2_X1 port map( A1 => n8288, A2 => n8289, ZN => n29720);
   U27079 : NAND2_X1 port map( A1 => n8293, A2 => n8292, ZN => n29721);
   U27094 : NAND2_X1 port map( A1 => n23758, A2 => n29131, ZN => n23475);
   U27108 : NAND2_X1 port map( A1 => n2437, A2 => n2439, ZN => n27253);
   U27166 : AOI21_X1 port map( B1 => n8214, B2 => n8215, A => n8213, ZN => 
                           n8220);
   U27167 : NAND2_X1 port map( A1 => n7625, A2 => n8216, ZN => n8214);
   U27177 : NAND2_X1 port map( A1 => n6855, A2 => n15398, ZN => n29290);
   U27199 : NAND2_X1 port map( A1 => n29723, A2 => n29722, ZN => n12026);
   U27200 : OAI21_X1 port map( B1 => n4650, B2 => n3882, A => n4649, ZN => 
                           n29723);
   U27225 : XNOR2_X1 port map( A => n29724, B => n4607, ZN => Ciphertext(112));
   U27252 : NAND3_X1 port map( A1 => n26147, A2 => n26148, A3 => n6952, ZN => 
                           n29724);
   U27273 : AOI22_X2 port map( A1 => n7874, A2 => n5360, B1 => n7875, B2 => 
                           n7959, ZN => n8116);
   U27331 : NAND3_X1 port map( A1 => n403, A2 => n29727, A3 => n29725, ZN => 
                           n24349);
   U27361 : NAND2_X1 port map( A1 => n29128, A2 => n29726, ZN => n29725);
   U27362 : NAND2_X1 port map( A1 => n14922, A2 => n14621, ZN => n14706);
   U27378 : NAND2_X1 port map( A1 => n29728, A2 => n28934, ZN => n7558);
   U27380 : NAND2_X1 port map( A1 => n28933, A2 => n29119, ZN => n29728);
   U27381 : NAND3_X1 port map( A1 => n29150, A2 => n11113, A3 => n10461, ZN => 
                           n2868);
   U27387 : NAND3_X1 port map( A1 => n382, A2 => n383, A3 => n19997, ZN => 
                           n6452);
   U27404 : NAND3_X1 port map( A1 => n7947, A2 => n8257, A3 => n8258, ZN => 
                           n7467);
   U27411 : NAND2_X1 port map( A1 => n22457, A2 => n29729, ZN => n24610);
   U27495 : AND2_X2 port map( A1 => n5342, A2 => n29730, ZN => n15311);
   U27499 : NAND2_X1 port map( A1 => n28273, A2 => n28351, ZN => n29730);
   U27514 : AND3_X2 port map( A1 => n14387, A2 => n14388, A3 => n14389, ZN => 
                           n16443);
   U27622 : NAND2_X2 port map( A1 => n29731, A2 => n5280, ZN => n12181);
   U27635 : NAND2_X1 port map( A1 => n5278, A2 => n5277, ZN => n29731);
   U27650 : OAI211_X2 port map( C1 => n24292, C2 => n24291, A => n24290, B => 
                           n24289, ZN => n25890);
   U27651 : OAI21_X1 port map( B1 => n13720, B2 => n13587, A => n29732, ZN => 
                           n13898);
   U27747 : NAND2_X1 port map( A1 => n13587, A2 => n28569, ZN => n29732);
   U27808 : AOI22_X1 port map( A1 => n21861, A2 => n23779, B1 => n23514, B2 => 
                           n21862, ZN => n29733);
   U27809 : NAND3_X1 port map( A1 => n11905, A2 => n12430, A3 => n29734, ZN => 
                           n11912);
   U27846 : NAND2_X1 port map( A1 => n12429, A2 => n29735, ZN => n29734);
   U27874 : NAND2_X1 port map( A1 => n8351, A2 => n8077, ZN => n8078);
   U27875 : OR2_X2 port map( A1 => n7799, A2 => n7798, ZN => n8077);
   U27904 : NAND3_X1 port map( A1 => n20330, A2 => n1881, A3 => n20623, ZN => 
                           n20331);
   U27910 : OAI22_X1 port map( A1 => n26616, A2 => n28228, B1 => n29736, B2 => 
                           n922, ZN => n26502);
   U27945 : NAND2_X1 port map( A1 => n28452, A2 => n26614, ZN => n29736);
   U28102 : NAND3_X1 port map( A1 => n28800, A2 => n17467, A3 => n29737, ZN => 
                           n3981);
   U28105 : NAND2_X1 port map( A1 => n968, A2 => n17018, ZN => n29738);
   U28108 : OR2_X1 port map( A1 => n23010, A2 => n29583, ZN => n23012);
   U28132 : NOR2_X2 port map( A1 => n10590, A2 => n10591, ZN => n12363);
   U28136 : NAND2_X1 port map( A1 => n23020, A2 => n24691, ZN => n23027);
   U28137 : NAND2_X1 port map( A1 => n20175, A2 => n20174, ZN => n29739);
   U28169 : NAND2_X1 port map( A1 => n29740, A2 => n18441, ZN => n17739);
   U28173 : NAND2_X1 port map( A1 => n18181, A2 => n18178, ZN => n29740);
   U28177 : NAND2_X1 port map( A1 => n29774, A2 => n29741, ZN => n18512);
   U28180 : NAND2_X1 port map( A1 => n4089, A2 => n17492, ZN => n29741);
   U28189 : NAND3_X1 port map( A1 => n596, A2 => n8984, A3 => n8983, ZN => 
                           n8985);
   U28190 : NAND2_X1 port map( A1 => n26129, A2 => n27178, ZN => n26264);
   U28193 : AND2_X2 port map( A1 => n29743, A2 => n29742, ZN => n22374);
   U28211 : NAND2_X1 port map( A1 => n21505, A2 => n21506, ZN => n29742);
   U28214 : NAND2_X1 port map( A1 => n21508, A2 => n29744, ZN => n29743);
   U28228 : NAND2_X1 port map( A1 => n21504, A2 => n28611, ZN => n29744);
   U28232 : OAI211_X1 port map( C1 => n24597, C2 => n24595, A => n24730, B => 
                           n29745, ZN => n5654);
   U28233 : NAND2_X1 port map( A1 => n29746, A2 => n24595, ZN => n29745);
   U28238 : INV_X1 port map( A => n24596, ZN => n29746);
   U28239 : NAND3_X2 port map( A1 => n28887, A2 => n10462, A3 => n4630, ZN => 
                           n11877);
   U28271 : NAND3_X1 port map( A1 => n14729, A2 => n14733, A3 => n14730, ZN => 
                           n14732);
   U28288 : XNOR2_X1 port map( A => n19575, B => n19016, ZN => n18855);
   U28295 : XNOR2_X1 port map( A => n19075, B => n19463, ZN => n19016);
   U28300 : NAND2_X1 port map( A1 => n29747, A2 => n530, ZN => n16877);
   U28301 : AND2_X1 port map( A1 => n29636, A2 => n28775, ZN => n29747);
   U28306 : NAND2_X1 port map( A1 => n491, A2 => n20933, ZN => n20762);
   U28309 : OAI21_X1 port map( B1 => n11617, B2 => n12507, A => n10864, ZN => 
                           n29748);
   U28310 : NAND3_X1 port map( A1 => n7309, A2 => n7601, A3 => n5149, ZN => 
                           n5361);
   U28311 : NAND2_X1 port map( A1 => n1697, A2 => n4294, ZN => n29008);
   U28312 : INV_X1 port map( A => n10723, ZN => n10612);
   U28313 : NAND2_X1 port map( A1 => n10976, A2 => n10948, ZN => n10723);
   U28314 : NAND2_X1 port map( A1 => n10648, A2 => n12337, ZN => n12346);
   U28315 : NAND2_X2 port map( A1 => n29749, A2 => n10480, ZN => n12337);
   U28316 : NAND2_X1 port map( A1 => n29752, A2 => n29750, ZN => n7125);
   U28317 : NAND2_X1 port map( A1 => n8139, A2 => n29751, ZN => n29750);
   U28318 : INV_X1 port map( A => n7560, ZN => n29751);
   U28319 : NAND2_X1 port map( A1 => n8041, A2 => n7560, ZN => n29752);
   U28320 : OAI21_X1 port map( B1 => n24667, B2 => n29754, A => n29753, ZN => 
                           n24384);
   U28321 : NAND2_X1 port map( A1 => n24667, A2 => n24383, ZN => n29753);
   U28322 : AND2_X1 port map( A1 => n23006, A2 => n23162, ZN => n23523);
   U28323 : NAND3_X1 port map( A1 => n18186, A2 => n18187, A3 => n29199, ZN => 
                           n2136);
   U28324 : NOR2_X1 port map( A1 => n29755, A2 => n26066, ZN => n26067);
   U28325 : INV_X1 port map( A => n26309, ZN => n29755);
   U28326 : NAND2_X1 port map( A1 => n26865, A2 => n29048, ZN => n26309);
   U28327 : OAI211_X2 port map( C1 => n8871, C2 => n8872, A => n8869, B => 
                           n8870, ZN => n10251);
   U28328 : NAND3_X1 port map( A1 => n28808, A2 => n8812, A3 => n8808, ZN => 
                           n8253);
   U28329 : OAI21_X1 port map( B1 => n11956, B2 => n571, A => n29757, ZN => 
                           n11200);
   U28330 : NAND2_X1 port map( A1 => n571, A2 => n12261, ZN => n29757);
   U28331 : NAND2_X1 port map( A1 => n11175, A2 => n11174, ZN => n11178);
   U28332 : NAND2_X1 port map( A1 => n3218, A2 => n29758, ZN => n15617);
   U28333 : NAND2_X1 port map( A1 => n2497, A2 => n2495, ZN => n29758);
   U28334 : NAND2_X1 port map( A1 => n29759, A2 => n17013, ZN => n6130);
   U28335 : NAND2_X1 port map( A1 => n16790, A2 => n5714, ZN => n29759);
   U28336 : NAND2_X1 port map( A1 => n13954, A2 => n29760, ZN => n13894);
   U28337 : NAND2_X1 port map( A1 => n14216, A2 => n14217, ZN => n13954);
   U28338 : OAI211_X2 port map( C1 => n4104, C2 => n20869, A => n28943, B => 
                           n29761, ZN => n22523);
   U28339 : NAND2_X1 port map( A1 => n20866, A2 => n4104, ZN => n29761);
   U28340 : NAND2_X1 port map( A1 => n514, A2 => n18343, ZN => n1480);
   U28341 : XNOR2_X1 port map( A => n29762, B => n1184, ZN => Ciphertext(116));
   U28342 : NAND3_X1 port map( A1 => n2792, A2 => n1216, A3 => n2793, ZN => 
                           n29762);
   U28343 : NAND2_X1 port map( A1 => n4035, A2 => n4036, ZN => n4034);
   U28344 : XNOR2_X1 port map( A => n22883, B => n22882, ZN => n29763);
   U28345 : XNOR2_X1 port map( A => n29764, B => n17697, ZN => n17726);
   U28346 : XNOR2_X1 port map( A => n17690, B => n18114, ZN => n29764);
   U28347 : NAND2_X1 port map( A1 => n5917, A2 => n10749, ZN => n3129);
   U28348 : XNOR2_X2 port map( A => n5002, B => n5003, ZN => n14414);
   U28349 : OAI211_X2 port map( C1 => n24807, C2 => n4335, A => n4334, B => 
                           n4333, ZN => n25515);
   U28350 : OAI21_X1 port map( B1 => n400, B2 => n27702, A => n29765, ZN => 
                           n28667);
   U28351 : INV_X1 port map( A => n2011, ZN => n29765);
   U28352 : OR3_X1 port map( A1 => n23357, A2 => n23355, A3 => n1837, ZN => 
                           n28924);
   U28353 : NAND3_X1 port map( A1 => n4306, A2 => n20603, A3 => n1915, ZN => 
                           n5252);
   U28354 : NAND2_X1 port map( A1 => n4914, A2 => n29766, ZN => n16855);
   U28355 : INV_X1 port map( A => n16850, ZN => n29766);
   U28356 : NAND2_X2 port map( A1 => n29768, A2 => n29767, ZN => n15464);
   U28357 : NAND3_X1 port map( A1 => n2344, A2 => n28804, A3 => n2346, ZN => 
                           n29767);
   U28358 : NAND2_X1 port map( A1 => n2607, A2 => n4012, ZN => n29768);
   U28359 : XNOR2_X1 port map( A => n29769, B => n19686, ZN => n4042);
   U28360 : AND2_X2 port map( A1 => n5163, A2 => n5162, ZN => n19484);
   U28361 : INV_X1 port map( A => n16574, ZN => n16009);
   U28362 : XNOR2_X1 port map( A => n16574, B => n16039, ZN => n16453);
   U28363 : NOR2_X2 port map( A1 => n15468, A2 => n15467, ZN => n16574);
   U28364 : NAND2_X1 port map( A1 => n29770, A2 => n7619, ZN => n7360);
   U28365 : OAI22_X1 port map( A1 => n8236, A2 => n7920, B1 => n8231, B2 => 
                           n7919, ZN => n29770);
   U28366 : NAND3_X1 port map( A1 => n19976, A2 => n6114, A3 => n504, ZN => 
                           n4889);
   U28367 : NAND2_X1 port map( A1 => n29002, A2 => n29003, ZN => n23240);
   U28368 : AND3_X2 port map( A1 => n24535, A2 => n132, A3 => n24537, ZN => 
                           n26080);
   U28369 : NAND2_X1 port map( A1 => n16866, A2 => n17824, ZN => n16867);
   U28370 : NAND2_X1 port map( A1 => n27666, A2 => n28373, ZN => n27670);
   U28371 : NAND2_X1 port map( A1 => n14285, A2 => n14084, ZN => n4451);
   U28372 : NAND2_X1 port map( A1 => n7843, A2 => n29772, ZN => n29771);
   U28373 : OR2_X1 port map( A1 => n10929, A2 => n10932, ZN => n9467);
   U28374 : OR2_X2 port map( A1 => n29773, A2 => n16545, ZN => n16611);
   U28375 : NAND2_X1 port map( A1 => n16542, A2 => n16543, ZN => n29773);
   U28376 : OR2_X2 port map( A1 => n10495, A2 => n10496, ZN => n11869);
   U28377 : OAI21_X1 port map( B1 => n16881, B2 => n17495, A => n17062, ZN => 
                           n29774);
   U28378 : NAND2_X1 port map( A1 => n29775, A2 => n23200, ZN => n24634);
   U28379 : OAI21_X1 port map( B1 => n28955, B2 => n28954, A => n23795, ZN => 
                           n29775);
   U28380 : INV_X1 port map( A => n23705, ZN => n3616);
   U28381 : NOR2_X1 port map( A1 => n23707, A2 => n29776, ZN => n23708);
   U28382 : NAND2_X1 port map( A1 => n29777, A2 => n23705, ZN => n29776);
   U28383 : NAND2_X1 port map( A1 => n23706, A2 => n29618, ZN => n23705);
   U28384 : INV_X1 port map( A => n22451, ZN => n29777);
   U28385 : INV_X1 port map( A => n22863, ZN => n5541);
   U28386 : NAND2_X1 port map( A1 => n23297, A2 => n23831, ZN => n22863);
   U28387 : NAND3_X2 port map( A1 => n1177, A2 => n1176, A3 => n6049, ZN => 
                           n24817);
   U28388 : NAND2_X1 port map( A1 => n29781, A2 => n29779, ZN => n1078);
   U28389 : NAND2_X1 port map( A1 => n29780, A2 => n21603, ZN => n29779);
   U28390 : NAND2_X1 port map( A1 => n21605, A2 => n20721, ZN => n29780);
   U28391 : NAND2_X1 port map( A1 => n29782, A2 => n20649, ZN => n29781);
   U28392 : INV_X1 port map( A => n21603, ZN => n29782);
   U28393 : NAND2_X1 port map( A1 => n24376, A2 => n1883, ZN => n23093);
   U28394 : NAND2_X2 port map( A1 => n23120, A2 => n23121, ZN => n25845);
   U28395 : OR2_X1 port map( A1 => n11490, A2 => n11431, ZN => n2302);
   U28396 : AOI22_X1 port map( A1 => n11429, A2 => n11428, B1 => n6482, B2 => 
                           n11794, ZN => n11490);
   U28397 : XNOR2_X1 port map( A => n16252, B => n16414, ZN => n15625);
   U28398 : OAI211_X2 port map( C1 => n15461, C2 => n15460, A => n1702, B => 
                           n1701, ZN => n16252);
   U28399 : AND2_X2 port map( A1 => n28363, A2 => n28364, ZN => n12232);
   U28400 : XNOR2_X1 port map( A => n29784, B => n29783, ZN => Ciphertext(35));
   U28401 : INV_X1 port map( A => n3516, ZN => n29783);
   U28402 : NAND2_X1 port map( A1 => n29786, A2 => n29785, ZN => n29784);
   U28403 : NAND2_X1 port map( A1 => n26706, A2 => n28592, ZN => n29785);
   U28404 : NAND2_X1 port map( A1 => n26705, A2 => n393, ZN => n29786);
   U28405 : NAND3_X1 port map( A1 => n23529, A2 => n23531, A3 => n28164, ZN => 
                           n23532);
   U28406 : XNOR2_X2 port map( A => n20061, B => n20062, ZN => n28164);
   U28407 : OAI211_X2 port map( C1 => n15051, C2 => n15052, A => n29787, B => 
                           n28872, ZN => n16480);
   U28408 : XNOR2_X1 port map( A => n15870, B => n28585, ZN => n15871);
   U28409 : OAI21_X2 port map( B1 => n15461, B2 => n14980, A => n14798, ZN => 
                           n28585);
   U28410 : NAND2_X1 port map( A1 => n29791, A2 => n29788, ZN => n26803);
   U28411 : NAND2_X1 port map( A1 => n29790, A2 => n29789, ZN => n29788);
   U28412 : NOR2_X1 port map( A1 => n26797, A2 => n26800, ZN => n29789);
   U28413 : NAND2_X1 port map( A1 => n26798, A2 => n26799, ZN => n29790);
   U28414 : NAND2_X1 port map( A1 => n26801, A2 => n26800, ZN => n29791);
   U28415 : NAND2_X1 port map( A1 => n5961, A2 => n8527, ZN => n5960);
   U28416 : NAND2_X1 port map( A1 => n906, A2 => n29328, ZN => n6602);
   U28417 : NAND2_X1 port map( A1 => n5639, A2 => n17436, ZN => n237);
   U28418 : OAI21_X1 port map( B1 => n1930, B2 => n29793, A => n29792, ZN => 
                           n20662);
   U28419 : NAND2_X1 port map( A1 => n1929, A2 => n29314, ZN => n29792);
   U28420 : INV_X1 port map( A => n21472, ZN => n29793);
   U28421 : AOI21_X1 port map( B1 => n7524, B2 => n7748, A => n7533, ZN => 
                           n29794);
   U28422 : NAND3_X1 port map( A1 => n29795, A2 => n10842, A3 => n10843, ZN => 
                           n10845);
   U28423 : NAND2_X1 port map( A1 => n1812, A2 => n11038, ZN => n29795);
   U28424 : OAI21_X2 port map( B1 => n8094, B2 => n9037, A => n29796, ZN => 
                           n9878);
   U28425 : NAND2_X1 port map( A1 => n6092, A2 => n8792, ZN => n29796);
   U28426 : NAND2_X1 port map( A1 => n23427, A2 => n28122, ZN => n23340);
   U28427 : NOR2_X1 port map( A1 => n17611, A2 => n29797, ZN => n18408);
   U28428 : XNOR2_X1 port map( A => n6270, B => n13542, ZN => n29798);
   U28429 : NAND2_X1 port map( A1 => n12511, A2 => n3653, ZN => n11994);
   U28430 : NOR2_X1 port map( A1 => n1746, A2 => n12507, ZN => n12511);
   U28431 : XNOR2_X1 port map( A => n29799, B => n2523, ZN => Ciphertext(164));
   U28432 : NAND2_X1 port map( A1 => n3064, A2 => n3063, ZN => n29799);
   U28433 : AOI21_X2 port map( B1 => n14219, B2 => n29800, A => n6231, ZN => 
                           n15333);
   U28434 : NAND2_X1 port map( A1 => n3045, A2 => n6466, ZN => n29800);
   U28435 : NAND3_X2 port map( A1 => n11525, A2 => n11526, A3 => n11523, ZN => 
                           n11982);
   U28436 : XNOR2_X1 port map( A => n29801, B => n10346, ZN => n9663);
   U28437 : XNOR2_X1 port map( A => n1891, B => n3501, ZN => n29801);
   U28438 : NOR2_X1 port map( A1 => n29570, A2 => n28783, ZN => n26633);
   U28439 : AOI22_X1 port map( A1 => n19990, A2 => n20166, B1 => n385, B2 => 
                           n19991, ZN => n1460);
   U28440 : NOR3_X1 port map( A1 => n18372, A2 => n18337, A3 => n18370, ZN => 
                           n17888);
   U28441 : XNOR2_X2 port map( A => n15157, B => n15158, ZN => n17421);
   U28442 : XNOR2_X2 port map( A => n15549, B => n15550, ZN => n17347);
   U28443 : NOR2_X2 port map( A1 => n26638, A2 => n26639, ZN => n29095);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Top is

   port( clk : in std_logic;  Plaintext, Key : in std_logic_vector (191 downto 
         0);  Ciphertext : out std_logic_vector (191 downto 0));

end SPEEDY_Top;

architecture SYN_Behavioral of SPEEDY_Top is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SPEEDY_Rounds7_0
      port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : 
            out std_logic_vector (191 downto 0));
   end component;
   
   signal reg_in_191_port, reg_in_190_port, reg_in_189_port, reg_in_188_port, 
      reg_in_187_port, reg_in_186_port, reg_in_185_port, reg_in_184_port, 
      reg_in_183_port, reg_in_182_port, reg_in_181_port, reg_in_180_port, 
      reg_in_179_port, reg_in_178_port, reg_in_177_port, reg_in_176_port, 
      reg_in_175_port, reg_in_174_port, reg_in_173_port, reg_in_172_port, 
      reg_in_171_port, reg_in_170_port, reg_in_169_port, reg_in_168_port, 
      reg_in_167_port, reg_in_166_port, reg_in_165_port, reg_in_164_port, 
      reg_in_163_port, reg_in_162_port, reg_in_161_port, reg_in_160_port, 
      reg_in_159_port, reg_in_158_port, reg_in_157_port, reg_in_156_port, 
      reg_in_155_port, reg_in_154_port, reg_in_153_port, reg_in_152_port, 
      reg_in_151_port, reg_in_150_port, reg_in_149_port, reg_in_148_port, 
      reg_in_147_port, reg_in_146_port, reg_in_145_port, reg_in_144_port, 
      reg_in_143_port, reg_in_142_port, reg_in_141_port, reg_in_140_port, 
      reg_in_139_port, reg_in_138_port, reg_in_137_port, reg_in_136_port, 
      reg_in_135_port, reg_in_134_port, reg_in_133_port, reg_in_132_port, 
      reg_in_131_port, reg_in_130_port, reg_in_129_port, reg_in_128_port, 
      reg_in_127_port, reg_in_126_port, reg_in_125_port, reg_in_124_port, 
      reg_in_123_port, reg_in_122_port, reg_in_121_port, reg_in_120_port, 
      reg_in_119_port, reg_in_118_port, reg_in_117_port, reg_in_116_port, 
      reg_in_115_port, reg_in_114_port, reg_in_113_port, reg_in_112_port, 
      reg_in_111_port, reg_in_110_port, reg_in_109_port, reg_in_108_port, 
      reg_in_107_port, reg_in_106_port, reg_in_105_port, reg_in_104_port, 
      reg_in_103_port, reg_in_102_port, reg_in_101_port, reg_in_100_port, 
      reg_in_99_port, reg_in_98_port, reg_in_97_port, reg_in_96_port, 
      reg_in_95_port, reg_in_94_port, reg_in_93_port, reg_in_92_port, 
      reg_in_91_port, reg_in_90_port, reg_in_89_port, reg_in_88_port, 
      reg_in_87_port, reg_in_86_port, reg_in_85_port, reg_in_84_port, 
      reg_in_83_port, reg_in_82_port, reg_in_81_port, reg_in_80_port, 
      reg_in_79_port, reg_in_78_port, reg_in_77_port, reg_in_76_port, 
      reg_in_75_port, reg_in_74_port, reg_in_73_port, reg_in_72_port, 
      reg_in_71_port, reg_in_70_port, reg_in_69_port, reg_in_68_port, 
      reg_in_67_port, reg_in_66_port, reg_in_65_port, reg_in_64_port, 
      reg_in_63_port, reg_in_62_port, reg_in_61_port, reg_in_60_port, 
      reg_in_59_port, reg_in_58_port, reg_in_57_port, reg_in_56_port, 
      reg_in_55_port, reg_in_54_port, reg_in_53_port, reg_in_52_port, 
      reg_in_51_port, reg_in_50_port, reg_in_49_port, reg_in_48_port, 
      reg_in_47_port, reg_in_46_port, reg_in_45_port, reg_in_44_port, 
      reg_in_43_port, reg_in_42_port, reg_in_41_port, reg_in_40_port, 
      reg_in_39_port, reg_in_38_port, reg_in_37_port, reg_in_36_port, 
      reg_in_35_port, reg_in_34_port, reg_in_33_port, reg_in_32_port, 
      reg_in_31_port, reg_in_30_port, reg_in_29_port, reg_in_28_port, 
      reg_in_27_port, reg_in_26_port, reg_in_25_port, reg_in_24_port, 
      reg_in_23_port, reg_in_22_port, reg_in_21_port, reg_in_20_port, 
      reg_in_19_port, reg_in_18_port, reg_in_17_port, reg_in_16_port, 
      reg_in_15_port, reg_in_14_port, reg_in_13_port, reg_in_12_port, 
      reg_in_11_port, reg_in_10_port, reg_in_9_port, reg_in_8_port, 
      reg_in_7_port, reg_in_6_port, reg_in_5_port, reg_in_4_port, reg_in_3_port
      , reg_in_2_port, reg_in_1_port, reg_in_0_port, reg_key_191_port, 
      reg_key_190_port, reg_key_189_port, reg_key_188_port, reg_key_187_port, 
      reg_key_186_port, reg_key_185_port, reg_key_184_port, reg_key_183_port, 
      reg_key_182_port, reg_key_181_port, reg_key_180_port, reg_key_179_port, 
      reg_key_178_port, reg_key_177_port, reg_key_176_port, reg_key_175_port, 
      reg_key_174_port, reg_key_173_port, reg_key_172_port, reg_key_171_port, 
      reg_key_170_port, reg_key_169_port, reg_key_168_port, reg_key_167_port, 
      reg_key_166_port, reg_key_165_port, reg_key_164_port, reg_key_163_port, 
      reg_key_162_port, reg_key_161_port, reg_key_160_port, reg_key_159_port, 
      reg_key_158_port, reg_key_157_port, reg_key_156_port, reg_key_155_port, 
      reg_key_154_port, reg_key_153_port, reg_key_152_port, reg_key_151_port, 
      reg_key_150_port, reg_key_149_port, reg_key_148_port, reg_key_147_port, 
      reg_key_146_port, reg_key_145_port, reg_key_144_port, reg_key_143_port, 
      reg_key_142_port, reg_key_141_port, reg_key_140_port, reg_key_139_port, 
      reg_key_138_port, reg_key_137_port, reg_key_136_port, reg_key_135_port, 
      reg_key_134_port, reg_key_133_port, reg_key_132_port, reg_key_131_port, 
      reg_key_130_port, reg_key_129_port, reg_key_128_port, reg_key_127_port, 
      reg_key_126_port, reg_key_125_port, reg_key_124_port, reg_key_123_port, 
      reg_key_122_port, reg_key_121_port, reg_key_120_port, reg_key_119_port, 
      reg_key_118_port, reg_key_117_port, reg_key_116_port, reg_key_115_port, 
      reg_key_114_port, reg_key_113_port, reg_key_112_port, reg_key_111_port, 
      reg_key_110_port, reg_key_109_port, reg_key_108_port, reg_key_107_port, 
      reg_key_106_port, reg_key_105_port, reg_key_104_port, reg_key_103_port, 
      reg_key_102_port, reg_key_101_port, reg_key_100_port, reg_key_99_port, 
      reg_key_98_port, reg_key_97_port, reg_key_96_port, reg_key_95_port, 
      reg_key_94_port, reg_key_93_port, reg_key_92_port, reg_key_91_port, 
      reg_key_90_port, reg_key_89_port, reg_key_88_port, reg_key_87_port, 
      reg_key_86_port, reg_key_85_port, reg_key_84_port, reg_key_83_port, 
      reg_key_82_port, reg_key_81_port, reg_key_80_port, reg_key_79_port, 
      reg_key_78_port, reg_key_77_port, reg_key_76_port, reg_key_75_port, 
      reg_key_74_port, reg_key_73_port, reg_key_72_port, reg_key_71_port, 
      reg_key_70_port, reg_key_69_port, reg_key_68_port, reg_key_67_port, 
      reg_key_66_port, reg_key_65_port, reg_key_64_port, reg_key_63_port, 
      reg_key_62_port, reg_key_61_port, reg_key_60_port, reg_key_59_port, 
      reg_key_58_port, reg_key_57_port, reg_key_56_port, reg_key_55_port, 
      reg_key_54_port, reg_key_53_port, reg_key_52_port, reg_key_51_port, 
      reg_key_50_port, reg_key_49_port, reg_key_48_port, reg_key_47_port, 
      reg_key_46_port, reg_key_45_port, reg_key_44_port, reg_key_43_port, 
      reg_key_42_port, reg_key_41_port, reg_key_40_port, reg_key_39_port, 
      reg_key_38_port, reg_key_37_port, reg_key_36_port, reg_key_35_port, 
      reg_key_34_port, reg_key_33_port, reg_key_32_port, reg_key_31_port, 
      reg_key_30_port, reg_key_29_port, reg_key_28_port, reg_key_27_port, 
      reg_key_26_port, reg_key_25_port, reg_key_24_port, reg_key_23_port, 
      reg_key_22_port, reg_key_21_port, reg_key_20_port, reg_key_19_port, 
      reg_key_18_port, reg_key_17_port, reg_key_16_port, reg_key_15_port, 
      reg_key_14_port, reg_key_13_port, reg_key_12_port, reg_key_11_port, 
      reg_key_10_port, reg_key_9_port, reg_key_8_port, reg_key_7_port, 
      reg_key_6_port, reg_key_5_port, reg_key_4_port, reg_key_3_port, 
      reg_key_2_port, reg_key_1_port, reg_key_0_port, reg_out_191_port, 
      reg_out_190_port, reg_out_189_port, reg_out_188_port, reg_out_187_port, 
      reg_out_186_port, reg_out_185_port, reg_out_184_port, reg_out_183_port, 
      reg_out_182_port, reg_out_181_port, reg_out_180_port, reg_out_179_port, 
      reg_out_178_port, reg_out_177_port, reg_out_176_port, reg_out_175_port, 
      reg_out_174_port, reg_out_173_port, reg_out_172_port, reg_out_171_port, 
      reg_out_170_port, reg_out_169_port, reg_out_168_port, reg_out_167_port, 
      reg_out_166_port, reg_out_165_port, reg_out_164_port, reg_out_163_port, 
      reg_out_162_port, reg_out_161_port, reg_out_160_port, reg_out_159_port, 
      reg_out_158_port, reg_out_157_port, reg_out_156_port, reg_out_155_port, 
      reg_out_154_port, reg_out_153_port, reg_out_152_port, reg_out_151_port, 
      reg_out_150_port, reg_out_149_port, reg_out_148_port, reg_out_147_port, 
      reg_out_146_port, reg_out_145_port, reg_out_144_port, reg_out_143_port, 
      reg_out_142_port, reg_out_141_port, reg_out_140_port, reg_out_139_port, 
      reg_out_138_port, reg_out_137_port, reg_out_136_port, reg_out_135_port, 
      reg_out_134_port, reg_out_133_port, reg_out_132_port, reg_out_131_port, 
      reg_out_130_port, reg_out_129_port, reg_out_128_port, reg_out_127_port, 
      reg_out_126_port, reg_out_125_port, reg_out_124_port, reg_out_123_port, 
      reg_out_122_port, reg_out_121_port, reg_out_120_port, reg_out_119_port, 
      reg_out_118_port, reg_out_117_port, reg_out_116_port, reg_out_115_port, 
      reg_out_114_port, reg_out_113_port, reg_out_112_port, reg_out_111_port, 
      reg_out_110_port, reg_out_109_port, reg_out_108_port, reg_out_107_port, 
      reg_out_106_port, reg_out_105_port, reg_out_104_port, reg_out_103_port, 
      reg_out_102_port, reg_out_101_port, reg_out_100_port, reg_out_99_port, 
      reg_out_98_port, reg_out_97_port, reg_out_96_port, reg_out_95_port, 
      reg_out_94_port, reg_out_93_port, reg_out_92_port, reg_out_91_port, 
      reg_out_90_port, reg_out_89_port, reg_out_88_port, reg_out_87_port, 
      reg_out_86_port, reg_out_85_port, reg_out_84_port, reg_out_83_port, 
      reg_out_82_port, reg_out_81_port, reg_out_80_port, reg_out_79_port, 
      reg_out_78_port, reg_out_77_port, reg_out_76_port, reg_out_75_port, 
      reg_out_74_port, reg_out_73_port, reg_out_72_port, reg_out_71_port, 
      reg_out_70_port, reg_out_69_port, reg_out_68_port, reg_out_67_port, 
      reg_out_66_port, reg_out_65_port, reg_out_64_port, reg_out_63_port, 
      reg_out_62_port, reg_out_61_port, reg_out_60_port, reg_out_59_port, 
      reg_out_58_port, reg_out_57_port, reg_out_56_port, reg_out_55_port, 
      reg_out_54_port, reg_out_53_port, reg_out_52_port, reg_out_51_port, 
      reg_out_50_port, reg_out_49_port, reg_out_48_port, reg_out_47_port, 
      reg_out_46_port, reg_out_45_port, reg_out_44_port, reg_out_43_port, 
      reg_out_42_port, reg_out_41_port, reg_out_40_port, reg_out_39_port, 
      reg_out_38_port, reg_out_37_port, reg_out_36_port, reg_out_35_port, 
      reg_out_34_port, reg_out_33_port, reg_out_32_port, reg_out_31_port, 
      reg_out_30_port, reg_out_29_port, reg_out_28_port, reg_out_27_port, 
      reg_out_26_port, reg_out_25_port, reg_out_24_port, reg_out_23_port, 
      reg_out_22_port, reg_out_21_port, reg_out_20_port, reg_out_19_port, 
      reg_out_18_port, reg_out_17_port, reg_out_16_port, reg_out_15_port, 
      reg_out_14_port, reg_out_13_port, reg_out_12_port, reg_out_11_port, 
      reg_out_10_port, reg_out_9_port, reg_out_8_port, reg_out_7_port, 
      reg_out_6_port, reg_out_5_port, reg_out_4_port, reg_out_3_port, 
      reg_out_2_port, reg_out_1_port, reg_out_0_port, n10, n12, n_1000, n_1001,
      n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575 : std_logic;

begin
   
   reg_in_regx191x : DFF_X1 port map( D => Plaintext(191), CK => clk, Q => 
                           reg_in_191_port, QN => n_1000);
   reg_in_regx190x : DFF_X1 port map( D => Plaintext(190), CK => clk, Q => 
                           reg_in_190_port, QN => n_1001);
   reg_in_regx189x : DFF_X1 port map( D => Plaintext(189), CK => clk, Q => 
                           reg_in_189_port, QN => n_1002);
   reg_in_regx188x : DFF_X1 port map( D => Plaintext(188), CK => clk, Q => 
                           reg_in_188_port, QN => n_1003);
   reg_in_regx187x : DFF_X1 port map( D => Plaintext(187), CK => clk, Q => 
                           reg_in_187_port, QN => n_1004);
   reg_in_regx186x : DFF_X1 port map( D => Plaintext(186), CK => clk, Q => 
                           reg_in_186_port, QN => n_1005);
   reg_in_regx185x : DFF_X1 port map( D => Plaintext(185), CK => clk, Q => 
                           reg_in_185_port, QN => n_1006);
   reg_in_regx184x : DFF_X1 port map( D => Plaintext(184), CK => clk, Q => 
                           reg_in_184_port, QN => n_1007);
   reg_in_regx183x : DFF_X1 port map( D => Plaintext(183), CK => clk, Q => 
                           reg_in_183_port, QN => n_1008);
   reg_in_regx182x : DFF_X1 port map( D => Plaintext(182), CK => clk, Q => 
                           reg_in_182_port, QN => n_1009);
   reg_in_regx181x : DFF_X1 port map( D => Plaintext(181), CK => clk, Q => 
                           reg_in_181_port, QN => n_1010);
   reg_in_regx180x : DFF_X1 port map( D => Plaintext(180), CK => clk, Q => 
                           reg_in_180_port, QN => n_1011);
   reg_in_regx179x : DFF_X1 port map( D => Plaintext(179), CK => clk, Q => 
                           reg_in_179_port, QN => n_1012);
   reg_in_regx178x : DFF_X1 port map( D => Plaintext(178), CK => clk, Q => 
                           reg_in_178_port, QN => n_1013);
   reg_in_regx177x : DFF_X1 port map( D => Plaintext(177), CK => clk, Q => 
                           reg_in_177_port, QN => n_1014);
   reg_in_regx176x : DFF_X1 port map( D => Plaintext(176), CK => clk, Q => 
                           reg_in_176_port, QN => n_1015);
   reg_in_regx175x : DFF_X1 port map( D => Plaintext(175), CK => clk, Q => 
                           reg_in_175_port, QN => n_1016);
   reg_in_regx174x : DFF_X1 port map( D => Plaintext(174), CK => clk, Q => 
                           reg_in_174_port, QN => n_1017);
   reg_in_regx173x : DFF_X1 port map( D => Plaintext(173), CK => clk, Q => 
                           reg_in_173_port, QN => n_1018);
   reg_in_regx172x : DFF_X1 port map( D => Plaintext(172), CK => clk, Q => 
                           reg_in_172_port, QN => n_1019);
   reg_in_regx171x : DFF_X1 port map( D => Plaintext(171), CK => clk, Q => 
                           reg_in_171_port, QN => n_1020);
   reg_in_regx170x : DFF_X1 port map( D => Plaintext(170), CK => clk, Q => 
                           reg_in_170_port, QN => n_1021);
   reg_in_regx169x : DFF_X1 port map( D => Plaintext(169), CK => clk, Q => 
                           reg_in_169_port, QN => n_1022);
   reg_in_regx168x : DFF_X1 port map( D => Plaintext(168), CK => clk, Q => 
                           reg_in_168_port, QN => n_1023);
   reg_in_regx167x : DFF_X1 port map( D => Plaintext(167), CK => clk, Q => 
                           reg_in_167_port, QN => n_1024);
   reg_in_regx166x : DFF_X1 port map( D => Plaintext(166), CK => clk, Q => 
                           reg_in_166_port, QN => n_1025);
   reg_in_regx165x : DFF_X1 port map( D => Plaintext(165), CK => clk, Q => 
                           reg_in_165_port, QN => n_1026);
   reg_in_regx164x : DFF_X1 port map( D => Plaintext(164), CK => clk, Q => 
                           reg_in_164_port, QN => n_1027);
   reg_in_regx163x : DFF_X1 port map( D => Plaintext(163), CK => clk, Q => 
                           reg_in_163_port, QN => n_1028);
   reg_in_regx162x : DFF_X1 port map( D => Plaintext(162), CK => clk, Q => 
                           reg_in_162_port, QN => n_1029);
   reg_in_regx161x : DFF_X1 port map( D => Plaintext(161), CK => clk, Q => 
                           reg_in_161_port, QN => n_1030);
   reg_in_regx160x : DFF_X1 port map( D => Plaintext(160), CK => clk, Q => 
                           reg_in_160_port, QN => n_1031);
   reg_in_regx159x : DFF_X1 port map( D => Plaintext(159), CK => clk, Q => 
                           reg_in_159_port, QN => n_1032);
   reg_in_regx158x : DFF_X1 port map( D => Plaintext(158), CK => clk, Q => 
                           reg_in_158_port, QN => n_1033);
   reg_in_regx157x : DFF_X1 port map( D => Plaintext(157), CK => clk, Q => 
                           reg_in_157_port, QN => n_1034);
   reg_in_regx156x : DFF_X1 port map( D => Plaintext(156), CK => clk, Q => 
                           reg_in_156_port, QN => n_1035);
   reg_in_regx155x : DFF_X1 port map( D => Plaintext(155), CK => clk, Q => 
                           reg_in_155_port, QN => n_1036);
   reg_in_regx154x : DFF_X1 port map( D => Plaintext(154), CK => clk, Q => 
                           reg_in_154_port, QN => n_1037);
   reg_in_regx153x : DFF_X1 port map( D => Plaintext(153), CK => clk, Q => 
                           reg_in_153_port, QN => n_1038);
   reg_in_regx152x : DFF_X1 port map( D => Plaintext(152), CK => clk, Q => 
                           reg_in_152_port, QN => n_1039);
   reg_in_regx151x : DFF_X1 port map( D => Plaintext(151), CK => clk, Q => 
                           reg_in_151_port, QN => n_1040);
   reg_in_regx150x : DFF_X1 port map( D => Plaintext(150), CK => clk, Q => 
                           reg_in_150_port, QN => n_1041);
   reg_in_regx149x : DFF_X1 port map( D => Plaintext(149), CK => clk, Q => 
                           reg_in_149_port, QN => n_1042);
   reg_in_regx148x : DFF_X1 port map( D => Plaintext(148), CK => clk, Q => 
                           reg_in_148_port, QN => n_1043);
   reg_in_regx147x : DFF_X1 port map( D => Plaintext(147), CK => clk, Q => 
                           reg_in_147_port, QN => n_1044);
   reg_in_regx146x : DFF_X1 port map( D => Plaintext(146), CK => clk, Q => 
                           reg_in_146_port, QN => n_1045);
   reg_in_regx145x : DFF_X1 port map( D => Plaintext(145), CK => clk, Q => 
                           reg_in_145_port, QN => n_1046);
   reg_in_regx144x : DFF_X1 port map( D => Plaintext(144), CK => clk, Q => 
                           reg_in_144_port, QN => n_1047);
   reg_in_regx143x : DFF_X1 port map( D => Plaintext(143), CK => clk, Q => 
                           reg_in_143_port, QN => n_1048);
   reg_in_regx142x : DFF_X1 port map( D => Plaintext(142), CK => clk, Q => 
                           reg_in_142_port, QN => n_1049);
   reg_in_regx141x : DFF_X1 port map( D => Plaintext(141), CK => clk, Q => 
                           reg_in_141_port, QN => n_1050);
   reg_in_regx140x : DFF_X1 port map( D => Plaintext(140), CK => clk, Q => 
                           reg_in_140_port, QN => n_1051);
   reg_in_regx139x : DFF_X1 port map( D => Plaintext(139), CK => clk, Q => 
                           reg_in_139_port, QN => n_1052);
   reg_in_regx138x : DFF_X1 port map( D => Plaintext(138), CK => clk, Q => 
                           reg_in_138_port, QN => n_1053);
   reg_in_regx137x : DFF_X1 port map( D => Plaintext(137), CK => clk, Q => 
                           reg_in_137_port, QN => n_1054);
   reg_in_regx136x : DFF_X1 port map( D => Plaintext(136), CK => clk, Q => 
                           reg_in_136_port, QN => n_1055);
   reg_in_regx135x : DFF_X1 port map( D => Plaintext(135), CK => clk, Q => 
                           reg_in_135_port, QN => n_1056);
   reg_in_regx134x : DFF_X1 port map( D => Plaintext(134), CK => clk, Q => 
                           reg_in_134_port, QN => n_1057);
   reg_in_regx133x : DFF_X1 port map( D => Plaintext(133), CK => clk, Q => 
                           reg_in_133_port, QN => n_1058);
   reg_in_regx132x : DFF_X1 port map( D => Plaintext(132), CK => clk, Q => 
                           reg_in_132_port, QN => n_1059);
   reg_in_regx131x : DFF_X1 port map( D => Plaintext(131), CK => clk, Q => 
                           reg_in_131_port, QN => n_1060);
   reg_in_regx130x : DFF_X1 port map( D => Plaintext(130), CK => clk, Q => 
                           reg_in_130_port, QN => n_1061);
   reg_in_regx129x : DFF_X1 port map( D => Plaintext(129), CK => clk, Q => 
                           reg_in_129_port, QN => n_1062);
   reg_in_regx128x : DFF_X1 port map( D => Plaintext(128), CK => clk, Q => 
                           reg_in_128_port, QN => n_1063);
   reg_in_regx127x : DFF_X1 port map( D => Plaintext(127), CK => clk, Q => 
                           reg_in_127_port, QN => n_1064);
   reg_in_regx126x : DFF_X1 port map( D => Plaintext(126), CK => clk, Q => 
                           reg_in_126_port, QN => n_1065);
   reg_in_regx125x : DFF_X1 port map( D => Plaintext(125), CK => clk, Q => 
                           reg_in_125_port, QN => n_1066);
   reg_in_regx124x : DFF_X1 port map( D => Plaintext(124), CK => clk, Q => 
                           reg_in_124_port, QN => n_1067);
   reg_in_regx123x : DFF_X1 port map( D => Plaintext(123), CK => clk, Q => 
                           reg_in_123_port, QN => n_1068);
   reg_in_regx122x : DFF_X1 port map( D => Plaintext(122), CK => clk, Q => 
                           reg_in_122_port, QN => n_1069);
   reg_in_regx121x : DFF_X1 port map( D => Plaintext(121), CK => clk, Q => 
                           reg_in_121_port, QN => n_1070);
   reg_in_regx120x : DFF_X1 port map( D => Plaintext(120), CK => clk, Q => 
                           reg_in_120_port, QN => n_1071);
   reg_in_regx119x : DFF_X1 port map( D => Plaintext(119), CK => clk, Q => 
                           reg_in_119_port, QN => n_1072);
   reg_in_regx118x : DFF_X1 port map( D => Plaintext(118), CK => clk, Q => 
                           reg_in_118_port, QN => n_1073);
   reg_in_regx117x : DFF_X1 port map( D => Plaintext(117), CK => clk, Q => 
                           reg_in_117_port, QN => n_1074);
   reg_in_regx116x : DFF_X1 port map( D => Plaintext(116), CK => clk, Q => 
                           reg_in_116_port, QN => n_1075);
   reg_in_regx115x : DFF_X1 port map( D => Plaintext(115), CK => clk, Q => 
                           reg_in_115_port, QN => n_1076);
   reg_in_regx114x : DFF_X1 port map( D => Plaintext(114), CK => clk, Q => 
                           reg_in_114_port, QN => n_1077);
   reg_in_regx113x : DFF_X1 port map( D => Plaintext(113), CK => clk, Q => 
                           reg_in_113_port, QN => n_1078);
   reg_in_regx112x : DFF_X1 port map( D => Plaintext(112), CK => clk, Q => 
                           reg_in_112_port, QN => n_1079);
   reg_in_regx111x : DFF_X1 port map( D => Plaintext(111), CK => clk, Q => 
                           reg_in_111_port, QN => n_1080);
   reg_in_regx110x : DFF_X1 port map( D => Plaintext(110), CK => clk, Q => 
                           reg_in_110_port, QN => n_1081);
   reg_in_regx109x : DFF_X1 port map( D => Plaintext(109), CK => clk, Q => 
                           reg_in_109_port, QN => n_1082);
   reg_in_regx108x : DFF_X1 port map( D => Plaintext(108), CK => clk, Q => 
                           reg_in_108_port, QN => n_1083);
   reg_in_regx107x : DFF_X1 port map( D => Plaintext(107), CK => clk, Q => 
                           reg_in_107_port, QN => n_1084);
   reg_in_regx106x : DFF_X1 port map( D => Plaintext(106), CK => clk, Q => 
                           reg_in_106_port, QN => n_1085);
   reg_in_regx105x : DFF_X1 port map( D => Plaintext(105), CK => clk, Q => 
                           reg_in_105_port, QN => n_1086);
   reg_in_regx104x : DFF_X1 port map( D => Plaintext(104), CK => clk, Q => 
                           reg_in_104_port, QN => n_1087);
   reg_in_regx103x : DFF_X1 port map( D => Plaintext(103), CK => clk, Q => 
                           reg_in_103_port, QN => n_1088);
   reg_in_regx102x : DFF_X1 port map( D => Plaintext(102), CK => clk, Q => 
                           reg_in_102_port, QN => n_1089);
   reg_in_regx101x : DFF_X1 port map( D => Plaintext(101), CK => clk, Q => 
                           reg_in_101_port, QN => n_1090);
   reg_in_regx100x : DFF_X1 port map( D => Plaintext(100), CK => clk, Q => 
                           reg_in_100_port, QN => n_1091);
   reg_in_regx99x : DFF_X1 port map( D => Plaintext(99), CK => clk, Q => 
                           reg_in_99_port, QN => n_1092);
   reg_in_regx98x : DFF_X1 port map( D => Plaintext(98), CK => clk, Q => 
                           reg_in_98_port, QN => n_1093);
   reg_in_regx97x : DFF_X1 port map( D => Plaintext(97), CK => clk, Q => 
                           reg_in_97_port, QN => n_1094);
   reg_in_regx96x : DFF_X1 port map( D => Plaintext(96), CK => clk, Q => 
                           reg_in_96_port, QN => n_1095);
   reg_in_regx95x : DFF_X1 port map( D => Plaintext(95), CK => clk, Q => 
                           reg_in_95_port, QN => n_1096);
   reg_in_regx94x : DFF_X1 port map( D => Plaintext(94), CK => clk, Q => 
                           reg_in_94_port, QN => n_1097);
   reg_in_regx93x : DFF_X1 port map( D => Plaintext(93), CK => clk, Q => 
                           reg_in_93_port, QN => n_1098);
   reg_in_regx92x : DFF_X1 port map( D => Plaintext(92), CK => clk, Q => 
                           reg_in_92_port, QN => n_1099);
   reg_in_regx91x : DFF_X1 port map( D => Plaintext(91), CK => clk, Q => 
                           reg_in_91_port, QN => n_1100);
   reg_in_regx90x : DFF_X1 port map( D => Plaintext(90), CK => clk, Q => 
                           reg_in_90_port, QN => n_1101);
   reg_in_regx89x : DFF_X1 port map( D => Plaintext(89), CK => clk, Q => 
                           reg_in_89_port, QN => n_1102);
   reg_in_regx88x : DFF_X1 port map( D => Plaintext(88), CK => clk, Q => 
                           reg_in_88_port, QN => n_1103);
   reg_in_regx87x : DFF_X1 port map( D => Plaintext(87), CK => clk, Q => 
                           reg_in_87_port, QN => n_1104);
   reg_in_regx86x : DFF_X1 port map( D => Plaintext(86), CK => clk, Q => 
                           reg_in_86_port, QN => n_1105);
   reg_in_regx85x : DFF_X1 port map( D => Plaintext(85), CK => clk, Q => 
                           reg_in_85_port, QN => n_1106);
   reg_in_regx84x : DFF_X1 port map( D => Plaintext(84), CK => clk, Q => 
                           reg_in_84_port, QN => n_1107);
   reg_in_regx83x : DFF_X1 port map( D => Plaintext(83), CK => clk, Q => 
                           reg_in_83_port, QN => n_1108);
   reg_in_regx82x : DFF_X1 port map( D => Plaintext(82), CK => clk, Q => 
                           reg_in_82_port, QN => n_1109);
   reg_in_regx81x : DFF_X1 port map( D => Plaintext(81), CK => clk, Q => 
                           reg_in_81_port, QN => n_1110);
   reg_in_regx80x : DFF_X1 port map( D => Plaintext(80), CK => clk, Q => 
                           reg_in_80_port, QN => n_1111);
   reg_in_regx79x : DFF_X1 port map( D => Plaintext(79), CK => clk, Q => 
                           reg_in_79_port, QN => n_1112);
   reg_in_regx78x : DFF_X1 port map( D => Plaintext(78), CK => clk, Q => 
                           reg_in_78_port, QN => n_1113);
   reg_in_regx77x : DFF_X1 port map( D => Plaintext(77), CK => clk, Q => 
                           reg_in_77_port, QN => n_1114);
   reg_in_regx76x : DFF_X1 port map( D => Plaintext(76), CK => clk, Q => 
                           reg_in_76_port, QN => n_1115);
   reg_in_regx75x : DFF_X1 port map( D => Plaintext(75), CK => clk, Q => 
                           reg_in_75_port, QN => n_1116);
   reg_in_regx74x : DFF_X1 port map( D => Plaintext(74), CK => clk, Q => 
                           reg_in_74_port, QN => n_1117);
   reg_in_regx73x : DFF_X1 port map( D => Plaintext(73), CK => clk, Q => 
                           reg_in_73_port, QN => n_1118);
   reg_in_regx72x : DFF_X1 port map( D => Plaintext(72), CK => clk, Q => 
                           reg_in_72_port, QN => n_1119);
   reg_in_regx71x : DFF_X1 port map( D => Plaintext(71), CK => clk, Q => 
                           reg_in_71_port, QN => n_1120);
   reg_in_regx70x : DFF_X1 port map( D => Plaintext(70), CK => clk, Q => 
                           reg_in_70_port, QN => n_1121);
   reg_in_regx69x : DFF_X1 port map( D => Plaintext(69), CK => clk, Q => 
                           reg_in_69_port, QN => n_1122);
   reg_in_regx68x : DFF_X1 port map( D => Plaintext(68), CK => clk, Q => 
                           reg_in_68_port, QN => n_1123);
   reg_in_regx67x : DFF_X1 port map( D => Plaintext(67), CK => clk, Q => 
                           reg_in_67_port, QN => n_1124);
   reg_in_regx66x : DFF_X1 port map( D => Plaintext(66), CK => clk, Q => 
                           reg_in_66_port, QN => n_1125);
   reg_in_regx65x : DFF_X1 port map( D => Plaintext(65), CK => clk, Q => 
                           reg_in_65_port, QN => n_1126);
   reg_in_regx64x : DFF_X1 port map( D => Plaintext(64), CK => clk, Q => 
                           reg_in_64_port, QN => n_1127);
   reg_in_regx63x : DFF_X1 port map( D => Plaintext(63), CK => clk, Q => 
                           reg_in_63_port, QN => n_1128);
   reg_in_regx62x : DFF_X1 port map( D => Plaintext(62), CK => clk, Q => 
                           reg_in_62_port, QN => n_1129);
   reg_in_regx61x : DFF_X1 port map( D => Plaintext(61), CK => clk, Q => 
                           reg_in_61_port, QN => n_1130);
   reg_in_regx60x : DFF_X1 port map( D => Plaintext(60), CK => clk, Q => 
                           reg_in_60_port, QN => n_1131);
   reg_in_regx59x : DFF_X1 port map( D => Plaintext(59), CK => clk, Q => 
                           reg_in_59_port, QN => n_1132);
   reg_in_regx58x : DFF_X1 port map( D => Plaintext(58), CK => clk, Q => 
                           reg_in_58_port, QN => n_1133);
   reg_in_regx57x : DFF_X1 port map( D => Plaintext(57), CK => clk, Q => 
                           reg_in_57_port, QN => n_1134);
   reg_in_regx56x : DFF_X1 port map( D => Plaintext(56), CK => clk, Q => 
                           reg_in_56_port, QN => n_1135);
   reg_in_regx55x : DFF_X1 port map( D => Plaintext(55), CK => clk, Q => 
                           reg_in_55_port, QN => n_1136);
   reg_in_regx54x : DFF_X1 port map( D => Plaintext(54), CK => clk, Q => 
                           reg_in_54_port, QN => n_1137);
   reg_in_regx53x : DFF_X1 port map( D => Plaintext(53), CK => clk, Q => 
                           reg_in_53_port, QN => n_1138);
   reg_in_regx52x : DFF_X1 port map( D => Plaintext(52), CK => clk, Q => 
                           reg_in_52_port, QN => n_1139);
   reg_in_regx51x : DFF_X1 port map( D => Plaintext(51), CK => clk, Q => 
                           reg_in_51_port, QN => n_1140);
   reg_in_regx50x : DFF_X1 port map( D => Plaintext(50), CK => clk, Q => 
                           reg_in_50_port, QN => n_1141);
   reg_in_regx49x : DFF_X1 port map( D => Plaintext(49), CK => clk, Q => 
                           reg_in_49_port, QN => n_1142);
   reg_in_regx48x : DFF_X1 port map( D => Plaintext(48), CK => clk, Q => 
                           reg_in_48_port, QN => n_1143);
   reg_in_regx47x : DFF_X1 port map( D => Plaintext(47), CK => clk, Q => 
                           reg_in_47_port, QN => n_1144);
   reg_in_regx46x : DFF_X1 port map( D => Plaintext(46), CK => clk, Q => 
                           reg_in_46_port, QN => n_1145);
   reg_in_regx45x : DFF_X1 port map( D => Plaintext(45), CK => clk, Q => 
                           reg_in_45_port, QN => n_1146);
   reg_in_regx44x : DFF_X1 port map( D => Plaintext(44), CK => clk, Q => 
                           reg_in_44_port, QN => n_1147);
   reg_in_regx43x : DFF_X1 port map( D => Plaintext(43), CK => clk, Q => 
                           reg_in_43_port, QN => n_1148);
   reg_in_regx42x : DFF_X1 port map( D => Plaintext(42), CK => clk, Q => 
                           reg_in_42_port, QN => n_1149);
   reg_in_regx41x : DFF_X1 port map( D => Plaintext(41), CK => clk, Q => 
                           reg_in_41_port, QN => n_1150);
   reg_in_regx40x : DFF_X1 port map( D => Plaintext(40), CK => clk, Q => 
                           reg_in_40_port, QN => n_1151);
   reg_in_regx39x : DFF_X1 port map( D => Plaintext(39), CK => clk, Q => 
                           reg_in_39_port, QN => n_1152);
   reg_in_regx38x : DFF_X1 port map( D => Plaintext(38), CK => clk, Q => 
                           reg_in_38_port, QN => n_1153);
   reg_in_regx37x : DFF_X1 port map( D => Plaintext(37), CK => clk, Q => 
                           reg_in_37_port, QN => n_1154);
   reg_in_regx36x : DFF_X1 port map( D => Plaintext(36), CK => clk, Q => 
                           reg_in_36_port, QN => n_1155);
   reg_in_regx35x : DFF_X1 port map( D => Plaintext(35), CK => clk, Q => 
                           reg_in_35_port, QN => n_1156);
   reg_in_regx34x : DFF_X1 port map( D => Plaintext(34), CK => clk, Q => 
                           reg_in_34_port, QN => n_1157);
   reg_in_regx33x : DFF_X1 port map( D => Plaintext(33), CK => clk, Q => 
                           reg_in_33_port, QN => n_1158);
   reg_in_regx32x : DFF_X1 port map( D => Plaintext(32), CK => clk, Q => 
                           reg_in_32_port, QN => n_1159);
   reg_in_regx31x : DFF_X1 port map( D => Plaintext(31), CK => clk, Q => 
                           reg_in_31_port, QN => n_1160);
   reg_in_regx30x : DFF_X1 port map( D => Plaintext(30), CK => clk, Q => 
                           reg_in_30_port, QN => n_1161);
   reg_in_regx29x : DFF_X1 port map( D => Plaintext(29), CK => clk, Q => 
                           reg_in_29_port, QN => n_1162);
   reg_in_regx28x : DFF_X1 port map( D => Plaintext(28), CK => clk, Q => 
                           reg_in_28_port, QN => n_1163);
   reg_in_regx27x : DFF_X1 port map( D => Plaintext(27), CK => clk, Q => 
                           reg_in_27_port, QN => n_1164);
   reg_in_regx26x : DFF_X1 port map( D => Plaintext(26), CK => clk, Q => 
                           reg_in_26_port, QN => n_1165);
   reg_in_regx25x : DFF_X1 port map( D => Plaintext(25), CK => clk, Q => 
                           reg_in_25_port, QN => n_1166);
   reg_in_regx24x : DFF_X1 port map( D => Plaintext(24), CK => clk, Q => 
                           reg_in_24_port, QN => n_1167);
   reg_in_regx23x : DFF_X1 port map( D => Plaintext(23), CK => clk, Q => 
                           reg_in_23_port, QN => n_1168);
   reg_in_regx22x : DFF_X1 port map( D => Plaintext(22), CK => clk, Q => 
                           reg_in_22_port, QN => n_1169);
   reg_in_regx21x : DFF_X1 port map( D => Plaintext(21), CK => clk, Q => 
                           reg_in_21_port, QN => n_1170);
   reg_in_regx20x : DFF_X1 port map( D => Plaintext(20), CK => clk, Q => 
                           reg_in_20_port, QN => n_1171);
   reg_in_regx19x : DFF_X1 port map( D => Plaintext(19), CK => clk, Q => 
                           reg_in_19_port, QN => n_1172);
   reg_in_regx18x : DFF_X1 port map( D => Plaintext(18), CK => clk, Q => 
                           reg_in_18_port, QN => n_1173);
   reg_in_regx17x : DFF_X1 port map( D => Plaintext(17), CK => clk, Q => 
                           reg_in_17_port, QN => n_1174);
   reg_in_regx16x : DFF_X1 port map( D => Plaintext(16), CK => clk, Q => 
                           reg_in_16_port, QN => n_1175);
   reg_in_regx15x : DFF_X1 port map( D => Plaintext(15), CK => clk, Q => 
                           reg_in_15_port, QN => n_1176);
   reg_in_regx14x : DFF_X1 port map( D => Plaintext(14), CK => clk, Q => 
                           reg_in_14_port, QN => n_1177);
   reg_in_regx13x : DFF_X1 port map( D => Plaintext(13), CK => clk, Q => 
                           reg_in_13_port, QN => n_1178);
   reg_in_regx12x : DFF_X1 port map( D => Plaintext(12), CK => clk, Q => 
                           reg_in_12_port, QN => n_1179);
   reg_in_regx11x : DFF_X1 port map( D => Plaintext(11), CK => clk, Q => 
                           reg_in_11_port, QN => n_1180);
   reg_in_regx10x : DFF_X1 port map( D => Plaintext(10), CK => clk, Q => 
                           reg_in_10_port, QN => n_1181);
   reg_in_regx9x : DFF_X1 port map( D => Plaintext(9), CK => clk, Q => 
                           reg_in_9_port, QN => n_1182);
   reg_in_regx8x : DFF_X1 port map( D => Plaintext(8), CK => clk, Q => 
                           reg_in_8_port, QN => n_1183);
   reg_in_regx7x : DFF_X1 port map( D => Plaintext(7), CK => clk, Q => 
                           reg_in_7_port, QN => n_1184);
   reg_in_regx6x : DFF_X1 port map( D => Plaintext(6), CK => clk, Q => 
                           reg_in_6_port, QN => n_1185);
   reg_in_regx5x : DFF_X1 port map( D => Plaintext(5), CK => clk, Q => 
                           reg_in_5_port, QN => n_1186);
   reg_in_regx4x : DFF_X1 port map( D => Plaintext(4), CK => clk, Q => 
                           reg_in_4_port, QN => n_1187);
   reg_in_regx3x : DFF_X1 port map( D => Plaintext(3), CK => clk, Q => 
                           reg_in_3_port, QN => n_1188);
   reg_in_regx2x : DFF_X1 port map( D => Plaintext(2), CK => clk, Q => 
                           reg_in_2_port, QN => n_1189);
   reg_in_regx1x : DFF_X1 port map( D => Plaintext(1), CK => clk, Q => 
                           reg_in_1_port, QN => n_1190);
   reg_in_regx0x : DFF_X1 port map( D => Plaintext(0), CK => clk, Q => 
                           reg_in_0_port, QN => n_1191);
   reg_key_regx190x : DFF_X1 port map( D => Key(190), CK => clk, Q => 
                           reg_key_190_port, QN => n_1192);
   reg_key_regx187x : DFF_X1 port map( D => Key(187), CK => clk, Q => 
                           reg_key_187_port, QN => n_1193);
   reg_key_regx179x : DFF_X1 port map( D => Key(179), CK => clk, Q => 
                           reg_key_179_port, QN => n_1194);
   reg_key_regx173x : DFF_X1 port map( D => Key(173), CK => clk, Q => 
                           reg_key_173_port, QN => n_1195);
   reg_key_regx168x : DFF_X1 port map( D => Key(168), CK => clk, Q => 
                           reg_key_168_port, QN => n_1196);
   reg_key_regx151x : DFF_X1 port map( D => Key(151), CK => clk, Q => 
                           reg_key_151_port, QN => n_1197);
   reg_key_regx148x : DFF_X1 port map( D => Key(148), CK => clk, Q => 
                           reg_key_148_port, QN => n_1198);
   reg_key_regx122x : DFF_X1 port map( D => Key(122), CK => clk, Q => 
                           reg_key_122_port, QN => n_1199);
   reg_key_regx104x : DFF_X1 port map( D => Key(104), CK => clk, Q => 
                           reg_key_104_port, QN => n_1200);
   reg_key_regx91x : DFF_X1 port map( D => Key(91), CK => clk, Q => 
                           reg_key_91_port, QN => n_1201);
   reg_key_regx83x : DFF_X1 port map( D => Key(83), CK => clk, Q => 
                           reg_key_83_port, QN => n_1202);
   reg_key_regx79x : DFF_X1 port map( D => Key(79), CK => clk, Q => 
                           reg_key_79_port, QN => n_1203);
   reg_key_regx74x : DFF_X1 port map( D => Key(74), CK => clk, Q => 
                           reg_key_74_port, QN => n_1204);
   reg_key_regx68x : DFF_X1 port map( D => Key(68), CK => clk, Q => 
                           reg_key_68_port, QN => n_1205);
   reg_key_regx66x : DFF_X1 port map( D => Key(66), CK => clk, Q => 
                           reg_key_66_port, QN => n_1206);
   reg_key_regx56x : DFF_X1 port map( D => Key(56), CK => clk, Q => 
                           reg_key_56_port, QN => n_1207);
   reg_key_regx53x : DFF_X1 port map( D => Key(53), CK => clk, Q => 
                           reg_key_53_port, QN => n_1208);
   reg_key_regx51x : DFF_X1 port map( D => Key(51), CK => clk, Q => 
                           reg_key_51_port, QN => n_1209);
   reg_key_regx40x : DFF_X1 port map( D => Key(40), CK => clk, Q => 
                           reg_key_40_port, QN => n_1210);
   reg_key_regx35x : DFF_X1 port map( D => Key(35), CK => clk, Q => 
                           reg_key_35_port, QN => n_1211);
   reg_key_regx19x : DFF_X1 port map( D => Key(19), CK => clk, Q => 
                           reg_key_19_port, QN => n_1212);
   reg_key_regx11x : DFF_X1 port map( D => Key(11), CK => clk, Q => 
                           reg_key_11_port, QN => n_1213);
   reg_key_regx9x : DFF_X1 port map( D => Key(9), CK => clk, Q => 
                           reg_key_9_port, QN => n_1214);
   reg_key_regx8x : DFF_X1 port map( D => Key(8), CK => clk, Q => 
                           reg_key_8_port, QN => n_1215);
   Ciphertext_regx191x : DFF_X1 port map( D => reg_out_191_port, CK => clk, Q 
                           => Ciphertext(191), QN => n_1216);
   Ciphertext_regx190x : DFF_X1 port map( D => reg_out_190_port, CK => clk, Q 
                           => Ciphertext(190), QN => n_1217);
   Ciphertext_regx189x : DFF_X1 port map( D => reg_out_189_port, CK => clk, Q 
                           => Ciphertext(189), QN => n_1218);
   Ciphertext_regx187x : DFF_X1 port map( D => reg_out_187_port, CK => clk, Q 
                           => Ciphertext(187), QN => n_1219);
   Ciphertext_regx186x : DFF_X1 port map( D => reg_out_186_port, CK => clk, Q 
                           => Ciphertext(186), QN => n_1220);
   Ciphertext_regx185x : DFF_X1 port map( D => reg_out_185_port, CK => clk, Q 
                           => Ciphertext(185), QN => n_1221);
   Ciphertext_regx184x : DFF_X1 port map( D => reg_out_184_port, CK => clk, Q 
                           => Ciphertext(184), QN => n_1222);
   Ciphertext_regx183x : DFF_X1 port map( D => reg_out_183_port, CK => clk, Q 
                           => Ciphertext(183), QN => n_1223);
   Ciphertext_regx182x : DFF_X1 port map( D => reg_out_182_port, CK => clk, Q 
                           => Ciphertext(182), QN => n_1224);
   Ciphertext_regx181x : DFF_X1 port map( D => reg_out_181_port, CK => clk, Q 
                           => Ciphertext(181), QN => n_1225);
   Ciphertext_regx180x : DFF_X1 port map( D => reg_out_180_port, CK => clk, Q 
                           => Ciphertext(180), QN => n_1226);
   Ciphertext_regx179x : DFF_X1 port map( D => reg_out_179_port, CK => clk, Q 
                           => Ciphertext(179), QN => n_1227);
   Ciphertext_regx178x : DFF_X1 port map( D => reg_out_178_port, CK => clk, Q 
                           => Ciphertext(178), QN => n_1228);
   Ciphertext_regx177x : DFF_X1 port map( D => reg_out_177_port, CK => clk, Q 
                           => Ciphertext(177), QN => n_1229);
   Ciphertext_regx176x : DFF_X1 port map( D => reg_out_176_port, CK => clk, Q 
                           => Ciphertext(176), QN => n_1230);
   Ciphertext_regx175x : DFF_X1 port map( D => reg_out_175_port, CK => clk, Q 
                           => Ciphertext(175), QN => n_1231);
   Ciphertext_regx174x : DFF_X1 port map( D => reg_out_174_port, CK => clk, Q 
                           => Ciphertext(174), QN => n_1232);
   Ciphertext_regx173x : DFF_X1 port map( D => reg_out_173_port, CK => clk, Q 
                           => Ciphertext(173), QN => n_1233);
   Ciphertext_regx172x : DFF_X1 port map( D => reg_out_172_port, CK => clk, Q 
                           => Ciphertext(172), QN => n_1234);
   Ciphertext_regx171x : DFF_X1 port map( D => reg_out_171_port, CK => clk, Q 
                           => Ciphertext(171), QN => n_1235);
   Ciphertext_regx170x : DFF_X1 port map( D => reg_out_170_port, CK => clk, Q 
                           => Ciphertext(170), QN => n_1236);
   Ciphertext_regx169x : DFF_X1 port map( D => reg_out_169_port, CK => clk, Q 
                           => Ciphertext(169), QN => n_1237);
   Ciphertext_regx167x : DFF_X1 port map( D => reg_out_167_port, CK => clk, Q 
                           => Ciphertext(167), QN => n_1238);
   Ciphertext_regx166x : DFF_X1 port map( D => reg_out_166_port, CK => clk, Q 
                           => Ciphertext(166), QN => n_1239);
   Ciphertext_regx165x : DFF_X1 port map( D => reg_out_165_port, CK => clk, Q 
                           => Ciphertext(165), QN => n_1240);
   Ciphertext_regx164x : DFF_X1 port map( D => reg_out_164_port, CK => clk, Q 
                           => Ciphertext(164), QN => n_1241);
   Ciphertext_regx163x : DFF_X1 port map( D => reg_out_163_port, CK => clk, Q 
                           => Ciphertext(163), QN => n_1242);
   Ciphertext_regx162x : DFF_X1 port map( D => reg_out_162_port, CK => clk, Q 
                           => Ciphertext(162), QN => n_1243);
   Ciphertext_regx161x : DFF_X1 port map( D => reg_out_161_port, CK => clk, Q 
                           => Ciphertext(161), QN => n_1244);
   Ciphertext_regx160x : DFF_X1 port map( D => reg_out_160_port, CK => clk, Q 
                           => Ciphertext(160), QN => n_1245);
   Ciphertext_regx159x : DFF_X1 port map( D => reg_out_159_port, CK => clk, Q 
                           => Ciphertext(159), QN => n_1246);
   Ciphertext_regx158x : DFF_X1 port map( D => reg_out_158_port, CK => clk, Q 
                           => Ciphertext(158), QN => n_1247);
   Ciphertext_regx157x : DFF_X1 port map( D => reg_out_157_port, CK => clk, Q 
                           => Ciphertext(157), QN => n_1248);
   Ciphertext_regx156x : DFF_X1 port map( D => reg_out_156_port, CK => clk, Q 
                           => Ciphertext(156), QN => n_1249);
   Ciphertext_regx155x : DFF_X1 port map( D => reg_out_155_port, CK => clk, Q 
                           => Ciphertext(155), QN => n_1250);
   Ciphertext_regx154x : DFF_X1 port map( D => reg_out_154_port, CK => clk, Q 
                           => Ciphertext(154), QN => n_1251);
   Ciphertext_regx153x : DFF_X1 port map( D => reg_out_153_port, CK => clk, Q 
                           => Ciphertext(153), QN => n_1252);
   Ciphertext_regx152x : DFF_X1 port map( D => reg_out_152_port, CK => clk, Q 
                           => Ciphertext(152), QN => n_1253);
   Ciphertext_regx150x : DFF_X1 port map( D => reg_out_150_port, CK => clk, Q 
                           => Ciphertext(150), QN => n_1254);
   Ciphertext_regx149x : DFF_X1 port map( D => reg_out_149_port, CK => clk, Q 
                           => Ciphertext(149), QN => n_1255);
   Ciphertext_regx147x : DFF_X1 port map( D => reg_out_147_port, CK => clk, Q 
                           => Ciphertext(147), QN => n_1256);
   Ciphertext_regx146x : DFF_X1 port map( D => reg_out_146_port, CK => clk, Q 
                           => Ciphertext(146), QN => n_1257);
   Ciphertext_regx145x : DFF_X1 port map( D => reg_out_145_port, CK => clk, Q 
                           => Ciphertext(145), QN => n_1258);
   Ciphertext_regx144x : DFF_X1 port map( D => reg_out_144_port, CK => clk, Q 
                           => Ciphertext(144), QN => n_1259);
   Ciphertext_regx143x : DFF_X1 port map( D => reg_out_143_port, CK => clk, Q 
                           => Ciphertext(143), QN => n_1260);
   Ciphertext_regx142x : DFF_X1 port map( D => reg_out_142_port, CK => clk, Q 
                           => Ciphertext(142), QN => n_1261);
   Ciphertext_regx141x : DFF_X1 port map( D => reg_out_141_port, CK => clk, Q 
                           => Ciphertext(141), QN => n_1262);
   Ciphertext_regx139x : DFF_X1 port map( D => reg_out_139_port, CK => clk, Q 
                           => Ciphertext(139), QN => n_1263);
   Ciphertext_regx138x : DFF_X1 port map( D => reg_out_138_port, CK => clk, Q 
                           => Ciphertext(138), QN => n_1264);
   Ciphertext_regx137x : DFF_X1 port map( D => reg_out_137_port, CK => clk, Q 
                           => Ciphertext(137), QN => n_1265);
   Ciphertext_regx136x : DFF_X1 port map( D => reg_out_136_port, CK => clk, Q 
                           => Ciphertext(136), QN => n_1266);
   Ciphertext_regx135x : DFF_X1 port map( D => reg_out_135_port, CK => clk, Q 
                           => Ciphertext(135), QN => n_1267);
   Ciphertext_regx134x : DFF_X1 port map( D => reg_out_134_port, CK => clk, Q 
                           => Ciphertext(134), QN => n_1268);
   Ciphertext_regx133x : DFF_X1 port map( D => reg_out_133_port, CK => clk, Q 
                           => Ciphertext(133), QN => n_1269);
   Ciphertext_regx132x : DFF_X1 port map( D => reg_out_132_port, CK => clk, Q 
                           => Ciphertext(132), QN => n_1270);
   Ciphertext_regx131x : DFF_X1 port map( D => reg_out_131_port, CK => clk, Q 
                           => Ciphertext(131), QN => n_1271);
   Ciphertext_regx130x : DFF_X1 port map( D => reg_out_130_port, CK => clk, Q 
                           => Ciphertext(130), QN => n_1272);
   Ciphertext_regx129x : DFF_X1 port map( D => reg_out_129_port, CK => clk, Q 
                           => Ciphertext(129), QN => n_1273);
   Ciphertext_regx128x : DFF_X1 port map( D => reg_out_128_port, CK => clk, Q 
                           => Ciphertext(128), QN => n_1274);
   Ciphertext_regx127x : DFF_X1 port map( D => reg_out_127_port, CK => clk, Q 
                           => Ciphertext(127), QN => n_1275);
   Ciphertext_regx126x : DFF_X1 port map( D => reg_out_126_port, CK => clk, Q 
                           => Ciphertext(126), QN => n_1276);
   Ciphertext_regx125x : DFF_X1 port map( D => reg_out_125_port, CK => clk, Q 
                           => Ciphertext(125), QN => n_1277);
   Ciphertext_regx124x : DFF_X1 port map( D => reg_out_124_port, CK => clk, Q 
                           => Ciphertext(124), QN => n_1278);
   Ciphertext_regx123x : DFF_X1 port map( D => reg_out_123_port, CK => clk, Q 
                           => Ciphertext(123), QN => n_1279);
   Ciphertext_regx122x : DFF_X1 port map( D => reg_out_122_port, CK => clk, Q 
                           => Ciphertext(122), QN => n_1280);
   Ciphertext_regx120x : DFF_X1 port map( D => reg_out_120_port, CK => clk, Q 
                           => Ciphertext(120), QN => n_1281);
   Ciphertext_regx119x : DFF_X1 port map( D => reg_out_119_port, CK => clk, Q 
                           => Ciphertext(119), QN => n_1282);
   Ciphertext_regx118x : DFF_X1 port map( D => reg_out_118_port, CK => clk, Q 
                           => Ciphertext(118), QN => n_1283);
   Ciphertext_regx117x : DFF_X1 port map( D => reg_out_117_port, CK => clk, Q 
                           => Ciphertext(117), QN => n_1284);
   Ciphertext_regx116x : DFF_X1 port map( D => reg_out_116_port, CK => clk, Q 
                           => Ciphertext(116), QN => n_1285);
   Ciphertext_regx115x : DFF_X1 port map( D => reg_out_115_port, CK => clk, Q 
                           => Ciphertext(115), QN => n_1286);
   Ciphertext_regx114x : DFF_X1 port map( D => reg_out_114_port, CK => clk, Q 
                           => Ciphertext(114), QN => n_1287);
   Ciphertext_regx113x : DFF_X1 port map( D => reg_out_113_port, CK => clk, Q 
                           => Ciphertext(113), QN => n_1288);
   Ciphertext_regx112x : DFF_X1 port map( D => reg_out_112_port, CK => clk, Q 
                           => Ciphertext(112), QN => n_1289);
   Ciphertext_regx110x : DFF_X1 port map( D => reg_out_110_port, CK => clk, Q 
                           => Ciphertext(110), QN => n_1290);
   Ciphertext_regx109x : DFF_X1 port map( D => reg_out_109_port, CK => clk, Q 
                           => Ciphertext(109), QN => n_1291);
   Ciphertext_regx107x : DFF_X1 port map( D => reg_out_107_port, CK => clk, Q 
                           => Ciphertext(107), QN => n_1292);
   Ciphertext_regx106x : DFF_X1 port map( D => reg_out_106_port, CK => clk, Q 
                           => Ciphertext(106), QN => n_1293);
   Ciphertext_regx104x : DFF_X1 port map( D => reg_out_104_port, CK => clk, Q 
                           => Ciphertext(104), QN => n_1294);
   Ciphertext_regx103x : DFF_X1 port map( D => reg_out_103_port, CK => clk, Q 
                           => Ciphertext(103), QN => n_1295);
   Ciphertext_regx101x : DFF_X1 port map( D => reg_out_101_port, CK => clk, Q 
                           => Ciphertext(101), QN => n_1296);
   Ciphertext_regx100x : DFF_X1 port map( D => reg_out_100_port, CK => clk, Q 
                           => Ciphertext(100), QN => n_1297);
   Ciphertext_regx99x : DFF_X1 port map( D => reg_out_99_port, CK => clk, Q => 
                           Ciphertext(99), QN => n_1298);
   Ciphertext_regx98x : DFF_X1 port map( D => reg_out_98_port, CK => clk, Q => 
                           Ciphertext(98), QN => n_1299);
   Ciphertext_regx97x : DFF_X1 port map( D => reg_out_97_port, CK => clk, Q => 
                           Ciphertext(97), QN => n_1300);
   Ciphertext_regx96x : DFF_X1 port map( D => reg_out_96_port, CK => clk, Q => 
                           Ciphertext(96), QN => n_1301);
   Ciphertext_regx95x : DFF_X1 port map( D => reg_out_95_port, CK => clk, Q => 
                           Ciphertext(95), QN => n_1302);
   Ciphertext_regx94x : DFF_X1 port map( D => reg_out_94_port, CK => clk, Q => 
                           Ciphertext(94), QN => n_1303);
   Ciphertext_regx93x : DFF_X1 port map( D => reg_out_93_port, CK => clk, Q => 
                           Ciphertext(93), QN => n_1304);
   Ciphertext_regx92x : DFF_X1 port map( D => reg_out_92_port, CK => clk, Q => 
                           Ciphertext(92), QN => n_1305);
   Ciphertext_regx91x : DFF_X1 port map( D => reg_out_91_port, CK => clk, Q => 
                           Ciphertext(91), QN => n_1306);
   Ciphertext_regx90x : DFF_X1 port map( D => reg_out_90_port, CK => clk, Q => 
                           Ciphertext(90), QN => n_1307);
   Ciphertext_regx89x : DFF_X1 port map( D => reg_out_89_port, CK => clk, Q => 
                           Ciphertext(89), QN => n_1308);
   Ciphertext_regx88x : DFF_X1 port map( D => reg_out_88_port, CK => clk, Q => 
                           Ciphertext(88), QN => n_1309);
   Ciphertext_regx87x : DFF_X1 port map( D => reg_out_87_port, CK => clk, Q => 
                           Ciphertext(87), QN => n_1310);
   Ciphertext_regx86x : DFF_X1 port map( D => reg_out_86_port, CK => clk, Q => 
                           Ciphertext(86), QN => n_1311);
   Ciphertext_regx85x : DFF_X1 port map( D => reg_out_85_port, CK => clk, Q => 
                           Ciphertext(85), QN => n_1312);
   Ciphertext_regx83x : DFF_X1 port map( D => reg_out_83_port, CK => clk, Q => 
                           Ciphertext(83), QN => n_1313);
   Ciphertext_regx82x : DFF_X1 port map( D => reg_out_82_port, CK => clk, Q => 
                           Ciphertext(82), QN => n_1314);
   Ciphertext_regx81x : DFF_X1 port map( D => reg_out_81_port, CK => clk, Q => 
                           Ciphertext(81), QN => n_1315);
   Ciphertext_regx80x : DFF_X1 port map( D => reg_out_80_port, CK => clk, Q => 
                           Ciphertext(80), QN => n_1316);
   Ciphertext_regx79x : DFF_X1 port map( D => reg_out_79_port, CK => clk, Q => 
                           Ciphertext(79), QN => n_1317);
   Ciphertext_regx78x : DFF_X1 port map( D => reg_out_78_port, CK => clk, Q => 
                           Ciphertext(78), QN => n_1318);
   Ciphertext_regx77x : DFF_X1 port map( D => reg_out_77_port, CK => clk, Q => 
                           Ciphertext(77), QN => n_1319);
   Ciphertext_regx76x : DFF_X1 port map( D => reg_out_76_port, CK => clk, Q => 
                           Ciphertext(76), QN => n_1320);
   Ciphertext_regx75x : DFF_X1 port map( D => reg_out_75_port, CK => clk, Q => 
                           Ciphertext(75), QN => n_1321);
   Ciphertext_regx74x : DFF_X1 port map( D => reg_out_74_port, CK => clk, Q => 
                           Ciphertext(74), QN => n_1322);
   Ciphertext_regx72x : DFF_X1 port map( D => reg_out_72_port, CK => clk, Q => 
                           Ciphertext(72), QN => n_1323);
   Ciphertext_regx71x : DFF_X1 port map( D => reg_out_71_port, CK => clk, Q => 
                           Ciphertext(71), QN => n_1324);
   Ciphertext_regx70x : DFF_X1 port map( D => reg_out_70_port, CK => clk, Q => 
                           Ciphertext(70), QN => n_1325);
   Ciphertext_regx69x : DFF_X1 port map( D => reg_out_69_port, CK => clk, Q => 
                           Ciphertext(69), QN => n_1326);
   Ciphertext_regx68x : DFF_X1 port map( D => reg_out_68_port, CK => clk, Q => 
                           Ciphertext(68), QN => n_1327);
   Ciphertext_regx67x : DFF_X1 port map( D => reg_out_67_port, CK => clk, Q => 
                           Ciphertext(67), QN => n_1328);
   Ciphertext_regx66x : DFF_X1 port map( D => reg_out_66_port, CK => clk, Q => 
                           Ciphertext(66), QN => n_1329);
   Ciphertext_regx65x : DFF_X1 port map( D => reg_out_65_port, CK => clk, Q => 
                           Ciphertext(65), QN => n_1330);
   Ciphertext_regx64x : DFF_X1 port map( D => reg_out_64_port, CK => clk, Q => 
                           Ciphertext(64), QN => n_1331);
   Ciphertext_regx63x : DFF_X1 port map( D => reg_out_63_port, CK => clk, Q => 
                           Ciphertext(63), QN => n_1332);
   Ciphertext_regx62x : DFF_X1 port map( D => reg_out_62_port, CK => clk, Q => 
                           Ciphertext(62), QN => n_1333);
   Ciphertext_regx61x : DFF_X1 port map( D => reg_out_61_port, CK => clk, Q => 
                           Ciphertext(61), QN => n_1334);
   Ciphertext_regx60x : DFF_X1 port map( D => reg_out_60_port, CK => clk, Q => 
                           Ciphertext(60), QN => n_1335);
   Ciphertext_regx59x : DFF_X1 port map( D => reg_out_59_port, CK => clk, Q => 
                           Ciphertext(59), QN => n_1336);
   Ciphertext_regx58x : DFF_X1 port map( D => reg_out_58_port, CK => clk, Q => 
                           Ciphertext(58), QN => n_1337);
   Ciphertext_regx57x : DFF_X1 port map( D => reg_out_57_port, CK => clk, Q => 
                           Ciphertext(57), QN => n_1338);
   Ciphertext_regx56x : DFF_X1 port map( D => reg_out_56_port, CK => clk, Q => 
                           Ciphertext(56), QN => n_1339);
   Ciphertext_regx55x : DFF_X1 port map( D => reg_out_55_port, CK => clk, Q => 
                           Ciphertext(55), QN => n_1340);
   Ciphertext_regx54x : DFF_X1 port map( D => reg_out_54_port, CK => clk, Q => 
                           Ciphertext(54), QN => n_1341);
   Ciphertext_regx53x : DFF_X1 port map( D => reg_out_53_port, CK => clk, Q => 
                           Ciphertext(53), QN => n_1342);
   Ciphertext_regx52x : DFF_X1 port map( D => reg_out_52_port, CK => clk, Q => 
                           Ciphertext(52), QN => n_1343);
   Ciphertext_regx49x : DFF_X1 port map( D => reg_out_49_port, CK => clk, Q => 
                           Ciphertext(49), QN => n_1344);
   Ciphertext_regx48x : DFF_X1 port map( D => reg_out_48_port, CK => clk, Q => 
                           Ciphertext(48), QN => n_1345);
   Ciphertext_regx47x : DFF_X1 port map( D => reg_out_47_port, CK => clk, Q => 
                           Ciphertext(47), QN => n_1346);
   Ciphertext_regx46x : DFF_X1 port map( D => reg_out_46_port, CK => clk, Q => 
                           Ciphertext(46), QN => n_1347);
   Ciphertext_regx45x : DFF_X1 port map( D => reg_out_45_port, CK => clk, Q => 
                           Ciphertext(45), QN => n_1348);
   Ciphertext_regx43x : DFF_X1 port map( D => reg_out_43_port, CK => clk, Q => 
                           Ciphertext(43), QN => n_1349);
   Ciphertext_regx42x : DFF_X1 port map( D => reg_out_42_port, CK => clk, Q => 
                           Ciphertext(42), QN => n_1350);
   Ciphertext_regx41x : DFF_X1 port map( D => reg_out_41_port, CK => clk, Q => 
                           Ciphertext(41), QN => n_1351);
   Ciphertext_regx39x : DFF_X1 port map( D => reg_out_39_port, CK => clk, Q => 
                           Ciphertext(39), QN => n_1352);
   Ciphertext_regx38x : DFF_X1 port map( D => reg_out_38_port, CK => clk, Q => 
                           Ciphertext(38), QN => n_1353);
   Ciphertext_regx37x : DFF_X1 port map( D => reg_out_37_port, CK => clk, Q => 
                           Ciphertext(37), QN => n_1354);
   Ciphertext_regx36x : DFF_X1 port map( D => reg_out_36_port, CK => clk, Q => 
                           Ciphertext(36), QN => n_1355);
   Ciphertext_regx35x : DFF_X1 port map( D => reg_out_35_port, CK => clk, Q => 
                           Ciphertext(35), QN => n_1356);
   Ciphertext_regx34x : DFF_X1 port map( D => reg_out_34_port, CK => clk, Q => 
                           Ciphertext(34), QN => n_1357);
   Ciphertext_regx33x : DFF_X1 port map( D => reg_out_33_port, CK => clk, Q => 
                           Ciphertext(33), QN => n_1358);
   Ciphertext_regx32x : DFF_X1 port map( D => reg_out_32_port, CK => clk, Q => 
                           Ciphertext(32), QN => n_1359);
   Ciphertext_regx31x : DFF_X1 port map( D => reg_out_31_port, CK => clk, Q => 
                           Ciphertext(31), QN => n_1360);
   Ciphertext_regx30x : DFF_X1 port map( D => reg_out_30_port, CK => clk, Q => 
                           Ciphertext(30), QN => n_1361);
   Ciphertext_regx29x : DFF_X1 port map( D => reg_out_29_port, CK => clk, Q => 
                           Ciphertext(29), QN => n_1362);
   Ciphertext_regx27x : DFF_X1 port map( D => reg_out_27_port, CK => clk, Q => 
                           Ciphertext(27), QN => n_1363);
   Ciphertext_regx26x : DFF_X1 port map( D => reg_out_26_port, CK => clk, Q => 
                           Ciphertext(26), QN => n_1364);
   Ciphertext_regx25x : DFF_X1 port map( D => reg_out_25_port, CK => clk, Q => 
                           Ciphertext(25), QN => n_1365);
   Ciphertext_regx24x : DFF_X1 port map( D => reg_out_24_port, CK => clk, Q => 
                           Ciphertext(24), QN => n_1366);
   Ciphertext_regx23x : DFF_X1 port map( D => reg_out_23_port, CK => clk, Q => 
                           Ciphertext(23), QN => n_1367);
   Ciphertext_regx22x : DFF_X1 port map( D => reg_out_22_port, CK => clk, Q => 
                           Ciphertext(22), QN => n_1368);
   Ciphertext_regx21x : DFF_X1 port map( D => reg_out_21_port, CK => clk, Q => 
                           Ciphertext(21), QN => n_1369);
   Ciphertext_regx20x : DFF_X1 port map( D => reg_out_20_port, CK => clk, Q => 
                           Ciphertext(20), QN => n_1370);
   Ciphertext_regx19x : DFF_X1 port map( D => reg_out_19_port, CK => clk, Q => 
                           Ciphertext(19), QN => n_1371);
   Ciphertext_regx18x : DFF_X1 port map( D => reg_out_18_port, CK => clk, Q => 
                           Ciphertext(18), QN => n_1372);
   Ciphertext_regx17x : DFF_X1 port map( D => reg_out_17_port, CK => clk, Q => 
                           Ciphertext(17), QN => n_1373);
   Ciphertext_regx16x : DFF_X1 port map( D => reg_out_16_port, CK => clk, Q => 
                           Ciphertext(16), QN => n_1374);
   Ciphertext_regx15x : DFF_X1 port map( D => reg_out_15_port, CK => clk, Q => 
                           Ciphertext(15), QN => n_1375);
   Ciphertext_regx14x : DFF_X1 port map( D => reg_out_14_port, CK => clk, Q => 
                           Ciphertext(14), QN => n_1376);
   Ciphertext_regx13x : DFF_X1 port map( D => reg_out_13_port, CK => clk, Q => 
                           Ciphertext(13), QN => n_1377);
   Ciphertext_regx12x : DFF_X1 port map( D => reg_out_12_port, CK => clk, Q => 
                           Ciphertext(12), QN => n_1378);
   Ciphertext_regx11x : DFF_X1 port map( D => reg_out_11_port, CK => clk, Q => 
                           Ciphertext(11), QN => n_1379);
   Ciphertext_regx10x : DFF_X1 port map( D => reg_out_10_port, CK => clk, Q => 
                           Ciphertext(10), QN => n_1380);
   Ciphertext_regx9x : DFF_X1 port map( D => reg_out_9_port, CK => clk, Q => 
                           Ciphertext(9), QN => n_1381);
   Ciphertext_regx8x : DFF_X1 port map( D => reg_out_8_port, CK => clk, Q => 
                           Ciphertext(8), QN => n_1382);
   Ciphertext_regx7x : DFF_X1 port map( D => reg_out_7_port, CK => clk, Q => 
                           Ciphertext(7), QN => n_1383);
   Ciphertext_regx6x : DFF_X1 port map( D => reg_out_6_port, CK => clk, Q => 
                           Ciphertext(6), QN => n_1384);
   Ciphertext_regx5x : DFF_X1 port map( D => reg_out_5_port, CK => clk, Q => 
                           Ciphertext(5), QN => n_1385);
   Ciphertext_regx4x : DFF_X1 port map( D => reg_out_4_port, CK => clk, Q => 
                           Ciphertext(4), QN => n_1386);
   Ciphertext_regx3x : DFF_X1 port map( D => reg_out_3_port, CK => clk, Q => 
                           Ciphertext(3), QN => n_1387);
   Ciphertext_regx2x : DFF_X1 port map( D => reg_out_2_port, CK => clk, Q => 
                           Ciphertext(2), QN => n_1388);
   Ciphertext_regx1x : DFF_X1 port map( D => reg_out_1_port, CK => clk, Q => 
                           Ciphertext(1), QN => n_1389);
   Ciphertext_regx40x : DFF_X1 port map( D => reg_out_40_port, CK => clk, Q => 
                           Ciphertext(40), QN => n_1390);
   reg_key_regx49x : DFF_X1 port map( D => Key(49), CK => clk, Q => 
                           reg_key_49_port, QN => n_1391);
   reg_key_regx147x : DFF_X1 port map( D => Key(147), CK => clk, Q => 
                           reg_key_147_port, QN => n_1392);
   Ciphertext_regx151x : DFF_X1 port map( D => reg_out_151_port, CK => clk, Q 
                           => Ciphertext(151), QN => n_1393);
   reg_key_regx1x : DFF_X1 port map( D => Key(1), CK => clk, Q => 
                           reg_key_1_port, QN => n_1394);
   reg_key_regx176x : DFF_X1 port map( D => Key(176), CK => clk, Q => 
                           reg_key_176_port, QN => n_1395);
   reg_key_regx159x : DFF_X1 port map( D => Key(159), CK => clk, Q => 
                           reg_key_159_port, QN => n_1396);
   reg_key_regx155x : DFF_X1 port map( D => Key(155), CK => clk, Q => 
                           reg_key_155_port, QN => n_1397);
   Ciphertext_regx51x : DFF_X1 port map( D => reg_out_51_port, CK => clk, Q => 
                           Ciphertext(51), QN => n_1398);
   reg_key_regx119x : DFF_X1 port map( D => Key(119), CK => clk, Q => 
                           reg_key_119_port, QN => n_1399);
   reg_key_regx44x : DFF_X1 port map( D => Key(44), CK => clk, Q => 
                           reg_key_44_port, QN => n_1400);
   reg_key_regx116x : DFF_X1 port map( D => Key(116), CK => clk, Q => 
                           reg_key_116_port, QN => n_1401);
   reg_key_regx137x : DFF_X1 port map( D => Key(137), CK => clk, Q => 
                           reg_key_137_port, QN => n_1402);
   reg_key_regx167x : DFF_X1 port map( D => Key(167), CK => clk, Q => 
                           reg_key_167_port, QN => n_1403);
   reg_key_regx50x : DFF_X1 port map( D => Key(50), CK => clk, Q => 
                           reg_key_50_port, QN => n_1404);
   reg_key_regx129x : DFF_X1 port map( D => Key(129), CK => clk, Q => 
                           reg_key_129_port, QN => n_1405);
   reg_key_regx111x : DFF_X1 port map( D => Key(111), CK => clk, Q => 
                           reg_key_111_port, QN => n_1406);
   reg_key_regx20x : DFF_X1 port map( D => Key(20), CK => clk, Q => 
                           reg_key_20_port, QN => n_1407);
   reg_key_regx33x : DFF_X1 port map( D => Key(33), CK => clk, Q => 
                           reg_key_33_port, QN => n_1408);
   reg_key_regx178x : DFF_X1 port map( D => Key(178), CK => clk, Q => 
                           reg_key_178_port, QN => n_1409);
   reg_key_regx135x : DFF_X1 port map( D => Key(135), CK => clk, Q => 
                           reg_key_135_port, QN => n_1410);
   reg_key_regx2x : DFF_X1 port map( D => Key(2), CK => clk, Q => 
                           reg_key_2_port, QN => n_1411);
   reg_key_regx77x : DFF_X1 port map( D => Key(77), CK => clk, Q => 
                           reg_key_77_port, QN => n_1412);
   reg_key_regx101x : DFF_X1 port map( D => Key(101), CK => clk, Q => 
                           reg_key_101_port, QN => n_1413);
   reg_key_regx125x : DFF_X1 port map( D => Key(125), CK => clk, Q => 
                           reg_key_125_port, QN => n_1414);
   reg_key_regx191x : DFF_X1 port map( D => Key(191), CK => clk, Q => 
                           reg_key_191_port, QN => n_1415);
   reg_key_regx175x : DFF_X1 port map( D => Key(175), CK => clk, Q => 
                           reg_key_175_port, QN => n_1416);
   reg_key_regx3x : DFF_X1 port map( D => Key(3), CK => clk, Q => 
                           reg_key_3_port, QN => n_1417);
   reg_key_regx153x : DFF_X1 port map( D => Key(153), CK => clk, Q => 
                           reg_key_153_port, QN => n_1418);
   reg_key_regx32x : DFF_X1 port map( D => Key(32), CK => clk, Q => 
                           reg_key_32_port, QN => n_1419);
   reg_key_regx112x : DFF_X1 port map( D => Key(112), CK => clk, Q => 
                           reg_key_112_port, QN => n_1420);
   reg_key_regx80x : DFF_X1 port map( D => Key(80), CK => clk, Q => 
                           reg_key_80_port, QN => n_1421);
   reg_key_regx150x : DFF_X1 port map( D => Key(150), CK => clk, Q => 
                           reg_key_150_port, QN => n_1422);
   reg_key_regx107x : DFF_X1 port map( D => Key(107), CK => clk, Q => 
                           reg_key_107_port, QN => n_1423);
   reg_key_regx98x : DFF_X1 port map( D => Key(98), CK => clk, Q => 
                           reg_key_98_port, QN => n_1424);
   reg_key_regx87x : DFF_X1 port map( D => Key(87), CK => clk, Q => 
                           reg_key_87_port, QN => n_1425);
   reg_key_regx189x : DFF_X1 port map( D => Key(189), CK => clk, Q => 
                           reg_key_189_port, QN => n_1426);
   reg_key_regx174x : DFF_X1 port map( D => Key(174), CK => clk, Q => 
                           reg_key_174_port, QN => n_1427);
   reg_key_regx28x : DFF_X1 port map( D => Key(28), CK => clk, Q => 
                           reg_key_28_port, QN => n_1428);
   reg_key_regx26x : DFF_X1 port map( D => Key(26), CK => clk, Q => 
                           reg_key_26_port, QN => n_1429);
   reg_key_regx134x : DFF_X1 port map( D => Key(134), CK => clk, Q => 
                           reg_key_134_port, QN => n_1430);
   reg_key_regx70x : DFF_X1 port map( D => Key(70), CK => clk, Q => 
                           reg_key_70_port, QN => n_1431);
   reg_key_regx177x : DFF_X1 port map( D => Key(177), CK => clk, Q => 
                           reg_key_177_port, QN => n_1432);
   reg_key_regx82x : DFF_X1 port map( D => Key(82), CK => clk, Q => 
                           reg_key_82_port, QN => n_1433);
   reg_key_regx92x : DFF_X1 port map( D => Key(92), CK => clk, Q => 
                           reg_key_92_port, QN => n_1434);
   reg_key_regx140x : DFF_X1 port map( D => Key(140), CK => clk, Q => 
                           reg_key_140_port, QN => n_1435);
   reg_key_regx57x : DFF_X1 port map( D => Key(57), CK => clk, Q => 
                           reg_key_57_port, QN => n_1436);
   reg_key_regx183x : DFF_X1 port map( D => Key(183), CK => clk, Q => 
                           reg_key_183_port, QN => n_1437);
   reg_key_regx171x : DFF_X1 port map( D => Key(171), CK => clk, Q => 
                           reg_key_171_port, QN => n_1438);
   reg_key_regx152x : DFF_X1 port map( D => Key(152), CK => clk, Q => 
                           reg_key_152_port, QN => n_1439);
   reg_key_regx108x : DFF_X1 port map( D => Key(108), CK => clk, Q => 
                           reg_key_108_port, QN => n_1440);
   reg_key_regx41x : DFF_X1 port map( D => Key(41), CK => clk, Q => 
                           reg_key_41_port, QN => n_1441);
   reg_key_regx130x : DFF_X1 port map( D => Key(130), CK => clk, Q => 
                           reg_key_130_port, QN => n_1442);
   reg_key_regx27x : DFF_X1 port map( D => Key(27), CK => clk, Q => 
                           reg_key_27_port, QN => n_1443);
   reg_key_regx23x : DFF_X1 port map( D => Key(23), CK => clk, Q => 
                           reg_key_23_port, QN => n_1444);
   reg_key_regx43x : DFF_X1 port map( D => Key(43), CK => clk, Q => 
                           reg_key_43_port, QN => n_1445);
   reg_key_regx169x : DFF_X1 port map( D => Key(169), CK => clk, Q => 
                           reg_key_169_port, QN => n_1446);
   reg_key_regx131x : DFF_X1 port map( D => Key(131), CK => clk, Q => 
                           reg_key_131_port, QN => n_1447);
   reg_key_regx185x : DFF_X1 port map( D => Key(185), CK => clk, Q => 
                           reg_key_185_port, QN => n_1448);
   reg_key_regx36x : DFF_X1 port map( D => Key(36), CK => clk, Q => 
                           reg_key_36_port, QN => n_1449);
   reg_key_regx86x : DFF_X1 port map( D => Key(86), CK => clk, Q => 
                           reg_key_86_port, QN => n_1450);
   reg_key_regx161x : DFF_X1 port map( D => Key(161), CK => clk, Q => 
                           reg_key_161_port, QN => n_1451);
   reg_key_regx71x : DFF_X1 port map( D => Key(71), CK => clk, Q => 
                           reg_key_71_port, QN => n_1452);
   reg_key_regx123x : DFF_X1 port map( D => Key(123), CK => clk, Q => 
                           reg_key_123_port, QN => n_1453);
   reg_key_regx157x : DFF_X1 port map( D => Key(157), CK => clk, Q => 
                           reg_key_157_port, QN => n_1454);
   reg_key_regx170x : DFF_X1 port map( D => Key(170), CK => clk, Q => 
                           reg_key_170_port, QN => n_1455);
   Ciphertext_regx44x : DFF_X1 port map( D => reg_out_44_port, CK => clk, Q => 
                           Ciphertext(44), QN => n_1456);
   Ciphertext_regx73x : DFF_X1 port map( D => reg_out_73_port, CK => clk, Q => 
                           Ciphertext(73), QN => n_1457);
   reg_key_regx22x : DFF_X1 port map( D => Key(22), CK => clk, Q => 
                           reg_key_22_port, QN => n_1458);
   reg_key_regx186x : DFF_X1 port map( D => Key(186), CK => clk, Q => 
                           reg_key_186_port, QN => n_1459);
   reg_key_regx76x : DFF_X1 port map( D => Key(76), CK => clk, Q => 
                           reg_key_76_port, QN => n_1460);
   reg_key_regx103x : DFF_X1 port map( D => Key(103), CK => clk, Q => 
                           reg_key_103_port, QN => n_1461);
   reg_key_regx48x : DFF_X1 port map( D => Key(48), CK => clk, Q => 
                           reg_key_48_port, QN => n_1462);
   reg_key_regx47x : DFF_X1 port map( D => Key(47), CK => clk, Q => 
                           reg_key_47_port, QN => n_1463);
   reg_key_regx184x : DFF_X1 port map( D => Key(184), CK => clk, Q => 
                           reg_key_184_port, QN => n_1464);
   reg_key_regx156x : DFF_X1 port map( D => Key(156), CK => clk, Q => 
                           reg_key_156_port, QN => n_1465);
   reg_key_regx46x : DFF_X1 port map( D => Key(46), CK => clk, Q => 
                           reg_key_46_port, QN => n_1466);
   reg_key_regx128x : DFF_X1 port map( D => Key(128), CK => clk, Q => 
                           reg_key_128_port, QN => n_1467);
   reg_key_regx73x : DFF_X1 port map( D => Key(73), CK => clk, Q => 
                           reg_key_73_port, QN => n_1468);
   reg_key_regx45x : DFF_X1 port map( D => Key(45), CK => clk, Q => 
                           reg_key_45_port, QN => n_1469);
   reg_key_regx17x : DFF_X1 port map( D => Key(17), CK => clk, Q => 
                           reg_key_17_port, QN => n_1470);
   reg_key_regx154x : DFF_X1 port map( D => Key(154), CK => clk, Q => 
                           reg_key_154_port, QN => n_1471);
   reg_key_regx180x : DFF_X1 port map( D => Key(180), CK => clk, Q => 
                           reg_key_180_port, QN => n_1472);
   reg_key_regx124x : DFF_X1 port map( D => Key(124), CK => clk, Q => 
                           reg_key_124_port, QN => n_1473);
   reg_key_regx96x : DFF_X1 port map( D => Key(96), CK => clk, Q => 
                           reg_key_96_port, QN => n_1474);
   reg_key_regx67x : DFF_X1 port map( D => Key(67), CK => clk, Q => 
                           reg_key_67_port, QN => n_1475);
   reg_key_regx149x : DFF_X1 port map( D => Key(149), CK => clk, Q => 
                           reg_key_149_port, QN => n_1476);
   reg_key_regx39x : DFF_X1 port map( D => Key(39), CK => clk, Q => 
                           reg_key_39_port, QN => n_1477);
   reg_key_regx146x : DFF_X1 port map( D => Key(146), CK => clk, Q => 
                           reg_key_146_port, QN => n_1478);
   reg_key_regx118x : DFF_X1 port map( D => Key(118), CK => clk, Q => 
                           reg_key_118_port, QN => n_1479);
   reg_key_regx63x : DFF_X1 port map( D => Key(63), CK => clk, Q => 
                           reg_key_63_port, QN => n_1480);
   reg_key_regx145x : DFF_X1 port map( D => Key(145), CK => clk, Q => 
                           reg_key_145_port, QN => n_1481);
   reg_key_regx90x : DFF_X1 port map( D => Key(90), CK => clk, Q => 
                           reg_key_90_port, QN => n_1482);
   reg_key_regx117x : DFF_X1 port map( D => Key(117), CK => clk, Q => 
                           reg_key_117_port, QN => n_1483);
   reg_key_regx62x : DFF_X1 port map( D => Key(62), CK => clk, Q => 
                           reg_key_62_port, QN => n_1484);
   reg_key_regx34x : DFF_X1 port map( D => Key(34), CK => clk, Q => 
                           reg_key_34_port, QN => n_1485);
   reg_key_regx143x : DFF_X1 port map( D => Key(143), CK => clk, Q => 
                           reg_key_143_port, QN => n_1486);
   reg_key_regx88x : DFF_X1 port map( D => Key(88), CK => clk, Q => 
                           reg_key_88_port, QN => n_1487);
   reg_key_regx115x : DFF_X1 port map( D => Key(115), CK => clk, Q => 
                           reg_key_115_port, QN => n_1488);
   reg_key_regx5x : DFF_X1 port map( D => Key(5), CK => clk, Q => 
                           reg_key_5_port, QN => n_1489);
   reg_key_regx142x : DFF_X1 port map( D => Key(142), CK => clk, Q => 
                           reg_key_142_port, QN => n_1490);
   reg_key_regx31x : DFF_X1 port map( D => Key(31), CK => clk, Q => 
                           reg_key_31_port, QN => n_1491);
   reg_key_regx113x : DFF_X1 port map( D => Key(113), CK => clk, Q => 
                           reg_key_113_port, QN => n_1492);
   reg_key_regx58x : DFF_X1 port map( D => Key(58), CK => clk, Q => 
                           reg_key_58_port, QN => n_1493);
   reg_key_regx30x : DFF_X1 port map( D => Key(30), CK => clk, Q => 
                           reg_key_30_port, QN => n_1494);
   reg_key_regx29x : DFF_X1 port map( D => Key(29), CK => clk, Q => 
                           reg_key_29_port, QN => n_1495);
   reg_key_regx138x : DFF_X1 port map( D => Key(138), CK => clk, Q => 
                           reg_key_138_port, QN => n_1496);
   reg_key_regx110x : DFF_X1 port map( D => Key(110), CK => clk, Q => 
                           reg_key_110_port, QN => n_1497);
   reg_key_regx55x : DFF_X1 port map( D => Key(55), CK => clk, Q => 
                           reg_key_55_port, QN => n_1498);
   reg_key_regx164x : DFF_X1 port map( D => Key(164), CK => clk, Q => 
                           reg_key_164_port, QN => n_1499);
   reg_key_regx109x : DFF_X1 port map( D => Key(109), CK => clk, Q => 
                           reg_key_109_port, QN => n_1500);
   reg_key_regx136x : DFF_X1 port map( D => Key(136), CK => clk, Q => 
                           reg_key_136_port, QN => n_1501);
   reg_key_regx81x : DFF_X1 port map( D => Key(81), CK => clk, Q => 
                           reg_key_81_port, QN => n_1502);
   reg_key_regx163x : DFF_X1 port map( D => Key(163), CK => clk, Q => 
                           reg_key_163_port, QN => n_1503);
   reg_key_regx162x : DFF_X1 port map( D => Key(162), CK => clk, Q => 
                           reg_key_162_port, QN => n_1504);
   reg_key_regx106x : DFF_X1 port map( D => Key(106), CK => clk, Q => 
                           reg_key_106_port, QN => n_1505);
   reg_key_regx133x : DFF_X1 port map( D => Key(133), CK => clk, Q => 
                           reg_key_133_port, QN => n_1506);
   reg_key_regx105x : DFF_X1 port map( D => Key(105), CK => clk, Q => 
                           reg_key_105_port, QN => n_1507);
   reg_key_regx165x : DFF_X1 port map( D => Key(165), CK => clk, Q => 
                           reg_key_165_port, QN => n_1508);
   reg_key_regx97x : DFF_X1 port map( D => Key(97), CK => clk, Q => 
                           reg_key_97_port, QN => n_1509);
   reg_key_regx158x : DFF_X1 port map( D => Key(158), CK => clk, Q => 
                           reg_key_158_port, QN => n_1510);
   reg_key_regx102x : DFF_X1 port map( D => Key(102), CK => clk, Q => 
                           reg_key_102_port, QN => n_1511);
   reg_key_regx18x : DFF_X1 port map( D => Key(18), CK => clk, Q => 
                           reg_key_18_port, QN => n_1512);
   reg_key_regx182x : DFF_X1 port map( D => Key(182), CK => clk, Q => 
                           reg_key_182_port, QN => n_1513);
   reg_key_regx72x : DFF_X1 port map( D => Key(72), CK => clk, Q => 
                           reg_key_72_port, QN => n_1514);
   reg_key_regx99x : DFF_X1 port map( D => Key(99), CK => clk, Q => 
                           reg_key_99_port, QN => n_1515);
   reg_key_regx181x : DFF_X1 port map( D => Key(181), CK => clk, Q => 
                           reg_key_181_port, QN => n_1516);
   reg_key_regx42x : DFF_X1 port map( D => Key(42), CK => clk, Q => 
                           reg_key_42_port, QN => n_1517);
   reg_key_regx14x : DFF_X1 port map( D => Key(14), CK => clk, Q => 
                           reg_key_14_port, QN => n_1518);
   reg_key_regx12x : DFF_X1 port map( D => Key(12), CK => clk, Q => 
                           reg_key_12_port, QN => n_1519);
   reg_key_regx38x : DFF_X1 port map( D => Key(38), CK => clk, Q => 
                           reg_key_38_port, QN => n_1520);
   reg_key_regx120x : DFF_X1 port map( D => Key(120), CK => clk, Q => 
                           reg_key_120_port, QN => n_1521);
   reg_key_regx10x : DFF_X1 port map( D => Key(10), CK => clk, Q => 
                           reg_key_10_port, QN => n_1522);
   reg_key_regx89x : DFF_X1 port map( D => Key(89), CK => clk, Q => 
                           reg_key_89_port, QN => n_1523);
   reg_key_regx59x : DFF_X1 port map( D => Key(59), CK => clk, Q => 
                           reg_key_59_port, QN => n_1524);
   reg_key_regx85x : DFF_X1 port map( D => Key(85), CK => clk, Q => 
                           reg_key_85_port, QN => n_1525);
   reg_key_regx139x : DFF_X1 port map( D => Key(139), CK => clk, Q => 
                           reg_key_139_port, QN => n_1526);
   reg_key_regx52x : DFF_X1 port map( D => Key(52), CK => clk, Q => 
                           reg_key_52_port, QN => n_1527);
   reg_key_regx132x : DFF_X1 port map( D => Key(132), CK => clk, Q => 
                           reg_key_132_port, QN => n_1528);
   reg_key_regx126x : DFF_X1 port map( D => Key(126), CK => clk, Q => 
                           reg_key_126_port, QN => n_1529);
   reg_key_regx75x : DFF_X1 port map( D => Key(75), CK => clk, Q => 
                           reg_key_75_port, QN => n_1530);
   reg_key_regx127x : DFF_X1 port map( D => Key(127), CK => clk, Q => 
                           reg_key_127_port, QN => n_1531);
   reg_key_regx69x : DFF_X1 port map( D => Key(69), CK => clk, Q => 
                           reg_key_69_port, QN => n_1532);
   reg_key_regx114x : DFF_X1 port map( D => Key(114), CK => clk, Q => 
                           reg_key_114_port, QN => n_1533);
   reg_key_regx141x : DFF_X1 port map( D => Key(141), CK => clk, Q => 
                           reg_key_141_port, QN => n_1534);
   reg_key_regx188x : DFF_X1 port map( D => Key(188), CK => clk, Q => 
                           reg_key_188_port, QN => n_1535);
   reg_key_regx60x : DFF_X1 port map( D => Key(60), CK => clk, Q => 
                           reg_key_60_port, QN => n_1536);
   reg_key_regx6x : DFF_X1 port map( D => Key(6), CK => clk, Q => 
                           reg_key_6_port, QN => n_1537);
   reg_key_regx4x : DFF_X1 port map( D => Key(4), CK => clk, Q => 
                           reg_key_4_port, QN => n_1538);
   reg_key_regx15x : DFF_X1 port map( D => Key(15), CK => clk, Q => 
                           reg_key_15_port, QN => n_1539);
   reg_key_regx24x : DFF_X1 port map( D => Key(24), CK => clk, Q => 
                           reg_key_24_port, QN => n_1540);
   reg_key_regx65x : DFF_X1 port map( D => Key(65), CK => clk, Q => 
                           reg_key_65_port, QN => n_1541);
   reg_key_regx16x : DFF_X1 port map( D => Key(16), CK => clk, Q => 
                           reg_key_16_port, QN => n_1542);
   reg_key_regx0x : DFF_X1 port map( D => Key(0), CK => clk, Q => 
                           reg_key_0_port, QN => n_1543);
   reg_key_regx13x : DFF_X1 port map( D => Key(13), CK => clk, Q => 
                           reg_key_13_port, QN => n_1544);
   reg_key_regx37x : DFF_X1 port map( D => Key(37), CK => clk, Q => 
                           reg_key_37_port, QN => n_1545);
   reg_key_regx93x : DFF_X1 port map( D => Key(93), CK => clk, Q => 
                           reg_key_93_port, QN => n_1546);
   reg_key_regx94x : DFF_X1 port map( D => Key(94), CK => clk, Q => 
                           reg_key_94_port, QN => n_1547);
   reg_key_regx21x : DFF_X1 port map( D => Key(21), CK => clk, Q => 
                           reg_key_21_port, QN => n_1548);
   reg_key_regx7x : DFF_X1 port map( D => Key(7), CK => clk, Q => 
                           reg_key_7_port, QN => n_1549);
   reg_key_regx95x : DFF_X1 port map( D => Key(95), CK => clk, Q => 
                           reg_key_95_port, QN => n_1550);
   reg_key_regx61x : DFF_X1 port map( D => Key(61), CK => clk, Q => 
                           reg_key_61_port, QN => n_1551);
   reg_key_regx121x : DFF_X1 port map( D => Key(121), CK => clk, Q => 
                           reg_key_121_port, QN => n_1552);
   reg_key_regx64x : DFF_X1 port map( D => Key(64), CK => clk, Q => 
                           reg_key_64_port, QN => n_1553);
   reg_key_regx166x : DFF_X1 port map( D => Key(166), CK => clk, Q => 
                           reg_key_166_port, QN => n_1554);
   reg_key_regx84x : DFF_X1 port map( D => Key(84), CK => clk, Q => 
                           reg_key_84_port, QN => n_1555);
   reg_key_regx54x : DFF_X1 port map( D => Key(54), CK => clk, Q => 
                           reg_key_54_port, QN => n_1556);
   reg_key_regx160x : DFF_X1 port map( D => Key(160), CK => clk, Q => 
                           reg_key_160_port, QN => n_1557);
   reg_key_regx25x : DFF_X1 port map( D => Key(25), CK => clk, Q => 
                           reg_key_25_port, QN => n_1558);
   reg_key_regx78x : DFF_X1 port map( D => Key(78), CK => clk, Q => 
                           reg_key_78_port, QN => n_1559);
   Ciphertext_regx105x : DFF_X2 port map( D => reg_out_105_port, CK => clk, Q 
                           => Ciphertext(105), QN => n_1560);
   Ciphertext_regx102x : DFF_X1 port map( D => reg_out_102_port, CK => clk, Q 
                           => Ciphertext(102), QN => n_1561);
   Ciphertext_regx28x : DFF_X2 port map( D => reg_out_28_port, CK => clk, Q => 
                           Ciphertext(28), QN => n_1562);
   reg_key_regx144x : DFF_X1 port map( D => Key(144), CK => clk, Q => 
                           reg_key_144_port, QN => n_1563);
   reg_key_regx172x : DFF_X1 port map( D => Key(172), CK => clk, Q => 
                           reg_key_172_port, QN => n_1564);
   Ciphertext_regx50x : DFFRS_X1 port map( D => reg_out_50_port, CK => clk, RN 
                           => n10, SN => n10, Q => Ciphertext(50), QN => n_1565
                           );
   Ciphertext_regx168x : DFF_X1 port map( D => reg_out_168_port, CK => clk, Q 
                           => Ciphertext(168), QN => n_1566);
   Ciphertext_regx140x : DFF_X1 port map( D => reg_out_140_port, CK => clk, Q 
                           => Ciphertext(140), QN => n_1567);
   reg_key_regx100x : DFF_X1 port map( D => Key(100), CK => clk, Q => 
                           reg_key_100_port, QN => n_1568);
   n10 <= '1';
   SPEEDY_instance : SPEEDY_Rounds7_0 port map( Plaintext(191) => 
                           reg_in_191_port, Plaintext(190) => reg_in_190_port, 
                           Plaintext(189) => reg_in_189_port, Plaintext(188) =>
                           reg_in_188_port, Plaintext(187) => reg_in_187_port, 
                           Plaintext(186) => reg_in_186_port, Plaintext(185) =>
                           reg_in_185_port, Plaintext(184) => reg_in_184_port, 
                           Plaintext(183) => reg_in_183_port, Plaintext(182) =>
                           reg_in_182_port, Plaintext(181) => reg_in_181_port, 
                           Plaintext(180) => reg_in_180_port, Plaintext(179) =>
                           reg_in_179_port, Plaintext(178) => reg_in_178_port, 
                           Plaintext(177) => reg_in_177_port, Plaintext(176) =>
                           reg_in_176_port, Plaintext(175) => reg_in_175_port, 
                           Plaintext(174) => reg_in_174_port, Plaintext(173) =>
                           reg_in_173_port, Plaintext(172) => reg_in_172_port, 
                           Plaintext(171) => reg_in_171_port, Plaintext(170) =>
                           reg_in_170_port, Plaintext(169) => reg_in_169_port, 
                           Plaintext(168) => reg_in_168_port, Plaintext(167) =>
                           reg_in_167_port, Plaintext(166) => reg_in_166_port, 
                           Plaintext(165) => reg_in_165_port, Plaintext(164) =>
                           reg_in_164_port, Plaintext(163) => reg_in_163_port, 
                           Plaintext(162) => reg_in_162_port, Plaintext(161) =>
                           reg_in_161_port, Plaintext(160) => reg_in_160_port, 
                           Plaintext(159) => reg_in_159_port, Plaintext(158) =>
                           reg_in_158_port, Plaintext(157) => reg_in_157_port, 
                           Plaintext(156) => reg_in_156_port, Plaintext(155) =>
                           reg_in_155_port, Plaintext(154) => reg_in_154_port, 
                           Plaintext(153) => reg_in_153_port, Plaintext(152) =>
                           reg_in_152_port, Plaintext(151) => reg_in_151_port, 
                           Plaintext(150) => reg_in_150_port, Plaintext(149) =>
                           reg_in_149_port, Plaintext(148) => reg_in_148_port, 
                           Plaintext(147) => reg_in_147_port, Plaintext(146) =>
                           reg_in_146_port, Plaintext(145) => reg_in_145_port, 
                           Plaintext(144) => reg_in_144_port, Plaintext(143) =>
                           reg_in_143_port, Plaintext(142) => reg_in_142_port, 
                           Plaintext(141) => reg_in_141_port, Plaintext(140) =>
                           reg_in_140_port, Plaintext(139) => reg_in_139_port, 
                           Plaintext(138) => reg_in_138_port, Plaintext(137) =>
                           reg_in_137_port, Plaintext(136) => reg_in_136_port, 
                           Plaintext(135) => reg_in_135_port, Plaintext(134) =>
                           reg_in_134_port, Plaintext(133) => reg_in_133_port, 
                           Plaintext(132) => reg_in_132_port, Plaintext(131) =>
                           reg_in_131_port, Plaintext(130) => reg_in_130_port, 
                           Plaintext(129) => reg_in_129_port, Plaintext(128) =>
                           reg_in_128_port, Plaintext(127) => reg_in_127_port, 
                           Plaintext(126) => reg_in_126_port, Plaintext(125) =>
                           reg_in_125_port, Plaintext(124) => reg_in_124_port, 
                           Plaintext(123) => reg_in_123_port, Plaintext(122) =>
                           reg_in_122_port, Plaintext(121) => reg_in_121_port, 
                           Plaintext(120) => reg_in_120_port, Plaintext(119) =>
                           reg_in_119_port, Plaintext(118) => reg_in_118_port, 
                           Plaintext(117) => reg_in_117_port, Plaintext(116) =>
                           reg_in_116_port, Plaintext(115) => reg_in_115_port, 
                           Plaintext(114) => reg_in_114_port, Plaintext(113) =>
                           reg_in_113_port, Plaintext(112) => reg_in_112_port, 
                           Plaintext(111) => reg_in_111_port, Plaintext(110) =>
                           reg_in_110_port, Plaintext(109) => reg_in_109_port, 
                           Plaintext(108) => reg_in_108_port, Plaintext(107) =>
                           reg_in_107_port, Plaintext(106) => reg_in_106_port, 
                           Plaintext(105) => reg_in_105_port, Plaintext(104) =>
                           reg_in_104_port, Plaintext(103) => reg_in_103_port, 
                           Plaintext(102) => reg_in_102_port, Plaintext(101) =>
                           reg_in_101_port, Plaintext(100) => reg_in_100_port, 
                           Plaintext(99) => reg_in_99_port, Plaintext(98) => 
                           reg_in_98_port, Plaintext(97) => reg_in_97_port, 
                           Plaintext(96) => reg_in_96_port, Plaintext(95) => 
                           reg_in_95_port, Plaintext(94) => reg_in_94_port, 
                           Plaintext(93) => reg_in_93_port, Plaintext(92) => 
                           reg_in_92_port, Plaintext(91) => reg_in_91_port, 
                           Plaintext(90) => reg_in_90_port, Plaintext(89) => 
                           reg_in_89_port, Plaintext(88) => reg_in_88_port, 
                           Plaintext(87) => reg_in_87_port, Plaintext(86) => 
                           reg_in_86_port, Plaintext(85) => reg_in_85_port, 
                           Plaintext(84) => reg_in_84_port, Plaintext(83) => 
                           reg_in_83_port, Plaintext(82) => reg_in_82_port, 
                           Plaintext(81) => reg_in_81_port, Plaintext(80) => 
                           reg_in_80_port, Plaintext(79) => reg_in_79_port, 
                           Plaintext(78) => reg_in_78_port, Plaintext(77) => 
                           reg_in_77_port, Plaintext(76) => reg_in_76_port, 
                           Plaintext(75) => reg_in_75_port, Plaintext(74) => 
                           reg_in_74_port, Plaintext(73) => reg_in_73_port, 
                           Plaintext(72) => reg_in_72_port, Plaintext(71) => 
                           reg_in_71_port, Plaintext(70) => reg_in_70_port, 
                           Plaintext(69) => reg_in_69_port, Plaintext(68) => 
                           reg_in_68_port, Plaintext(67) => reg_in_67_port, 
                           Plaintext(66) => reg_in_66_port, Plaintext(65) => 
                           reg_in_65_port, Plaintext(64) => reg_in_64_port, 
                           Plaintext(63) => reg_in_63_port, Plaintext(62) => 
                           reg_in_62_port, Plaintext(61) => reg_in_61_port, 
                           Plaintext(60) => reg_in_60_port, Plaintext(59) => 
                           reg_in_59_port, Plaintext(58) => reg_in_58_port, 
                           Plaintext(57) => reg_in_57_port, Plaintext(56) => 
                           reg_in_56_port, Plaintext(55) => reg_in_55_port, 
                           Plaintext(54) => reg_in_54_port, Plaintext(53) => 
                           reg_in_53_port, Plaintext(52) => reg_in_52_port, 
                           Plaintext(51) => reg_in_51_port, Plaintext(50) => 
                           reg_in_50_port, Plaintext(49) => reg_in_49_port, 
                           Plaintext(48) => reg_in_48_port, Plaintext(47) => 
                           reg_in_47_port, Plaintext(46) => reg_in_46_port, 
                           Plaintext(45) => reg_in_45_port, Plaintext(44) => 
                           reg_in_44_port, Plaintext(43) => reg_in_43_port, 
                           Plaintext(42) => reg_in_42_port, Plaintext(41) => 
                           reg_in_41_port, Plaintext(40) => reg_in_40_port, 
                           Plaintext(39) => reg_in_39_port, Plaintext(38) => 
                           reg_in_38_port, Plaintext(37) => reg_in_37_port, 
                           Plaintext(36) => reg_in_36_port, Plaintext(35) => 
                           reg_in_35_port, Plaintext(34) => reg_in_34_port, 
                           Plaintext(33) => reg_in_33_port, Plaintext(32) => 
                           reg_in_32_port, Plaintext(31) => reg_in_31_port, 
                           Plaintext(30) => reg_in_30_port, Plaintext(29) => 
                           reg_in_29_port, Plaintext(28) => reg_in_28_port, 
                           Plaintext(27) => reg_in_27_port, Plaintext(26) => 
                           reg_in_26_port, Plaintext(25) => reg_in_25_port, 
                           Plaintext(24) => reg_in_24_port, Plaintext(23) => 
                           reg_in_23_port, Plaintext(22) => reg_in_22_port, 
                           Plaintext(21) => reg_in_21_port, Plaintext(20) => 
                           reg_in_20_port, Plaintext(19) => reg_in_19_port, 
                           Plaintext(18) => reg_in_18_port, Plaintext(17) => 
                           reg_in_17_port, Plaintext(16) => reg_in_16_port, 
                           Plaintext(15) => reg_in_15_port, Plaintext(14) => 
                           reg_in_14_port, Plaintext(13) => reg_in_13_port, 
                           Plaintext(12) => reg_in_12_port, Plaintext(11) => 
                           reg_in_11_port, Plaintext(10) => reg_in_10_port, 
                           Plaintext(9) => reg_in_9_port, Plaintext(8) => 
                           reg_in_8_port, Plaintext(7) => reg_in_7_port, 
                           Plaintext(6) => reg_in_6_port, Plaintext(5) => 
                           reg_in_5_port, Plaintext(4) => reg_in_4_port, 
                           Plaintext(3) => reg_in_3_port, Plaintext(2) => 
                           reg_in_2_port, Plaintext(1) => reg_in_1_port, 
                           Plaintext(0) => reg_in_0_port, Key(191) => 
                           reg_key_191_port, Key(190) => reg_key_190_port, 
                           Key(189) => reg_key_189_port, Key(188) => 
                           reg_key_188_port, Key(187) => reg_key_187_port, 
                           Key(186) => reg_key_186_port, Key(185) => 
                           reg_key_185_port, Key(184) => reg_key_184_port, 
                           Key(183) => reg_key_183_port, Key(182) => 
                           reg_key_182_port, Key(181) => reg_key_181_port, 
                           Key(180) => reg_key_180_port, Key(179) => 
                           reg_key_179_port, Key(178) => reg_key_178_port, 
                           Key(177) => reg_key_177_port, Key(176) => 
                           reg_key_176_port, Key(175) => reg_key_175_port, 
                           Key(174) => reg_key_174_port, Key(173) => 
                           reg_key_173_port, Key(172) => reg_key_172_port, 
                           Key(171) => reg_key_171_port, Key(170) => 
                           reg_key_170_port, Key(169) => reg_key_169_port, 
                           Key(168) => reg_key_168_port, Key(167) => 
                           reg_key_167_port, Key(166) => reg_key_166_port, 
                           Key(165) => reg_key_165_port, Key(164) => 
                           reg_key_164_port, Key(163) => reg_key_163_port, 
                           Key(162) => reg_key_162_port, Key(161) => 
                           reg_key_161_port, Key(160) => reg_key_160_port, 
                           Key(159) => reg_key_159_port, Key(158) => 
                           reg_key_158_port, Key(157) => reg_key_157_port, 
                           Key(156) => reg_key_156_port, Key(155) => 
                           reg_key_155_port, Key(154) => reg_key_154_port, 
                           Key(153) => reg_key_153_port, Key(152) => 
                           reg_key_152_port, Key(151) => reg_key_151_port, 
                           Key(150) => reg_key_150_port, Key(149) => 
                           reg_key_149_port, Key(148) => reg_key_148_port, 
                           Key(147) => reg_key_147_port, Key(146) => 
                           reg_key_146_port, Key(145) => reg_key_145_port, 
                           Key(144) => reg_key_144_port, Key(143) => 
                           reg_key_143_port, Key(142) => reg_key_142_port, 
                           Key(141) => reg_key_141_port, Key(140) => 
                           reg_key_140_port, Key(139) => reg_key_139_port, 
                           Key(138) => reg_key_138_port, Key(137) => 
                           reg_key_137_port, Key(136) => reg_key_136_port, 
                           Key(135) => reg_key_135_port, Key(134) => 
                           reg_key_134_port, Key(133) => reg_key_133_port, 
                           Key(132) => reg_key_132_port, Key(131) => 
                           reg_key_131_port, Key(130) => reg_key_130_port, 
                           Key(129) => reg_key_129_port, Key(128) => 
                           reg_key_128_port, Key(127) => reg_key_127_port, 
                           Key(126) => reg_key_126_port, Key(125) => 
                           reg_key_125_port, Key(124) => reg_key_124_port, 
                           Key(123) => reg_key_123_port, Key(122) => 
                           reg_key_122_port, Key(121) => reg_key_121_port, 
                           Key(120) => reg_key_120_port, Key(119) => 
                           reg_key_119_port, Key(118) => reg_key_118_port, 
                           Key(117) => reg_key_117_port, Key(116) => 
                           reg_key_116_port, Key(115) => reg_key_115_port, 
                           Key(114) => reg_key_114_port, Key(113) => 
                           reg_key_113_port, Key(112) => reg_key_112_port, 
                           Key(111) => reg_key_111_port, Key(110) => 
                           reg_key_110_port, Key(109) => reg_key_109_port, 
                           Key(108) => reg_key_108_port, Key(107) => 
                           reg_key_107_port, Key(106) => reg_key_106_port, 
                           Key(105) => reg_key_105_port, Key(104) => 
                           reg_key_104_port, Key(103) => reg_key_103_port, 
                           Key(102) => reg_key_102_port, Key(101) => 
                           reg_key_101_port, Key(100) => reg_key_100_port, 
                           Key(99) => reg_key_99_port, Key(98) => 
                           reg_key_98_port, Key(97) => reg_key_97_port, Key(96)
                           => reg_key_96_port, Key(95) => reg_key_95_port, 
                           Key(94) => reg_key_94_port, Key(93) => 
                           reg_key_93_port, Key(92) => reg_key_92_port, Key(91)
                           => reg_key_91_port, Key(90) => reg_key_90_port, 
                           Key(89) => reg_key_89_port, Key(88) => 
                           reg_key_88_port, Key(87) => reg_key_87_port, Key(86)
                           => reg_key_86_port, Key(85) => reg_key_85_port, 
                           Key(84) => reg_key_84_port, Key(83) => 
                           reg_key_83_port, Key(82) => reg_key_82_port, Key(81)
                           => reg_key_81_port, Key(80) => reg_key_80_port, 
                           Key(79) => reg_key_79_port, Key(78) => 
                           reg_key_78_port, Key(77) => reg_key_77_port, Key(76)
                           => reg_key_76_port, Key(75) => reg_key_75_port, 
                           Key(74) => reg_key_74_port, Key(73) => 
                           reg_key_73_port, Key(72) => reg_key_72_port, Key(71)
                           => reg_key_71_port, Key(70) => reg_key_70_port, 
                           Key(69) => reg_key_69_port, Key(68) => 
                           reg_key_68_port, Key(67) => reg_key_67_port, Key(66)
                           => reg_key_66_port, Key(65) => reg_key_65_port, 
                           Key(64) => reg_key_64_port, Key(63) => 
                           reg_key_63_port, Key(62) => reg_key_62_port, Key(61)
                           => reg_key_61_port, Key(60) => reg_key_60_port, 
                           Key(59) => reg_key_59_port, Key(58) => 
                           reg_key_58_port, Key(57) => reg_key_57_port, Key(56)
                           => reg_key_56_port, Key(55) => reg_key_55_port, 
                           Key(54) => reg_key_54_port, Key(53) => 
                           reg_key_53_port, Key(52) => reg_key_52_port, Key(51)
                           => reg_key_51_port, Key(50) => reg_key_50_port, 
                           Key(49) => reg_key_49_port, Key(48) => 
                           reg_key_48_port, Key(47) => reg_key_47_port, Key(46)
                           => reg_key_46_port, Key(45) => reg_key_45_port, 
                           Key(44) => reg_key_44_port, Key(43) => 
                           reg_key_43_port, Key(42) => reg_key_42_port, Key(41)
                           => reg_key_41_port, Key(40) => reg_key_40_port, 
                           Key(39) => reg_key_39_port, Key(38) => 
                           reg_key_38_port, Key(37) => reg_key_37_port, Key(36)
                           => reg_key_36_port, Key(35) => reg_key_35_port, 
                           Key(34) => reg_key_34_port, Key(33) => 
                           reg_key_33_port, Key(32) => reg_key_32_port, Key(31)
                           => reg_key_31_port, Key(30) => reg_key_30_port, 
                           Key(29) => reg_key_29_port, Key(28) => 
                           reg_key_28_port, Key(27) => reg_key_27_port, Key(26)
                           => reg_key_26_port, Key(25) => reg_key_25_port, 
                           Key(24) => reg_key_24_port, Key(23) => 
                           reg_key_23_port, Key(22) => reg_key_22_port, Key(21)
                           => reg_key_21_port, Key(20) => reg_key_20_port, 
                           Key(19) => reg_key_19_port, Key(18) => 
                           reg_key_18_port, Key(17) => reg_key_17_port, Key(16)
                           => reg_key_16_port, Key(15) => reg_key_15_port, 
                           Key(14) => reg_key_14_port, Key(13) => 
                           reg_key_13_port, Key(12) => reg_key_12_port, Key(11)
                           => reg_key_11_port, Key(10) => reg_key_10_port, 
                           Key(9) => reg_key_9_port, Key(8) => reg_key_8_port, 
                           Key(7) => reg_key_7_port, Key(6) => reg_key_6_port, 
                           Key(5) => reg_key_5_port, Key(4) => reg_key_4_port, 
                           Key(3) => reg_key_3_port, Key(2) => reg_key_2_port, 
                           Key(1) => reg_key_1_port, Key(0) => reg_key_0_port, 
                           Ciphertext(191) => reg_out_191_port, Ciphertext(190)
                           => reg_out_190_port, Ciphertext(189) => 
                           reg_out_189_port, Ciphertext(188) => 
                           reg_out_188_port, Ciphertext(187) => 
                           reg_out_187_port, Ciphertext(186) => 
                           reg_out_186_port, Ciphertext(185) => 
                           reg_out_185_port, Ciphertext(184) => 
                           reg_out_184_port, Ciphertext(183) => 
                           reg_out_183_port, Ciphertext(182) => 
                           reg_out_182_port, Ciphertext(181) => 
                           reg_out_181_port, Ciphertext(180) => 
                           reg_out_180_port, Ciphertext(179) => 
                           reg_out_179_port, Ciphertext(178) => 
                           reg_out_178_port, Ciphertext(177) => 
                           reg_out_177_port, Ciphertext(176) => 
                           reg_out_176_port, Ciphertext(175) => 
                           reg_out_175_port, Ciphertext(174) => 
                           reg_out_174_port, Ciphertext(173) => 
                           reg_out_173_port, Ciphertext(172) => 
                           reg_out_172_port, Ciphertext(171) => 
                           reg_out_171_port, Ciphertext(170) => 
                           reg_out_170_port, Ciphertext(169) => 
                           reg_out_169_port, Ciphertext(168) => 
                           reg_out_168_port, Ciphertext(167) => 
                           reg_out_167_port, Ciphertext(166) => 
                           reg_out_166_port, Ciphertext(165) => 
                           reg_out_165_port, Ciphertext(164) => 
                           reg_out_164_port, Ciphertext(163) => 
                           reg_out_163_port, Ciphertext(162) => 
                           reg_out_162_port, Ciphertext(161) => 
                           reg_out_161_port, Ciphertext(160) => 
                           reg_out_160_port, Ciphertext(159) => 
                           reg_out_159_port, Ciphertext(158) => 
                           reg_out_158_port, Ciphertext(157) => 
                           reg_out_157_port, Ciphertext(156) => 
                           reg_out_156_port, Ciphertext(155) => 
                           reg_out_155_port, Ciphertext(154) => 
                           reg_out_154_port, Ciphertext(153) => 
                           reg_out_153_port, Ciphertext(152) => 
                           reg_out_152_port, Ciphertext(151) => 
                           reg_out_151_port, Ciphertext(150) => 
                           reg_out_150_port, Ciphertext(149) => 
                           reg_out_149_port, Ciphertext(148) => 
                           reg_out_148_port, Ciphertext(147) => 
                           reg_out_147_port, Ciphertext(146) => 
                           reg_out_146_port, Ciphertext(145) => 
                           reg_out_145_port, Ciphertext(144) => 
                           reg_out_144_port, Ciphertext(143) => 
                           reg_out_143_port, Ciphertext(142) => 
                           reg_out_142_port, Ciphertext(141) => 
                           reg_out_141_port, Ciphertext(140) => 
                           reg_out_140_port, Ciphertext(139) => 
                           reg_out_139_port, Ciphertext(138) => 
                           reg_out_138_port, Ciphertext(137) => 
                           reg_out_137_port, Ciphertext(136) => 
                           reg_out_136_port, Ciphertext(135) => 
                           reg_out_135_port, Ciphertext(134) => 
                           reg_out_134_port, Ciphertext(133) => 
                           reg_out_133_port, Ciphertext(132) => 
                           reg_out_132_port, Ciphertext(131) => 
                           reg_out_131_port, Ciphertext(130) => 
                           reg_out_130_port, Ciphertext(129) => 
                           reg_out_129_port, Ciphertext(128) => 
                           reg_out_128_port, Ciphertext(127) => 
                           reg_out_127_port, Ciphertext(126) => 
                           reg_out_126_port, Ciphertext(125) => 
                           reg_out_125_port, Ciphertext(124) => 
                           reg_out_124_port, Ciphertext(123) => 
                           reg_out_123_port, Ciphertext(122) => 
                           reg_out_122_port, Ciphertext(121) => 
                           reg_out_121_port, Ciphertext(120) => 
                           reg_out_120_port, Ciphertext(119) => 
                           reg_out_119_port, Ciphertext(118) => 
                           reg_out_118_port, Ciphertext(117) => 
                           reg_out_117_port, Ciphertext(116) => 
                           reg_out_116_port, Ciphertext(115) => 
                           reg_out_115_port, Ciphertext(114) => 
                           reg_out_114_port, Ciphertext(113) => 
                           reg_out_113_port, Ciphertext(112) => 
                           reg_out_112_port, Ciphertext(111) => 
                           reg_out_111_port, Ciphertext(110) => 
                           reg_out_110_port, Ciphertext(109) => 
                           reg_out_109_port, Ciphertext(108) => 
                           reg_out_108_port, Ciphertext(107) => 
                           reg_out_107_port, Ciphertext(106) => 
                           reg_out_106_port, Ciphertext(105) => 
                           reg_out_105_port, Ciphertext(104) => 
                           reg_out_104_port, Ciphertext(103) => 
                           reg_out_103_port, Ciphertext(102) => 
                           reg_out_102_port, Ciphertext(101) => 
                           reg_out_101_port, Ciphertext(100) => 
                           reg_out_100_port, Ciphertext(99) => reg_out_99_port,
                           Ciphertext(98) => reg_out_98_port, Ciphertext(97) =>
                           reg_out_97_port, Ciphertext(96) => reg_out_96_port, 
                           Ciphertext(95) => reg_out_95_port, Ciphertext(94) =>
                           reg_out_94_port, Ciphertext(93) => reg_out_93_port, 
                           Ciphertext(92) => reg_out_92_port, Ciphertext(91) =>
                           reg_out_91_port, Ciphertext(90) => reg_out_90_port, 
                           Ciphertext(89) => reg_out_89_port, Ciphertext(88) =>
                           reg_out_88_port, Ciphertext(87) => reg_out_87_port, 
                           Ciphertext(86) => reg_out_86_port, Ciphertext(85) =>
                           reg_out_85_port, Ciphertext(84) => reg_out_84_port, 
                           Ciphertext(83) => reg_out_83_port, Ciphertext(82) =>
                           reg_out_82_port, Ciphertext(81) => reg_out_81_port, 
                           Ciphertext(80) => reg_out_80_port, Ciphertext(79) =>
                           reg_out_79_port, Ciphertext(78) => reg_out_78_port, 
                           Ciphertext(77) => reg_out_77_port, Ciphertext(76) =>
                           reg_out_76_port, Ciphertext(75) => reg_out_75_port, 
                           Ciphertext(74) => reg_out_74_port, Ciphertext(73) =>
                           reg_out_73_port, Ciphertext(72) => reg_out_72_port, 
                           Ciphertext(71) => reg_out_71_port, Ciphertext(70) =>
                           reg_out_70_port, Ciphertext(69) => reg_out_69_port, 
                           Ciphertext(68) => reg_out_68_port, Ciphertext(67) =>
                           reg_out_67_port, Ciphertext(66) => reg_out_66_port, 
                           Ciphertext(65) => reg_out_65_port, Ciphertext(64) =>
                           reg_out_64_port, Ciphertext(63) => reg_out_63_port, 
                           Ciphertext(62) => reg_out_62_port, Ciphertext(61) =>
                           reg_out_61_port, Ciphertext(60) => reg_out_60_port, 
                           Ciphertext(59) => reg_out_59_port, Ciphertext(58) =>
                           reg_out_58_port, Ciphertext(57) => reg_out_57_port, 
                           Ciphertext(56) => reg_out_56_port, Ciphertext(55) =>
                           reg_out_55_port, Ciphertext(54) => reg_out_54_port, 
                           Ciphertext(53) => reg_out_53_port, Ciphertext(52) =>
                           reg_out_52_port, Ciphertext(51) => reg_out_51_port, 
                           Ciphertext(50) => reg_out_50_port, Ciphertext(49) =>
                           reg_out_49_port, Ciphertext(48) => reg_out_48_port, 
                           Ciphertext(47) => reg_out_47_port, Ciphertext(46) =>
                           reg_out_46_port, Ciphertext(45) => reg_out_45_port, 
                           Ciphertext(44) => reg_out_44_port, Ciphertext(43) =>
                           reg_out_43_port, Ciphertext(42) => reg_out_42_port, 
                           Ciphertext(41) => reg_out_41_port, Ciphertext(40) =>
                           reg_out_40_port, Ciphertext(39) => reg_out_39_port, 
                           Ciphertext(38) => reg_out_38_port, Ciphertext(37) =>
                           reg_out_37_port, Ciphertext(36) => reg_out_36_port, 
                           Ciphertext(35) => reg_out_35_port, Ciphertext(34) =>
                           reg_out_34_port, Ciphertext(33) => reg_out_33_port, 
                           Ciphertext(32) => reg_out_32_port, Ciphertext(31) =>
                           reg_out_31_port, Ciphertext(30) => reg_out_30_port, 
                           Ciphertext(29) => reg_out_29_port, Ciphertext(28) =>
                           reg_out_28_port, Ciphertext(27) => reg_out_27_port, 
                           Ciphertext(26) => reg_out_26_port, Ciphertext(25) =>
                           reg_out_25_port, Ciphertext(24) => reg_out_24_port, 
                           Ciphertext(23) => reg_out_23_port, Ciphertext(22) =>
                           reg_out_22_port, Ciphertext(21) => reg_out_21_port, 
                           Ciphertext(20) => reg_out_20_port, Ciphertext(19) =>
                           reg_out_19_port, Ciphertext(18) => reg_out_18_port, 
                           Ciphertext(17) => reg_out_17_port, Ciphertext(16) =>
                           reg_out_16_port, Ciphertext(15) => reg_out_15_port, 
                           Ciphertext(14) => reg_out_14_port, Ciphertext(13) =>
                           reg_out_13_port, Ciphertext(12) => reg_out_12_port, 
                           Ciphertext(11) => reg_out_11_port, Ciphertext(10) =>
                           reg_out_10_port, Ciphertext(9) => reg_out_9_port, 
                           Ciphertext(8) => reg_out_8_port, Ciphertext(7) => 
                           reg_out_7_port, Ciphertext(6) => reg_out_6_port, 
                           Ciphertext(5) => reg_out_5_port, Ciphertext(4) => 
                           reg_out_4_port, Ciphertext(3) => reg_out_3_port, 
                           Ciphertext(2) => reg_out_2_port, Ciphertext(1) => 
                           reg_out_1_port, Ciphertext(0) => reg_out_0_port);
   Ciphertext_regx111x : DFF_X2 port map( D => reg_out_111_port, CK => clk, Q 
                           => Ciphertext(111), QN => n_1569);
   Ciphertext_regx108x : DFF_X2 port map( D => reg_out_108_port, CK => clk, Q 
                           => Ciphertext(108), QN => n_1570);
   Ciphertext_regx121x : DFFRS_X1 port map( D => reg_out_121_port, CK => clk, 
                           RN => n12, SN => n12, Q => Ciphertext(121), QN => 
                           n_1571);
   Ciphertext_regx84x : DFF_X2 port map( D => reg_out_84_port, CK => clk, Q => 
                           Ciphertext(84), QN => n_1572);
   Ciphertext_regx188x : DFF_X2 port map( D => reg_out_188_port, CK => clk, Q 
                           => Ciphertext(188), QN => n_1573);
   Ciphertext_regx0x : DFF_X1 port map( D => reg_out_0_port, CK => clk, Q => 
                           Ciphertext(0), QN => n_1574);
   Ciphertext_regx148x : DFF_X1 port map( D => reg_out_148_port, CK => clk, Q 
                           => Ciphertext(148), QN => n_1575);
   n12 <= '1';

end SYN_Behavioral;
