module SPEEDY_Rounds5_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   \RI1[1][191] , \RI1[1][190] , \RI1[1][189] , \RI1[1][188] ,
         \RI1[1][187] , \RI1[1][186] , \RI1[1][185] , \RI1[1][184] ,
         \RI1[1][183] , \RI1[1][182] , \RI1[1][181] , \RI1[1][180] ,
         \RI1[1][179] , \RI1[1][178] , \RI1[1][177] , \RI1[1][176] ,
         \RI1[1][175] , \RI1[1][174] , \RI1[1][173] , \RI1[1][172] ,
         \RI1[1][171] , \RI1[1][170] , \RI1[1][169] , \RI1[1][168] ,
         \RI1[1][167] , \RI1[1][166] , \RI1[1][165] , \RI1[1][164] ,
         \RI1[1][163] , \RI1[1][162] , \RI1[1][161] , \RI1[1][160] ,
         \RI1[1][159] , \RI1[1][158] , \RI1[1][157] , \RI1[1][156] ,
         \RI1[1][155] , \RI1[1][154] , \RI1[1][153] , \RI1[1][152] ,
         \RI1[1][151] , \RI1[1][150] , \RI1[1][149] , \RI1[1][148] ,
         \RI1[1][147] , \RI1[1][146] , \RI1[1][145] , \RI1[1][144] ,
         \RI1[1][143] , \RI1[1][142] , \RI1[1][141] , \RI1[1][140] ,
         \RI1[1][139] , \RI1[1][138] , \RI1[1][137] , \RI1[1][136] ,
         \RI1[1][135] , \RI1[1][134] , \RI1[1][133] , \RI1[1][132] ,
         \RI1[1][131] , \RI1[1][130] , \RI1[1][129] , \RI1[1][128] ,
         \RI1[1][127] , \RI1[1][126] , \RI1[1][125] , \RI1[1][124] ,
         \RI1[1][123] , \RI1[1][122] , \RI1[1][121] , \RI1[1][120] ,
         \RI1[1][119] , \RI1[1][118] , \RI1[1][117] , \RI1[1][116] ,
         \RI1[1][115] , \RI1[1][114] , \RI1[1][113] , \RI1[1][112] ,
         \RI1[1][111] , \RI1[1][110] , \RI1[1][109] , \RI1[1][108] ,
         \RI1[1][107] , \RI1[1][106] , \RI1[1][105] , \RI1[1][104] ,
         \RI1[1][103] , \RI1[1][102] , \RI1[1][101] , \RI1[1][100] ,
         \RI1[1][99] , \RI1[1][98] , \RI1[1][97] , \RI1[1][96] , \RI1[1][95] ,
         \RI1[1][94] , \RI1[1][93] , \RI1[1][92] , \RI1[1][91] , \RI1[1][90] ,
         \RI1[1][89] , \RI1[1][88] , \RI1[1][87] , \RI1[1][86] , \RI1[1][85] ,
         \RI1[1][84] , \RI1[1][83] , \RI1[1][82] , \RI1[1][81] , \RI1[1][80] ,
         \RI1[1][79] , \RI1[1][78] , \RI1[1][77] , \RI1[1][76] , \RI1[1][75] ,
         \RI1[1][74] , \RI1[1][73] , \RI1[1][72] , \RI1[1][71] , \RI1[1][70] ,
         \RI1[1][69] , \RI1[1][68] , \RI1[1][67] , \RI1[1][66] , \RI1[1][65] ,
         \RI1[1][64] , \RI1[1][63] , \RI1[1][62] , \RI1[1][61] , \RI1[1][60] ,
         \RI1[1][59] , \RI1[1][58] , \RI1[1][57] , \RI1[1][56] , \RI1[1][55] ,
         \RI1[1][54] , \RI1[1][53] , \RI1[1][52] , \RI1[1][51] , \RI1[1][50] ,
         \RI1[1][49] , \RI1[1][48] , \RI1[1][47] , \RI1[1][46] , \RI1[1][45] ,
         \RI1[1][44] , \RI1[1][43] , \RI1[1][42] , \RI1[1][41] , \RI1[1][40] ,
         \RI1[1][39] , \RI1[1][38] , \RI1[1][37] , \RI1[1][36] , \RI1[1][35] ,
         \RI1[1][34] , \RI1[1][33] , \RI1[1][32] , \RI1[1][31] , \RI1[1][30] ,
         \RI1[1][29] , \RI1[1][28] , \RI1[1][27] , \RI1[1][26] , \RI1[1][25] ,
         \RI1[1][24] , \RI1[1][23] , \RI1[1][22] , \RI1[1][21] , \RI1[1][20] ,
         \RI1[1][19] , \RI1[1][18] , \RI1[1][17] , \RI1[1][16] , \RI1[1][15] ,
         \RI1[1][14] , \RI1[1][13] , \RI1[1][12] , \RI1[1][11] , \RI1[1][10] ,
         \RI1[1][9] , \RI1[1][8] , \RI1[1][7] , \RI1[1][6] , \RI1[1][5] ,
         \RI1[1][4] , \RI1[1][3] , \RI1[1][2] , \RI1[1][1] , \RI1[1][0] ,
         \RI1[2][191] , \RI1[2][190] , \RI1[2][189] , \RI1[2][188] ,
         \RI1[2][187] , \RI1[2][186] , \RI1[2][185] , \RI1[2][184] ,
         \RI1[2][183] , \RI1[2][182] , \RI1[2][181] , \RI1[2][180] ,
         \RI1[2][179] , \RI1[2][178] , \RI1[2][177] , \RI1[2][176] ,
         \RI1[2][175] , \RI1[2][174] , \RI1[2][173] , \RI1[2][172] ,
         \RI1[2][171] , \RI1[2][170] , \RI1[2][169] , \RI1[2][168] ,
         \RI1[2][167] , \RI1[2][166] , \RI1[2][165] , \RI1[2][164] ,
         \RI1[2][163] , \RI1[2][162] , \RI1[2][161] , \RI1[2][160] ,
         \RI1[2][159] , \RI1[2][158] , \RI1[2][157] , \RI1[2][156] ,
         \RI1[2][155] , \RI1[2][154] , \RI1[2][153] , \RI1[2][152] ,
         \RI1[2][151] , \RI1[2][150] , \RI1[2][149] , \RI1[2][148] ,
         \RI1[2][147] , \RI1[2][146] , \RI1[2][145] , \RI1[2][144] ,
         \RI1[2][143] , \RI1[2][142] , \RI1[2][141] , \RI1[2][140] ,
         \RI1[2][139] , \RI1[2][138] , \RI1[2][137] , \RI1[2][136] ,
         \RI1[2][135] , \RI1[2][134] , \RI1[2][133] , \RI1[2][132] ,
         \RI1[2][131] , \RI1[2][130] , \RI1[2][129] , \RI1[2][128] ,
         \RI1[2][127] , \RI1[2][126] , \RI1[2][125] , \RI1[2][124] ,
         \RI1[2][123] , \RI1[2][122] , \RI1[2][121] , \RI1[2][120] ,
         \RI1[2][119] , \RI1[2][118] , \RI1[2][117] , \RI1[2][116] ,
         \RI1[2][115] , \RI1[2][114] , \RI1[2][113] , \RI1[2][112] ,
         \RI1[2][111] , \RI1[2][110] , \RI1[2][109] , \RI1[2][108] ,
         \RI1[2][107] , \RI1[2][106] , \RI1[2][105] , \RI1[2][104] ,
         \RI1[2][103] , \RI1[2][102] , \RI1[2][101] , \RI1[2][100] ,
         \RI1[2][99] , \RI1[2][98] , \RI1[2][97] , \RI1[2][96] , \RI1[2][95] ,
         \RI1[2][94] , \RI1[2][93] , \RI1[2][92] , \RI1[2][91] , \RI1[2][90] ,
         \RI1[2][89] , \RI1[2][88] , \RI1[2][87] , \RI1[2][86] , \RI1[2][85] ,
         \RI1[2][84] , \RI1[2][83] , \RI1[2][82] , \RI1[2][81] , \RI1[2][80] ,
         \RI1[2][79] , \RI1[2][78] , \RI1[2][77] , \RI1[2][76] , \RI1[2][75] ,
         \RI1[2][74] , \RI1[2][73] , \RI1[2][72] , \RI1[2][71] , \RI1[2][70] ,
         \RI1[2][69] , \RI1[2][68] , \RI1[2][67] , \RI1[2][66] , \RI1[2][65] ,
         \RI1[2][64] , \RI1[2][63] , \RI1[2][62] , \RI1[2][61] , \RI1[2][60] ,
         \RI1[2][59] , \RI1[2][58] , \RI1[2][57] , \RI1[2][56] , \RI1[2][55] ,
         \RI1[2][54] , \RI1[2][53] , \RI1[2][52] , \RI1[2][51] , \RI1[2][50] ,
         \RI1[2][49] , \RI1[2][48] , \RI1[2][47] , \RI1[2][46] , \RI1[2][45] ,
         \RI1[2][44] , \RI1[2][43] , \RI1[2][42] , \RI1[2][41] , \RI1[2][40] ,
         \RI1[2][39] , \RI1[2][38] , \RI1[2][37] , \RI1[2][36] , \RI1[2][35] ,
         \RI1[2][34] , \RI1[2][33] , \RI1[2][32] , \RI1[2][31] , \RI1[2][30] ,
         \RI1[2][29] , \RI1[2][28] , \RI1[2][27] , \RI1[2][26] , \RI1[2][25] ,
         \RI1[2][24] , \RI1[2][23] , \RI1[2][22] , \RI1[2][21] , \RI1[2][20] ,
         \RI1[2][19] , \RI1[2][18] , \RI1[2][17] , \RI1[2][16] , \RI1[2][15] ,
         \RI1[2][14] , \RI1[2][13] , \RI1[2][12] , \RI1[2][11] , \RI1[2][10] ,
         \RI1[2][9] , \RI1[2][8] , \RI1[2][7] , \RI1[2][6] , \RI1[2][5] ,
         \RI1[2][4] , \RI1[2][3] , \RI1[2][2] , \RI1[2][1] , \RI1[2][0] ,
         \RI1[3][191] , \RI1[3][190] , \RI1[3][189] , \RI1[3][188] ,
         \RI1[3][187] , \RI1[3][186] , \RI1[3][185] , \RI1[3][184] ,
         \RI1[3][183] , \RI1[3][182] , \RI1[3][181] , \RI1[3][180] ,
         \RI1[3][179] , \RI1[3][178] , \RI1[3][177] , \RI1[3][176] ,
         \RI1[3][175] , \RI1[3][174] , \RI1[3][173] , \RI1[3][172] ,
         \RI1[3][171] , \RI1[3][170] , \RI1[3][169] , \RI1[3][168] ,
         \RI1[3][167] , \RI1[3][166] , \RI1[3][165] , \RI1[3][164] ,
         \RI1[3][163] , \RI1[3][162] , \RI1[3][161] , \RI1[3][160] ,
         \RI1[3][159] , \RI1[3][158] , \RI1[3][157] , \RI1[3][156] ,
         \RI1[3][155] , \RI1[3][154] , \RI1[3][153] , \RI1[3][152] ,
         \RI1[3][151] , \RI1[3][150] , \RI1[3][149] , \RI1[3][148] ,
         \RI1[3][147] , \RI1[3][146] , \RI1[3][145] , \RI1[3][144] ,
         \RI1[3][143] , \RI1[3][142] , \RI1[3][141] , \RI1[3][140] ,
         \RI1[3][139] , \RI1[3][138] , \RI1[3][137] , \RI1[3][136] ,
         \RI1[3][135] , \RI1[3][134] , \RI1[3][133] , \RI1[3][132] ,
         \RI1[3][131] , \RI1[3][130] , \RI1[3][129] , \RI1[3][128] ,
         \RI1[3][127] , \RI1[3][126] , \RI1[3][125] , \RI1[3][124] ,
         \RI1[3][123] , \RI1[3][122] , \RI1[3][121] , \RI1[3][120] ,
         \RI1[3][119] , \RI1[3][118] , \RI1[3][117] , \RI1[3][116] ,
         \RI1[3][115] , \RI1[3][114] , \RI1[3][113] , \RI1[3][112] ,
         \RI1[3][111] , \RI1[3][110] , \RI1[3][109] , \RI1[3][108] ,
         \RI1[3][107] , \RI1[3][106] , \RI1[3][105] , \RI1[3][104] ,
         \RI1[3][103] , \RI1[3][102] , \RI1[3][101] , \RI1[3][100] ,
         \RI1[3][99] , \RI1[3][98] , \RI1[3][97] , \RI1[3][96] , \RI1[3][95] ,
         \RI1[3][94] , \RI1[3][93] , \RI1[3][92] , \RI1[3][91] , \RI1[3][90] ,
         \RI1[3][89] , \RI1[3][88] , \RI1[3][87] , \RI1[3][86] , \RI1[3][85] ,
         \RI1[3][84] , \RI1[3][83] , \RI1[3][82] , \RI1[3][81] , \RI1[3][80] ,
         \RI1[3][79] , \RI1[3][78] , \RI1[3][77] , \RI1[3][76] , \RI1[3][75] ,
         \RI1[3][74] , \RI1[3][73] , \RI1[3][72] , \RI1[3][71] , \RI1[3][70] ,
         \RI1[3][69] , \RI1[3][68] , \RI1[3][67] , \RI1[3][66] , \RI1[3][65] ,
         \RI1[3][64] , \RI1[3][63] , \RI1[3][62] , \RI1[3][61] , \RI1[3][60] ,
         \RI1[3][59] , \RI1[3][58] , \RI1[3][57] , \RI1[3][56] , \RI1[3][55] ,
         \RI1[3][54] , \RI1[3][53] , \RI1[3][52] , \RI1[3][51] , \RI1[3][50] ,
         \RI1[3][49] , \RI1[3][48] , \RI1[3][47] , \RI1[3][46] , \RI1[3][45] ,
         \RI1[3][44] , \RI1[3][43] , \RI1[3][42] , \RI1[3][41] , \RI1[3][40] ,
         \RI1[3][39] , \RI1[3][38] , \RI1[3][37] , \RI1[3][36] , \RI1[3][35] ,
         \RI1[3][34] , \RI1[3][33] , \RI1[3][32] , \RI1[3][31] , \RI1[3][30] ,
         \RI1[3][29] , \RI1[3][28] , \RI1[3][27] , \RI1[3][26] , \RI1[3][25] ,
         \RI1[3][24] , \RI1[3][23] , \RI1[3][22] , \RI1[3][21] , \RI1[3][20] ,
         \RI1[3][19] , \RI1[3][18] , \RI1[3][17] , \RI1[3][16] , \RI1[3][15] ,
         \RI1[3][14] , \RI1[3][13] , \RI1[3][12] , \RI1[3][11] , \RI1[3][10] ,
         \RI1[3][9] , \RI1[3][8] , \RI1[3][7] , \RI1[3][6] , \RI1[3][5] ,
         \RI1[3][4] , \RI1[3][3] , \RI1[3][2] , \RI1[3][1] , \RI1[3][0] ,
         \RI1[4][191] , \RI1[4][190] , \RI1[4][189] , \RI1[4][188] ,
         \RI1[4][187] , \RI1[4][186] , \RI1[4][185] , \RI1[4][184] ,
         \RI1[4][183] , \RI1[4][182] , \RI1[4][181] , \RI1[4][180] ,
         \RI1[4][179] , \RI1[4][178] , \RI1[4][177] , \RI1[4][176] ,
         \RI1[4][175] , \RI1[4][174] , \RI1[4][173] , \RI1[4][172] ,
         \RI1[4][171] , \RI1[4][170] , \RI1[4][169] , \RI1[4][168] ,
         \RI1[4][167] , \RI1[4][166] , \RI1[4][165] , \RI1[4][164] ,
         \RI1[4][163] , \RI1[4][162] , \RI1[4][161] , \RI1[4][160] ,
         \RI1[4][159] , \RI1[4][158] , \RI1[4][157] , \RI1[4][156] ,
         \RI1[4][155] , \RI1[4][154] , \RI1[4][153] , \RI1[4][152] ,
         \RI1[4][151] , \RI1[4][150] , \RI1[4][149] , \RI1[4][148] ,
         \RI1[4][147] , \RI1[4][146] , \RI1[4][145] , \RI1[4][144] ,
         \RI1[4][143] , \RI1[4][142] , \RI1[4][141] , \RI1[4][140] ,
         \RI1[4][139] , \RI1[4][138] , \RI1[4][137] , \RI1[4][136] ,
         \RI1[4][135] , \RI1[4][134] , \RI1[4][133] , \RI1[4][132] ,
         \RI1[4][131] , \RI1[4][130] , \RI1[4][129] , \RI1[4][128] ,
         \RI1[4][127] , \RI1[4][126] , \RI1[4][125] , \RI1[4][124] ,
         \RI1[4][123] , \RI1[4][122] , \RI1[4][121] , \RI1[4][120] ,
         \RI1[4][119] , \RI1[4][118] , \RI1[4][117] , \RI1[4][116] ,
         \RI1[4][115] , \RI1[4][114] , \RI1[4][113] , \RI1[4][112] ,
         \RI1[4][111] , \RI1[4][110] , \RI1[4][109] , \RI1[4][108] ,
         \RI1[4][107] , \RI1[4][106] , \RI1[4][105] , \RI1[4][104] ,
         \RI1[4][103] , \RI1[4][102] , \RI1[4][101] , \RI1[4][100] ,
         \RI1[4][99] , \RI1[4][98] , \RI1[4][97] , \RI1[4][96] , \RI1[4][95] ,
         \RI1[4][94] , \RI1[4][93] , \RI1[4][92] , \RI1[4][91] , \RI1[4][90] ,
         \RI1[4][89] , \RI1[4][88] , \RI1[4][87] , \RI1[4][86] , \RI1[4][85] ,
         \RI1[4][84] , \RI1[4][83] , \RI1[4][82] , \RI1[4][81] , \RI1[4][80] ,
         \RI1[4][79] , \RI1[4][78] , \RI1[4][77] , \RI1[4][76] , \RI1[4][75] ,
         \RI1[4][74] , \RI1[4][73] , \RI1[4][72] , \RI1[4][71] , \RI1[4][70] ,
         \RI1[4][69] , \RI1[4][68] , \RI1[4][67] , \RI1[4][66] , \RI1[4][65] ,
         \RI1[4][64] , \RI1[4][63] , \RI1[4][62] , \RI1[4][61] , \RI1[4][60] ,
         \RI1[4][59] , \RI1[4][58] , \RI1[4][57] , \RI1[4][56] , \RI1[4][55] ,
         \RI1[4][54] , \RI1[4][53] , \RI1[4][52] , \RI1[4][51] , \RI1[4][50] ,
         \RI1[4][49] , \RI1[4][48] , \RI1[4][47] , \RI1[4][46] , \RI1[4][45] ,
         \RI1[4][44] , \RI1[4][43] , \RI1[4][42] , \RI1[4][41] , \RI1[4][40] ,
         \RI1[4][39] , \RI1[4][38] , \RI1[4][37] , \RI1[4][36] , \RI1[4][35] ,
         \RI1[4][34] , \RI1[4][33] , \RI1[4][32] , \RI1[4][31] , \RI1[4][30] ,
         \RI1[4][29] , \RI1[4][28] , \RI1[4][27] , \RI1[4][26] , \RI1[4][25] ,
         \RI1[4][24] , \RI1[4][23] , \RI1[4][22] , \RI1[4][21] , \RI1[4][20] ,
         \RI1[4][19] , \RI1[4][18] , \RI1[4][17] , \RI1[4][16] , \RI1[4][15] ,
         \RI1[4][14] , \RI1[4][13] , \RI1[4][12] , \RI1[4][11] , \RI1[4][10] ,
         \RI1[4][9] , \RI1[4][8] , \RI1[4][7] , \RI1[4][6] , \RI1[4][5] ,
         \RI1[4][4] , \RI1[4][3] , \RI1[4][2] , \RI1[4][1] , \RI1[4][0] ,
         \RI3[0][191] , \RI3[0][190] , \RI3[0][189] , \RI3[0][188] ,
         \RI3[0][187] , \RI3[0][186] , \RI3[0][185] , \RI3[0][184] ,
         \RI3[0][183] , \RI3[0][182] , \RI3[0][181] , \RI3[0][180] ,
         \RI3[0][179] , \RI3[0][178] , \RI3[0][177] , \RI3[0][176] ,
         \RI3[0][175] , \RI3[0][174] , \RI3[0][173] , \RI3[0][171] ,
         \RI3[0][170] , \RI3[0][169] , \RI3[0][168] , \RI3[0][167] ,
         \RI3[0][166] , \RI3[0][165] , \RI3[0][164] , \RI3[0][163] ,
         \RI3[0][162] , \RI3[0][161] , \RI3[0][160] , \RI3[0][159] ,
         \RI3[0][158] , \RI3[0][157] , \RI3[0][156] , \RI3[0][155] ,
         \RI3[0][154] , \RI3[0][153] , \RI3[0][152] , \RI3[0][151] ,
         \RI3[0][150] , \RI3[0][149] , \RI3[0][148] , \RI3[0][147] ,
         \RI3[0][146] , \RI3[0][145] , \RI3[0][144] , \RI3[0][143] ,
         \RI3[0][142] , \RI3[0][141] , \RI3[0][140] , \RI3[0][139] ,
         \RI3[0][138] , \RI3[0][137] , \RI3[0][136] , \RI3[0][135] ,
         \RI3[0][134] , \RI3[0][133] , \RI3[0][132] , \RI3[0][131] ,
         \RI3[0][130] , \RI3[0][129] , \RI3[0][128] , \RI3[0][127] ,
         \RI3[0][126] , \RI3[0][125] , \RI3[0][124] , \RI3[0][123] ,
         \RI3[0][122] , \RI3[0][121] , \RI3[0][120] , \RI3[0][119] ,
         \RI3[0][118] , \RI3[0][117] , \RI3[0][116] , \RI3[0][115] ,
         \RI3[0][114] , \RI3[0][113] , \RI3[0][112] , \RI3[0][111] ,
         \RI3[0][110] , \RI3[0][109] , \RI3[0][108] , \RI3[0][107] ,
         \RI3[0][106] , \RI3[0][105] , \RI3[0][104] , \RI3[0][103] ,
         \RI3[0][102] , \RI3[0][101] , \RI3[0][99] , \RI3[0][98] ,
         \RI3[0][97] , \RI3[0][96] , \RI3[0][95] , \RI3[0][94] , \RI3[0][93] ,
         \RI3[0][92] , \RI3[0][91] , \RI3[0][90] , \RI3[0][89] , \RI3[0][88] ,
         \RI3[0][87] , \RI3[0][86] , \RI3[0][85] , \RI3[0][84] , \RI3[0][83] ,
         \RI3[0][82] , \RI3[0][81] , \RI3[0][80] , \RI3[0][79] , \RI3[0][78] ,
         \RI3[0][77] , \RI3[0][76] , \RI3[0][75] , \RI3[0][74] , \RI3[0][73] ,
         \RI3[0][72] , \RI3[0][71] , \RI3[0][70] , \RI3[0][69] , \RI3[0][68] ,
         \RI3[0][67] , \RI3[0][66] , \RI3[0][65] , \RI3[0][64] , \RI3[0][63] ,
         \RI3[0][62] , \RI3[0][61] , \RI3[0][60] , \RI3[0][59] , \RI3[0][58] ,
         \RI3[0][57] , \RI3[0][56] , \RI3[0][55] , \RI3[0][54] , \RI3[0][53] ,
         \RI3[0][51] , \RI3[0][50] , \RI3[0][49] , \RI3[0][48] , \RI3[0][47] ,
         \RI3[0][46] , \RI3[0][45] , \RI3[0][44] , \RI3[0][43] , \RI3[0][42] ,
         \RI3[0][41] , \RI3[0][40] , \RI3[0][39] , \RI3[0][38] , \RI3[0][37] ,
         \RI3[0][36] , \RI3[0][35] , \RI3[0][34] , \RI3[0][33] , \RI3[0][32] ,
         \RI3[0][31] , \RI3[0][30] , \RI3[0][29] , \RI3[0][28] , \RI3[0][27] ,
         \RI3[0][26] , \RI3[0][25] , \RI3[0][24] , \RI3[0][23] , \RI3[0][22] ,
         \RI3[0][21] , \RI3[0][20] , \RI3[0][19] , \RI3[0][18] , \RI3[0][17] ,
         \RI3[0][16] , \RI3[0][15] , \RI3[0][14] , \RI3[0][13] , \RI3[0][12] ,
         \RI3[0][11] , \RI3[0][10] , \RI3[0][9] , \RI3[0][8] , \RI3[0][7] ,
         \RI3[0][6] , \RI3[0][5] , \RI3[0][4] , \RI3[0][3] , \RI3[0][2] ,
         \RI3[0][1] , \RI3[0][0] , \RI3[1][191] , \RI3[1][190] , \RI3[1][189] ,
         \RI3[1][188] , \RI3[1][187] , \RI3[1][186] , \RI3[1][185] ,
         \RI3[1][184] , \RI3[1][183] , \RI3[1][182] , \RI3[1][181] ,
         \RI3[1][180] , \RI3[1][179] , \RI3[1][178] , \RI3[1][177] ,
         \RI3[1][176] , \RI3[1][175] , \RI3[1][174] , \RI3[1][173] ,
         \RI3[1][172] , \RI3[1][171] , \RI3[1][170] , \RI3[1][169] ,
         \RI3[1][168] , \RI3[1][167] , \RI3[1][166] , \RI3[1][165] ,
         \RI3[1][164] , \RI3[1][163] , \RI3[1][162] , \RI3[1][161] ,
         \RI3[1][160] , \RI3[1][159] , \RI3[1][158] , \RI3[1][157] ,
         \RI3[1][156] , \RI3[1][155] , \RI3[1][154] , \RI3[1][153] ,
         \RI3[1][152] , \RI3[1][151] , \RI3[1][150] , \RI3[1][149] ,
         \RI3[1][147] , \RI3[1][146] , \RI3[1][145] , \RI3[1][144] ,
         \RI3[1][143] , \RI3[1][142] , \RI3[1][141] , \RI3[1][140] ,
         \RI3[1][139] , \RI3[1][138] , \RI3[1][137] , \RI3[1][136] ,
         \RI3[1][135] , \RI3[1][134] , \RI3[1][133] , \RI3[1][132] ,
         \RI3[1][131] , \RI3[1][130] , \RI3[1][129] , \RI3[1][128] ,
         \RI3[1][127] , \RI3[1][126] , \RI3[1][125] , \RI3[1][124] ,
         \RI3[1][123] , \RI3[1][122] , \RI3[1][121] , \RI3[1][120] ,
         \RI3[1][119] , \RI3[1][118] , \RI3[1][117] , \RI3[1][116] ,
         \RI3[1][115] , \RI3[1][114] , \RI3[1][113] , \RI3[1][112] ,
         \RI3[1][111] , \RI3[1][110] , \RI3[1][109] , \RI3[1][108] ,
         \RI3[1][107] , \RI3[1][106] , \RI3[1][105] , \RI3[1][104] ,
         \RI3[1][103] , \RI3[1][102] , \RI3[1][101] , \RI3[1][100] ,
         \RI3[1][99] , \RI3[1][98] , \RI3[1][97] , \RI3[1][96] , \RI3[1][95] ,
         \RI3[1][94] , \RI3[1][93] , \RI3[1][92] , \RI3[1][91] , \RI3[1][90] ,
         \RI3[1][89] , \RI3[1][88] , \RI3[1][87] , \RI3[1][86] , \RI3[1][85] ,
         \RI3[1][84] , \RI3[1][83] , \RI3[1][82] , \RI3[1][81] , \RI3[1][80] ,
         \RI3[1][79] , \RI3[1][78] , \RI3[1][77] , \RI3[1][76] , \RI3[1][75] ,
         \RI3[1][74] , \RI3[1][73] , \RI3[1][72] , \RI3[1][71] , \RI3[1][70] ,
         \RI3[1][69] , \RI3[1][68] , \RI3[1][67] , \RI3[1][66] , \RI3[1][65] ,
         \RI3[1][64] , \RI3[1][63] , \RI3[1][62] , \RI3[1][61] , \RI3[1][60] ,
         \RI3[1][59] , \RI3[1][58] , \RI3[1][57] , \RI3[1][56] , \RI3[1][55] ,
         \RI3[1][54] , \RI3[1][53] , \RI3[1][52] , \RI3[1][51] , \RI3[1][50] ,
         \RI3[1][49] , \RI3[1][48] , \RI3[1][47] , \RI3[1][46] , \RI3[1][45] ,
         \RI3[1][44] , \RI3[1][43] , \RI3[1][42] , \RI3[1][41] , \RI3[1][40] ,
         \RI3[1][39] , \RI3[1][38] , \RI3[1][37] , \RI3[1][36] , \RI3[1][35] ,
         \RI3[1][34] , \RI3[1][33] , \RI3[1][32] , \RI3[1][31] , \RI3[1][30] ,
         \RI3[1][29] , \RI3[1][28] , \RI3[1][27] , \RI3[1][26] , \RI3[1][25] ,
         \RI3[1][24] , \RI3[1][23] , \RI3[1][22] , \RI3[1][21] , \RI3[1][20] ,
         \RI3[1][19] , \RI3[1][18] , \RI3[1][17] , \RI3[1][16] , \RI3[1][15] ,
         \RI3[1][14] , \RI3[1][13] , \RI3[1][12] , \RI3[1][11] , \RI3[1][10] ,
         \RI3[1][9] , \RI3[1][8] , \RI3[1][7] , \RI3[1][6] , \RI3[1][5] ,
         \RI3[1][4] , \RI3[1][3] , \RI3[1][2] , \RI3[1][1] , \RI3[1][0] ,
         \RI3[2][191] , \RI3[2][190] , \RI3[2][189] , \RI3[2][188] ,
         \RI3[2][187] , \RI3[2][186] , \RI3[2][185] , \RI3[2][184] ,
         \RI3[2][183] , \RI3[2][182] , \RI3[2][181] , \RI3[2][180] ,
         \RI3[2][179] , \RI3[2][178] , \RI3[2][177] , \RI3[2][176] ,
         \RI3[2][175] , \RI3[2][174] , \RI3[2][173] , \RI3[2][172] ,
         \RI3[2][171] , \RI3[2][170] , \RI3[2][169] , \RI3[2][168] ,
         \RI3[2][167] , \RI3[2][166] , \RI3[2][165] , \RI3[2][164] ,
         \RI3[2][163] , \RI3[2][162] , \RI3[2][161] , \RI3[2][160] ,
         \RI3[2][159] , \RI3[2][158] , \RI3[2][157] , \RI3[2][156] ,
         \RI3[2][155] , \RI3[2][154] , \RI3[2][153] , \RI3[2][152] ,
         \RI3[2][151] , \RI3[2][150] , \RI3[2][149] , \RI3[2][148] ,
         \RI3[2][147] , \RI3[2][146] , \RI3[2][145] , \RI3[2][144] ,
         \RI3[2][143] , \RI3[2][142] , \RI3[2][141] , \RI3[2][140] ,
         \RI3[2][139] , \RI3[2][138] , \RI3[2][137] , \RI3[2][136] ,
         \RI3[2][135] , \RI3[2][134] , \RI3[2][133] , \RI3[2][132] ,
         \RI3[2][131] , \RI3[2][130] , \RI3[2][129] , \RI3[2][128] ,
         \RI3[2][127] , \RI3[2][126] , \RI3[2][125] , \RI3[2][124] ,
         \RI3[2][123] , \RI3[2][122] , \RI3[2][121] , \RI3[2][120] ,
         \RI3[2][119] , \RI3[2][118] , \RI3[2][117] , \RI3[2][116] ,
         \RI3[2][115] , \RI3[2][114] , \RI3[2][113] , \RI3[2][112] ,
         \RI3[2][111] , \RI3[2][110] , \RI3[2][109] , \RI3[2][108] ,
         \RI3[2][107] , \RI3[2][106] , \RI3[2][105] , \RI3[2][104] ,
         \RI3[2][103] , \RI3[2][102] , \RI3[2][101] , \RI3[2][100] ,
         \RI3[2][99] , \RI3[2][98] , \RI3[2][97] , \RI3[2][96] , \RI3[2][95] ,
         \RI3[2][94] , \RI3[2][93] , \RI3[2][92] , \RI3[2][91] , \RI3[2][90] ,
         \RI3[2][89] , \RI3[2][88] , \RI3[2][87] , \RI3[2][86] , \RI3[2][85] ,
         \RI3[2][84] , \RI3[2][83] , \RI3[2][82] , \RI3[2][81] , \RI3[2][80] ,
         \RI3[2][79] , \RI3[2][78] , \RI3[2][77] , \RI3[2][76] , \RI3[2][75] ,
         \RI3[2][74] , \RI3[2][73] , \RI3[2][72] , \RI3[2][71] , \RI3[2][70] ,
         \RI3[2][69] , \RI3[2][68] , \RI3[2][67] , \RI3[2][66] , \RI3[2][65] ,
         \RI3[2][64] , \RI3[2][63] , \RI3[2][62] , \RI3[2][61] , \RI3[2][60] ,
         \RI3[2][59] , \RI3[2][58] , \RI3[2][57] , \RI3[2][56] , \RI3[2][55] ,
         \RI3[2][54] , \RI3[2][53] , \RI3[2][52] , \RI3[2][51] , \RI3[2][50] ,
         \RI3[2][49] , \RI3[2][48] , \RI3[2][47] , \RI3[2][46] , \RI3[2][45] ,
         \RI3[2][44] , \RI3[2][43] , \RI3[2][42] , \RI3[2][41] , \RI3[2][40] ,
         \RI3[2][39] , \RI3[2][38] , \RI3[2][37] , \RI3[2][36] , \RI3[2][35] ,
         \RI3[2][34] , \RI3[2][33] , \RI3[2][32] , \RI3[2][31] , \RI3[2][30] ,
         \RI3[2][29] , \RI3[2][28] , \RI3[2][27] , \RI3[2][26] , \RI3[2][25] ,
         \RI3[2][24] , \RI3[2][23] , \RI3[2][22] , \RI3[2][21] , \RI3[2][20] ,
         \RI3[2][19] , \RI3[2][18] , \RI3[2][17] , \RI3[2][16] , \RI3[2][15] ,
         \RI3[2][14] , \RI3[2][13] , \RI3[2][12] , \RI3[2][11] , \RI3[2][10] ,
         \RI3[2][9] , \RI3[2][8] , \RI3[2][7] , \RI3[2][6] , \RI3[2][5] ,
         \RI3[2][4] , \RI3[2][3] , \RI3[2][2] , \RI3[2][1] , \RI3[2][0] ,
         \RI3[3][191] , \RI3[3][190] , \RI3[3][189] , \RI3[3][188] ,
         \RI3[3][187] , \RI3[3][186] , \RI3[3][185] , \RI3[3][184] ,
         \RI3[3][183] , \RI3[3][182] , \RI3[3][181] , \RI3[3][180] ,
         \RI3[3][179] , \RI3[3][178] , \RI3[3][177] , \RI3[3][176] ,
         \RI3[3][175] , \RI3[3][174] , \RI3[3][173] , \RI3[3][172] ,
         \RI3[3][171] , \RI3[3][170] , \RI3[3][169] , \RI3[3][168] ,
         \RI3[3][167] , \RI3[3][165] , \RI3[3][164] , \RI3[3][163] ,
         \RI3[3][162] , \RI3[3][161] , \RI3[3][159] , \RI3[3][158] ,
         \RI3[3][157] , \RI3[3][156] , \RI3[3][155] , \RI3[3][154] ,
         \RI3[3][153] , \RI3[3][152] , \RI3[3][151] , \RI3[3][150] ,
         \RI3[3][149] , \RI3[3][148] , \RI3[3][147] , \RI3[3][146] ,
         \RI3[3][145] , \RI3[3][144] , \RI3[3][143] , \RI3[3][141] ,
         \RI3[3][140] , \RI3[3][139] , \RI3[3][138] , \RI3[3][137] ,
         \RI3[3][136] , \RI3[3][135] , \RI3[3][134] , \RI3[3][133] ,
         \RI3[3][132] , \RI3[3][131] , \RI3[3][130] , \RI3[3][129] ,
         \RI3[3][128] , \RI3[3][127] , \RI3[3][126] , \RI3[3][125] ,
         \RI3[3][124] , \RI3[3][123] , \RI3[3][122] , \RI3[3][121] ,
         \RI3[3][120] , \RI3[3][119] , \RI3[3][118] , \RI3[3][117] ,
         \RI3[3][116] , \RI3[3][115] , \RI3[3][114] , \RI3[3][113] ,
         \RI3[3][111] , \RI3[3][110] , \RI3[3][109] , \RI3[3][108] ,
         \RI3[3][107] , \RI3[3][106] , \RI3[3][105] , \RI3[3][104] ,
         \RI3[3][103] , \RI3[3][102] , \RI3[3][101] , \RI3[3][99] ,
         \RI3[3][98] , \RI3[3][96] , \RI3[3][95] , \RI3[3][94] , \RI3[3][93] ,
         \RI3[3][92] , \RI3[3][91] , \RI3[3][90] , \RI3[3][89] , \RI3[3][88] ,
         \RI3[3][87] , \RI3[3][86] , \RI3[3][85] , \RI3[3][84] , \RI3[3][83] ,
         \RI3[3][81] , \RI3[3][80] , \RI3[3][79] , \RI3[3][78] , \RI3[3][77] ,
         \RI3[3][76] , \RI3[3][75] , \RI3[3][74] , \RI3[3][73] , \RI3[3][72] ,
         \RI3[3][71] , \RI3[3][69] , \RI3[3][68] , \RI3[3][67] , \RI3[3][66] ,
         \RI3[3][65] , \RI3[3][64] , \RI3[3][63] , \RI3[3][62] , \RI3[3][61] ,
         \RI3[3][60] , \RI3[3][59] , \RI3[3][57] , \RI3[3][56] , \RI3[3][55] ,
         \RI3[3][54] , \RI3[3][53] , \RI3[3][51] , \RI3[3][50] , \RI3[3][49] ,
         \RI3[3][48] , \RI3[3][47] , \RI3[3][46] , \RI3[3][45] , \RI3[3][44] ,
         \RI3[3][43] , \RI3[3][42] , \RI3[3][41] , \RI3[3][39] , \RI3[3][38] ,
         \RI3[3][37] , \RI3[3][36] , \RI3[3][35] , \RI3[3][33] , \RI3[3][32] ,
         \RI3[3][31] , \RI3[3][30] , \RI3[3][29] , \RI3[3][28] , \RI3[3][27] ,
         \RI3[3][26] , \RI3[3][25] , \RI3[3][24] , \RI3[3][23] , \RI3[3][21] ,
         \RI3[3][20] , \RI3[3][19] , \RI3[3][18] , \RI3[3][17] , \RI3[3][16] ,
         \RI3[3][15] , \RI3[3][14] , \RI3[3][13] , \RI3[3][12] , \RI3[3][11] ,
         \RI3[3][10] , \RI3[3][9] , \RI3[3][8] , \RI3[3][7] , \RI3[3][6] ,
         \RI3[3][5] , \RI3[3][3] , \RI3[3][2] , \RI3[3][1] , \RI3[3][0] ,
         \RI3[4][191] , \RI3[4][190] , \RI3[4][189] , \RI3[4][188] ,
         \RI3[4][187] , \RI3[4][186] , \RI3[4][185] , \RI3[4][184] ,
         \RI3[4][183] , \RI3[4][182] , \RI3[4][181] , \RI3[4][180] ,
         \RI3[4][179] , \RI3[4][178] , \RI3[4][177] , \RI3[4][176] ,
         \RI3[4][175] , \RI3[4][173] , \RI3[4][172] , \RI3[4][171] ,
         \RI3[4][170] , \RI3[4][169] , \RI3[4][168] , \RI3[4][167] ,
         \RI3[4][166] , \RI3[4][165] , \RI3[4][164] , \RI3[4][163] ,
         \RI3[4][162] , \RI3[4][161] , \RI3[4][159] , \RI3[4][158] ,
         \RI3[4][157] , \RI3[4][156] , \RI3[4][155] , \RI3[4][154] ,
         \RI3[4][153] , \RI3[4][152] , \RI3[4][151] , \RI3[4][150] ,
         \RI3[4][149] , \RI3[4][148] , \RI3[4][147] , \RI3[4][146] ,
         \RI3[4][145] , \RI3[4][144] , \RI3[4][143] , \RI3[4][141] ,
         \RI3[4][140] , \RI3[4][139] , \RI3[4][138] , \RI3[4][137] ,
         \RI3[4][136] , \RI3[4][135] , \RI3[4][134] , \RI3[4][133] ,
         \RI3[4][132] , \RI3[4][131] , \RI3[4][130] , \RI3[4][129] ,
         \RI3[4][128] , \RI3[4][127] , \RI3[4][126] , \RI3[4][125] ,
         \RI3[4][123] , \RI3[4][122] , \RI3[4][121] , \RI3[4][120] ,
         \RI3[4][119] , \RI3[4][118] , \RI3[4][117] , \RI3[4][116] ,
         \RI3[4][115] , \RI3[4][114] , \RI3[4][113] , \RI3[4][112] ,
         \RI3[4][111] , \RI3[4][110] , \RI3[4][109] , \RI3[4][108] ,
         \RI3[4][107] , \RI3[4][105] , \RI3[4][104] , \RI3[4][103] ,
         \RI3[4][102] , \RI3[4][101] , \RI3[4][100] , \RI3[4][99] ,
         \RI3[4][98] , \RI3[4][97] , \RI3[4][96] , \RI3[4][95] , \RI3[4][94] ,
         \RI3[4][93] , \RI3[4][92] , \RI3[4][91] , \RI3[4][90] , \RI3[4][89] ,
         \RI3[4][88] , \RI3[4][87] , \RI3[4][86] , \RI3[4][85] , \RI3[4][84] ,
         \RI3[4][83] , \RI3[4][82] , \RI3[4][81] , \RI3[4][80] , \RI3[4][79] ,
         \RI3[4][78] , \RI3[4][77] , \RI3[4][76] , \RI3[4][75] , \RI3[4][74] ,
         \RI3[4][73] , \RI3[4][72] , \RI3[4][71] , \RI3[4][69] , \RI3[4][68] ,
         \RI3[4][67] , \RI3[4][66] , \RI3[4][65] , \RI3[4][64] , \RI3[4][63] ,
         \RI3[4][62] , \RI3[4][61] , \RI3[4][60] , \RI3[4][59] , \RI3[4][58] ,
         \RI3[4][57] , \RI3[4][56] , \RI3[4][55] , \RI3[4][53] , \RI3[4][52] ,
         \RI3[4][51] , \RI3[4][50] , \RI3[4][49] , \RI3[4][48] , \RI3[4][47] ,
         \RI3[4][46] , \RI3[4][45] , \RI3[4][44] , \RI3[4][43] , \RI3[4][42] ,
         \RI3[4][41] , \RI3[4][40] , \RI3[4][39] , \RI3[4][38] , \RI3[4][37] ,
         \RI3[4][36] , \RI3[4][35] , \RI3[4][34] , \RI3[4][33] , \RI3[4][32] ,
         \RI3[4][31] , \RI3[4][30] , \RI3[4][29] , \RI3[4][27] , \RI3[4][26] ,
         \RI3[4][25] , \RI3[4][24] , \RI3[4][23] , \RI3[4][22] , \RI3[4][21] ,
         \RI3[4][20] , \RI3[4][19] , \RI3[4][18] , \RI3[4][17] , \RI3[4][15] ,
         \RI3[4][14] , \RI3[4][11] , \RI3[4][10] , \RI3[4][9] , \RI3[4][8] ,
         \RI3[4][7] , \RI3[4][6] , \RI3[4][4] , \RI3[4][3] , \RI3[4][2] ,
         \RI3[4][1] , \RI3[4][0] , \RI4[4][187] , \RI4[4][183] , \RI4[4][159] ,
         \RI4[4][141] , \RI4[4][105] , \RI4[4][81] , \RI4[4][75] ,
         \RI4[4][51] , \RI4[4][45] , \RI4[4][33] , \RI4[4][3] , \RI5[0][190] ,
         \RI5[0][187] , \RI5[0][186] , \RI5[0][184] , \RI5[0][181] ,
         \RI5[0][180] , \RI5[0][178] , \RI5[0][176] , \RI5[0][175] ,
         \RI5[0][174] , \RI5[0][172] , \RI5[0][171] , \RI5[0][170] ,
         \RI5[0][169] , \RI5[0][168] , \RI5[0][166] , \RI5[0][165] ,
         \RI5[0][163] , \RI5[0][162] , \RI5[0][160] , \RI5[0][157] ,
         \RI5[0][156] , \RI5[0][152] , \RI5[0][151] , \RI5[0][150] ,
         \RI5[0][148] , \RI5[0][144] , \RI5[0][142] , \RI5[0][139] ,
         \RI5[0][138] , \RI5[0][136] , \RI5[0][134] , \RI5[0][133] ,
         \RI5[0][132] , \RI5[0][130] , \RI5[0][129] , \RI5[0][128] ,
         \RI5[0][127] , \RI5[0][124] , \RI5[0][123] , \RI5[0][122] ,
         \RI5[0][121] , \RI5[0][120] , \RI5[0][118] , \RI5[0][115] ,
         \RI5[0][114] , \RI5[0][112] , \RI5[0][109] , \RI5[0][108] ,
         \RI5[0][106] , \RI5[0][104] , \RI5[0][103] , \RI5[0][102] ,
         \RI5[0][99] , \RI5[0][98] , \RI5[0][97] , \RI5[0][96] , \RI5[0][94] ,
         \RI5[0][93] , \RI5[0][92] , \RI5[0][91] , \RI5[0][90] , \RI5[0][88] ,
         \RI5[0][87] , \RI5[0][84] , \RI5[0][82] , \RI5[0][80] , \RI5[0][79] ,
         \RI5[0][76] , \RI5[0][73] , \RI5[0][72] , \RI5[0][68] , \RI5[0][67] ,
         \RI5[0][66] , \RI5[0][64] , \RI5[0][63] , \RI5[0][62] , \RI5[0][61] ,
         \RI5[0][60] , \RI5[0][58] , \RI5[0][55] , \RI5[0][54] , \RI5[0][52] ,
         \RI5[0][49] , \RI5[0][48] , \RI5[0][46] , \RI5[0][45] , \RI5[0][43] ,
         \RI5[0][42] , \RI5[0][38] , \RI5[0][37] , \RI5[0][36] , \RI5[0][33] ,
         \RI5[0][32] , \RI5[0][31] , \RI5[0][30] , \RI5[0][28] , \RI5[0][27] ,
         \RI5[0][25] , \RI5[0][24] , \RI5[0][22] , \RI5[0][19] , \RI5[0][18] ,
         \RI5[0][14] , \RI5[0][13] , \RI5[0][12] , \RI5[0][9] , \RI5[0][8] ,
         \RI5[0][7] , \RI5[0][4] , \RI5[0][3] , \RI5[0][2] , \RI5[0][1] ,
         \RI5[0][0] , \RI5[1][190] , \RI5[1][189] , \RI5[1][187] ,
         \RI5[1][186] , \RI5[1][184] , \RI5[1][183] , \RI5[1][182] ,
         \RI5[1][181] , \RI5[1][180] , \RI5[1][179] , \RI5[1][177] ,
         \RI5[1][175] , \RI5[1][172] , \RI5[1][171] , \RI5[1][170] ,
         \RI5[1][169] , \RI5[1][168] , \RI5[1][166] , \RI5[1][165] ,
         \RI5[1][163] , \RI5[1][162] , \RI5[1][160] , \RI5[1][158] ,
         \RI5[1][157] , \RI5[1][156] , \RI5[1][152] , \RI5[1][151] ,
         \RI5[1][150] , \RI5[1][147] , \RI5[1][145] , \RI5[1][144] ,
         \RI5[1][142] , \RI5[1][141] , \RI5[1][140] , \RI5[1][139] ,
         \RI5[1][138] , \RI5[1][136] , \RI5[1][135] , \RI5[1][134] ,
         \RI5[1][133] , \RI5[1][132] , \RI5[1][130] , \RI5[1][129] ,
         \RI5[1][128] , \RI5[1][127] , \RI5[1][126] , \RI5[1][124] ,
         \RI5[1][123] , \RI5[1][122] , \RI5[1][121] , \RI5[1][120] ,
         \RI5[1][118] , \RI5[1][117] , \RI5[1][115] , \RI5[1][114] ,
         \RI5[1][112] , \RI5[1][111] , \RI5[1][109] , \RI5[1][108] ,
         \RI5[1][106] , \RI5[1][104] , \RI5[1][103] , \RI5[1][102] ,
         \RI5[1][100] , \RI5[1][97] , \RI5[1][96] , \RI5[1][94] , \RI5[1][93] ,
         \RI5[1][91] , \RI5[1][90] , \RI5[1][89] , \RI5[1][88] , \RI5[1][87] ,
         \RI5[1][86] , \RI5[1][85] , \RI5[1][84] , \RI5[1][81] , \RI5[1][79] ,
         \RI5[1][78] , \RI5[1][76] , \RI5[1][75] , \RI5[1][74] , \RI5[1][73] ,
         \RI5[1][72] , \RI5[1][70] , \RI5[1][68] , \RI5[1][67] , \RI5[1][66] ,
         \RI5[1][64] , \RI5[1][63] , \RI5[1][62] , \RI5[1][61] , \RI5[1][60] ,
         \RI5[1][58] , \RI5[1][57] , \RI5[1][56] , \RI5[1][55] , \RI5[1][54] ,
         \RI5[1][52] , \RI5[1][51] , \RI5[1][49] , \RI5[1][48] , \RI5[1][46] ,
         \RI5[1][45] , \RI5[1][44] , \RI5[1][43] , \RI5[1][42] , \RI5[1][40] ,
         \RI5[1][39] , \RI5[1][38] , \RI5[1][37] , \RI5[1][36] , \RI5[1][34] ,
         \RI5[1][33] , \RI5[1][32] , \RI5[1][31] , \RI5[1][30] , \RI5[1][28] ,
         \RI5[1][26] , \RI5[1][25] , \RI5[1][24] , \RI5[1][22] , \RI5[1][21] ,
         \RI5[1][19] , \RI5[1][18] , \RI5[1][16] , \RI5[1][14] , \RI5[1][13] ,
         \RI5[1][12] , \RI5[1][10] , \RI5[1][9] , \RI5[1][7] , \RI5[1][6] ,
         \RI5[1][4] , \RI5[1][3] , \RI5[1][2] , \RI5[1][1] , \RI5[1][0] ,
         \RI5[2][190] , \RI5[2][188] , \RI5[2][187] , \RI5[2][186] ,
         \RI5[2][183] , \RI5[2][182] , \RI5[2][181] , \RI5[2][180] ,
         \RI5[2][178] , \RI5[2][177] , \RI5[2][175] , \RI5[2][174] ,
         \RI5[2][172] , \RI5[2][171] , \RI5[2][170] , \RI5[2][169] ,
         \RI5[2][168] , \RI5[2][166] , \RI5[2][165] , \RI5[2][164] ,
         \RI5[2][163] , \RI5[2][162] , \RI5[2][160] , \RI5[2][159] ,
         \RI5[2][158] , \RI5[2][157] , \RI5[2][156] , \RI5[2][154] ,
         \RI5[2][152] , \RI5[2][151] , \RI5[2][150] , \RI5[2][148] ,
         \RI5[2][147] , \RI5[2][146] , \RI5[2][145] , \RI5[2][144] ,
         \RI5[2][142] , \RI5[2][141] , \RI5[2][140] , \RI5[2][139] ,
         \RI5[2][138] , \RI5[2][135] , \RI5[2][134] , \RI5[2][133] ,
         \RI5[2][132] , \RI5[2][130] , \RI5[2][129] , \RI5[2][128] ,
         \RI5[2][127] , \RI5[2][126] , \RI5[2][124] , \RI5[2][123] ,
         \RI5[2][122] , \RI5[2][121] , \RI5[2][120] , \RI5[2][117] ,
         \RI5[2][116] , \RI5[2][115] , \RI5[2][114] , \RI5[2][112] ,
         \RI5[2][111] , \RI5[2][110] , \RI5[2][109] , \RI5[2][108] ,
         \RI5[2][106] , \RI5[2][105] , \RI5[2][103] , \RI5[2][102] ,
         \RI5[2][100] , \RI5[2][99] , \RI5[2][98] , \RI5[2][97] , \RI5[2][96] ,
         \RI5[2][94] , \RI5[2][93] , \RI5[2][92] , \RI5[2][91] , \RI5[2][90] ,
         \RI5[2][88] , \RI5[2][87] , \RI5[2][86] , \RI5[2][85] , \RI5[2][84] ,
         \RI5[2][82] , \RI5[2][81] , \RI5[2][79] , \RI5[2][78] , \RI5[2][76] ,
         \RI5[2][75] , \RI5[2][74] , \RI5[2][73] , \RI5[2][72] , \RI5[2][70] ,
         \RI5[2][69] , \RI5[2][67] , \RI5[2][66] , \RI5[2][64] , \RI5[2][62] ,
         \RI5[2][61] , \RI5[2][60] , \RI5[2][56] , \RI5[2][55] , \RI5[2][54] ,
         \RI5[2][52] , \RI5[2][51] , \RI5[2][50] , \RI5[2][49] , \RI5[2][48] ,
         \RI5[2][46] , \RI5[2][45] , \RI5[2][44] , \RI5[2][43] , \RI5[2][42] ,
         \RI5[2][40] , \RI5[2][39] , \RI5[2][37] , \RI5[2][36] , \RI5[2][34] ,
         \RI5[2][33] , \RI5[2][32] , \RI5[2][30] , \RI5[2][26] , \RI5[2][25] ,
         \RI5[2][24] , \RI5[2][22] , \RI5[2][21] , \RI5[2][19] , \RI5[2][18] ,
         \RI5[2][16] , \RI5[2][14] , \RI5[2][13] , \RI5[2][12] , \RI5[2][10] ,
         \RI5[2][9] , \RI5[2][7] , \RI5[2][6] , \RI5[2][4] , \RI5[2][3] ,
         \RI5[2][2] , \RI5[2][1] , \RI5[2][0] , \RI5[3][190] , \RI5[3][189] ,
         \RI5[3][188] , \RI5[3][187] , \RI5[3][186] , \RI5[3][185] ,
         \RI5[3][184] , \RI5[3][181] , \RI5[3][180] , \RI5[3][177] ,
         \RI5[3][175] , \RI5[3][174] , \RI5[3][172] , \RI5[3][171] ,
         \RI5[3][170] , \RI5[3][169] , \RI5[3][168] , \RI5[3][165] ,
         \RI5[3][164] , \RI5[3][163] , \RI5[3][162] , \RI5[3][160] ,
         \RI5[3][159] , \RI5[3][158] , \RI5[3][157] , \RI5[3][156] ,
         \RI5[3][154] , \RI5[3][153] , \RI5[3][152] , \RI5[3][151] ,
         \RI5[3][150] , \RI5[3][149] , \RI5[3][148] , \RI5[3][147] ,
         \RI5[3][145] , \RI5[3][144] , \RI5[3][141] , \RI5[3][140] ,
         \RI5[3][139] , \RI5[3][138] , \RI5[3][136] , \RI5[3][135] ,
         \RI5[3][134] , \RI5[3][133] , \RI5[3][132] , \RI5[3][131] ,
         \RI5[3][130] , \RI5[3][129] , \RI5[3][127] , \RI5[3][126] ,
         \RI5[3][123] , \RI5[3][121] , \RI5[3][120] , \RI5[3][118] ,
         \RI5[3][117] , \RI5[3][116] , \RI5[3][115] , \RI5[3][114] ,
         \RI5[3][113] , \RI5[3][111] , \RI5[3][109] , \RI5[3][108] ,
         \RI5[3][106] , \RI5[3][105] , \RI5[3][103] , \RI5[3][102] ,
         \RI5[3][101] , \RI5[3][99] , \RI5[3][98] , \RI5[3][97] , \RI5[3][96] ,
         \RI5[3][94] , \RI5[3][93] , \RI5[3][92] , \RI5[3][90] , \RI5[3][89] ,
         \RI5[3][88] , \RI5[3][87] , \RI5[3][86] , \RI5[3][85] , \RI5[3][84] ,
         \RI5[3][82] , \RI5[3][81] , \RI5[3][80] , \RI5[3][79] , \RI5[3][78] ,
         \RI5[3][76] , \RI5[3][75] , \RI5[3][73] , \RI5[3][72] , \RI5[3][71] ,
         \RI5[3][69] , \RI5[3][68] , \RI5[3][67] , \RI5[3][66] , \RI5[3][64] ,
         \RI5[3][63] , \RI5[3][61] , \RI5[3][60] , \RI5[3][58] , \RI5[3][57] ,
         \RI5[3][56] , \RI5[3][55] , \RI5[3][54] , \RI5[3][51] , \RI5[3][50] ,
         \RI5[3][49] , \RI5[3][48] , \RI5[3][47] , \RI5[3][46] , \RI5[3][45] ,
         \RI5[3][44] , \RI5[3][43] , \RI5[3][42] , \RI5[3][41] , \RI5[3][40] ,
         \RI5[3][39] , \RI5[3][38] , \RI5[3][37] , \RI5[3][36] , \RI5[3][33] ,
         \RI5[3][31] , \RI5[3][30] , \RI5[3][28] , \RI5[3][27] , \RI5[3][26] ,
         \RI5[3][25] , \RI5[3][24] , \RI5[3][23] , \RI5[3][21] , \RI5[3][19] ,
         \RI5[3][18] , \RI5[3][17] , \RI5[3][16] , \RI5[3][15] , \RI5[3][14] ,
         \RI5[3][13] , \RI5[3][12] , \RI5[3][11] , \RI5[3][9] , \RI5[3][8] ,
         \RI5[3][7] , \RI5[3][6] , \RI5[3][5] , \RI5[3][3] , \RI5[3][2] ,
         \RI5[3][1] , \RI5[3][0] , \MC_ARK_ARC_1_0/temp6[190] ,
         \MC_ARK_ARC_1_0/temp6[188] , \MC_ARK_ARC_1_0/temp6[187] ,
         \MC_ARK_ARC_1_0/temp6[186] , \MC_ARK_ARC_1_0/temp6[184] ,
         \MC_ARK_ARC_1_0/temp6[183] , \MC_ARK_ARC_1_0/temp6[182] ,
         \MC_ARK_ARC_1_0/temp6[181] , \MC_ARK_ARC_1_0/temp6[180] ,
         \MC_ARK_ARC_1_0/temp6[178] , \MC_ARK_ARC_1_0/temp6[176] ,
         \MC_ARK_ARC_1_0/temp6[175] , \MC_ARK_ARC_1_0/temp6[174] ,
         \MC_ARK_ARC_1_0/temp6[172] , \MC_ARK_ARC_1_0/temp6[171] ,
         \MC_ARK_ARC_1_0/temp6[170] , \MC_ARK_ARC_1_0/temp6[169] ,
         \MC_ARK_ARC_1_0/temp6[168] , \MC_ARK_ARC_1_0/temp6[166] ,
         \MC_ARK_ARC_1_0/temp6[165] , \MC_ARK_ARC_1_0/temp6[164] ,
         \MC_ARK_ARC_1_0/temp6[163] , \MC_ARK_ARC_1_0/temp6[162] ,
         \MC_ARK_ARC_1_0/temp6[160] , \MC_ARK_ARC_1_0/temp6[159] ,
         \MC_ARK_ARC_1_0/temp6[157] , \MC_ARK_ARC_1_0/temp6[156] ,
         \MC_ARK_ARC_1_0/temp6[155] , \MC_ARK_ARC_1_0/temp6[154] ,
         \MC_ARK_ARC_1_0/temp6[153] , \MC_ARK_ARC_1_0/temp6[152] ,
         \MC_ARK_ARC_1_0/temp6[151] , \MC_ARK_ARC_1_0/temp6[150] ,
         \MC_ARK_ARC_1_0/temp6[148] , \MC_ARK_ARC_1_0/temp6[147] ,
         \MC_ARK_ARC_1_0/temp6[145] , \MC_ARK_ARC_1_0/temp6[144] ,
         \MC_ARK_ARC_1_0/temp6[143] , \MC_ARK_ARC_1_0/temp6[142] ,
         \MC_ARK_ARC_1_0/temp6[141] , \MC_ARK_ARC_1_0/temp6[140] ,
         \MC_ARK_ARC_1_0/temp6[139] , \MC_ARK_ARC_1_0/temp6[138] ,
         \MC_ARK_ARC_1_0/temp6[137] , \MC_ARK_ARC_1_0/temp6[136] ,
         \MC_ARK_ARC_1_0/temp6[135] , \MC_ARK_ARC_1_0/temp6[134] ,
         \MC_ARK_ARC_1_0/temp6[133] , \MC_ARK_ARC_1_0/temp6[132] ,
         \MC_ARK_ARC_1_0/temp6[131] , \MC_ARK_ARC_1_0/temp6[130] ,
         \MC_ARK_ARC_1_0/temp6[129] , \MC_ARK_ARC_1_0/temp6[128] ,
         \MC_ARK_ARC_1_0/temp6[127] , \MC_ARK_ARC_1_0/temp6[126] ,
         \MC_ARK_ARC_1_0/temp6[124] , \MC_ARK_ARC_1_0/temp6[123] ,
         \MC_ARK_ARC_1_0/temp6[122] , \MC_ARK_ARC_1_0/temp6[121] ,
         \MC_ARK_ARC_1_0/temp6[120] , \MC_ARK_ARC_1_0/temp6[118] ,
         \MC_ARK_ARC_1_0/temp6[117] , \MC_ARK_ARC_1_0/temp6[116] ,
         \MC_ARK_ARC_1_0/temp6[115] , \MC_ARK_ARC_1_0/temp6[114] ,
         \MC_ARK_ARC_1_0/temp6[112] , \MC_ARK_ARC_1_0/temp6[111] ,
         \MC_ARK_ARC_1_0/temp6[110] , \MC_ARK_ARC_1_0/temp6[109] ,
         \MC_ARK_ARC_1_0/temp6[108] , \MC_ARK_ARC_1_0/temp6[107] ,
         \MC_ARK_ARC_1_0/temp6[106] , \MC_ARK_ARC_1_0/temp6[105] ,
         \MC_ARK_ARC_1_0/temp6[104] , \MC_ARK_ARC_1_0/temp6[103] ,
         \MC_ARK_ARC_1_0/temp6[102] , \MC_ARK_ARC_1_0/temp6[101] ,
         \MC_ARK_ARC_1_0/temp6[100] , \MC_ARK_ARC_1_0/temp6[99] ,
         \MC_ARK_ARC_1_0/temp6[98] , \MC_ARK_ARC_1_0/temp6[97] ,
         \MC_ARK_ARC_1_0/temp6[96] , \MC_ARK_ARC_1_0/temp6[94] ,
         \MC_ARK_ARC_1_0/temp6[93] , \MC_ARK_ARC_1_0/temp6[92] ,
         \MC_ARK_ARC_1_0/temp6[91] , \MC_ARK_ARC_1_0/temp6[90] ,
         \MC_ARK_ARC_1_0/temp6[88] , \MC_ARK_ARC_1_0/temp6[87] ,
         \MC_ARK_ARC_1_0/temp6[86] , \MC_ARK_ARC_1_0/temp6[85] ,
         \MC_ARK_ARC_1_0/temp6[84] , \MC_ARK_ARC_1_0/temp6[82] ,
         \MC_ARK_ARC_1_0/temp6[81] , \MC_ARK_ARC_1_0/temp6[80] ,
         \MC_ARK_ARC_1_0/temp6[79] , \MC_ARK_ARC_1_0/temp6[78] ,
         \MC_ARK_ARC_1_0/temp6[76] , \MC_ARK_ARC_1_0/temp6[75] ,
         \MC_ARK_ARC_1_0/temp6[73] , \MC_ARK_ARC_1_0/temp6[72] ,
         \MC_ARK_ARC_1_0/temp6[70] , \MC_ARK_ARC_1_0/temp6[69] ,
         \MC_ARK_ARC_1_0/temp6[68] , \MC_ARK_ARC_1_0/temp6[67] ,
         \MC_ARK_ARC_1_0/temp6[66] , \MC_ARK_ARC_1_0/temp6[65] ,
         \MC_ARK_ARC_1_0/temp6[64] , \MC_ARK_ARC_1_0/temp6[63] ,
         \MC_ARK_ARC_1_0/temp6[62] , \MC_ARK_ARC_1_0/temp6[61] ,
         \MC_ARK_ARC_1_0/temp6[60] , \MC_ARK_ARC_1_0/temp6[58] ,
         \MC_ARK_ARC_1_0/temp6[57] , \MC_ARK_ARC_1_0/temp6[56] ,
         \MC_ARK_ARC_1_0/temp6[55] , \MC_ARK_ARC_1_0/temp6[54] ,
         \MC_ARK_ARC_1_0/temp6[52] , \MC_ARK_ARC_1_0/temp6[51] ,
         \MC_ARK_ARC_1_0/temp6[50] , \MC_ARK_ARC_1_0/temp6[49] ,
         \MC_ARK_ARC_1_0/temp6[48] , \MC_ARK_ARC_1_0/temp6[46] ,
         \MC_ARK_ARC_1_0/temp6[45] , \MC_ARK_ARC_1_0/temp6[43] ,
         \MC_ARK_ARC_1_0/temp6[42] , \MC_ARK_ARC_1_0/temp6[40] ,
         \MC_ARK_ARC_1_0/temp6[39] , \MC_ARK_ARC_1_0/temp6[37] ,
         \MC_ARK_ARC_1_0/temp6[36] , \MC_ARK_ARC_1_0/temp6[34] ,
         \MC_ARK_ARC_1_0/temp6[33] , \MC_ARK_ARC_1_0/temp6[32] ,
         \MC_ARK_ARC_1_0/temp6[31] , \MC_ARK_ARC_1_0/temp6[30] ,
         \MC_ARK_ARC_1_0/temp6[29] , \MC_ARK_ARC_1_0/temp6[28] ,
         \MC_ARK_ARC_1_0/temp6[26] , \MC_ARK_ARC_1_0/temp6[25] ,
         \MC_ARK_ARC_1_0/temp6[24] , \MC_ARK_ARC_1_0/temp6[22] ,
         \MC_ARK_ARC_1_0/temp6[21] , \MC_ARK_ARC_1_0/temp6[20] ,
         \MC_ARK_ARC_1_0/temp6[19] , \MC_ARK_ARC_1_0/temp6[18] ,
         \MC_ARK_ARC_1_0/temp6[16] , \MC_ARK_ARC_1_0/temp6[15] ,
         \MC_ARK_ARC_1_0/temp6[14] , \MC_ARK_ARC_1_0/temp6[13] ,
         \MC_ARK_ARC_1_0/temp6[12] , \MC_ARK_ARC_1_0/temp6[10] ,
         \MC_ARK_ARC_1_0/temp6[9] , \MC_ARK_ARC_1_0/temp6[8] ,
         \MC_ARK_ARC_1_0/temp6[7] , \MC_ARK_ARC_1_0/temp6[6] ,
         \MC_ARK_ARC_1_0/temp6[4] , \MC_ARK_ARC_1_0/temp6[3] ,
         \MC_ARK_ARC_1_0/temp6[2] , \MC_ARK_ARC_1_0/temp6[1] ,
         \MC_ARK_ARC_1_0/temp6[0] , \MC_ARK_ARC_1_0/temp5[190] ,
         \MC_ARK_ARC_1_0/temp5[188] , \MC_ARK_ARC_1_0/temp5[187] ,
         \MC_ARK_ARC_1_0/temp5[186] , \MC_ARK_ARC_1_0/temp5[185] ,
         \MC_ARK_ARC_1_0/temp5[184] , \MC_ARK_ARC_1_0/temp5[183] ,
         \MC_ARK_ARC_1_0/temp5[182] , \MC_ARK_ARC_1_0/temp5[181] ,
         \MC_ARK_ARC_1_0/temp5[180] , \MC_ARK_ARC_1_0/temp5[179] ,
         \MC_ARK_ARC_1_0/temp5[178] , \MC_ARK_ARC_1_0/temp5[177] ,
         \MC_ARK_ARC_1_0/temp5[176] , \MC_ARK_ARC_1_0/temp5[175] ,
         \MC_ARK_ARC_1_0/temp5[174] , \MC_ARK_ARC_1_0/temp5[173] ,
         \MC_ARK_ARC_1_0/temp5[172] , \MC_ARK_ARC_1_0/temp5[171] ,
         \MC_ARK_ARC_1_0/temp5[170] , \MC_ARK_ARC_1_0/temp5[169] ,
         \MC_ARK_ARC_1_0/temp5[168] , \MC_ARK_ARC_1_0/temp5[166] ,
         \MC_ARK_ARC_1_0/temp5[165] , \MC_ARK_ARC_1_0/temp5[164] ,
         \MC_ARK_ARC_1_0/temp5[163] , \MC_ARK_ARC_1_0/temp5[162] ,
         \MC_ARK_ARC_1_0/temp5[160] , \MC_ARK_ARC_1_0/temp5[159] ,
         \MC_ARK_ARC_1_0/temp5[158] , \MC_ARK_ARC_1_0/temp5[157] ,
         \MC_ARK_ARC_1_0/temp5[156] , \MC_ARK_ARC_1_0/temp5[155] ,
         \MC_ARK_ARC_1_0/temp5[154] , \MC_ARK_ARC_1_0/temp5[153] ,
         \MC_ARK_ARC_1_0/temp5[151] , \MC_ARK_ARC_1_0/temp5[150] ,
         \MC_ARK_ARC_1_0/temp5[149] , \MC_ARK_ARC_1_0/temp5[148] ,
         \MC_ARK_ARC_1_0/temp5[147] , \MC_ARK_ARC_1_0/temp5[145] ,
         \MC_ARK_ARC_1_0/temp5[144] , \MC_ARK_ARC_1_0/temp5[143] ,
         \MC_ARK_ARC_1_0/temp5[142] , \MC_ARK_ARC_1_0/temp5[141] ,
         \MC_ARK_ARC_1_0/temp5[140] , \MC_ARK_ARC_1_0/temp5[139] ,
         \MC_ARK_ARC_1_0/temp5[138] , \MC_ARK_ARC_1_0/temp5[137] ,
         \MC_ARK_ARC_1_0/temp5[136] , \MC_ARK_ARC_1_0/temp5[135] ,
         \MC_ARK_ARC_1_0/temp5[134] , \MC_ARK_ARC_1_0/temp5[133] ,
         \MC_ARK_ARC_1_0/temp5[132] , \MC_ARK_ARC_1_0/temp5[131] ,
         \MC_ARK_ARC_1_0/temp5[130] , \MC_ARK_ARC_1_0/temp5[129] ,
         \MC_ARK_ARC_1_0/temp5[128] , \MC_ARK_ARC_1_0/temp5[127] ,
         \MC_ARK_ARC_1_0/temp5[126] , \MC_ARK_ARC_1_0/temp5[125] ,
         \MC_ARK_ARC_1_0/temp5[124] , \MC_ARK_ARC_1_0/temp5[123] ,
         \MC_ARK_ARC_1_0/temp5[122] , \MC_ARK_ARC_1_0/temp5[121] ,
         \MC_ARK_ARC_1_0/temp5[120] , \MC_ARK_ARC_1_0/temp5[119] ,
         \MC_ARK_ARC_1_0/temp5[116] , \MC_ARK_ARC_1_0/temp5[115] ,
         \MC_ARK_ARC_1_0/temp5[114] , \MC_ARK_ARC_1_0/temp5[112] ,
         \MC_ARK_ARC_1_0/temp5[111] , \MC_ARK_ARC_1_0/temp5[110] ,
         \MC_ARK_ARC_1_0/temp5[109] , \MC_ARK_ARC_1_0/temp5[108] ,
         \MC_ARK_ARC_1_0/temp5[107] , \MC_ARK_ARC_1_0/temp5[106] ,
         \MC_ARK_ARC_1_0/temp5[105] , \MC_ARK_ARC_1_0/temp5[104] ,
         \MC_ARK_ARC_1_0/temp5[103] , \MC_ARK_ARC_1_0/temp5[102] ,
         \MC_ARK_ARC_1_0/temp5[101] , \MC_ARK_ARC_1_0/temp5[100] ,
         \MC_ARK_ARC_1_0/temp5[99] , \MC_ARK_ARC_1_0/temp5[98] ,
         \MC_ARK_ARC_1_0/temp5[97] , \MC_ARK_ARC_1_0/temp5[96] ,
         \MC_ARK_ARC_1_0/temp5[94] , \MC_ARK_ARC_1_0/temp5[93] ,
         \MC_ARK_ARC_1_0/temp5[92] , \MC_ARK_ARC_1_0/temp5[91] ,
         \MC_ARK_ARC_1_0/temp5[90] , \MC_ARK_ARC_1_0/temp5[88] ,
         \MC_ARK_ARC_1_0/temp5[87] , \MC_ARK_ARC_1_0/temp5[86] ,
         \MC_ARK_ARC_1_0/temp5[85] , \MC_ARK_ARC_1_0/temp5[84] ,
         \MC_ARK_ARC_1_0/temp5[82] , \MC_ARK_ARC_1_0/temp5[81] ,
         \MC_ARK_ARC_1_0/temp5[80] , \MC_ARK_ARC_1_0/temp5[79] ,
         \MC_ARK_ARC_1_0/temp5[78] , \MC_ARK_ARC_1_0/temp5[76] ,
         \MC_ARK_ARC_1_0/temp5[75] , \MC_ARK_ARC_1_0/temp5[73] ,
         \MC_ARK_ARC_1_0/temp5[72] , \MC_ARK_ARC_1_0/temp5[70] ,
         \MC_ARK_ARC_1_0/temp5[69] , \MC_ARK_ARC_1_0/temp5[68] ,
         \MC_ARK_ARC_1_0/temp5[67] , \MC_ARK_ARC_1_0/temp5[66] ,
         \MC_ARK_ARC_1_0/temp5[65] , \MC_ARK_ARC_1_0/temp5[64] ,
         \MC_ARK_ARC_1_0/temp5[63] , \MC_ARK_ARC_1_0/temp5[62] ,
         \MC_ARK_ARC_1_0/temp5[61] , \MC_ARK_ARC_1_0/temp5[60] ,
         \MC_ARK_ARC_1_0/temp5[58] , \MC_ARK_ARC_1_0/temp5[57] ,
         \MC_ARK_ARC_1_0/temp5[56] , \MC_ARK_ARC_1_0/temp5[55] ,
         \MC_ARK_ARC_1_0/temp5[54] , \MC_ARK_ARC_1_0/temp5[52] ,
         \MC_ARK_ARC_1_0/temp5[51] , \MC_ARK_ARC_1_0/temp5[50] ,
         \MC_ARK_ARC_1_0/temp5[49] , \MC_ARK_ARC_1_0/temp5[48] ,
         \MC_ARK_ARC_1_0/temp5[46] , \MC_ARK_ARC_1_0/temp5[45] ,
         \MC_ARK_ARC_1_0/temp5[43] , \MC_ARK_ARC_1_0/temp5[42] ,
         \MC_ARK_ARC_1_0/temp5[40] , \MC_ARK_ARC_1_0/temp5[39] ,
         \MC_ARK_ARC_1_0/temp5[37] , \MC_ARK_ARC_1_0/temp5[36] ,
         \MC_ARK_ARC_1_0/temp5[34] , \MC_ARK_ARC_1_0/temp5[33] ,
         \MC_ARK_ARC_1_0/temp5[32] , \MC_ARK_ARC_1_0/temp5[31] ,
         \MC_ARK_ARC_1_0/temp5[30] , \MC_ARK_ARC_1_0/temp5[29] ,
         \MC_ARK_ARC_1_0/temp5[28] , \MC_ARK_ARC_1_0/temp5[26] ,
         \MC_ARK_ARC_1_0/temp5[25] , \MC_ARK_ARC_1_0/temp5[24] ,
         \MC_ARK_ARC_1_0/temp5[22] , \MC_ARK_ARC_1_0/temp5[21] ,
         \MC_ARK_ARC_1_0/temp5[20] , \MC_ARK_ARC_1_0/temp5[19] ,
         \MC_ARK_ARC_1_0/temp5[18] , \MC_ARK_ARC_1_0/temp5[16] ,
         \MC_ARK_ARC_1_0/temp5[15] , \MC_ARK_ARC_1_0/temp5[14] ,
         \MC_ARK_ARC_1_0/temp5[13] , \MC_ARK_ARC_1_0/temp5[12] ,
         \MC_ARK_ARC_1_0/temp5[10] , \MC_ARK_ARC_1_0/temp5[9] ,
         \MC_ARK_ARC_1_0/temp5[8] , \MC_ARK_ARC_1_0/temp5[7] ,
         \MC_ARK_ARC_1_0/temp5[6] , \MC_ARK_ARC_1_0/temp5[4] ,
         \MC_ARK_ARC_1_0/temp5[3] , \MC_ARK_ARC_1_0/temp5[2] ,
         \MC_ARK_ARC_1_0/temp5[1] , \MC_ARK_ARC_1_0/temp5[0] ,
         \MC_ARK_ARC_1_0/temp4[191] , \MC_ARK_ARC_1_0/temp4[190] ,
         \MC_ARK_ARC_1_0/temp4[189] , \MC_ARK_ARC_1_0/temp4[188] ,
         \MC_ARK_ARC_1_0/temp4[187] , \MC_ARK_ARC_1_0/temp4[186] ,
         \MC_ARK_ARC_1_0/temp4[185] , \MC_ARK_ARC_1_0/temp4[184] ,
         \MC_ARK_ARC_1_0/temp4[183] , \MC_ARK_ARC_1_0/temp4[182] ,
         \MC_ARK_ARC_1_0/temp4[181] , \MC_ARK_ARC_1_0/temp4[180] ,
         \MC_ARK_ARC_1_0/temp4[179] , \MC_ARK_ARC_1_0/temp4[178] ,
         \MC_ARK_ARC_1_0/temp4[177] , \MC_ARK_ARC_1_0/temp4[176] ,
         \MC_ARK_ARC_1_0/temp4[175] , \MC_ARK_ARC_1_0/temp4[174] ,
         \MC_ARK_ARC_1_0/temp4[173] , \MC_ARK_ARC_1_0/temp4[172] ,
         \MC_ARK_ARC_1_0/temp4[171] , \MC_ARK_ARC_1_0/temp4[170] ,
         \MC_ARK_ARC_1_0/temp4[169] , \MC_ARK_ARC_1_0/temp4[168] ,
         \MC_ARK_ARC_1_0/temp4[167] , \MC_ARK_ARC_1_0/temp4[166] ,
         \MC_ARK_ARC_1_0/temp4[165] , \MC_ARK_ARC_1_0/temp4[164] ,
         \MC_ARK_ARC_1_0/temp4[163] , \MC_ARK_ARC_1_0/temp4[162] ,
         \MC_ARK_ARC_1_0/temp4[161] , \MC_ARK_ARC_1_0/temp4[160] ,
         \MC_ARK_ARC_1_0/temp4[159] , \MC_ARK_ARC_1_0/temp4[158] ,
         \MC_ARK_ARC_1_0/temp4[157] , \MC_ARK_ARC_1_0/temp4[156] ,
         \MC_ARK_ARC_1_0/temp4[155] , \MC_ARK_ARC_1_0/temp4[154] ,
         \MC_ARK_ARC_1_0/temp4[153] , \MC_ARK_ARC_1_0/temp4[152] ,
         \MC_ARK_ARC_1_0/temp4[151] , \MC_ARK_ARC_1_0/temp4[150] ,
         \MC_ARK_ARC_1_0/temp4[149] , \MC_ARK_ARC_1_0/temp4[148] ,
         \MC_ARK_ARC_1_0/temp4[147] , \MC_ARK_ARC_1_0/temp4[146] ,
         \MC_ARK_ARC_1_0/temp4[145] , \MC_ARK_ARC_1_0/temp4[144] ,
         \MC_ARK_ARC_1_0/temp4[143] , \MC_ARK_ARC_1_0/temp4[142] ,
         \MC_ARK_ARC_1_0/temp4[141] , \MC_ARK_ARC_1_0/temp4[140] ,
         \MC_ARK_ARC_1_0/temp4[139] , \MC_ARK_ARC_1_0/temp4[138] ,
         \MC_ARK_ARC_1_0/temp4[137] , \MC_ARK_ARC_1_0/temp4[136] ,
         \MC_ARK_ARC_1_0/temp4[135] , \MC_ARK_ARC_1_0/temp4[134] ,
         \MC_ARK_ARC_1_0/temp4[133] , \MC_ARK_ARC_1_0/temp4[132] ,
         \MC_ARK_ARC_1_0/temp4[131] , \MC_ARK_ARC_1_0/temp4[130] ,
         \MC_ARK_ARC_1_0/temp4[129] , \MC_ARK_ARC_1_0/temp4[128] ,
         \MC_ARK_ARC_1_0/temp4[127] , \MC_ARK_ARC_1_0/temp4[126] ,
         \MC_ARK_ARC_1_0/temp4[125] , \MC_ARK_ARC_1_0/temp4[124] ,
         \MC_ARK_ARC_1_0/temp4[123] , \MC_ARK_ARC_1_0/temp4[122] ,
         \MC_ARK_ARC_1_0/temp4[121] , \MC_ARK_ARC_1_0/temp4[120] ,
         \MC_ARK_ARC_1_0/temp4[119] , \MC_ARK_ARC_1_0/temp4[118] ,
         \MC_ARK_ARC_1_0/temp4[117] , \MC_ARK_ARC_1_0/temp4[116] ,
         \MC_ARK_ARC_1_0/temp4[115] , \MC_ARK_ARC_1_0/temp4[114] ,
         \MC_ARK_ARC_1_0/temp4[113] , \MC_ARK_ARC_1_0/temp4[112] ,
         \MC_ARK_ARC_1_0/temp4[111] , \MC_ARK_ARC_1_0/temp4[110] ,
         \MC_ARK_ARC_1_0/temp4[109] , \MC_ARK_ARC_1_0/temp4[108] ,
         \MC_ARK_ARC_1_0/temp4[107] , \MC_ARK_ARC_1_0/temp4[106] ,
         \MC_ARK_ARC_1_0/temp4[105] , \MC_ARK_ARC_1_0/temp4[104] ,
         \MC_ARK_ARC_1_0/temp4[103] , \MC_ARK_ARC_1_0/temp4[102] ,
         \MC_ARK_ARC_1_0/temp4[101] , \MC_ARK_ARC_1_0/temp4[100] ,
         \MC_ARK_ARC_1_0/temp4[99] , \MC_ARK_ARC_1_0/temp4[98] ,
         \MC_ARK_ARC_1_0/temp4[97] , \MC_ARK_ARC_1_0/temp4[96] ,
         \MC_ARK_ARC_1_0/temp4[95] , \MC_ARK_ARC_1_0/temp4[94] ,
         \MC_ARK_ARC_1_0/temp4[93] , \MC_ARK_ARC_1_0/temp4[92] ,
         \MC_ARK_ARC_1_0/temp4[91] , \MC_ARK_ARC_1_0/temp4[90] ,
         \MC_ARK_ARC_1_0/temp4[89] , \MC_ARK_ARC_1_0/temp4[88] ,
         \MC_ARK_ARC_1_0/temp4[87] , \MC_ARK_ARC_1_0/temp4[86] ,
         \MC_ARK_ARC_1_0/temp4[85] , \MC_ARK_ARC_1_0/temp4[84] ,
         \MC_ARK_ARC_1_0/temp4[83] , \MC_ARK_ARC_1_0/temp4[82] ,
         \MC_ARK_ARC_1_0/temp4[81] , \MC_ARK_ARC_1_0/temp4[80] ,
         \MC_ARK_ARC_1_0/temp4[79] , \MC_ARK_ARC_1_0/temp4[78] ,
         \MC_ARK_ARC_1_0/temp4[77] , \MC_ARK_ARC_1_0/temp4[76] ,
         \MC_ARK_ARC_1_0/temp4[75] , \MC_ARK_ARC_1_0/temp4[74] ,
         \MC_ARK_ARC_1_0/temp4[73] , \MC_ARK_ARC_1_0/temp4[72] ,
         \MC_ARK_ARC_1_0/temp4[71] , \MC_ARK_ARC_1_0/temp4[70] ,
         \MC_ARK_ARC_1_0/temp4[69] , \MC_ARK_ARC_1_0/temp4[68] ,
         \MC_ARK_ARC_1_0/temp4[67] , \MC_ARK_ARC_1_0/temp4[66] ,
         \MC_ARK_ARC_1_0/temp4[65] , \MC_ARK_ARC_1_0/temp4[64] ,
         \MC_ARK_ARC_1_0/temp4[63] , \MC_ARK_ARC_1_0/temp4[62] ,
         \MC_ARK_ARC_1_0/temp4[61] , \MC_ARK_ARC_1_0/temp4[60] ,
         \MC_ARK_ARC_1_0/temp4[59] , \MC_ARK_ARC_1_0/temp4[58] ,
         \MC_ARK_ARC_1_0/temp4[57] , \MC_ARK_ARC_1_0/temp4[56] ,
         \MC_ARK_ARC_1_0/temp4[55] , \MC_ARK_ARC_1_0/temp4[54] ,
         \MC_ARK_ARC_1_0/temp4[53] , \MC_ARK_ARC_1_0/temp4[52] ,
         \MC_ARK_ARC_1_0/temp4[51] , \MC_ARK_ARC_1_0/temp4[50] ,
         \MC_ARK_ARC_1_0/temp4[49] , \MC_ARK_ARC_1_0/temp4[48] ,
         \MC_ARK_ARC_1_0/temp4[47] , \MC_ARK_ARC_1_0/temp4[46] ,
         \MC_ARK_ARC_1_0/temp4[45] , \MC_ARK_ARC_1_0/temp4[44] ,
         \MC_ARK_ARC_1_0/temp4[43] , \MC_ARK_ARC_1_0/temp4[42] ,
         \MC_ARK_ARC_1_0/temp4[41] , \MC_ARK_ARC_1_0/temp4[40] ,
         \MC_ARK_ARC_1_0/temp4[39] , \MC_ARK_ARC_1_0/temp4[38] ,
         \MC_ARK_ARC_1_0/temp4[37] , \MC_ARK_ARC_1_0/temp4[36] ,
         \MC_ARK_ARC_1_0/temp4[35] , \MC_ARK_ARC_1_0/temp4[34] ,
         \MC_ARK_ARC_1_0/temp4[33] , \MC_ARK_ARC_1_0/temp4[32] ,
         \MC_ARK_ARC_1_0/temp4[31] , \MC_ARK_ARC_1_0/temp4[30] ,
         \MC_ARK_ARC_1_0/temp4[29] , \MC_ARK_ARC_1_0/temp4[28] ,
         \MC_ARK_ARC_1_0/temp4[27] , \MC_ARK_ARC_1_0/temp4[26] ,
         \MC_ARK_ARC_1_0/temp4[25] , \MC_ARK_ARC_1_0/temp4[24] ,
         \MC_ARK_ARC_1_0/temp4[23] , \MC_ARK_ARC_1_0/temp4[22] ,
         \MC_ARK_ARC_1_0/temp4[21] , \MC_ARK_ARC_1_0/temp4[20] ,
         \MC_ARK_ARC_1_0/temp4[19] , \MC_ARK_ARC_1_0/temp4[18] ,
         \MC_ARK_ARC_1_0/temp4[17] , \MC_ARK_ARC_1_0/temp4[16] ,
         \MC_ARK_ARC_1_0/temp4[15] , \MC_ARK_ARC_1_0/temp4[14] ,
         \MC_ARK_ARC_1_0/temp4[13] , \MC_ARK_ARC_1_0/temp4[12] ,
         \MC_ARK_ARC_1_0/temp4[11] , \MC_ARK_ARC_1_0/temp4[10] ,
         \MC_ARK_ARC_1_0/temp4[9] , \MC_ARK_ARC_1_0/temp4[8] ,
         \MC_ARK_ARC_1_0/temp4[7] , \MC_ARK_ARC_1_0/temp4[6] ,
         \MC_ARK_ARC_1_0/temp4[5] , \MC_ARK_ARC_1_0/temp4[4] ,
         \MC_ARK_ARC_1_0/temp4[3] , \MC_ARK_ARC_1_0/temp4[2] ,
         \MC_ARK_ARC_1_0/temp4[1] , \MC_ARK_ARC_1_0/temp4[0] ,
         \MC_ARK_ARC_1_0/temp3[191] , \MC_ARK_ARC_1_0/temp3[190] ,
         \MC_ARK_ARC_1_0/temp3[189] , \MC_ARK_ARC_1_0/temp3[188] ,
         \MC_ARK_ARC_1_0/temp3[187] , \MC_ARK_ARC_1_0/temp3[186] ,
         \MC_ARK_ARC_1_0/temp3[185] , \MC_ARK_ARC_1_0/temp3[184] ,
         \MC_ARK_ARC_1_0/temp3[183] , \MC_ARK_ARC_1_0/temp3[182] ,
         \MC_ARK_ARC_1_0/temp3[181] , \MC_ARK_ARC_1_0/temp3[180] ,
         \MC_ARK_ARC_1_0/temp3[179] , \MC_ARK_ARC_1_0/temp3[178] ,
         \MC_ARK_ARC_1_0/temp3[177] , \MC_ARK_ARC_1_0/temp3[176] ,
         \MC_ARK_ARC_1_0/temp3[175] , \MC_ARK_ARC_1_0/temp3[174] ,
         \MC_ARK_ARC_1_0/temp3[173] , \MC_ARK_ARC_1_0/temp3[172] ,
         \MC_ARK_ARC_1_0/temp3[171] , \MC_ARK_ARC_1_0/temp3[170] ,
         \MC_ARK_ARC_1_0/temp3[169] , \MC_ARK_ARC_1_0/temp3[168] ,
         \MC_ARK_ARC_1_0/temp3[167] , \MC_ARK_ARC_1_0/temp3[166] ,
         \MC_ARK_ARC_1_0/temp3[165] , \MC_ARK_ARC_1_0/temp3[164] ,
         \MC_ARK_ARC_1_0/temp3[163] , \MC_ARK_ARC_1_0/temp3[162] ,
         \MC_ARK_ARC_1_0/temp3[161] , \MC_ARK_ARC_1_0/temp3[160] ,
         \MC_ARK_ARC_1_0/temp3[159] , \MC_ARK_ARC_1_0/temp3[158] ,
         \MC_ARK_ARC_1_0/temp3[157] , \MC_ARK_ARC_1_0/temp3[156] ,
         \MC_ARK_ARC_1_0/temp3[155] , \MC_ARK_ARC_1_0/temp3[154] ,
         \MC_ARK_ARC_1_0/temp3[153] , \MC_ARK_ARC_1_0/temp3[152] ,
         \MC_ARK_ARC_1_0/temp3[151] , \MC_ARK_ARC_1_0/temp3[150] ,
         \MC_ARK_ARC_1_0/temp3[149] , \MC_ARK_ARC_1_0/temp3[148] ,
         \MC_ARK_ARC_1_0/temp3[147] , \MC_ARK_ARC_1_0/temp3[146] ,
         \MC_ARK_ARC_1_0/temp3[145] , \MC_ARK_ARC_1_0/temp3[144] ,
         \MC_ARK_ARC_1_0/temp3[143] , \MC_ARK_ARC_1_0/temp3[142] ,
         \MC_ARK_ARC_1_0/temp3[141] , \MC_ARK_ARC_1_0/temp3[140] ,
         \MC_ARK_ARC_1_0/temp3[139] , \MC_ARK_ARC_1_0/temp3[138] ,
         \MC_ARK_ARC_1_0/temp3[137] , \MC_ARK_ARC_1_0/temp3[136] ,
         \MC_ARK_ARC_1_0/temp3[135] , \MC_ARK_ARC_1_0/temp3[134] ,
         \MC_ARK_ARC_1_0/temp3[133] , \MC_ARK_ARC_1_0/temp3[132] ,
         \MC_ARK_ARC_1_0/temp3[131] , \MC_ARK_ARC_1_0/temp3[130] ,
         \MC_ARK_ARC_1_0/temp3[129] , \MC_ARK_ARC_1_0/temp3[128] ,
         \MC_ARK_ARC_1_0/temp3[127] , \MC_ARK_ARC_1_0/temp3[126] ,
         \MC_ARK_ARC_1_0/temp3[125] , \MC_ARK_ARC_1_0/temp3[124] ,
         \MC_ARK_ARC_1_0/temp3[123] , \MC_ARK_ARC_1_0/temp3[122] ,
         \MC_ARK_ARC_1_0/temp3[121] , \MC_ARK_ARC_1_0/temp3[120] ,
         \MC_ARK_ARC_1_0/temp3[119] , \MC_ARK_ARC_1_0/temp3[118] ,
         \MC_ARK_ARC_1_0/temp3[117] , \MC_ARK_ARC_1_0/temp3[116] ,
         \MC_ARK_ARC_1_0/temp3[115] , \MC_ARK_ARC_1_0/temp3[114] ,
         \MC_ARK_ARC_1_0/temp3[113] , \MC_ARK_ARC_1_0/temp3[112] ,
         \MC_ARK_ARC_1_0/temp3[111] , \MC_ARK_ARC_1_0/temp3[110] ,
         \MC_ARK_ARC_1_0/temp3[109] , \MC_ARK_ARC_1_0/temp3[108] ,
         \MC_ARK_ARC_1_0/temp3[107] , \MC_ARK_ARC_1_0/temp3[106] ,
         \MC_ARK_ARC_1_0/temp3[105] , \MC_ARK_ARC_1_0/temp3[104] ,
         \MC_ARK_ARC_1_0/temp3[103] , \MC_ARK_ARC_1_0/temp3[102] ,
         \MC_ARK_ARC_1_0/temp3[101] , \MC_ARK_ARC_1_0/temp3[100] ,
         \MC_ARK_ARC_1_0/temp3[99] , \MC_ARK_ARC_1_0/temp3[98] ,
         \MC_ARK_ARC_1_0/temp3[97] , \MC_ARK_ARC_1_0/temp3[96] ,
         \MC_ARK_ARC_1_0/temp3[95] , \MC_ARK_ARC_1_0/temp3[94] ,
         \MC_ARK_ARC_1_0/temp3[93] , \MC_ARK_ARC_1_0/temp3[92] ,
         \MC_ARK_ARC_1_0/temp3[91] , \MC_ARK_ARC_1_0/temp3[90] ,
         \MC_ARK_ARC_1_0/temp3[89] , \MC_ARK_ARC_1_0/temp3[88] ,
         \MC_ARK_ARC_1_0/temp3[87] , \MC_ARK_ARC_1_0/temp3[86] ,
         \MC_ARK_ARC_1_0/temp3[85] , \MC_ARK_ARC_1_0/temp3[84] ,
         \MC_ARK_ARC_1_0/temp3[83] , \MC_ARK_ARC_1_0/temp3[82] ,
         \MC_ARK_ARC_1_0/temp3[81] , \MC_ARK_ARC_1_0/temp3[80] ,
         \MC_ARK_ARC_1_0/temp3[79] , \MC_ARK_ARC_1_0/temp3[78] ,
         \MC_ARK_ARC_1_0/temp3[77] , \MC_ARK_ARC_1_0/temp3[76] ,
         \MC_ARK_ARC_1_0/temp3[75] , \MC_ARK_ARC_1_0/temp3[74] ,
         \MC_ARK_ARC_1_0/temp3[73] , \MC_ARK_ARC_1_0/temp3[72] ,
         \MC_ARK_ARC_1_0/temp3[71] , \MC_ARK_ARC_1_0/temp3[70] ,
         \MC_ARK_ARC_1_0/temp3[69] , \MC_ARK_ARC_1_0/temp3[68] ,
         \MC_ARK_ARC_1_0/temp3[67] , \MC_ARK_ARC_1_0/temp3[66] ,
         \MC_ARK_ARC_1_0/temp3[65] , \MC_ARK_ARC_1_0/temp3[64] ,
         \MC_ARK_ARC_1_0/temp3[63] , \MC_ARK_ARC_1_0/temp3[62] ,
         \MC_ARK_ARC_1_0/temp3[61] , \MC_ARK_ARC_1_0/temp3[60] ,
         \MC_ARK_ARC_1_0/temp3[59] , \MC_ARK_ARC_1_0/temp3[58] ,
         \MC_ARK_ARC_1_0/temp3[57] , \MC_ARK_ARC_1_0/temp3[56] ,
         \MC_ARK_ARC_1_0/temp3[55] , \MC_ARK_ARC_1_0/temp3[54] ,
         \MC_ARK_ARC_1_0/temp3[53] , \MC_ARK_ARC_1_0/temp3[52] ,
         \MC_ARK_ARC_1_0/temp3[51] , \MC_ARK_ARC_1_0/temp3[50] ,
         \MC_ARK_ARC_1_0/temp3[49] , \MC_ARK_ARC_1_0/temp3[48] ,
         \MC_ARK_ARC_1_0/temp3[47] , \MC_ARK_ARC_1_0/temp3[46] ,
         \MC_ARK_ARC_1_0/temp3[45] , \MC_ARK_ARC_1_0/temp3[44] ,
         \MC_ARK_ARC_1_0/temp3[43] , \MC_ARK_ARC_1_0/temp3[42] ,
         \MC_ARK_ARC_1_0/temp3[41] , \MC_ARK_ARC_1_0/temp3[40] ,
         \MC_ARK_ARC_1_0/temp3[39] , \MC_ARK_ARC_1_0/temp3[38] ,
         \MC_ARK_ARC_1_0/temp3[37] , \MC_ARK_ARC_1_0/temp3[36] ,
         \MC_ARK_ARC_1_0/temp3[35] , \MC_ARK_ARC_1_0/temp3[34] ,
         \MC_ARK_ARC_1_0/temp3[33] , \MC_ARK_ARC_1_0/temp3[32] ,
         \MC_ARK_ARC_1_0/temp3[31] , \MC_ARK_ARC_1_0/temp3[30] ,
         \MC_ARK_ARC_1_0/temp3[29] , \MC_ARK_ARC_1_0/temp3[28] ,
         \MC_ARK_ARC_1_0/temp3[27] , \MC_ARK_ARC_1_0/temp3[26] ,
         \MC_ARK_ARC_1_0/temp3[25] , \MC_ARK_ARC_1_0/temp3[24] ,
         \MC_ARK_ARC_1_0/temp3[23] , \MC_ARK_ARC_1_0/temp3[22] ,
         \MC_ARK_ARC_1_0/temp3[21] , \MC_ARK_ARC_1_0/temp3[20] ,
         \MC_ARK_ARC_1_0/temp3[19] , \MC_ARK_ARC_1_0/temp3[18] ,
         \MC_ARK_ARC_1_0/temp3[17] , \MC_ARK_ARC_1_0/temp3[16] ,
         \MC_ARK_ARC_1_0/temp3[15] , \MC_ARK_ARC_1_0/temp3[14] ,
         \MC_ARK_ARC_1_0/temp3[13] , \MC_ARK_ARC_1_0/temp3[12] ,
         \MC_ARK_ARC_1_0/temp3[11] , \MC_ARK_ARC_1_0/temp3[10] ,
         \MC_ARK_ARC_1_0/temp3[9] , \MC_ARK_ARC_1_0/temp3[8] ,
         \MC_ARK_ARC_1_0/temp3[7] , \MC_ARK_ARC_1_0/temp3[6] ,
         \MC_ARK_ARC_1_0/temp3[5] , \MC_ARK_ARC_1_0/temp3[4] ,
         \MC_ARK_ARC_1_0/temp3[3] , \MC_ARK_ARC_1_0/temp3[2] ,
         \MC_ARK_ARC_1_0/temp3[1] , \MC_ARK_ARC_1_0/temp3[0] ,
         \MC_ARK_ARC_1_0/temp2[191] , \MC_ARK_ARC_1_0/temp2[190] ,
         \MC_ARK_ARC_1_0/temp2[189] , \MC_ARK_ARC_1_0/temp2[188] ,
         \MC_ARK_ARC_1_0/temp2[187] , \MC_ARK_ARC_1_0/temp2[186] ,
         \MC_ARK_ARC_1_0/temp2[185] , \MC_ARK_ARC_1_0/temp2[184] ,
         \MC_ARK_ARC_1_0/temp2[183] , \MC_ARK_ARC_1_0/temp2[182] ,
         \MC_ARK_ARC_1_0/temp2[181] , \MC_ARK_ARC_1_0/temp2[180] ,
         \MC_ARK_ARC_1_0/temp2[179] , \MC_ARK_ARC_1_0/temp2[178] ,
         \MC_ARK_ARC_1_0/temp2[177] , \MC_ARK_ARC_1_0/temp2[176] ,
         \MC_ARK_ARC_1_0/temp2[175] , \MC_ARK_ARC_1_0/temp2[174] ,
         \MC_ARK_ARC_1_0/temp2[173] , \MC_ARK_ARC_1_0/temp2[172] ,
         \MC_ARK_ARC_1_0/temp2[171] , \MC_ARK_ARC_1_0/temp2[170] ,
         \MC_ARK_ARC_1_0/temp2[169] , \MC_ARK_ARC_1_0/temp2[168] ,
         \MC_ARK_ARC_1_0/temp2[167] , \MC_ARK_ARC_1_0/temp2[166] ,
         \MC_ARK_ARC_1_0/temp2[165] , \MC_ARK_ARC_1_0/temp2[164] ,
         \MC_ARK_ARC_1_0/temp2[163] , \MC_ARK_ARC_1_0/temp2[162] ,
         \MC_ARK_ARC_1_0/temp2[161] , \MC_ARK_ARC_1_0/temp2[160] ,
         \MC_ARK_ARC_1_0/temp2[159] , \MC_ARK_ARC_1_0/temp2[158] ,
         \MC_ARK_ARC_1_0/temp2[157] , \MC_ARK_ARC_1_0/temp2[156] ,
         \MC_ARK_ARC_1_0/temp2[155] , \MC_ARK_ARC_1_0/temp2[154] ,
         \MC_ARK_ARC_1_0/temp2[153] , \MC_ARK_ARC_1_0/temp2[152] ,
         \MC_ARK_ARC_1_0/temp2[151] , \MC_ARK_ARC_1_0/temp2[150] ,
         \MC_ARK_ARC_1_0/temp2[149] , \MC_ARK_ARC_1_0/temp2[148] ,
         \MC_ARK_ARC_1_0/temp2[147] , \MC_ARK_ARC_1_0/temp2[146] ,
         \MC_ARK_ARC_1_0/temp2[145] , \MC_ARK_ARC_1_0/temp2[144] ,
         \MC_ARK_ARC_1_0/temp2[143] , \MC_ARK_ARC_1_0/temp2[142] ,
         \MC_ARK_ARC_1_0/temp2[141] , \MC_ARK_ARC_1_0/temp2[140] ,
         \MC_ARK_ARC_1_0/temp2[139] , \MC_ARK_ARC_1_0/temp2[138] ,
         \MC_ARK_ARC_1_0/temp2[137] , \MC_ARK_ARC_1_0/temp2[136] ,
         \MC_ARK_ARC_1_0/temp2[135] , \MC_ARK_ARC_1_0/temp2[134] ,
         \MC_ARK_ARC_1_0/temp2[133] , \MC_ARK_ARC_1_0/temp2[132] ,
         \MC_ARK_ARC_1_0/temp2[131] , \MC_ARK_ARC_1_0/temp2[130] ,
         \MC_ARK_ARC_1_0/temp2[129] , \MC_ARK_ARC_1_0/temp2[128] ,
         \MC_ARK_ARC_1_0/temp2[127] , \MC_ARK_ARC_1_0/temp2[126] ,
         \MC_ARK_ARC_1_0/temp2[125] , \MC_ARK_ARC_1_0/temp2[124] ,
         \MC_ARK_ARC_1_0/temp2[123] , \MC_ARK_ARC_1_0/temp2[122] ,
         \MC_ARK_ARC_1_0/temp2[121] , \MC_ARK_ARC_1_0/temp2[120] ,
         \MC_ARK_ARC_1_0/temp2[119] , \MC_ARK_ARC_1_0/temp2[118] ,
         \MC_ARK_ARC_1_0/temp2[117] , \MC_ARK_ARC_1_0/temp2[116] ,
         \MC_ARK_ARC_1_0/temp2[115] , \MC_ARK_ARC_1_0/temp2[114] ,
         \MC_ARK_ARC_1_0/temp2[113] , \MC_ARK_ARC_1_0/temp2[112] ,
         \MC_ARK_ARC_1_0/temp2[111] , \MC_ARK_ARC_1_0/temp2[110] ,
         \MC_ARK_ARC_1_0/temp2[109] , \MC_ARK_ARC_1_0/temp2[108] ,
         \MC_ARK_ARC_1_0/temp2[107] , \MC_ARK_ARC_1_0/temp2[106] ,
         \MC_ARK_ARC_1_0/temp2[105] , \MC_ARK_ARC_1_0/temp2[104] ,
         \MC_ARK_ARC_1_0/temp2[103] , \MC_ARK_ARC_1_0/temp2[102] ,
         \MC_ARK_ARC_1_0/temp2[101] , \MC_ARK_ARC_1_0/temp2[100] ,
         \MC_ARK_ARC_1_0/temp2[99] , \MC_ARK_ARC_1_0/temp2[98] ,
         \MC_ARK_ARC_1_0/temp2[97] , \MC_ARK_ARC_1_0/temp2[96] ,
         \MC_ARK_ARC_1_0/temp2[95] , \MC_ARK_ARC_1_0/temp2[94] ,
         \MC_ARK_ARC_1_0/temp2[93] , \MC_ARK_ARC_1_0/temp2[92] ,
         \MC_ARK_ARC_1_0/temp2[91] , \MC_ARK_ARC_1_0/temp2[90] ,
         \MC_ARK_ARC_1_0/temp2[89] , \MC_ARK_ARC_1_0/temp2[88] ,
         \MC_ARK_ARC_1_0/temp2[87] , \MC_ARK_ARC_1_0/temp2[86] ,
         \MC_ARK_ARC_1_0/temp2[85] , \MC_ARK_ARC_1_0/temp2[84] ,
         \MC_ARK_ARC_1_0/temp2[83] , \MC_ARK_ARC_1_0/temp2[82] ,
         \MC_ARK_ARC_1_0/temp2[81] , \MC_ARK_ARC_1_0/temp2[80] ,
         \MC_ARK_ARC_1_0/temp2[79] , \MC_ARK_ARC_1_0/temp2[78] ,
         \MC_ARK_ARC_1_0/temp2[77] , \MC_ARK_ARC_1_0/temp2[76] ,
         \MC_ARK_ARC_1_0/temp2[75] , \MC_ARK_ARC_1_0/temp2[74] ,
         \MC_ARK_ARC_1_0/temp2[73] , \MC_ARK_ARC_1_0/temp2[72] ,
         \MC_ARK_ARC_1_0/temp2[71] , \MC_ARK_ARC_1_0/temp2[70] ,
         \MC_ARK_ARC_1_0/temp2[69] , \MC_ARK_ARC_1_0/temp2[68] ,
         \MC_ARK_ARC_1_0/temp2[67] , \MC_ARK_ARC_1_0/temp2[66] ,
         \MC_ARK_ARC_1_0/temp2[65] , \MC_ARK_ARC_1_0/temp2[64] ,
         \MC_ARK_ARC_1_0/temp2[63] , \MC_ARK_ARC_1_0/temp2[62] ,
         \MC_ARK_ARC_1_0/temp2[61] , \MC_ARK_ARC_1_0/temp2[60] ,
         \MC_ARK_ARC_1_0/temp2[59] , \MC_ARK_ARC_1_0/temp2[58] ,
         \MC_ARK_ARC_1_0/temp2[57] , \MC_ARK_ARC_1_0/temp2[56] ,
         \MC_ARK_ARC_1_0/temp2[55] , \MC_ARK_ARC_1_0/temp2[54] ,
         \MC_ARK_ARC_1_0/temp2[53] , \MC_ARK_ARC_1_0/temp2[52] ,
         \MC_ARK_ARC_1_0/temp2[51] , \MC_ARK_ARC_1_0/temp2[50] ,
         \MC_ARK_ARC_1_0/temp2[49] , \MC_ARK_ARC_1_0/temp2[48] ,
         \MC_ARK_ARC_1_0/temp2[47] , \MC_ARK_ARC_1_0/temp2[46] ,
         \MC_ARK_ARC_1_0/temp2[45] , \MC_ARK_ARC_1_0/temp2[44] ,
         \MC_ARK_ARC_1_0/temp2[43] , \MC_ARK_ARC_1_0/temp2[42] ,
         \MC_ARK_ARC_1_0/temp2[41] , \MC_ARK_ARC_1_0/temp2[40] ,
         \MC_ARK_ARC_1_0/temp2[39] , \MC_ARK_ARC_1_0/temp2[38] ,
         \MC_ARK_ARC_1_0/temp2[37] , \MC_ARK_ARC_1_0/temp2[36] ,
         \MC_ARK_ARC_1_0/temp2[35] , \MC_ARK_ARC_1_0/temp2[34] ,
         \MC_ARK_ARC_1_0/temp2[33] , \MC_ARK_ARC_1_0/temp2[32] ,
         \MC_ARK_ARC_1_0/temp2[31] , \MC_ARK_ARC_1_0/temp2[30] ,
         \MC_ARK_ARC_1_0/temp2[29] , \MC_ARK_ARC_1_0/temp2[28] ,
         \MC_ARK_ARC_1_0/temp2[27] , \MC_ARK_ARC_1_0/temp2[26] ,
         \MC_ARK_ARC_1_0/temp2[25] , \MC_ARK_ARC_1_0/temp2[24] ,
         \MC_ARK_ARC_1_0/temp2[23] , \MC_ARK_ARC_1_0/temp2[22] ,
         \MC_ARK_ARC_1_0/temp2[21] , \MC_ARK_ARC_1_0/temp2[20] ,
         \MC_ARK_ARC_1_0/temp2[19] , \MC_ARK_ARC_1_0/temp2[18] ,
         \MC_ARK_ARC_1_0/temp2[17] , \MC_ARK_ARC_1_0/temp2[16] ,
         \MC_ARK_ARC_1_0/temp2[15] , \MC_ARK_ARC_1_0/temp2[14] ,
         \MC_ARK_ARC_1_0/temp2[13] , \MC_ARK_ARC_1_0/temp2[12] ,
         \MC_ARK_ARC_1_0/temp2[11] , \MC_ARK_ARC_1_0/temp2[10] ,
         \MC_ARK_ARC_1_0/temp2[9] , \MC_ARK_ARC_1_0/temp2[8] ,
         \MC_ARK_ARC_1_0/temp2[7] , \MC_ARK_ARC_1_0/temp2[6] ,
         \MC_ARK_ARC_1_0/temp2[5] , \MC_ARK_ARC_1_0/temp2[4] ,
         \MC_ARK_ARC_1_0/temp2[3] , \MC_ARK_ARC_1_0/temp2[2] ,
         \MC_ARK_ARC_1_0/temp2[1] , \MC_ARK_ARC_1_0/temp2[0] ,
         \MC_ARK_ARC_1_0/temp1[191] , \MC_ARK_ARC_1_0/temp1[190] ,
         \MC_ARK_ARC_1_0/temp1[189] , \MC_ARK_ARC_1_0/temp1[188] ,
         \MC_ARK_ARC_1_0/temp1[187] , \MC_ARK_ARC_1_0/temp1[186] ,
         \MC_ARK_ARC_1_0/temp1[185] , \MC_ARK_ARC_1_0/temp1[184] ,
         \MC_ARK_ARC_1_0/temp1[183] , \MC_ARK_ARC_1_0/temp1[182] ,
         \MC_ARK_ARC_1_0/temp1[181] , \MC_ARK_ARC_1_0/temp1[180] ,
         \MC_ARK_ARC_1_0/temp1[179] , \MC_ARK_ARC_1_0/temp1[178] ,
         \MC_ARK_ARC_1_0/temp1[177] , \MC_ARK_ARC_1_0/temp1[176] ,
         \MC_ARK_ARC_1_0/temp1[175] , \MC_ARK_ARC_1_0/temp1[174] ,
         \MC_ARK_ARC_1_0/temp1[173] , \MC_ARK_ARC_1_0/temp1[172] ,
         \MC_ARK_ARC_1_0/temp1[171] , \MC_ARK_ARC_1_0/temp1[170] ,
         \MC_ARK_ARC_1_0/temp1[169] , \MC_ARK_ARC_1_0/temp1[168] ,
         \MC_ARK_ARC_1_0/temp1[167] , \MC_ARK_ARC_1_0/temp1[166] ,
         \MC_ARK_ARC_1_0/temp1[165] , \MC_ARK_ARC_1_0/temp1[164] ,
         \MC_ARK_ARC_1_0/temp1[163] , \MC_ARK_ARC_1_0/temp1[162] ,
         \MC_ARK_ARC_1_0/temp1[161] , \MC_ARK_ARC_1_0/temp1[160] ,
         \MC_ARK_ARC_1_0/temp1[159] , \MC_ARK_ARC_1_0/temp1[158] ,
         \MC_ARK_ARC_1_0/temp1[157] , \MC_ARK_ARC_1_0/temp1[156] ,
         \MC_ARK_ARC_1_0/temp1[155] , \MC_ARK_ARC_1_0/temp1[154] ,
         \MC_ARK_ARC_1_0/temp1[153] , \MC_ARK_ARC_1_0/temp1[152] ,
         \MC_ARK_ARC_1_0/temp1[151] , \MC_ARK_ARC_1_0/temp1[150] ,
         \MC_ARK_ARC_1_0/temp1[149] , \MC_ARK_ARC_1_0/temp1[148] ,
         \MC_ARK_ARC_1_0/temp1[147] , \MC_ARK_ARC_1_0/temp1[146] ,
         \MC_ARK_ARC_1_0/temp1[145] , \MC_ARK_ARC_1_0/temp1[144] ,
         \MC_ARK_ARC_1_0/temp1[143] , \MC_ARK_ARC_1_0/temp1[142] ,
         \MC_ARK_ARC_1_0/temp1[141] , \MC_ARK_ARC_1_0/temp1[140] ,
         \MC_ARK_ARC_1_0/temp1[139] , \MC_ARK_ARC_1_0/temp1[138] ,
         \MC_ARK_ARC_1_0/temp1[137] , \MC_ARK_ARC_1_0/temp1[136] ,
         \MC_ARK_ARC_1_0/temp1[135] , \MC_ARK_ARC_1_0/temp1[134] ,
         \MC_ARK_ARC_1_0/temp1[133] , \MC_ARK_ARC_1_0/temp1[132] ,
         \MC_ARK_ARC_1_0/temp1[131] , \MC_ARK_ARC_1_0/temp1[130] ,
         \MC_ARK_ARC_1_0/temp1[129] , \MC_ARK_ARC_1_0/temp1[128] ,
         \MC_ARK_ARC_1_0/temp1[127] , \MC_ARK_ARC_1_0/temp1[126] ,
         \MC_ARK_ARC_1_0/temp1[125] , \MC_ARK_ARC_1_0/temp1[124] ,
         \MC_ARK_ARC_1_0/temp1[123] , \MC_ARK_ARC_1_0/temp1[122] ,
         \MC_ARK_ARC_1_0/temp1[121] , \MC_ARK_ARC_1_0/temp1[120] ,
         \MC_ARK_ARC_1_0/temp1[119] , \MC_ARK_ARC_1_0/temp1[118] ,
         \MC_ARK_ARC_1_0/temp1[117] , \MC_ARK_ARC_1_0/temp1[116] ,
         \MC_ARK_ARC_1_0/temp1[115] , \MC_ARK_ARC_1_0/temp1[114] ,
         \MC_ARK_ARC_1_0/temp1[113] , \MC_ARK_ARC_1_0/temp1[112] ,
         \MC_ARK_ARC_1_0/temp1[111] , \MC_ARK_ARC_1_0/temp1[110] ,
         \MC_ARK_ARC_1_0/temp1[109] , \MC_ARK_ARC_1_0/temp1[108] ,
         \MC_ARK_ARC_1_0/temp1[107] , \MC_ARK_ARC_1_0/temp1[106] ,
         \MC_ARK_ARC_1_0/temp1[105] , \MC_ARK_ARC_1_0/temp1[104] ,
         \MC_ARK_ARC_1_0/temp1[103] , \MC_ARK_ARC_1_0/temp1[102] ,
         \MC_ARK_ARC_1_0/temp1[101] , \MC_ARK_ARC_1_0/temp1[100] ,
         \MC_ARK_ARC_1_0/temp1[99] , \MC_ARK_ARC_1_0/temp1[98] ,
         \MC_ARK_ARC_1_0/temp1[97] , \MC_ARK_ARC_1_0/temp1[96] ,
         \MC_ARK_ARC_1_0/temp1[95] , \MC_ARK_ARC_1_0/temp1[94] ,
         \MC_ARK_ARC_1_0/temp1[93] , \MC_ARK_ARC_1_0/temp1[92] ,
         \MC_ARK_ARC_1_0/temp1[91] , \MC_ARK_ARC_1_0/temp1[90] ,
         \MC_ARK_ARC_1_0/temp1[89] , \MC_ARK_ARC_1_0/temp1[88] ,
         \MC_ARK_ARC_1_0/temp1[87] , \MC_ARK_ARC_1_0/temp1[86] ,
         \MC_ARK_ARC_1_0/temp1[85] , \MC_ARK_ARC_1_0/temp1[84] ,
         \MC_ARK_ARC_1_0/temp1[83] , \MC_ARK_ARC_1_0/temp1[82] ,
         \MC_ARK_ARC_1_0/temp1[81] , \MC_ARK_ARC_1_0/temp1[80] ,
         \MC_ARK_ARC_1_0/temp1[79] , \MC_ARK_ARC_1_0/temp1[78] ,
         \MC_ARK_ARC_1_0/temp1[77] , \MC_ARK_ARC_1_0/temp1[76] ,
         \MC_ARK_ARC_1_0/temp1[75] , \MC_ARK_ARC_1_0/temp1[74] ,
         \MC_ARK_ARC_1_0/temp1[73] , \MC_ARK_ARC_1_0/temp1[72] ,
         \MC_ARK_ARC_1_0/temp1[71] , \MC_ARK_ARC_1_0/temp1[70] ,
         \MC_ARK_ARC_1_0/temp1[69] , \MC_ARK_ARC_1_0/temp1[68] ,
         \MC_ARK_ARC_1_0/temp1[67] , \MC_ARK_ARC_1_0/temp1[66] ,
         \MC_ARK_ARC_1_0/temp1[65] , \MC_ARK_ARC_1_0/temp1[64] ,
         \MC_ARK_ARC_1_0/temp1[63] , \MC_ARK_ARC_1_0/temp1[62] ,
         \MC_ARK_ARC_1_0/temp1[61] , \MC_ARK_ARC_1_0/temp1[60] ,
         \MC_ARK_ARC_1_0/temp1[59] , \MC_ARK_ARC_1_0/temp1[58] ,
         \MC_ARK_ARC_1_0/temp1[57] , \MC_ARK_ARC_1_0/temp1[56] ,
         \MC_ARK_ARC_1_0/temp1[55] , \MC_ARK_ARC_1_0/temp1[54] ,
         \MC_ARK_ARC_1_0/temp1[53] , \MC_ARK_ARC_1_0/temp1[52] ,
         \MC_ARK_ARC_1_0/temp1[51] , \MC_ARK_ARC_1_0/temp1[50] ,
         \MC_ARK_ARC_1_0/temp1[49] , \MC_ARK_ARC_1_0/temp1[48] ,
         \MC_ARK_ARC_1_0/temp1[47] , \MC_ARK_ARC_1_0/temp1[46] ,
         \MC_ARK_ARC_1_0/temp1[45] , \MC_ARK_ARC_1_0/temp1[44] ,
         \MC_ARK_ARC_1_0/temp1[43] , \MC_ARK_ARC_1_0/temp1[42] ,
         \MC_ARK_ARC_1_0/temp1[41] , \MC_ARK_ARC_1_0/temp1[40] ,
         \MC_ARK_ARC_1_0/temp1[39] , \MC_ARK_ARC_1_0/temp1[38] ,
         \MC_ARK_ARC_1_0/temp1[37] , \MC_ARK_ARC_1_0/temp1[36] ,
         \MC_ARK_ARC_1_0/temp1[35] , \MC_ARK_ARC_1_0/temp1[34] ,
         \MC_ARK_ARC_1_0/temp1[33] , \MC_ARK_ARC_1_0/temp1[32] ,
         \MC_ARK_ARC_1_0/temp1[31] , \MC_ARK_ARC_1_0/temp1[30] ,
         \MC_ARK_ARC_1_0/temp1[29] , \MC_ARK_ARC_1_0/temp1[28] ,
         \MC_ARK_ARC_1_0/temp1[27] , \MC_ARK_ARC_1_0/temp1[26] ,
         \MC_ARK_ARC_1_0/temp1[25] , \MC_ARK_ARC_1_0/temp1[24] ,
         \MC_ARK_ARC_1_0/temp1[23] , \MC_ARK_ARC_1_0/temp1[22] ,
         \MC_ARK_ARC_1_0/temp1[21] , \MC_ARK_ARC_1_0/temp1[20] ,
         \MC_ARK_ARC_1_0/temp1[19] , \MC_ARK_ARC_1_0/temp1[18] ,
         \MC_ARK_ARC_1_0/temp1[17] , \MC_ARK_ARC_1_0/temp1[16] ,
         \MC_ARK_ARC_1_0/temp1[15] , \MC_ARK_ARC_1_0/temp1[14] ,
         \MC_ARK_ARC_1_0/temp1[13] , \MC_ARK_ARC_1_0/temp1[12] ,
         \MC_ARK_ARC_1_0/temp1[11] , \MC_ARK_ARC_1_0/temp1[10] ,
         \MC_ARK_ARC_1_0/temp1[9] , \MC_ARK_ARC_1_0/temp1[8] ,
         \MC_ARK_ARC_1_0/temp1[7] , \MC_ARK_ARC_1_0/temp1[6] ,
         \MC_ARK_ARC_1_0/temp1[5] , \MC_ARK_ARC_1_0/temp1[4] ,
         \MC_ARK_ARC_1_0/temp1[3] , \MC_ARK_ARC_1_0/temp1[2] ,
         \MC_ARK_ARC_1_0/temp1[1] , \MC_ARK_ARC_1_0/temp1[0] ,
         \MC_ARK_ARC_1_0/buf_keyinput[187] ,
         \MC_ARK_ARC_1_0/buf_keyinput[158] ,
         \MC_ARK_ARC_1_0/buf_keyinput[136] , \MC_ARK_ARC_1_0/buf_keyinput[95] ,
         \MC_ARK_ARC_1_0/buf_keyinput[80] , \MC_ARK_ARC_1_0/buf_keyinput[40] ,
         \MC_ARK_ARC_1_0/buf_keyinput[11] ,
         \MC_ARK_ARC_1_0/buf_datainput[191] ,
         \MC_ARK_ARC_1_0/buf_datainput[190] ,
         \MC_ARK_ARC_1_0/buf_datainput[189] ,
         \MC_ARK_ARC_1_0/buf_datainput[188] ,
         \MC_ARK_ARC_1_0/buf_datainput[187] ,
         \MC_ARK_ARC_1_0/buf_datainput[186] ,
         \MC_ARK_ARC_1_0/buf_datainput[185] ,
         \MC_ARK_ARC_1_0/buf_datainput[183] ,
         \MC_ARK_ARC_1_0/buf_datainput[182] ,
         \MC_ARK_ARC_1_0/buf_datainput[181] ,
         \MC_ARK_ARC_1_0/buf_datainput[180] ,
         \MC_ARK_ARC_1_0/buf_datainput[179] ,
         \MC_ARK_ARC_1_0/buf_datainput[177] ,
         \MC_ARK_ARC_1_0/buf_datainput[176] ,
         \MC_ARK_ARC_1_0/buf_datainput[175] ,
         \MC_ARK_ARC_1_0/buf_datainput[173] ,
         \MC_ARK_ARC_1_0/buf_datainput[172] ,
         \MC_ARK_ARC_1_0/buf_datainput[171] ,
         \MC_ARK_ARC_1_0/buf_datainput[168] ,
         \MC_ARK_ARC_1_0/buf_datainput[167] ,
         \MC_ARK_ARC_1_0/buf_datainput[166] ,
         \MC_ARK_ARC_1_0/buf_datainput[164] ,
         \MC_ARK_ARC_1_0/buf_datainput[162] ,
         \MC_ARK_ARC_1_0/buf_datainput[161] ,
         \MC_ARK_ARC_1_0/buf_datainput[160] ,
         \MC_ARK_ARC_1_0/buf_datainput[159] ,
         \MC_ARK_ARC_1_0/buf_datainput[158] ,
         \MC_ARK_ARC_1_0/buf_datainput[155] ,
         \MC_ARK_ARC_1_0/buf_datainput[154] ,
         \MC_ARK_ARC_1_0/buf_datainput[153] ,
         \MC_ARK_ARC_1_0/buf_datainput[151] ,
         \MC_ARK_ARC_1_0/buf_datainput[149] ,
         \MC_ARK_ARC_1_0/buf_datainput[148] ,
         \MC_ARK_ARC_1_0/buf_datainput[147] ,
         \MC_ARK_ARC_1_0/buf_datainput[146] ,
         \MC_ARK_ARC_1_0/buf_datainput[145] ,
         \MC_ARK_ARC_1_0/buf_datainput[144] ,
         \MC_ARK_ARC_1_0/buf_datainput[143] ,
         \MC_ARK_ARC_1_0/buf_datainput[142] ,
         \MC_ARK_ARC_1_0/buf_datainput[141] ,
         \MC_ARK_ARC_1_0/buf_datainput[140] ,
         \MC_ARK_ARC_1_0/buf_datainput[139] ,
         \MC_ARK_ARC_1_0/buf_datainput[138] ,
         \MC_ARK_ARC_1_0/buf_datainput[137] ,
         \MC_ARK_ARC_1_0/buf_datainput[136] ,
         \MC_ARK_ARC_1_0/buf_datainput[135] ,
         \MC_ARK_ARC_1_0/buf_datainput[134] ,
         \MC_ARK_ARC_1_0/buf_datainput[133] ,
         \MC_ARK_ARC_1_0/buf_datainput[132] ,
         \MC_ARK_ARC_1_0/buf_datainput[131] ,
         \MC_ARK_ARC_1_0/buf_datainput[130] ,
         \MC_ARK_ARC_1_0/buf_datainput[129] ,
         \MC_ARK_ARC_1_0/buf_datainput[128] ,
         \MC_ARK_ARC_1_0/buf_datainput[127] ,
         \MC_ARK_ARC_1_0/buf_datainput[126] ,
         \MC_ARK_ARC_1_0/buf_datainput[125] ,
         \MC_ARK_ARC_1_0/buf_datainput[124] ,
         \MC_ARK_ARC_1_0/buf_datainput[122] ,
         \MC_ARK_ARC_1_0/buf_datainput[121] ,
         \MC_ARK_ARC_1_0/buf_datainput[120] ,
         \MC_ARK_ARC_1_0/buf_datainput[119] ,
         \MC_ARK_ARC_1_0/buf_datainput[118] ,
         \MC_ARK_ARC_1_0/buf_datainput[117] ,
         \MC_ARK_ARC_1_0/buf_datainput[116] ,
         \MC_ARK_ARC_1_0/buf_datainput[115] ,
         \MC_ARK_ARC_1_0/buf_datainput[114] ,
         \MC_ARK_ARC_1_0/buf_datainput[113] ,
         \MC_ARK_ARC_1_0/buf_datainput[111] ,
         \MC_ARK_ARC_1_0/buf_datainput[110] ,
         \MC_ARK_ARC_1_0/buf_datainput[109] ,
         \MC_ARK_ARC_1_0/buf_datainput[108] ,
         \MC_ARK_ARC_1_0/buf_datainput[107] ,
         \MC_ARK_ARC_1_0/buf_datainput[106] ,
         \MC_ARK_ARC_1_0/buf_datainput[105] ,
         \MC_ARK_ARC_1_0/buf_datainput[104] ,
         \MC_ARK_ARC_1_0/buf_datainput[103] ,
         \MC_ARK_ARC_1_0/buf_datainput[102] ,
         \MC_ARK_ARC_1_0/buf_datainput[101] ,
         \MC_ARK_ARC_1_0/buf_datainput[100] ,
         \MC_ARK_ARC_1_0/buf_datainput[99] ,
         \MC_ARK_ARC_1_0/buf_datainput[98] ,
         \MC_ARK_ARC_1_0/buf_datainput[97] ,
         \MC_ARK_ARC_1_0/buf_datainput[96] ,
         \MC_ARK_ARC_1_0/buf_datainput[95] ,
         \MC_ARK_ARC_1_0/buf_datainput[94] ,
         \MC_ARK_ARC_1_0/buf_datainput[93] ,
         \MC_ARK_ARC_1_0/buf_datainput[92] ,
         \MC_ARK_ARC_1_0/buf_datainput[91] ,
         \MC_ARK_ARC_1_0/buf_datainput[90] ,
         \MC_ARK_ARC_1_0/buf_datainput[89] ,
         \MC_ARK_ARC_1_0/buf_datainput[88] ,
         \MC_ARK_ARC_1_0/buf_datainput[87] ,
         \MC_ARK_ARC_1_0/buf_datainput[86] ,
         \MC_ARK_ARC_1_0/buf_datainput[85] ,
         \MC_ARK_ARC_1_0/buf_datainput[84] ,
         \MC_ARK_ARC_1_0/buf_datainput[83] ,
         \MC_ARK_ARC_1_0/buf_datainput[82] ,
         \MC_ARK_ARC_1_0/buf_datainput[81] ,
         \MC_ARK_ARC_1_0/buf_datainput[80] ,
         \MC_ARK_ARC_1_0/buf_datainput[79] ,
         \MC_ARK_ARC_1_0/buf_datainput[78] ,
         \MC_ARK_ARC_1_0/buf_datainput[77] ,
         \MC_ARK_ARC_1_0/buf_datainput[75] ,
         \MC_ARK_ARC_1_0/buf_datainput[74] ,
         \MC_ARK_ARC_1_0/buf_datainput[73] ,
         \MC_ARK_ARC_1_0/buf_datainput[72] ,
         \MC_ARK_ARC_1_0/buf_datainput[71] ,
         \MC_ARK_ARC_1_0/buf_datainput[70] ,
         \MC_ARK_ARC_1_0/buf_datainput[69] ,
         \MC_ARK_ARC_1_0/buf_datainput[68] ,
         \MC_ARK_ARC_1_0/buf_datainput[67] ,
         \MC_ARK_ARC_1_0/buf_datainput[66] ,
         \MC_ARK_ARC_1_0/buf_datainput[65] ,
         \MC_ARK_ARC_1_0/buf_datainput[64] ,
         \MC_ARK_ARC_1_0/buf_datainput[61] ,
         \MC_ARK_ARC_1_0/buf_datainput[59] ,
         \MC_ARK_ARC_1_0/buf_datainput[58] ,
         \MC_ARK_ARC_1_0/buf_datainput[57] ,
         \MC_ARK_ARC_1_0/buf_datainput[56] ,
         \MC_ARK_ARC_1_0/buf_datainput[55] ,
         \MC_ARK_ARC_1_0/buf_datainput[54] ,
         \MC_ARK_ARC_1_0/buf_datainput[53] ,
         \MC_ARK_ARC_1_0/buf_datainput[52] ,
         \MC_ARK_ARC_1_0/buf_datainput[51] ,
         \MC_ARK_ARC_1_0/buf_datainput[50] ,
         \MC_ARK_ARC_1_0/buf_datainput[49] ,
         \MC_ARK_ARC_1_0/buf_datainput[48] ,
         \MC_ARK_ARC_1_0/buf_datainput[47] ,
         \MC_ARK_ARC_1_0/buf_datainput[46] ,
         \MC_ARK_ARC_1_0/buf_datainput[44] ,
         \MC_ARK_ARC_1_0/buf_datainput[43] ,
         \MC_ARK_ARC_1_0/buf_datainput[42] ,
         \MC_ARK_ARC_1_0/buf_datainput[41] ,
         \MC_ARK_ARC_1_0/buf_datainput[40] ,
         \MC_ARK_ARC_1_0/buf_datainput[39] ,
         \MC_ARK_ARC_1_0/buf_datainput[38] ,
         \MC_ARK_ARC_1_0/buf_datainput[37] ,
         \MC_ARK_ARC_1_0/buf_datainput[36] ,
         \MC_ARK_ARC_1_0/buf_datainput[35] ,
         \MC_ARK_ARC_1_0/buf_datainput[34] ,
         \MC_ARK_ARC_1_0/buf_datainput[33] ,
         \MC_ARK_ARC_1_0/buf_datainput[32] ,
         \MC_ARK_ARC_1_0/buf_datainput[31] ,
         \MC_ARK_ARC_1_0/buf_datainput[30] ,
         \MC_ARK_ARC_1_0/buf_datainput[29] ,
         \MC_ARK_ARC_1_0/buf_datainput[28] ,
         \MC_ARK_ARC_1_0/buf_datainput[27] ,
         \MC_ARK_ARC_1_0/buf_datainput[26] ,
         \MC_ARK_ARC_1_0/buf_datainput[25] ,
         \MC_ARK_ARC_1_0/buf_datainput[24] ,
         \MC_ARK_ARC_1_0/buf_datainput[23] ,
         \MC_ARK_ARC_1_0/buf_datainput[22] ,
         \MC_ARK_ARC_1_0/buf_datainput[21] ,
         \MC_ARK_ARC_1_0/buf_datainput[20] ,
         \MC_ARK_ARC_1_0/buf_datainput[19] ,
         \MC_ARK_ARC_1_0/buf_datainput[18] ,
         \MC_ARK_ARC_1_0/buf_datainput[17] ,
         \MC_ARK_ARC_1_0/buf_datainput[16] ,
         \MC_ARK_ARC_1_0/buf_datainput[15] ,
         \MC_ARK_ARC_1_0/buf_datainput[14] ,
         \MC_ARK_ARC_1_0/buf_datainput[13] ,
         \MC_ARK_ARC_1_0/buf_datainput[12] ,
         \MC_ARK_ARC_1_0/buf_datainput[11] ,
         \MC_ARK_ARC_1_0/buf_datainput[10] , \MC_ARK_ARC_1_0/buf_datainput[9] ,
         \MC_ARK_ARC_1_0/buf_datainput[8] , \MC_ARK_ARC_1_0/buf_datainput[7] ,
         \MC_ARK_ARC_1_0/buf_datainput[6] , \MC_ARK_ARC_1_0/buf_datainput[5] ,
         \MC_ARK_ARC_1_0/buf_datainput[4] , \MC_ARK_ARC_1_0/buf_datainput[3] ,
         \MC_ARK_ARC_1_0/buf_datainput[0] , \MC_ARK_ARC_1_1/temp6[190] ,
         \MC_ARK_ARC_1_1/temp6[187] , \MC_ARK_ARC_1_1/temp6[186] ,
         \MC_ARK_ARC_1_1/temp6[184] , \MC_ARK_ARC_1_1/temp6[183] ,
         \MC_ARK_ARC_1_1/temp6[182] , \MC_ARK_ARC_1_1/temp6[181] ,
         \MC_ARK_ARC_1_1/temp6[180] , \MC_ARK_ARC_1_1/temp6[178] ,
         \MC_ARK_ARC_1_1/temp6[176] , \MC_ARK_ARC_1_1/temp6[175] ,
         \MC_ARK_ARC_1_1/temp6[174] , \MC_ARK_ARC_1_1/temp6[173] ,
         \MC_ARK_ARC_1_1/temp6[172] , \MC_ARK_ARC_1_1/temp6[171] ,
         \MC_ARK_ARC_1_1/temp6[170] , \MC_ARK_ARC_1_1/temp6[169] ,
         \MC_ARK_ARC_1_1/temp6[168] , \MC_ARK_ARC_1_1/temp6[167] ,
         \MC_ARK_ARC_1_1/temp6[166] , \MC_ARK_ARC_1_1/temp6[165] ,
         \MC_ARK_ARC_1_1/temp6[164] , \MC_ARK_ARC_1_1/temp6[163] ,
         \MC_ARK_ARC_1_1/temp6[162] , \MC_ARK_ARC_1_1/temp6[161] ,
         \MC_ARK_ARC_1_1/temp6[160] , \MC_ARK_ARC_1_1/temp6[158] ,
         \MC_ARK_ARC_1_1/temp6[157] , \MC_ARK_ARC_1_1/temp6[156] ,
         \MC_ARK_ARC_1_1/temp6[154] , \MC_ARK_ARC_1_1/temp6[153] ,
         \MC_ARK_ARC_1_1/temp6[152] , \MC_ARK_ARC_1_1/temp6[151] ,
         \MC_ARK_ARC_1_1/temp6[150] , \MC_ARK_ARC_1_1/temp6[148] ,
         \MC_ARK_ARC_1_1/temp6[147] , \MC_ARK_ARC_1_1/temp6[146] ,
         \MC_ARK_ARC_1_1/temp6[145] , \MC_ARK_ARC_1_1/temp6[144] ,
         \MC_ARK_ARC_1_1/temp6[142] , \MC_ARK_ARC_1_1/temp6[141] ,
         \MC_ARK_ARC_1_1/temp6[140] , \MC_ARK_ARC_1_1/temp6[139] ,
         \MC_ARK_ARC_1_1/temp6[138] , \MC_ARK_ARC_1_1/temp6[137] ,
         \MC_ARK_ARC_1_1/temp6[136] , \MC_ARK_ARC_1_1/temp6[135] ,
         \MC_ARK_ARC_1_1/temp6[133] , \MC_ARK_ARC_1_1/temp6[132] ,
         \MC_ARK_ARC_1_1/temp6[131] , \MC_ARK_ARC_1_1/temp6[130] ,
         \MC_ARK_ARC_1_1/temp6[129] , \MC_ARK_ARC_1_1/temp6[128] ,
         \MC_ARK_ARC_1_1/temp6[127] , \MC_ARK_ARC_1_1/temp6[126] ,
         \MC_ARK_ARC_1_1/temp6[125] , \MC_ARK_ARC_1_1/temp6[124] ,
         \MC_ARK_ARC_1_1/temp6[123] , \MC_ARK_ARC_1_1/temp6[122] ,
         \MC_ARK_ARC_1_1/temp6[121] , \MC_ARK_ARC_1_1/temp6[120] ,
         \MC_ARK_ARC_1_1/temp6[119] , \MC_ARK_ARC_1_1/temp6[118] ,
         \MC_ARK_ARC_1_1/temp6[117] , \MC_ARK_ARC_1_1/temp6[116] ,
         \MC_ARK_ARC_1_1/temp6[115] , \MC_ARK_ARC_1_1/temp6[114] ,
         \MC_ARK_ARC_1_1/temp6[113] , \MC_ARK_ARC_1_1/temp6[112] ,
         \MC_ARK_ARC_1_1/temp6[111] , \MC_ARK_ARC_1_1/temp6[109] ,
         \MC_ARK_ARC_1_1/temp6[108] , \MC_ARK_ARC_1_1/temp6[106] ,
         \MC_ARK_ARC_1_1/temp6[103] , \MC_ARK_ARC_1_1/temp6[102] ,
         \MC_ARK_ARC_1_1/temp6[101] , \MC_ARK_ARC_1_1/temp6[100] ,
         \MC_ARK_ARC_1_1/temp6[99] , \MC_ARK_ARC_1_1/temp6[98] ,
         \MC_ARK_ARC_1_1/temp6[97] , \MC_ARK_ARC_1_1/temp6[96] ,
         \MC_ARK_ARC_1_1/temp6[95] , \MC_ARK_ARC_1_1/temp6[93] ,
         \MC_ARK_ARC_1_1/temp6[92] , \MC_ARK_ARC_1_1/temp6[91] ,
         \MC_ARK_ARC_1_1/temp6[90] , \MC_ARK_ARC_1_1/temp6[88] ,
         \MC_ARK_ARC_1_1/temp6[87] , \MC_ARK_ARC_1_1/temp6[86] ,
         \MC_ARK_ARC_1_1/temp6[85] , \MC_ARK_ARC_1_1/temp6[84] ,
         \MC_ARK_ARC_1_1/temp6[82] , \MC_ARK_ARC_1_1/temp6[81] ,
         \MC_ARK_ARC_1_1/temp6[80] , \MC_ARK_ARC_1_1/temp6[79] ,
         \MC_ARK_ARC_1_1/temp6[78] , \MC_ARK_ARC_1_1/temp6[76] ,
         \MC_ARK_ARC_1_1/temp6[75] , \MC_ARK_ARC_1_1/temp6[74] ,
         \MC_ARK_ARC_1_1/temp6[73] , \MC_ARK_ARC_1_1/temp6[72] ,
         \MC_ARK_ARC_1_1/temp6[70] , \MC_ARK_ARC_1_1/temp6[69] ,
         \MC_ARK_ARC_1_1/temp6[68] , \MC_ARK_ARC_1_1/temp6[67] ,
         \MC_ARK_ARC_1_1/temp6[66] , \MC_ARK_ARC_1_1/temp6[64] ,
         \MC_ARK_ARC_1_1/temp6[63] , \MC_ARK_ARC_1_1/temp6[62] ,
         \MC_ARK_ARC_1_1/temp6[61] , \MC_ARK_ARC_1_1/temp6[60] ,
         \MC_ARK_ARC_1_1/temp6[59] , \MC_ARK_ARC_1_1/temp6[57] ,
         \MC_ARK_ARC_1_1/temp6[56] , \MC_ARK_ARC_1_1/temp6[55] ,
         \MC_ARK_ARC_1_1/temp6[54] , \MC_ARK_ARC_1_1/temp6[52] ,
         \MC_ARK_ARC_1_1/temp6[51] , \MC_ARK_ARC_1_1/temp6[50] ,
         \MC_ARK_ARC_1_1/temp6[49] , \MC_ARK_ARC_1_1/temp6[48] ,
         \MC_ARK_ARC_1_1/temp6[47] , \MC_ARK_ARC_1_1/temp6[46] ,
         \MC_ARK_ARC_1_1/temp6[45] , \MC_ARK_ARC_1_1/temp6[44] ,
         \MC_ARK_ARC_1_1/temp6[43] , \MC_ARK_ARC_1_1/temp6[42] ,
         \MC_ARK_ARC_1_1/temp6[41] , \MC_ARK_ARC_1_1/temp6[40] ,
         \MC_ARK_ARC_1_1/temp6[38] , \MC_ARK_ARC_1_1/temp6[37] ,
         \MC_ARK_ARC_1_1/temp6[36] , \MC_ARK_ARC_1_1/temp6[34] ,
         \MC_ARK_ARC_1_1/temp6[33] , \MC_ARK_ARC_1_1/temp6[32] ,
         \MC_ARK_ARC_1_1/temp6[31] , \MC_ARK_ARC_1_1/temp6[30] ,
         \MC_ARK_ARC_1_1/temp6[28] , \MC_ARK_ARC_1_1/temp6[27] ,
         \MC_ARK_ARC_1_1/temp6[26] , \MC_ARK_ARC_1_1/temp6[25] ,
         \MC_ARK_ARC_1_1/temp6[24] , \MC_ARK_ARC_1_1/temp6[23] ,
         \MC_ARK_ARC_1_1/temp6[22] , \MC_ARK_ARC_1_1/temp6[20] ,
         \MC_ARK_ARC_1_1/temp6[19] , \MC_ARK_ARC_1_1/temp6[18] ,
         \MC_ARK_ARC_1_1/temp6[16] , \MC_ARK_ARC_1_1/temp6[15] ,
         \MC_ARK_ARC_1_1/temp6[14] , \MC_ARK_ARC_1_1/temp6[13] ,
         \MC_ARK_ARC_1_1/temp6[12] , \MC_ARK_ARC_1_1/temp6[11] ,
         \MC_ARK_ARC_1_1/temp6[10] , \MC_ARK_ARC_1_1/temp6[9] ,
         \MC_ARK_ARC_1_1/temp6[8] , \MC_ARK_ARC_1_1/temp6[7] ,
         \MC_ARK_ARC_1_1/temp6[6] , \MC_ARK_ARC_1_1/temp6[5] ,
         \MC_ARK_ARC_1_1/temp6[4] , \MC_ARK_ARC_1_1/temp6[3] ,
         \MC_ARK_ARC_1_1/temp6[2] , \MC_ARK_ARC_1_1/temp6[1] ,
         \MC_ARK_ARC_1_1/temp6[0] , \MC_ARK_ARC_1_1/temp5[190] ,
         \MC_ARK_ARC_1_1/temp5[188] , \MC_ARK_ARC_1_1/temp5[187] ,
         \MC_ARK_ARC_1_1/temp5[186] , \MC_ARK_ARC_1_1/temp5[184] ,
         \MC_ARK_ARC_1_1/temp5[183] , \MC_ARK_ARC_1_1/temp5[182] ,
         \MC_ARK_ARC_1_1/temp5[181] , \MC_ARK_ARC_1_1/temp5[180] ,
         \MC_ARK_ARC_1_1/temp5[178] , \MC_ARK_ARC_1_1/temp5[176] ,
         \MC_ARK_ARC_1_1/temp5[175] , \MC_ARK_ARC_1_1/temp5[174] ,
         \MC_ARK_ARC_1_1/temp5[173] , \MC_ARK_ARC_1_1/temp5[172] ,
         \MC_ARK_ARC_1_1/temp5[171] , \MC_ARK_ARC_1_1/temp5[170] ,
         \MC_ARK_ARC_1_1/temp5[169] , \MC_ARK_ARC_1_1/temp5[168] ,
         \MC_ARK_ARC_1_1/temp5[167] , \MC_ARK_ARC_1_1/temp5[166] ,
         \MC_ARK_ARC_1_1/temp5[165] , \MC_ARK_ARC_1_1/temp5[164] ,
         \MC_ARK_ARC_1_1/temp5[163] , \MC_ARK_ARC_1_1/temp5[162] ,
         \MC_ARK_ARC_1_1/temp5[161] , \MC_ARK_ARC_1_1/temp5[160] ,
         \MC_ARK_ARC_1_1/temp5[159] , \MC_ARK_ARC_1_1/temp5[157] ,
         \MC_ARK_ARC_1_1/temp5[156] , \MC_ARK_ARC_1_1/temp5[154] ,
         \MC_ARK_ARC_1_1/temp5[153] , \MC_ARK_ARC_1_1/temp5[152] ,
         \MC_ARK_ARC_1_1/temp5[151] , \MC_ARK_ARC_1_1/temp5[150] ,
         \MC_ARK_ARC_1_1/temp5[148] , \MC_ARK_ARC_1_1/temp5[147] ,
         \MC_ARK_ARC_1_1/temp5[146] , \MC_ARK_ARC_1_1/temp5[145] ,
         \MC_ARK_ARC_1_1/temp5[144] , \MC_ARK_ARC_1_1/temp5[142] ,
         \MC_ARK_ARC_1_1/temp5[141] , \MC_ARK_ARC_1_1/temp5[140] ,
         \MC_ARK_ARC_1_1/temp5[139] , \MC_ARK_ARC_1_1/temp5[138] ,
         \MC_ARK_ARC_1_1/temp5[137] , \MC_ARK_ARC_1_1/temp5[136] ,
         \MC_ARK_ARC_1_1/temp5[135] , \MC_ARK_ARC_1_1/temp5[134] ,
         \MC_ARK_ARC_1_1/temp5[133] , \MC_ARK_ARC_1_1/temp5[132] ,
         \MC_ARK_ARC_1_1/temp5[131] , \MC_ARK_ARC_1_1/temp5[130] ,
         \MC_ARK_ARC_1_1/temp5[129] , \MC_ARK_ARC_1_1/temp5[127] ,
         \MC_ARK_ARC_1_1/temp5[126] , \MC_ARK_ARC_1_1/temp5[124] ,
         \MC_ARK_ARC_1_1/temp5[123] , \MC_ARK_ARC_1_1/temp5[122] ,
         \MC_ARK_ARC_1_1/temp5[121] , \MC_ARK_ARC_1_1/temp5[120] ,
         \MC_ARK_ARC_1_1/temp5[119] , \MC_ARK_ARC_1_1/temp5[118] ,
         \MC_ARK_ARC_1_1/temp5[117] , \MC_ARK_ARC_1_1/temp5[116] ,
         \MC_ARK_ARC_1_1/temp5[115] , \MC_ARK_ARC_1_1/temp5[114] ,
         \MC_ARK_ARC_1_1/temp5[113] , \MC_ARK_ARC_1_1/temp5[112] ,
         \MC_ARK_ARC_1_1/temp5[111] , \MC_ARK_ARC_1_1/temp5[110] ,
         \MC_ARK_ARC_1_1/temp5[109] , \MC_ARK_ARC_1_1/temp5[108] ,
         \MC_ARK_ARC_1_1/temp5[106] , \MC_ARK_ARC_1_1/temp5[105] ,
         \MC_ARK_ARC_1_1/temp5[103] , \MC_ARK_ARC_1_1/temp5[102] ,
         \MC_ARK_ARC_1_1/temp5[101] , \MC_ARK_ARC_1_1/temp5[100] ,
         \MC_ARK_ARC_1_1/temp5[99] , \MC_ARK_ARC_1_1/temp5[98] ,
         \MC_ARK_ARC_1_1/temp5[97] , \MC_ARK_ARC_1_1/temp5[96] ,
         \MC_ARK_ARC_1_1/temp5[95] , \MC_ARK_ARC_1_1/temp5[94] ,
         \MC_ARK_ARC_1_1/temp5[93] , \MC_ARK_ARC_1_1/temp5[92] ,
         \MC_ARK_ARC_1_1/temp5[91] , \MC_ARK_ARC_1_1/temp5[90] ,
         \MC_ARK_ARC_1_1/temp5[88] , \MC_ARK_ARC_1_1/temp5[87] ,
         \MC_ARK_ARC_1_1/temp5[86] , \MC_ARK_ARC_1_1/temp5[85] ,
         \MC_ARK_ARC_1_1/temp5[84] , \MC_ARK_ARC_1_1/temp5[82] ,
         \MC_ARK_ARC_1_1/temp5[81] , \MC_ARK_ARC_1_1/temp5[80] ,
         \MC_ARK_ARC_1_1/temp5[79] , \MC_ARK_ARC_1_1/temp5[78] ,
         \MC_ARK_ARC_1_1/temp5[76] , \MC_ARK_ARC_1_1/temp5[75] ,
         \MC_ARK_ARC_1_1/temp5[74] , \MC_ARK_ARC_1_1/temp5[73] ,
         \MC_ARK_ARC_1_1/temp5[72] , \MC_ARK_ARC_1_1/temp5[70] ,
         \MC_ARK_ARC_1_1/temp5[69] , \MC_ARK_ARC_1_1/temp5[68] ,
         \MC_ARK_ARC_1_1/temp5[67] , \MC_ARK_ARC_1_1/temp5[66] ,
         \MC_ARK_ARC_1_1/temp5[64] , \MC_ARK_ARC_1_1/temp5[62] ,
         \MC_ARK_ARC_1_1/temp5[61] , \MC_ARK_ARC_1_1/temp5[60] ,
         \MC_ARK_ARC_1_1/temp5[57] , \MC_ARK_ARC_1_1/temp5[56] ,
         \MC_ARK_ARC_1_1/temp5[55] , \MC_ARK_ARC_1_1/temp5[54] ,
         \MC_ARK_ARC_1_1/temp5[52] , \MC_ARK_ARC_1_1/temp5[50] ,
         \MC_ARK_ARC_1_1/temp5[49] , \MC_ARK_ARC_1_1/temp5[48] ,
         \MC_ARK_ARC_1_1/temp5[47] , \MC_ARK_ARC_1_1/temp5[46] ,
         \MC_ARK_ARC_1_1/temp5[45] , \MC_ARK_ARC_1_1/temp5[44] ,
         \MC_ARK_ARC_1_1/temp5[43] , \MC_ARK_ARC_1_1/temp5[42] ,
         \MC_ARK_ARC_1_1/temp5[41] , \MC_ARK_ARC_1_1/temp5[40] ,
         \MC_ARK_ARC_1_1/temp5[39] , \MC_ARK_ARC_1_1/temp5[38] ,
         \MC_ARK_ARC_1_1/temp5[37] , \MC_ARK_ARC_1_1/temp5[36] ,
         \MC_ARK_ARC_1_1/temp5[34] , \MC_ARK_ARC_1_1/temp5[33] ,
         \MC_ARK_ARC_1_1/temp5[32] , \MC_ARK_ARC_1_1/temp5[31] ,
         \MC_ARK_ARC_1_1/temp5[30] , \MC_ARK_ARC_1_1/temp5[28] ,
         \MC_ARK_ARC_1_1/temp5[27] , \MC_ARK_ARC_1_1/temp5[26] ,
         \MC_ARK_ARC_1_1/temp5[25] , \MC_ARK_ARC_1_1/temp5[24] ,
         \MC_ARK_ARC_1_1/temp5[23] , \MC_ARK_ARC_1_1/temp5[22] ,
         \MC_ARK_ARC_1_1/temp5[21] , \MC_ARK_ARC_1_1/temp5[20] ,
         \MC_ARK_ARC_1_1/temp5[19] , \MC_ARK_ARC_1_1/temp5[18] ,
         \MC_ARK_ARC_1_1/temp5[16] , \MC_ARK_ARC_1_1/temp5[15] ,
         \MC_ARK_ARC_1_1/temp5[14] , \MC_ARK_ARC_1_1/temp5[13] ,
         \MC_ARK_ARC_1_1/temp5[12] , \MC_ARK_ARC_1_1/temp5[11] ,
         \MC_ARK_ARC_1_1/temp5[10] , \MC_ARK_ARC_1_1/temp5[9] ,
         \MC_ARK_ARC_1_1/temp5[8] , \MC_ARK_ARC_1_1/temp5[7] ,
         \MC_ARK_ARC_1_1/temp5[6] , \MC_ARK_ARC_1_1/temp5[5] ,
         \MC_ARK_ARC_1_1/temp5[4] , \MC_ARK_ARC_1_1/temp5[3] ,
         \MC_ARK_ARC_1_1/temp5[2] , \MC_ARK_ARC_1_1/temp5[1] ,
         \MC_ARK_ARC_1_1/temp5[0] , \MC_ARK_ARC_1_1/temp4[191] ,
         \MC_ARK_ARC_1_1/temp4[190] , \MC_ARK_ARC_1_1/temp4[189] ,
         \MC_ARK_ARC_1_1/temp4[188] , \MC_ARK_ARC_1_1/temp4[187] ,
         \MC_ARK_ARC_1_1/temp4[186] , \MC_ARK_ARC_1_1/temp4[185] ,
         \MC_ARK_ARC_1_1/temp4[184] , \MC_ARK_ARC_1_1/temp4[183] ,
         \MC_ARK_ARC_1_1/temp4[182] , \MC_ARK_ARC_1_1/temp4[181] ,
         \MC_ARK_ARC_1_1/temp4[180] , \MC_ARK_ARC_1_1/temp4[179] ,
         \MC_ARK_ARC_1_1/temp4[178] , \MC_ARK_ARC_1_1/temp4[177] ,
         \MC_ARK_ARC_1_1/temp4[176] , \MC_ARK_ARC_1_1/temp4[175] ,
         \MC_ARK_ARC_1_1/temp4[174] , \MC_ARK_ARC_1_1/temp4[173] ,
         \MC_ARK_ARC_1_1/temp4[172] , \MC_ARK_ARC_1_1/temp4[171] ,
         \MC_ARK_ARC_1_1/temp4[170] , \MC_ARK_ARC_1_1/temp4[169] ,
         \MC_ARK_ARC_1_1/temp4[168] , \MC_ARK_ARC_1_1/temp4[167] ,
         \MC_ARK_ARC_1_1/temp4[166] , \MC_ARK_ARC_1_1/temp4[165] ,
         \MC_ARK_ARC_1_1/temp4[164] , \MC_ARK_ARC_1_1/temp4[163] ,
         \MC_ARK_ARC_1_1/temp4[162] , \MC_ARK_ARC_1_1/temp4[161] ,
         \MC_ARK_ARC_1_1/temp4[160] , \MC_ARK_ARC_1_1/temp4[159] ,
         \MC_ARK_ARC_1_1/temp4[158] , \MC_ARK_ARC_1_1/temp4[157] ,
         \MC_ARK_ARC_1_1/temp4[156] , \MC_ARK_ARC_1_1/temp4[155] ,
         \MC_ARK_ARC_1_1/temp4[154] , \MC_ARK_ARC_1_1/temp4[153] ,
         \MC_ARK_ARC_1_1/temp4[152] , \MC_ARK_ARC_1_1/temp4[151] ,
         \MC_ARK_ARC_1_1/temp4[150] , \MC_ARK_ARC_1_1/temp4[149] ,
         \MC_ARK_ARC_1_1/temp4[148] , \MC_ARK_ARC_1_1/temp4[147] ,
         \MC_ARK_ARC_1_1/temp4[146] , \MC_ARK_ARC_1_1/temp4[145] ,
         \MC_ARK_ARC_1_1/temp4[144] , \MC_ARK_ARC_1_1/temp4[143] ,
         \MC_ARK_ARC_1_1/temp4[142] , \MC_ARK_ARC_1_1/temp4[141] ,
         \MC_ARK_ARC_1_1/temp4[140] , \MC_ARK_ARC_1_1/temp4[139] ,
         \MC_ARK_ARC_1_1/temp4[138] , \MC_ARK_ARC_1_1/temp4[137] ,
         \MC_ARK_ARC_1_1/temp4[136] , \MC_ARK_ARC_1_1/temp4[135] ,
         \MC_ARK_ARC_1_1/temp4[134] , \MC_ARK_ARC_1_1/temp4[133] ,
         \MC_ARK_ARC_1_1/temp4[132] , \MC_ARK_ARC_1_1/temp4[131] ,
         \MC_ARK_ARC_1_1/temp4[130] , \MC_ARK_ARC_1_1/temp4[129] ,
         \MC_ARK_ARC_1_1/temp4[128] , \MC_ARK_ARC_1_1/temp4[127] ,
         \MC_ARK_ARC_1_1/temp4[126] , \MC_ARK_ARC_1_1/temp4[125] ,
         \MC_ARK_ARC_1_1/temp4[124] , \MC_ARK_ARC_1_1/temp4[123] ,
         \MC_ARK_ARC_1_1/temp4[122] , \MC_ARK_ARC_1_1/temp4[121] ,
         \MC_ARK_ARC_1_1/temp4[120] , \MC_ARK_ARC_1_1/temp4[119] ,
         \MC_ARK_ARC_1_1/temp4[118] , \MC_ARK_ARC_1_1/temp4[117] ,
         \MC_ARK_ARC_1_1/temp4[116] , \MC_ARK_ARC_1_1/temp4[115] ,
         \MC_ARK_ARC_1_1/temp4[114] , \MC_ARK_ARC_1_1/temp4[113] ,
         \MC_ARK_ARC_1_1/temp4[112] , \MC_ARK_ARC_1_1/temp4[111] ,
         \MC_ARK_ARC_1_1/temp4[110] , \MC_ARK_ARC_1_1/temp4[109] ,
         \MC_ARK_ARC_1_1/temp4[108] , \MC_ARK_ARC_1_1/temp4[107] ,
         \MC_ARK_ARC_1_1/temp4[106] , \MC_ARK_ARC_1_1/temp4[105] ,
         \MC_ARK_ARC_1_1/temp4[104] , \MC_ARK_ARC_1_1/temp4[103] ,
         \MC_ARK_ARC_1_1/temp4[102] , \MC_ARK_ARC_1_1/temp4[101] ,
         \MC_ARK_ARC_1_1/temp4[100] , \MC_ARK_ARC_1_1/temp4[99] ,
         \MC_ARK_ARC_1_1/temp4[98] , \MC_ARK_ARC_1_1/temp4[97] ,
         \MC_ARK_ARC_1_1/temp4[96] , \MC_ARK_ARC_1_1/temp4[95] ,
         \MC_ARK_ARC_1_1/temp4[94] , \MC_ARK_ARC_1_1/temp4[93] ,
         \MC_ARK_ARC_1_1/temp4[92] , \MC_ARK_ARC_1_1/temp4[91] ,
         \MC_ARK_ARC_1_1/temp4[90] , \MC_ARK_ARC_1_1/temp4[89] ,
         \MC_ARK_ARC_1_1/temp4[88] , \MC_ARK_ARC_1_1/temp4[87] ,
         \MC_ARK_ARC_1_1/temp4[86] , \MC_ARK_ARC_1_1/temp4[85] ,
         \MC_ARK_ARC_1_1/temp4[84] , \MC_ARK_ARC_1_1/temp4[83] ,
         \MC_ARK_ARC_1_1/temp4[82] , \MC_ARK_ARC_1_1/temp4[81] ,
         \MC_ARK_ARC_1_1/temp4[80] , \MC_ARK_ARC_1_1/temp4[79] ,
         \MC_ARK_ARC_1_1/temp4[78] , \MC_ARK_ARC_1_1/temp4[77] ,
         \MC_ARK_ARC_1_1/temp4[76] , \MC_ARK_ARC_1_1/temp4[75] ,
         \MC_ARK_ARC_1_1/temp4[74] , \MC_ARK_ARC_1_1/temp4[73] ,
         \MC_ARK_ARC_1_1/temp4[72] , \MC_ARK_ARC_1_1/temp4[71] ,
         \MC_ARK_ARC_1_1/temp4[70] , \MC_ARK_ARC_1_1/temp4[69] ,
         \MC_ARK_ARC_1_1/temp4[68] , \MC_ARK_ARC_1_1/temp4[67] ,
         \MC_ARK_ARC_1_1/temp4[66] , \MC_ARK_ARC_1_1/temp4[65] ,
         \MC_ARK_ARC_1_1/temp4[64] , \MC_ARK_ARC_1_1/temp4[63] ,
         \MC_ARK_ARC_1_1/temp4[62] , \MC_ARK_ARC_1_1/temp4[61] ,
         \MC_ARK_ARC_1_1/temp4[60] , \MC_ARK_ARC_1_1/temp4[59] ,
         \MC_ARK_ARC_1_1/temp4[58] , \MC_ARK_ARC_1_1/temp4[57] ,
         \MC_ARK_ARC_1_1/temp4[56] , \MC_ARK_ARC_1_1/temp4[55] ,
         \MC_ARK_ARC_1_1/temp4[54] , \MC_ARK_ARC_1_1/temp4[53] ,
         \MC_ARK_ARC_1_1/temp4[52] , \MC_ARK_ARC_1_1/temp4[51] ,
         \MC_ARK_ARC_1_1/temp4[50] , \MC_ARK_ARC_1_1/temp4[49] ,
         \MC_ARK_ARC_1_1/temp4[48] , \MC_ARK_ARC_1_1/temp4[47] ,
         \MC_ARK_ARC_1_1/temp4[46] , \MC_ARK_ARC_1_1/temp4[45] ,
         \MC_ARK_ARC_1_1/temp4[44] , \MC_ARK_ARC_1_1/temp4[43] ,
         \MC_ARK_ARC_1_1/temp4[42] , \MC_ARK_ARC_1_1/temp4[41] ,
         \MC_ARK_ARC_1_1/temp4[40] , \MC_ARK_ARC_1_1/temp4[39] ,
         \MC_ARK_ARC_1_1/temp4[38] , \MC_ARK_ARC_1_1/temp4[37] ,
         \MC_ARK_ARC_1_1/temp4[36] , \MC_ARK_ARC_1_1/temp4[35] ,
         \MC_ARK_ARC_1_1/temp4[34] , \MC_ARK_ARC_1_1/temp4[33] ,
         \MC_ARK_ARC_1_1/temp4[32] , \MC_ARK_ARC_1_1/temp4[31] ,
         \MC_ARK_ARC_1_1/temp4[30] , \MC_ARK_ARC_1_1/temp4[29] ,
         \MC_ARK_ARC_1_1/temp4[28] , \MC_ARK_ARC_1_1/temp4[27] ,
         \MC_ARK_ARC_1_1/temp4[26] , \MC_ARK_ARC_1_1/temp4[25] ,
         \MC_ARK_ARC_1_1/temp4[24] , \MC_ARK_ARC_1_1/temp4[23] ,
         \MC_ARK_ARC_1_1/temp4[22] , \MC_ARK_ARC_1_1/temp4[21] ,
         \MC_ARK_ARC_1_1/temp4[20] , \MC_ARK_ARC_1_1/temp4[19] ,
         \MC_ARK_ARC_1_1/temp4[18] , \MC_ARK_ARC_1_1/temp4[17] ,
         \MC_ARK_ARC_1_1/temp4[16] , \MC_ARK_ARC_1_1/temp4[15] ,
         \MC_ARK_ARC_1_1/temp4[14] , \MC_ARK_ARC_1_1/temp4[13] ,
         \MC_ARK_ARC_1_1/temp4[12] , \MC_ARK_ARC_1_1/temp4[11] ,
         \MC_ARK_ARC_1_1/temp4[10] , \MC_ARK_ARC_1_1/temp4[9] ,
         \MC_ARK_ARC_1_1/temp4[8] , \MC_ARK_ARC_1_1/temp4[7] ,
         \MC_ARK_ARC_1_1/temp4[6] , \MC_ARK_ARC_1_1/temp4[5] ,
         \MC_ARK_ARC_1_1/temp4[4] , \MC_ARK_ARC_1_1/temp4[3] ,
         \MC_ARK_ARC_1_1/temp4[2] , \MC_ARK_ARC_1_1/temp4[1] ,
         \MC_ARK_ARC_1_1/temp4[0] , \MC_ARK_ARC_1_1/temp3[191] ,
         \MC_ARK_ARC_1_1/temp3[190] , \MC_ARK_ARC_1_1/temp3[189] ,
         \MC_ARK_ARC_1_1/temp3[188] , \MC_ARK_ARC_1_1/temp3[187] ,
         \MC_ARK_ARC_1_1/temp3[186] , \MC_ARK_ARC_1_1/temp3[185] ,
         \MC_ARK_ARC_1_1/temp3[184] , \MC_ARK_ARC_1_1/temp3[183] ,
         \MC_ARK_ARC_1_1/temp3[182] , \MC_ARK_ARC_1_1/temp3[181] ,
         \MC_ARK_ARC_1_1/temp3[180] , \MC_ARK_ARC_1_1/temp3[179] ,
         \MC_ARK_ARC_1_1/temp3[178] , \MC_ARK_ARC_1_1/temp3[177] ,
         \MC_ARK_ARC_1_1/temp3[176] , \MC_ARK_ARC_1_1/temp3[175] ,
         \MC_ARK_ARC_1_1/temp3[174] , \MC_ARK_ARC_1_1/temp3[173] ,
         \MC_ARK_ARC_1_1/temp3[172] , \MC_ARK_ARC_1_1/temp3[171] ,
         \MC_ARK_ARC_1_1/temp3[170] , \MC_ARK_ARC_1_1/temp3[169] ,
         \MC_ARK_ARC_1_1/temp3[168] , \MC_ARK_ARC_1_1/temp3[167] ,
         \MC_ARK_ARC_1_1/temp3[166] , \MC_ARK_ARC_1_1/temp3[165] ,
         \MC_ARK_ARC_1_1/temp3[164] , \MC_ARK_ARC_1_1/temp3[163] ,
         \MC_ARK_ARC_1_1/temp3[162] , \MC_ARK_ARC_1_1/temp3[161] ,
         \MC_ARK_ARC_1_1/temp3[160] , \MC_ARK_ARC_1_1/temp3[159] ,
         \MC_ARK_ARC_1_1/temp3[158] , \MC_ARK_ARC_1_1/temp3[157] ,
         \MC_ARK_ARC_1_1/temp3[156] , \MC_ARK_ARC_1_1/temp3[155] ,
         \MC_ARK_ARC_1_1/temp3[154] , \MC_ARK_ARC_1_1/temp3[153] ,
         \MC_ARK_ARC_1_1/temp3[152] , \MC_ARK_ARC_1_1/temp3[151] ,
         \MC_ARK_ARC_1_1/temp3[150] , \MC_ARK_ARC_1_1/temp3[149] ,
         \MC_ARK_ARC_1_1/temp3[148] , \MC_ARK_ARC_1_1/temp3[147] ,
         \MC_ARK_ARC_1_1/temp3[146] , \MC_ARK_ARC_1_1/temp3[145] ,
         \MC_ARK_ARC_1_1/temp3[144] , \MC_ARK_ARC_1_1/temp3[143] ,
         \MC_ARK_ARC_1_1/temp3[142] , \MC_ARK_ARC_1_1/temp3[141] ,
         \MC_ARK_ARC_1_1/temp3[140] , \MC_ARK_ARC_1_1/temp3[139] ,
         \MC_ARK_ARC_1_1/temp3[138] , \MC_ARK_ARC_1_1/temp3[137] ,
         \MC_ARK_ARC_1_1/temp3[136] , \MC_ARK_ARC_1_1/temp3[135] ,
         \MC_ARK_ARC_1_1/temp3[134] , \MC_ARK_ARC_1_1/temp3[133] ,
         \MC_ARK_ARC_1_1/temp3[132] , \MC_ARK_ARC_1_1/temp3[131] ,
         \MC_ARK_ARC_1_1/temp3[130] , \MC_ARK_ARC_1_1/temp3[129] ,
         \MC_ARK_ARC_1_1/temp3[128] , \MC_ARK_ARC_1_1/temp3[127] ,
         \MC_ARK_ARC_1_1/temp3[126] , \MC_ARK_ARC_1_1/temp3[125] ,
         \MC_ARK_ARC_1_1/temp3[124] , \MC_ARK_ARC_1_1/temp3[123] ,
         \MC_ARK_ARC_1_1/temp3[122] , \MC_ARK_ARC_1_1/temp3[121] ,
         \MC_ARK_ARC_1_1/temp3[120] , \MC_ARK_ARC_1_1/temp3[119] ,
         \MC_ARK_ARC_1_1/temp3[118] , \MC_ARK_ARC_1_1/temp3[117] ,
         \MC_ARK_ARC_1_1/temp3[116] , \MC_ARK_ARC_1_1/temp3[115] ,
         \MC_ARK_ARC_1_1/temp3[114] , \MC_ARK_ARC_1_1/temp3[113] ,
         \MC_ARK_ARC_1_1/temp3[112] , \MC_ARK_ARC_1_1/temp3[111] ,
         \MC_ARK_ARC_1_1/temp3[110] , \MC_ARK_ARC_1_1/temp3[109] ,
         \MC_ARK_ARC_1_1/temp3[108] , \MC_ARK_ARC_1_1/temp3[107] ,
         \MC_ARK_ARC_1_1/temp3[106] , \MC_ARK_ARC_1_1/temp3[105] ,
         \MC_ARK_ARC_1_1/temp3[104] , \MC_ARK_ARC_1_1/temp3[103] ,
         \MC_ARK_ARC_1_1/temp3[102] , \MC_ARK_ARC_1_1/temp3[101] ,
         \MC_ARK_ARC_1_1/temp3[100] , \MC_ARK_ARC_1_1/temp3[99] ,
         \MC_ARK_ARC_1_1/temp3[98] , \MC_ARK_ARC_1_1/temp3[97] ,
         \MC_ARK_ARC_1_1/temp3[96] , \MC_ARK_ARC_1_1/temp3[95] ,
         \MC_ARK_ARC_1_1/temp3[94] , \MC_ARK_ARC_1_1/temp3[93] ,
         \MC_ARK_ARC_1_1/temp3[92] , \MC_ARK_ARC_1_1/temp3[91] ,
         \MC_ARK_ARC_1_1/temp3[90] , \MC_ARK_ARC_1_1/temp3[89] ,
         \MC_ARK_ARC_1_1/temp3[88] , \MC_ARK_ARC_1_1/temp3[87] ,
         \MC_ARK_ARC_1_1/temp3[86] , \MC_ARK_ARC_1_1/temp3[85] ,
         \MC_ARK_ARC_1_1/temp3[84] , \MC_ARK_ARC_1_1/temp3[83] ,
         \MC_ARK_ARC_1_1/temp3[82] , \MC_ARK_ARC_1_1/temp3[81] ,
         \MC_ARK_ARC_1_1/temp3[80] , \MC_ARK_ARC_1_1/temp3[79] ,
         \MC_ARK_ARC_1_1/temp3[78] , \MC_ARK_ARC_1_1/temp3[77] ,
         \MC_ARK_ARC_1_1/temp3[76] , \MC_ARK_ARC_1_1/temp3[75] ,
         \MC_ARK_ARC_1_1/temp3[74] , \MC_ARK_ARC_1_1/temp3[73] ,
         \MC_ARK_ARC_1_1/temp3[72] , \MC_ARK_ARC_1_1/temp3[71] ,
         \MC_ARK_ARC_1_1/temp3[70] , \MC_ARK_ARC_1_1/temp3[69] ,
         \MC_ARK_ARC_1_1/temp3[68] , \MC_ARK_ARC_1_1/temp3[67] ,
         \MC_ARK_ARC_1_1/temp3[66] , \MC_ARK_ARC_1_1/temp3[65] ,
         \MC_ARK_ARC_1_1/temp3[64] , \MC_ARK_ARC_1_1/temp3[63] ,
         \MC_ARK_ARC_1_1/temp3[62] , \MC_ARK_ARC_1_1/temp3[61] ,
         \MC_ARK_ARC_1_1/temp3[60] , \MC_ARK_ARC_1_1/temp3[59] ,
         \MC_ARK_ARC_1_1/temp3[58] , \MC_ARK_ARC_1_1/temp3[57] ,
         \MC_ARK_ARC_1_1/temp3[56] , \MC_ARK_ARC_1_1/temp3[55] ,
         \MC_ARK_ARC_1_1/temp3[54] , \MC_ARK_ARC_1_1/temp3[53] ,
         \MC_ARK_ARC_1_1/temp3[52] , \MC_ARK_ARC_1_1/temp3[51] ,
         \MC_ARK_ARC_1_1/temp3[50] , \MC_ARK_ARC_1_1/temp3[49] ,
         \MC_ARK_ARC_1_1/temp3[48] , \MC_ARK_ARC_1_1/temp3[47] ,
         \MC_ARK_ARC_1_1/temp3[46] , \MC_ARK_ARC_1_1/temp3[45] ,
         \MC_ARK_ARC_1_1/temp3[44] , \MC_ARK_ARC_1_1/temp3[43] ,
         \MC_ARK_ARC_1_1/temp3[42] , \MC_ARK_ARC_1_1/temp3[41] ,
         \MC_ARK_ARC_1_1/temp3[40] , \MC_ARK_ARC_1_1/temp3[39] ,
         \MC_ARK_ARC_1_1/temp3[38] , \MC_ARK_ARC_1_1/temp3[37] ,
         \MC_ARK_ARC_1_1/temp3[36] , \MC_ARK_ARC_1_1/temp3[35] ,
         \MC_ARK_ARC_1_1/temp3[34] , \MC_ARK_ARC_1_1/temp3[33] ,
         \MC_ARK_ARC_1_1/temp3[32] , \MC_ARK_ARC_1_1/temp3[31] ,
         \MC_ARK_ARC_1_1/temp3[30] , \MC_ARK_ARC_1_1/temp3[29] ,
         \MC_ARK_ARC_1_1/temp3[28] , \MC_ARK_ARC_1_1/temp3[27] ,
         \MC_ARK_ARC_1_1/temp3[26] , \MC_ARK_ARC_1_1/temp3[25] ,
         \MC_ARK_ARC_1_1/temp3[24] , \MC_ARK_ARC_1_1/temp3[23] ,
         \MC_ARK_ARC_1_1/temp3[22] , \MC_ARK_ARC_1_1/temp3[21] ,
         \MC_ARK_ARC_1_1/temp3[20] , \MC_ARK_ARC_1_1/temp3[19] ,
         \MC_ARK_ARC_1_1/temp3[18] , \MC_ARK_ARC_1_1/temp3[17] ,
         \MC_ARK_ARC_1_1/temp3[16] , \MC_ARK_ARC_1_1/temp3[15] ,
         \MC_ARK_ARC_1_1/temp3[14] , \MC_ARK_ARC_1_1/temp3[13] ,
         \MC_ARK_ARC_1_1/temp3[12] , \MC_ARK_ARC_1_1/temp3[10] ,
         \MC_ARK_ARC_1_1/temp3[9] , \MC_ARK_ARC_1_1/temp3[8] ,
         \MC_ARK_ARC_1_1/temp3[7] , \MC_ARK_ARC_1_1/temp3[6] ,
         \MC_ARK_ARC_1_1/temp3[5] , \MC_ARK_ARC_1_1/temp3[4] ,
         \MC_ARK_ARC_1_1/temp3[3] , \MC_ARK_ARC_1_1/temp3[2] ,
         \MC_ARK_ARC_1_1/temp3[1] , \MC_ARK_ARC_1_1/temp3[0] ,
         \MC_ARK_ARC_1_1/temp2[191] , \MC_ARK_ARC_1_1/temp2[190] ,
         \MC_ARK_ARC_1_1/temp2[189] , \MC_ARK_ARC_1_1/temp2[188] ,
         \MC_ARK_ARC_1_1/temp2[187] , \MC_ARK_ARC_1_1/temp2[186] ,
         \MC_ARK_ARC_1_1/temp2[185] , \MC_ARK_ARC_1_1/temp2[184] ,
         \MC_ARK_ARC_1_1/temp2[183] , \MC_ARK_ARC_1_1/temp2[182] ,
         \MC_ARK_ARC_1_1/temp2[181] , \MC_ARK_ARC_1_1/temp2[180] ,
         \MC_ARK_ARC_1_1/temp2[179] , \MC_ARK_ARC_1_1/temp2[178] ,
         \MC_ARK_ARC_1_1/temp2[177] , \MC_ARK_ARC_1_1/temp2[176] ,
         \MC_ARK_ARC_1_1/temp2[175] , \MC_ARK_ARC_1_1/temp2[174] ,
         \MC_ARK_ARC_1_1/temp2[173] , \MC_ARK_ARC_1_1/temp2[172] ,
         \MC_ARK_ARC_1_1/temp2[171] , \MC_ARK_ARC_1_1/temp2[170] ,
         \MC_ARK_ARC_1_1/temp2[169] , \MC_ARK_ARC_1_1/temp2[168] ,
         \MC_ARK_ARC_1_1/temp2[167] , \MC_ARK_ARC_1_1/temp2[166] ,
         \MC_ARK_ARC_1_1/temp2[165] , \MC_ARK_ARC_1_1/temp2[164] ,
         \MC_ARK_ARC_1_1/temp2[163] , \MC_ARK_ARC_1_1/temp2[162] ,
         \MC_ARK_ARC_1_1/temp2[161] , \MC_ARK_ARC_1_1/temp2[160] ,
         \MC_ARK_ARC_1_1/temp2[159] , \MC_ARK_ARC_1_1/temp2[158] ,
         \MC_ARK_ARC_1_1/temp2[157] , \MC_ARK_ARC_1_1/temp2[156] ,
         \MC_ARK_ARC_1_1/temp2[155] , \MC_ARK_ARC_1_1/temp2[154] ,
         \MC_ARK_ARC_1_1/temp2[153] , \MC_ARK_ARC_1_1/temp2[152] ,
         \MC_ARK_ARC_1_1/temp2[151] , \MC_ARK_ARC_1_1/temp2[150] ,
         \MC_ARK_ARC_1_1/temp2[149] , \MC_ARK_ARC_1_1/temp2[148] ,
         \MC_ARK_ARC_1_1/temp2[147] , \MC_ARK_ARC_1_1/temp2[146] ,
         \MC_ARK_ARC_1_1/temp2[145] , \MC_ARK_ARC_1_1/temp2[144] ,
         \MC_ARK_ARC_1_1/temp2[143] , \MC_ARK_ARC_1_1/temp2[142] ,
         \MC_ARK_ARC_1_1/temp2[141] , \MC_ARK_ARC_1_1/temp2[140] ,
         \MC_ARK_ARC_1_1/temp2[139] , \MC_ARK_ARC_1_1/temp2[138] ,
         \MC_ARK_ARC_1_1/temp2[137] , \MC_ARK_ARC_1_1/temp2[136] ,
         \MC_ARK_ARC_1_1/temp2[135] , \MC_ARK_ARC_1_1/temp2[134] ,
         \MC_ARK_ARC_1_1/temp2[133] , \MC_ARK_ARC_1_1/temp2[132] ,
         \MC_ARK_ARC_1_1/temp2[131] , \MC_ARK_ARC_1_1/temp2[130] ,
         \MC_ARK_ARC_1_1/temp2[129] , \MC_ARK_ARC_1_1/temp2[128] ,
         \MC_ARK_ARC_1_1/temp2[127] , \MC_ARK_ARC_1_1/temp2[126] ,
         \MC_ARK_ARC_1_1/temp2[125] , \MC_ARK_ARC_1_1/temp2[124] ,
         \MC_ARK_ARC_1_1/temp2[123] , \MC_ARK_ARC_1_1/temp2[122] ,
         \MC_ARK_ARC_1_1/temp2[121] , \MC_ARK_ARC_1_1/temp2[120] ,
         \MC_ARK_ARC_1_1/temp2[119] , \MC_ARK_ARC_1_1/temp2[118] ,
         \MC_ARK_ARC_1_1/temp2[117] , \MC_ARK_ARC_1_1/temp2[116] ,
         \MC_ARK_ARC_1_1/temp2[115] , \MC_ARK_ARC_1_1/temp2[114] ,
         \MC_ARK_ARC_1_1/temp2[113] , \MC_ARK_ARC_1_1/temp2[112] ,
         \MC_ARK_ARC_1_1/temp2[111] , \MC_ARK_ARC_1_1/temp2[110] ,
         \MC_ARK_ARC_1_1/temp2[109] , \MC_ARK_ARC_1_1/temp2[108] ,
         \MC_ARK_ARC_1_1/temp2[107] , \MC_ARK_ARC_1_1/temp2[106] ,
         \MC_ARK_ARC_1_1/temp2[105] , \MC_ARK_ARC_1_1/temp2[104] ,
         \MC_ARK_ARC_1_1/temp2[103] , \MC_ARK_ARC_1_1/temp2[102] ,
         \MC_ARK_ARC_1_1/temp2[101] , \MC_ARK_ARC_1_1/temp2[100] ,
         \MC_ARK_ARC_1_1/temp2[99] , \MC_ARK_ARC_1_1/temp2[98] ,
         \MC_ARK_ARC_1_1/temp2[97] , \MC_ARK_ARC_1_1/temp2[96] ,
         \MC_ARK_ARC_1_1/temp2[95] , \MC_ARK_ARC_1_1/temp2[94] ,
         \MC_ARK_ARC_1_1/temp2[93] , \MC_ARK_ARC_1_1/temp2[92] ,
         \MC_ARK_ARC_1_1/temp2[91] , \MC_ARK_ARC_1_1/temp2[90] ,
         \MC_ARK_ARC_1_1/temp2[89] , \MC_ARK_ARC_1_1/temp2[88] ,
         \MC_ARK_ARC_1_1/temp2[87] , \MC_ARK_ARC_1_1/temp2[86] ,
         \MC_ARK_ARC_1_1/temp2[85] , \MC_ARK_ARC_1_1/temp2[84] ,
         \MC_ARK_ARC_1_1/temp2[83] , \MC_ARK_ARC_1_1/temp2[82] ,
         \MC_ARK_ARC_1_1/temp2[81] , \MC_ARK_ARC_1_1/temp2[80] ,
         \MC_ARK_ARC_1_1/temp2[79] , \MC_ARK_ARC_1_1/temp2[78] ,
         \MC_ARK_ARC_1_1/temp2[77] , \MC_ARK_ARC_1_1/temp2[76] ,
         \MC_ARK_ARC_1_1/temp2[75] , \MC_ARK_ARC_1_1/temp2[74] ,
         \MC_ARK_ARC_1_1/temp2[73] , \MC_ARK_ARC_1_1/temp2[72] ,
         \MC_ARK_ARC_1_1/temp2[71] , \MC_ARK_ARC_1_1/temp2[70] ,
         \MC_ARK_ARC_1_1/temp2[69] , \MC_ARK_ARC_1_1/temp2[68] ,
         \MC_ARK_ARC_1_1/temp2[67] , \MC_ARK_ARC_1_1/temp2[66] ,
         \MC_ARK_ARC_1_1/temp2[65] , \MC_ARK_ARC_1_1/temp2[64] ,
         \MC_ARK_ARC_1_1/temp2[63] , \MC_ARK_ARC_1_1/temp2[62] ,
         \MC_ARK_ARC_1_1/temp2[61] , \MC_ARK_ARC_1_1/temp2[60] ,
         \MC_ARK_ARC_1_1/temp2[59] , \MC_ARK_ARC_1_1/temp2[58] ,
         \MC_ARK_ARC_1_1/temp2[57] , \MC_ARK_ARC_1_1/temp2[56] ,
         \MC_ARK_ARC_1_1/temp2[55] , \MC_ARK_ARC_1_1/temp2[54] ,
         \MC_ARK_ARC_1_1/temp2[53] , \MC_ARK_ARC_1_1/temp2[52] ,
         \MC_ARK_ARC_1_1/temp2[51] , \MC_ARK_ARC_1_1/temp2[50] ,
         \MC_ARK_ARC_1_1/temp2[49] , \MC_ARK_ARC_1_1/temp2[48] ,
         \MC_ARK_ARC_1_1/temp2[47] , \MC_ARK_ARC_1_1/temp2[46] ,
         \MC_ARK_ARC_1_1/temp2[45] , \MC_ARK_ARC_1_1/temp2[44] ,
         \MC_ARK_ARC_1_1/temp2[43] , \MC_ARK_ARC_1_1/temp2[42] ,
         \MC_ARK_ARC_1_1/temp2[41] , \MC_ARK_ARC_1_1/temp2[40] ,
         \MC_ARK_ARC_1_1/temp2[39] , \MC_ARK_ARC_1_1/temp2[38] ,
         \MC_ARK_ARC_1_1/temp2[37] , \MC_ARK_ARC_1_1/temp2[36] ,
         \MC_ARK_ARC_1_1/temp2[35] , \MC_ARK_ARC_1_1/temp2[34] ,
         \MC_ARK_ARC_1_1/temp2[33] , \MC_ARK_ARC_1_1/temp2[32] ,
         \MC_ARK_ARC_1_1/temp2[31] , \MC_ARK_ARC_1_1/temp2[30] ,
         \MC_ARK_ARC_1_1/temp2[29] , \MC_ARK_ARC_1_1/temp2[28] ,
         \MC_ARK_ARC_1_1/temp2[27] , \MC_ARK_ARC_1_1/temp2[26] ,
         \MC_ARK_ARC_1_1/temp2[25] , \MC_ARK_ARC_1_1/temp2[24] ,
         \MC_ARK_ARC_1_1/temp2[23] , \MC_ARK_ARC_1_1/temp2[22] ,
         \MC_ARK_ARC_1_1/temp2[21] , \MC_ARK_ARC_1_1/temp2[20] ,
         \MC_ARK_ARC_1_1/temp2[19] , \MC_ARK_ARC_1_1/temp2[18] ,
         \MC_ARK_ARC_1_1/temp2[17] , \MC_ARK_ARC_1_1/temp2[16] ,
         \MC_ARK_ARC_1_1/temp2[15] , \MC_ARK_ARC_1_1/temp2[14] ,
         \MC_ARK_ARC_1_1/temp2[13] , \MC_ARK_ARC_1_1/temp2[12] ,
         \MC_ARK_ARC_1_1/temp2[11] , \MC_ARK_ARC_1_1/temp2[10] ,
         \MC_ARK_ARC_1_1/temp2[9] , \MC_ARK_ARC_1_1/temp2[8] ,
         \MC_ARK_ARC_1_1/temp2[7] , \MC_ARK_ARC_1_1/temp2[6] ,
         \MC_ARK_ARC_1_1/temp2[5] , \MC_ARK_ARC_1_1/temp2[4] ,
         \MC_ARK_ARC_1_1/temp2[3] , \MC_ARK_ARC_1_1/temp2[2] ,
         \MC_ARK_ARC_1_1/temp2[1] , \MC_ARK_ARC_1_1/temp2[0] ,
         \MC_ARK_ARC_1_1/temp1[191] , \MC_ARK_ARC_1_1/temp1[190] ,
         \MC_ARK_ARC_1_1/temp1[189] , \MC_ARK_ARC_1_1/temp1[188] ,
         \MC_ARK_ARC_1_1/temp1[187] , \MC_ARK_ARC_1_1/temp1[186] ,
         \MC_ARK_ARC_1_1/temp1[185] , \MC_ARK_ARC_1_1/temp1[184] ,
         \MC_ARK_ARC_1_1/temp1[183] , \MC_ARK_ARC_1_1/temp1[182] ,
         \MC_ARK_ARC_1_1/temp1[181] , \MC_ARK_ARC_1_1/temp1[180] ,
         \MC_ARK_ARC_1_1/temp1[179] , \MC_ARK_ARC_1_1/temp1[178] ,
         \MC_ARK_ARC_1_1/temp1[177] , \MC_ARK_ARC_1_1/temp1[176] ,
         \MC_ARK_ARC_1_1/temp1[175] , \MC_ARK_ARC_1_1/temp1[174] ,
         \MC_ARK_ARC_1_1/temp1[173] , \MC_ARK_ARC_1_1/temp1[172] ,
         \MC_ARK_ARC_1_1/temp1[171] , \MC_ARK_ARC_1_1/temp1[170] ,
         \MC_ARK_ARC_1_1/temp1[169] , \MC_ARK_ARC_1_1/temp1[168] ,
         \MC_ARK_ARC_1_1/temp1[167] , \MC_ARK_ARC_1_1/temp1[166] ,
         \MC_ARK_ARC_1_1/temp1[165] , \MC_ARK_ARC_1_1/temp1[164] ,
         \MC_ARK_ARC_1_1/temp1[163] , \MC_ARK_ARC_1_1/temp1[162] ,
         \MC_ARK_ARC_1_1/temp1[161] , \MC_ARK_ARC_1_1/temp1[160] ,
         \MC_ARK_ARC_1_1/temp1[159] , \MC_ARK_ARC_1_1/temp1[158] ,
         \MC_ARK_ARC_1_1/temp1[157] , \MC_ARK_ARC_1_1/temp1[156] ,
         \MC_ARK_ARC_1_1/temp1[155] , \MC_ARK_ARC_1_1/temp1[154] ,
         \MC_ARK_ARC_1_1/temp1[153] , \MC_ARK_ARC_1_1/temp1[152] ,
         \MC_ARK_ARC_1_1/temp1[151] , \MC_ARK_ARC_1_1/temp1[150] ,
         \MC_ARK_ARC_1_1/temp1[149] , \MC_ARK_ARC_1_1/temp1[148] ,
         \MC_ARK_ARC_1_1/temp1[147] , \MC_ARK_ARC_1_1/temp1[146] ,
         \MC_ARK_ARC_1_1/temp1[145] , \MC_ARK_ARC_1_1/temp1[144] ,
         \MC_ARK_ARC_1_1/temp1[143] , \MC_ARK_ARC_1_1/temp1[142] ,
         \MC_ARK_ARC_1_1/temp1[141] , \MC_ARK_ARC_1_1/temp1[140] ,
         \MC_ARK_ARC_1_1/temp1[139] , \MC_ARK_ARC_1_1/temp1[138] ,
         \MC_ARK_ARC_1_1/temp1[137] , \MC_ARK_ARC_1_1/temp1[136] ,
         \MC_ARK_ARC_1_1/temp1[135] , \MC_ARK_ARC_1_1/temp1[134] ,
         \MC_ARK_ARC_1_1/temp1[133] , \MC_ARK_ARC_1_1/temp1[132] ,
         \MC_ARK_ARC_1_1/temp1[131] , \MC_ARK_ARC_1_1/temp1[130] ,
         \MC_ARK_ARC_1_1/temp1[129] , \MC_ARK_ARC_1_1/temp1[128] ,
         \MC_ARK_ARC_1_1/temp1[127] , \MC_ARK_ARC_1_1/temp1[126] ,
         \MC_ARK_ARC_1_1/temp1[125] , \MC_ARK_ARC_1_1/temp1[124] ,
         \MC_ARK_ARC_1_1/temp1[123] , \MC_ARK_ARC_1_1/temp1[122] ,
         \MC_ARK_ARC_1_1/temp1[121] , \MC_ARK_ARC_1_1/temp1[120] ,
         \MC_ARK_ARC_1_1/temp1[119] , \MC_ARK_ARC_1_1/temp1[118] ,
         \MC_ARK_ARC_1_1/temp1[117] , \MC_ARK_ARC_1_1/temp1[116] ,
         \MC_ARK_ARC_1_1/temp1[115] , \MC_ARK_ARC_1_1/temp1[114] ,
         \MC_ARK_ARC_1_1/temp1[113] , \MC_ARK_ARC_1_1/temp1[112] ,
         \MC_ARK_ARC_1_1/temp1[111] , \MC_ARK_ARC_1_1/temp1[110] ,
         \MC_ARK_ARC_1_1/temp1[109] , \MC_ARK_ARC_1_1/temp1[108] ,
         \MC_ARK_ARC_1_1/temp1[107] , \MC_ARK_ARC_1_1/temp1[106] ,
         \MC_ARK_ARC_1_1/temp1[105] , \MC_ARK_ARC_1_1/temp1[104] ,
         \MC_ARK_ARC_1_1/temp1[103] , \MC_ARK_ARC_1_1/temp1[102] ,
         \MC_ARK_ARC_1_1/temp1[101] , \MC_ARK_ARC_1_1/temp1[100] ,
         \MC_ARK_ARC_1_1/temp1[99] , \MC_ARK_ARC_1_1/temp1[98] ,
         \MC_ARK_ARC_1_1/temp1[97] , \MC_ARK_ARC_1_1/temp1[96] ,
         \MC_ARK_ARC_1_1/temp1[95] , \MC_ARK_ARC_1_1/temp1[94] ,
         \MC_ARK_ARC_1_1/temp1[93] , \MC_ARK_ARC_1_1/temp1[92] ,
         \MC_ARK_ARC_1_1/temp1[91] , \MC_ARK_ARC_1_1/temp1[90] ,
         \MC_ARK_ARC_1_1/temp1[89] , \MC_ARK_ARC_1_1/temp1[88] ,
         \MC_ARK_ARC_1_1/temp1[87] , \MC_ARK_ARC_1_1/temp1[86] ,
         \MC_ARK_ARC_1_1/temp1[85] , \MC_ARK_ARC_1_1/temp1[84] ,
         \MC_ARK_ARC_1_1/temp1[83] , \MC_ARK_ARC_1_1/temp1[82] ,
         \MC_ARK_ARC_1_1/temp1[81] , \MC_ARK_ARC_1_1/temp1[80] ,
         \MC_ARK_ARC_1_1/temp1[79] , \MC_ARK_ARC_1_1/temp1[78] ,
         \MC_ARK_ARC_1_1/temp1[77] , \MC_ARK_ARC_1_1/temp1[76] ,
         \MC_ARK_ARC_1_1/temp1[75] , \MC_ARK_ARC_1_1/temp1[74] ,
         \MC_ARK_ARC_1_1/temp1[73] , \MC_ARK_ARC_1_1/temp1[72] ,
         \MC_ARK_ARC_1_1/temp1[71] , \MC_ARK_ARC_1_1/temp1[70] ,
         \MC_ARK_ARC_1_1/temp1[69] , \MC_ARK_ARC_1_1/temp1[68] ,
         \MC_ARK_ARC_1_1/temp1[67] , \MC_ARK_ARC_1_1/temp1[66] ,
         \MC_ARK_ARC_1_1/temp1[65] , \MC_ARK_ARC_1_1/temp1[64] ,
         \MC_ARK_ARC_1_1/temp1[63] , \MC_ARK_ARC_1_1/temp1[62] ,
         \MC_ARK_ARC_1_1/temp1[61] , \MC_ARK_ARC_1_1/temp1[60] ,
         \MC_ARK_ARC_1_1/temp1[59] , \MC_ARK_ARC_1_1/temp1[58] ,
         \MC_ARK_ARC_1_1/temp1[57] , \MC_ARK_ARC_1_1/temp1[56] ,
         \MC_ARK_ARC_1_1/temp1[55] , \MC_ARK_ARC_1_1/temp1[54] ,
         \MC_ARK_ARC_1_1/temp1[53] , \MC_ARK_ARC_1_1/temp1[52] ,
         \MC_ARK_ARC_1_1/temp1[51] , \MC_ARK_ARC_1_1/temp1[50] ,
         \MC_ARK_ARC_1_1/temp1[49] , \MC_ARK_ARC_1_1/temp1[48] ,
         \MC_ARK_ARC_1_1/temp1[47] , \MC_ARK_ARC_1_1/temp1[46] ,
         \MC_ARK_ARC_1_1/temp1[45] , \MC_ARK_ARC_1_1/temp1[44] ,
         \MC_ARK_ARC_1_1/temp1[43] , \MC_ARK_ARC_1_1/temp1[42] ,
         \MC_ARK_ARC_1_1/temp1[41] , \MC_ARK_ARC_1_1/temp1[40] ,
         \MC_ARK_ARC_1_1/temp1[39] , \MC_ARK_ARC_1_1/temp1[38] ,
         \MC_ARK_ARC_1_1/temp1[37] , \MC_ARK_ARC_1_1/temp1[36] ,
         \MC_ARK_ARC_1_1/temp1[35] , \MC_ARK_ARC_1_1/temp1[34] ,
         \MC_ARK_ARC_1_1/temp1[33] , \MC_ARK_ARC_1_1/temp1[32] ,
         \MC_ARK_ARC_1_1/temp1[31] , \MC_ARK_ARC_1_1/temp1[30] ,
         \MC_ARK_ARC_1_1/temp1[29] , \MC_ARK_ARC_1_1/temp1[28] ,
         \MC_ARK_ARC_1_1/temp1[27] , \MC_ARK_ARC_1_1/temp1[26] ,
         \MC_ARK_ARC_1_1/temp1[25] , \MC_ARK_ARC_1_1/temp1[24] ,
         \MC_ARK_ARC_1_1/temp1[23] , \MC_ARK_ARC_1_1/temp1[22] ,
         \MC_ARK_ARC_1_1/temp1[21] , \MC_ARK_ARC_1_1/temp1[20] ,
         \MC_ARK_ARC_1_1/temp1[19] , \MC_ARK_ARC_1_1/temp1[18] ,
         \MC_ARK_ARC_1_1/temp1[17] , \MC_ARK_ARC_1_1/temp1[16] ,
         \MC_ARK_ARC_1_1/temp1[15] , \MC_ARK_ARC_1_1/temp1[14] ,
         \MC_ARK_ARC_1_1/temp1[13] , \MC_ARK_ARC_1_1/temp1[12] ,
         \MC_ARK_ARC_1_1/temp1[11] , \MC_ARK_ARC_1_1/temp1[10] ,
         \MC_ARK_ARC_1_1/temp1[9] , \MC_ARK_ARC_1_1/temp1[8] ,
         \MC_ARK_ARC_1_1/temp1[7] , \MC_ARK_ARC_1_1/temp1[6] ,
         \MC_ARK_ARC_1_1/temp1[5] , \MC_ARK_ARC_1_1/temp1[4] ,
         \MC_ARK_ARC_1_1/temp1[3] , \MC_ARK_ARC_1_1/temp1[2] ,
         \MC_ARK_ARC_1_1/temp1[1] , \MC_ARK_ARC_1_1/temp1[0] ,
         \MC_ARK_ARC_1_1/buf_keyinput[189] ,
         \MC_ARK_ARC_1_1/buf_keyinput[183] ,
         \MC_ARK_ARC_1_1/buf_keyinput[176] ,
         \MC_ARK_ARC_1_1/buf_keyinput[170] ,
         \MC_ARK_ARC_1_1/buf_keyinput[165] ,
         \MC_ARK_ARC_1_1/buf_keyinput[152] ,
         \MC_ARK_ARC_1_1/buf_keyinput[134] ,
         \MC_ARK_ARC_1_1/buf_keyinput[129] ,
         \MC_ARK_ARC_1_1/buf_keyinput[125] ,
         \MC_ARK_ARC_1_1/buf_keyinput[123] ,
         \MC_ARK_ARC_1_1/buf_keyinput[107] ,
         \MC_ARK_ARC_1_1/buf_keyinput[106] ,
         \MC_ARK_ARC_1_1/buf_keyinput[105] , \MC_ARK_ARC_1_1/buf_keyinput[74] ,
         \MC_ARK_ARC_1_1/buf_keyinput[62] , \MC_ARK_ARC_1_1/buf_keyinput[27] ,
         \MC_ARK_ARC_1_1/buf_keyinput[8] , \MC_ARK_ARC_1_1/buf_datainput[191] ,
         \MC_ARK_ARC_1_1/buf_datainput[190] ,
         \MC_ARK_ARC_1_1/buf_datainput[188] ,
         \MC_ARK_ARC_1_1/buf_datainput[187] ,
         \MC_ARK_ARC_1_1/buf_datainput[186] ,
         \MC_ARK_ARC_1_1/buf_datainput[185] ,
         \MC_ARK_ARC_1_1/buf_datainput[184] ,
         \MC_ARK_ARC_1_1/buf_datainput[182] ,
         \MC_ARK_ARC_1_1/buf_datainput[181] ,
         \MC_ARK_ARC_1_1/buf_datainput[180] ,
         \MC_ARK_ARC_1_1/buf_datainput[179] ,
         \MC_ARK_ARC_1_1/buf_datainput[178] ,
         \MC_ARK_ARC_1_1/buf_datainput[176] ,
         \MC_ARK_ARC_1_1/buf_datainput[175] ,
         \MC_ARK_ARC_1_1/buf_datainput[174] ,
         \MC_ARK_ARC_1_1/buf_datainput[173] ,
         \MC_ARK_ARC_1_1/buf_datainput[172] ,
         \MC_ARK_ARC_1_1/buf_datainput[170] ,
         \MC_ARK_ARC_1_1/buf_datainput[169] ,
         \MC_ARK_ARC_1_1/buf_datainput[168] ,
         \MC_ARK_ARC_1_1/buf_datainput[167] ,
         \MC_ARK_ARC_1_1/buf_datainput[166] ,
         \MC_ARK_ARC_1_1/buf_datainput[165] ,
         \MC_ARK_ARC_1_1/buf_datainput[163] ,
         \MC_ARK_ARC_1_1/buf_datainput[162] ,
         \MC_ARK_ARC_1_1/buf_datainput[161] ,
         \MC_ARK_ARC_1_1/buf_datainput[160] ,
         \MC_ARK_ARC_1_1/buf_datainput[159] ,
         \MC_ARK_ARC_1_1/buf_datainput[158] ,
         \MC_ARK_ARC_1_1/buf_datainput[157] ,
         \MC_ARK_ARC_1_1/buf_datainput[156] ,
         \MC_ARK_ARC_1_1/buf_datainput[155] ,
         \MC_ARK_ARC_1_1/buf_datainput[154] ,
         \MC_ARK_ARC_1_1/buf_datainput[153] ,
         \MC_ARK_ARC_1_1/buf_datainput[152] ,
         \MC_ARK_ARC_1_1/buf_datainput[151] ,
         \MC_ARK_ARC_1_1/buf_datainput[150] ,
         \MC_ARK_ARC_1_1/buf_datainput[149] ,
         \MC_ARK_ARC_1_1/buf_datainput[148] ,
         \MC_ARK_ARC_1_1/buf_datainput[146] ,
         \MC_ARK_ARC_1_1/buf_datainput[145] ,
         \MC_ARK_ARC_1_1/buf_datainput[144] ,
         \MC_ARK_ARC_1_1/buf_datainput[143] ,
         \MC_ARK_ARC_1_1/buf_datainput[142] ,
         \MC_ARK_ARC_1_1/buf_datainput[140] ,
         \MC_ARK_ARC_1_1/buf_datainput[139] ,
         \MC_ARK_ARC_1_1/buf_datainput[137] ,
         \MC_ARK_ARC_1_1/buf_datainput[136] ,
         \MC_ARK_ARC_1_1/buf_datainput[134] ,
         \MC_ARK_ARC_1_1/buf_datainput[133] ,
         \MC_ARK_ARC_1_1/buf_datainput[131] ,
         \MC_ARK_ARC_1_1/buf_datainput[130] ,
         \MC_ARK_ARC_1_1/buf_datainput[128] ,
         \MC_ARK_ARC_1_1/buf_datainput[127] ,
         \MC_ARK_ARC_1_1/buf_datainput[126] ,
         \MC_ARK_ARC_1_1/buf_datainput[125] ,
         \MC_ARK_ARC_1_1/buf_datainput[124] ,
         \MC_ARK_ARC_1_1/buf_datainput[122] ,
         \MC_ARK_ARC_1_1/buf_datainput[121] ,
         \MC_ARK_ARC_1_1/buf_datainput[120] ,
         \MC_ARK_ARC_1_1/buf_datainput[119] ,
         \MC_ARK_ARC_1_1/buf_datainput[118] ,
         \MC_ARK_ARC_1_1/buf_datainput[116] ,
         \MC_ARK_ARC_1_1/buf_datainput[115] ,
         \MC_ARK_ARC_1_1/buf_datainput[114] ,
         \MC_ARK_ARC_1_1/buf_datainput[112] ,
         \MC_ARK_ARC_1_1/buf_datainput[111] ,
         \MC_ARK_ARC_1_1/buf_datainput[110] ,
         \MC_ARK_ARC_1_1/buf_datainput[109] ,
         \MC_ARK_ARC_1_1/buf_datainput[108] ,
         \MC_ARK_ARC_1_1/buf_datainput[107] ,
         \MC_ARK_ARC_1_1/buf_datainput[106] ,
         \MC_ARK_ARC_1_1/buf_datainput[105] ,
         \MC_ARK_ARC_1_1/buf_datainput[104] ,
         \MC_ARK_ARC_1_1/buf_datainput[103] ,
         \MC_ARK_ARC_1_1/buf_datainput[102] ,
         \MC_ARK_ARC_1_1/buf_datainput[101] ,
         \MC_ARK_ARC_1_1/buf_datainput[100] ,
         \MC_ARK_ARC_1_1/buf_datainput[99] ,
         \MC_ARK_ARC_1_1/buf_datainput[98] ,
         \MC_ARK_ARC_1_1/buf_datainput[97] ,
         \MC_ARK_ARC_1_1/buf_datainput[96] ,
         \MC_ARK_ARC_1_1/buf_datainput[95] ,
         \MC_ARK_ARC_1_1/buf_datainput[94] ,
         \MC_ARK_ARC_1_1/buf_datainput[92] ,
         \MC_ARK_ARC_1_1/buf_datainput[91] ,
         \MC_ARK_ARC_1_1/buf_datainput[90] ,
         \MC_ARK_ARC_1_1/buf_datainput[89] ,
         \MC_ARK_ARC_1_1/buf_datainput[88] ,
         \MC_ARK_ARC_1_1/buf_datainput[87] ,
         \MC_ARK_ARC_1_1/buf_datainput[86] ,
         \MC_ARK_ARC_1_1/buf_datainput[85] ,
         \MC_ARK_ARC_1_1/buf_datainput[84] ,
         \MC_ARK_ARC_1_1/buf_datainput[83] ,
         \MC_ARK_ARC_1_1/buf_datainput[82] ,
         \MC_ARK_ARC_1_1/buf_datainput[80] ,
         \MC_ARK_ARC_1_1/buf_datainput[79] ,
         \MC_ARK_ARC_1_1/buf_datainput[78] ,
         \MC_ARK_ARC_1_1/buf_datainput[77] ,
         \MC_ARK_ARC_1_1/buf_datainput[76] ,
         \MC_ARK_ARC_1_1/buf_datainput[74] ,
         \MC_ARK_ARC_1_1/buf_datainput[73] ,
         \MC_ARK_ARC_1_1/buf_datainput[72] ,
         \MC_ARK_ARC_1_1/buf_datainput[71] ,
         \MC_ARK_ARC_1_1/buf_datainput[70] ,
         \MC_ARK_ARC_1_1/buf_datainput[69] ,
         \MC_ARK_ARC_1_1/buf_datainput[68] ,
         \MC_ARK_ARC_1_1/buf_datainput[67] ,
         \MC_ARK_ARC_1_1/buf_datainput[66] ,
         \MC_ARK_ARC_1_1/buf_datainput[65] ,
         \MC_ARK_ARC_1_1/buf_datainput[64] ,
         \MC_ARK_ARC_1_1/buf_datainput[63] ,
         \MC_ARK_ARC_1_1/buf_datainput[62] ,
         \MC_ARK_ARC_1_1/buf_datainput[61] ,
         \MC_ARK_ARC_1_1/buf_datainput[60] ,
         \MC_ARK_ARC_1_1/buf_datainput[59] ,
         \MC_ARK_ARC_1_1/buf_datainput[58] ,
         \MC_ARK_ARC_1_1/buf_datainput[55] ,
         \MC_ARK_ARC_1_1/buf_datainput[54] ,
         \MC_ARK_ARC_1_1/buf_datainput[52] ,
         \MC_ARK_ARC_1_1/buf_datainput[50] ,
         \MC_ARK_ARC_1_1/buf_datainput[49] ,
         \MC_ARK_ARC_1_1/buf_datainput[48] ,
         \MC_ARK_ARC_1_1/buf_datainput[47] ,
         \MC_ARK_ARC_1_1/buf_datainput[46] ,
         \MC_ARK_ARC_1_1/buf_datainput[45] ,
         \MC_ARK_ARC_1_1/buf_datainput[44] ,
         \MC_ARK_ARC_1_1/buf_datainput[43] ,
         \MC_ARK_ARC_1_1/buf_datainput[42] ,
         \MC_ARK_ARC_1_1/buf_datainput[41] ,
         \MC_ARK_ARC_1_1/buf_datainput[40] ,
         \MC_ARK_ARC_1_1/buf_datainput[39] ,
         \MC_ARK_ARC_1_1/buf_datainput[38] ,
         \MC_ARK_ARC_1_1/buf_datainput[37] ,
         \MC_ARK_ARC_1_1/buf_datainput[36] ,
         \MC_ARK_ARC_1_1/buf_datainput[35] ,
         \MC_ARK_ARC_1_1/buf_datainput[34] ,
         \MC_ARK_ARC_1_1/buf_datainput[33] ,
         \MC_ARK_ARC_1_1/buf_datainput[32] ,
         \MC_ARK_ARC_1_1/buf_datainput[31] ,
         \MC_ARK_ARC_1_1/buf_datainput[30] ,
         \MC_ARK_ARC_1_1/buf_datainput[29] ,
         \MC_ARK_ARC_1_1/buf_datainput[28] ,
         \MC_ARK_ARC_1_1/buf_datainput[27] ,
         \MC_ARK_ARC_1_1/buf_datainput[26] ,
         \MC_ARK_ARC_1_1/buf_datainput[25] ,
         \MC_ARK_ARC_1_1/buf_datainput[24] ,
         \MC_ARK_ARC_1_1/buf_datainput[23] ,
         \MC_ARK_ARC_1_1/buf_datainput[22] ,
         \MC_ARK_ARC_1_1/buf_datainput[21] ,
         \MC_ARK_ARC_1_1/buf_datainput[20] ,
         \MC_ARK_ARC_1_1/buf_datainput[19] ,
         \MC_ARK_ARC_1_1/buf_datainput[18] ,
         \MC_ARK_ARC_1_1/buf_datainput[17] ,
         \MC_ARK_ARC_1_1/buf_datainput[16] ,
         \MC_ARK_ARC_1_1/buf_datainput[15] ,
         \MC_ARK_ARC_1_1/buf_datainput[14] ,
         \MC_ARK_ARC_1_1/buf_datainput[13] ,
         \MC_ARK_ARC_1_1/buf_datainput[12] ,
         \MC_ARK_ARC_1_1/buf_datainput[10] , \MC_ARK_ARC_1_1/buf_datainput[8] ,
         \MC_ARK_ARC_1_1/buf_datainput[7] , \MC_ARK_ARC_1_1/buf_datainput[6] ,
         \MC_ARK_ARC_1_1/buf_datainput[5] , \MC_ARK_ARC_1_1/buf_datainput[4] ,
         \MC_ARK_ARC_1_1/buf_datainput[3] , \MC_ARK_ARC_1_1/buf_datainput[2] ,
         \MC_ARK_ARC_1_1/buf_datainput[1] , \MC_ARK_ARC_1_1/buf_datainput[0] ,
         \MC_ARK_ARC_1_2/temp6[190] , \MC_ARK_ARC_1_2/temp6[189] ,
         \MC_ARK_ARC_1_2/temp6[188] , \MC_ARK_ARC_1_2/temp6[187] ,
         \MC_ARK_ARC_1_2/temp6[186] , \MC_ARK_ARC_1_2/temp6[185] ,
         \MC_ARK_ARC_1_2/temp6[184] , \MC_ARK_ARC_1_2/temp6[183] ,
         \MC_ARK_ARC_1_2/temp6[182] , \MC_ARK_ARC_1_2/temp6[181] ,
         \MC_ARK_ARC_1_2/temp6[180] , \MC_ARK_ARC_1_2/temp6[179] ,
         \MC_ARK_ARC_1_2/temp6[178] , \MC_ARK_ARC_1_2/temp6[177] ,
         \MC_ARK_ARC_1_2/temp6[176] , \MC_ARK_ARC_1_2/temp6[174] ,
         \MC_ARK_ARC_1_2/temp6[172] , \MC_ARK_ARC_1_2/temp6[171] ,
         \MC_ARK_ARC_1_2/temp6[170] , \MC_ARK_ARC_1_2/temp6[169] ,
         \MC_ARK_ARC_1_2/temp6[168] , \MC_ARK_ARC_1_2/temp6[166] ,
         \MC_ARK_ARC_1_2/temp6[165] , \MC_ARK_ARC_1_2/temp6[164] ,
         \MC_ARK_ARC_1_2/temp6[163] , \MC_ARK_ARC_1_2/temp6[162] ,
         \MC_ARK_ARC_1_2/temp6[160] , \MC_ARK_ARC_1_2/temp6[159] ,
         \MC_ARK_ARC_1_2/temp6[158] , \MC_ARK_ARC_1_2/temp6[157] ,
         \MC_ARK_ARC_1_2/temp6[156] , \MC_ARK_ARC_1_2/temp6[154] ,
         \MC_ARK_ARC_1_2/temp6[153] , \MC_ARK_ARC_1_2/temp6[152] ,
         \MC_ARK_ARC_1_2/temp6[151] , \MC_ARK_ARC_1_2/temp6[150] ,
         \MC_ARK_ARC_1_2/temp6[148] , \MC_ARK_ARC_1_2/temp6[147] ,
         \MC_ARK_ARC_1_2/temp6[146] , \MC_ARK_ARC_1_2/temp6[145] ,
         \MC_ARK_ARC_1_2/temp6[144] , \MC_ARK_ARC_1_2/temp6[143] ,
         \MC_ARK_ARC_1_2/temp6[142] , \MC_ARK_ARC_1_2/temp6[141] ,
         \MC_ARK_ARC_1_2/temp6[140] , \MC_ARK_ARC_1_2/temp6[139] ,
         \MC_ARK_ARC_1_2/temp6[138] , \MC_ARK_ARC_1_2/temp6[137] ,
         \MC_ARK_ARC_1_2/temp6[136] , \MC_ARK_ARC_1_2/temp6[135] ,
         \MC_ARK_ARC_1_2/temp6[134] , \MC_ARK_ARC_1_2/temp6[133] ,
         \MC_ARK_ARC_1_2/temp6[132] , \MC_ARK_ARC_1_2/temp6[130] ,
         \MC_ARK_ARC_1_2/temp6[128] , \MC_ARK_ARC_1_2/temp6[127] ,
         \MC_ARK_ARC_1_2/temp6[126] , \MC_ARK_ARC_1_2/temp6[124] ,
         \MC_ARK_ARC_1_2/temp6[121] , \MC_ARK_ARC_1_2/temp6[120] ,
         \MC_ARK_ARC_1_2/temp6[119] , \MC_ARK_ARC_1_2/temp6[118] ,
         \MC_ARK_ARC_1_2/temp6[117] , \MC_ARK_ARC_1_2/temp6[116] ,
         \MC_ARK_ARC_1_2/temp6[115] , \MC_ARK_ARC_1_2/temp6[114] ,
         \MC_ARK_ARC_1_2/temp6[113] , \MC_ARK_ARC_1_2/temp6[112] ,
         \MC_ARK_ARC_1_2/temp6[111] , \MC_ARK_ARC_1_2/temp6[110] ,
         \MC_ARK_ARC_1_2/temp6[109] , \MC_ARK_ARC_1_2/temp6[108] ,
         \MC_ARK_ARC_1_2/temp6[107] , \MC_ARK_ARC_1_2/temp6[106] ,
         \MC_ARK_ARC_1_2/temp6[105] , \MC_ARK_ARC_1_2/temp6[104] ,
         \MC_ARK_ARC_1_2/temp6[103] , \MC_ARK_ARC_1_2/temp6[102] ,
         \MC_ARK_ARC_1_2/temp6[100] , \MC_ARK_ARC_1_2/temp6[99] ,
         \MC_ARK_ARC_1_2/temp6[98] , \MC_ARK_ARC_1_2/temp6[97] ,
         \MC_ARK_ARC_1_2/temp6[96] , \MC_ARK_ARC_1_2/temp6[95] ,
         \MC_ARK_ARC_1_2/temp6[93] , \MC_ARK_ARC_1_2/temp6[91] ,
         \MC_ARK_ARC_1_2/temp6[90] , \MC_ARK_ARC_1_2/temp6[88] ,
         \MC_ARK_ARC_1_2/temp6[87] , \MC_ARK_ARC_1_2/temp6[86] ,
         \MC_ARK_ARC_1_2/temp6[85] , \MC_ARK_ARC_1_2/temp6[84] ,
         \MC_ARK_ARC_1_2/temp6[83] , \MC_ARK_ARC_1_2/temp6[82] ,
         \MC_ARK_ARC_1_2/temp6[81] , \MC_ARK_ARC_1_2/temp6[79] ,
         \MC_ARK_ARC_1_2/temp6[78] , \MC_ARK_ARC_1_2/temp6[76] ,
         \MC_ARK_ARC_1_2/temp6[74] , \MC_ARK_ARC_1_2/temp6[73] ,
         \MC_ARK_ARC_1_2/temp6[72] , \MC_ARK_ARC_1_2/temp6[70] ,
         \MC_ARK_ARC_1_2/temp6[68] , \MC_ARK_ARC_1_2/temp6[67] ,
         \MC_ARK_ARC_1_2/temp6[66] , \MC_ARK_ARC_1_2/temp6[65] ,
         \MC_ARK_ARC_1_2/temp6[64] , \MC_ARK_ARC_1_2/temp6[61] ,
         \MC_ARK_ARC_1_2/temp6[60] , \MC_ARK_ARC_1_2/temp6[58] ,
         \MC_ARK_ARC_1_2/temp6[57] , \MC_ARK_ARC_1_2/temp6[55] ,
         \MC_ARK_ARC_1_2/temp6[54] , \MC_ARK_ARC_1_2/temp6[53] ,
         \MC_ARK_ARC_1_2/temp6[52] , \MC_ARK_ARC_1_2/temp6[51] ,
         \MC_ARK_ARC_1_2/temp6[49] , \MC_ARK_ARC_1_2/temp6[48] ,
         \MC_ARK_ARC_1_2/temp6[47] , \MC_ARK_ARC_1_2/temp6[46] ,
         \MC_ARK_ARC_1_2/temp6[45] , \MC_ARK_ARC_1_2/temp6[44] ,
         \MC_ARK_ARC_1_2/temp6[43] , \MC_ARK_ARC_1_2/temp6[42] ,
         \MC_ARK_ARC_1_2/temp6[40] , \MC_ARK_ARC_1_2/temp6[38] ,
         \MC_ARK_ARC_1_2/temp6[37] , \MC_ARK_ARC_1_2/temp6[36] ,
         \MC_ARK_ARC_1_2/temp6[35] , \MC_ARK_ARC_1_2/temp6[34] ,
         \MC_ARK_ARC_1_2/temp6[33] , \MC_ARK_ARC_1_2/temp6[32] ,
         \MC_ARK_ARC_1_2/temp6[31] , \MC_ARK_ARC_1_2/temp6[30] ,
         \MC_ARK_ARC_1_2/temp6[28] , \MC_ARK_ARC_1_2/temp6[27] ,
         \MC_ARK_ARC_1_2/temp6[26] , \MC_ARK_ARC_1_2/temp6[25] ,
         \MC_ARK_ARC_1_2/temp6[24] , \MC_ARK_ARC_1_2/temp6[22] ,
         \MC_ARK_ARC_1_2/temp6[21] , \MC_ARK_ARC_1_2/temp6[19] ,
         \MC_ARK_ARC_1_2/temp6[18] , \MC_ARK_ARC_1_2/temp6[16] ,
         \MC_ARK_ARC_1_2/temp6[15] , \MC_ARK_ARC_1_2/temp6[13] ,
         \MC_ARK_ARC_1_2/temp6[12] , \MC_ARK_ARC_1_2/temp6[11] ,
         \MC_ARK_ARC_1_2/temp6[10] , \MC_ARK_ARC_1_2/temp6[9] ,
         \MC_ARK_ARC_1_2/temp6[8] , \MC_ARK_ARC_1_2/temp6[7] ,
         \MC_ARK_ARC_1_2/temp6[6] , \MC_ARK_ARC_1_2/temp6[5] ,
         \MC_ARK_ARC_1_2/temp6[4] , \MC_ARK_ARC_1_2/temp6[3] ,
         \MC_ARK_ARC_1_2/temp6[2] , \MC_ARK_ARC_1_2/temp6[1] ,
         \MC_ARK_ARC_1_2/temp6[0] , \MC_ARK_ARC_1_2/temp5[190] ,
         \MC_ARK_ARC_1_2/temp5[189] , \MC_ARK_ARC_1_2/temp5[188] ,
         \MC_ARK_ARC_1_2/temp5[187] , \MC_ARK_ARC_1_2/temp5[186] ,
         \MC_ARK_ARC_1_2/temp5[185] , \MC_ARK_ARC_1_2/temp5[184] ,
         \MC_ARK_ARC_1_2/temp5[183] , \MC_ARK_ARC_1_2/temp5[182] ,
         \MC_ARK_ARC_1_2/temp5[181] , \MC_ARK_ARC_1_2/temp5[180] ,
         \MC_ARK_ARC_1_2/temp5[179] , \MC_ARK_ARC_1_2/temp5[178] ,
         \MC_ARK_ARC_1_2/temp5[177] , \MC_ARK_ARC_1_2/temp5[176] ,
         \MC_ARK_ARC_1_2/temp5[175] , \MC_ARK_ARC_1_2/temp5[174] ,
         \MC_ARK_ARC_1_2/temp5[172] , \MC_ARK_ARC_1_2/temp5[171] ,
         \MC_ARK_ARC_1_2/temp5[170] , \MC_ARK_ARC_1_2/temp5[169] ,
         \MC_ARK_ARC_1_2/temp5[168] , \MC_ARK_ARC_1_2/temp5[166] ,
         \MC_ARK_ARC_1_2/temp5[165] , \MC_ARK_ARC_1_2/temp5[164] ,
         \MC_ARK_ARC_1_2/temp5[163] , \MC_ARK_ARC_1_2/temp5[162] ,
         \MC_ARK_ARC_1_2/temp5[160] , \MC_ARK_ARC_1_2/temp5[159] ,
         \MC_ARK_ARC_1_2/temp5[158] , \MC_ARK_ARC_1_2/temp5[157] ,
         \MC_ARK_ARC_1_2/temp5[156] , \MC_ARK_ARC_1_2/temp5[154] ,
         \MC_ARK_ARC_1_2/temp5[153] , \MC_ARK_ARC_1_2/temp5[152] ,
         \MC_ARK_ARC_1_2/temp5[151] , \MC_ARK_ARC_1_2/temp5[150] ,
         \MC_ARK_ARC_1_2/temp5[148] , \MC_ARK_ARC_1_2/temp5[147] ,
         \MC_ARK_ARC_1_2/temp5[146] , \MC_ARK_ARC_1_2/temp5[145] ,
         \MC_ARK_ARC_1_2/temp5[144] , \MC_ARK_ARC_1_2/temp5[143] ,
         \MC_ARK_ARC_1_2/temp5[142] , \MC_ARK_ARC_1_2/temp5[141] ,
         \MC_ARK_ARC_1_2/temp5[140] , \MC_ARK_ARC_1_2/temp5[139] ,
         \MC_ARK_ARC_1_2/temp5[138] , \MC_ARK_ARC_1_2/temp5[137] ,
         \MC_ARK_ARC_1_2/temp5[136] , \MC_ARK_ARC_1_2/temp5[135] ,
         \MC_ARK_ARC_1_2/temp5[134] , \MC_ARK_ARC_1_2/temp5[133] ,
         \MC_ARK_ARC_1_2/temp5[132] , \MC_ARK_ARC_1_2/temp5[131] ,
         \MC_ARK_ARC_1_2/temp5[130] , \MC_ARK_ARC_1_2/temp5[128] ,
         \MC_ARK_ARC_1_2/temp5[127] , \MC_ARK_ARC_1_2/temp5[126] ,
         \MC_ARK_ARC_1_2/temp5[124] , \MC_ARK_ARC_1_2/temp5[121] ,
         \MC_ARK_ARC_1_2/temp5[120] , \MC_ARK_ARC_1_2/temp5[119] ,
         \MC_ARK_ARC_1_2/temp5[118] , \MC_ARK_ARC_1_2/temp5[117] ,
         \MC_ARK_ARC_1_2/temp5[116] , \MC_ARK_ARC_1_2/temp5[115] ,
         \MC_ARK_ARC_1_2/temp5[114] , \MC_ARK_ARC_1_2/temp5[113] ,
         \MC_ARK_ARC_1_2/temp5[112] , \MC_ARK_ARC_1_2/temp5[111] ,
         \MC_ARK_ARC_1_2/temp5[110] , \MC_ARK_ARC_1_2/temp5[109] ,
         \MC_ARK_ARC_1_2/temp5[108] , \MC_ARK_ARC_1_2/temp5[107] ,
         \MC_ARK_ARC_1_2/temp5[106] , \MC_ARK_ARC_1_2/temp5[105] ,
         \MC_ARK_ARC_1_2/temp5[104] , \MC_ARK_ARC_1_2/temp5[103] ,
         \MC_ARK_ARC_1_2/temp5[102] , \MC_ARK_ARC_1_2/temp5[100] ,
         \MC_ARK_ARC_1_2/temp5[99] , \MC_ARK_ARC_1_2/temp5[98] ,
         \MC_ARK_ARC_1_2/temp5[97] , \MC_ARK_ARC_1_2/temp5[96] ,
         \MC_ARK_ARC_1_2/temp5[95] , \MC_ARK_ARC_1_2/temp5[93] ,
         \MC_ARK_ARC_1_2/temp5[92] , \MC_ARK_ARC_1_2/temp5[91] ,
         \MC_ARK_ARC_1_2/temp5[90] , \MC_ARK_ARC_1_2/temp5[88] ,
         \MC_ARK_ARC_1_2/temp5[87] , \MC_ARK_ARC_1_2/temp5[86] ,
         \MC_ARK_ARC_1_2/temp5[85] , \MC_ARK_ARC_1_2/temp5[84] ,
         \MC_ARK_ARC_1_2/temp5[83] , \MC_ARK_ARC_1_2/temp5[82] ,
         \MC_ARK_ARC_1_2/temp5[79] , \MC_ARK_ARC_1_2/temp5[78] ,
         \MC_ARK_ARC_1_2/temp5[76] , \MC_ARK_ARC_1_2/temp5[75] ,
         \MC_ARK_ARC_1_2/temp5[74] , \MC_ARK_ARC_1_2/temp5[73] ,
         \MC_ARK_ARC_1_2/temp5[72] , \MC_ARK_ARC_1_2/temp5[71] ,
         \MC_ARK_ARC_1_2/temp5[70] , \MC_ARK_ARC_1_2/temp5[69] ,
         \MC_ARK_ARC_1_2/temp5[68] , \MC_ARK_ARC_1_2/temp5[67] ,
         \MC_ARK_ARC_1_2/temp5[66] , \MC_ARK_ARC_1_2/temp5[65] ,
         \MC_ARK_ARC_1_2/temp5[64] , \MC_ARK_ARC_1_2/temp5[63] ,
         \MC_ARK_ARC_1_2/temp5[62] , \MC_ARK_ARC_1_2/temp5[61] ,
         \MC_ARK_ARC_1_2/temp5[60] , \MC_ARK_ARC_1_2/temp5[59] ,
         \MC_ARK_ARC_1_2/temp5[58] , \MC_ARK_ARC_1_2/temp5[57] ,
         \MC_ARK_ARC_1_2/temp5[56] , \MC_ARK_ARC_1_2/temp5[55] ,
         \MC_ARK_ARC_1_2/temp5[54] , \MC_ARK_ARC_1_2/temp5[53] ,
         \MC_ARK_ARC_1_2/temp5[52] , \MC_ARK_ARC_1_2/temp5[51] ,
         \MC_ARK_ARC_1_2/temp5[50] , \MC_ARK_ARC_1_2/temp5[49] ,
         \MC_ARK_ARC_1_2/temp5[48] , \MC_ARK_ARC_1_2/temp5[47] ,
         \MC_ARK_ARC_1_2/temp5[46] , \MC_ARK_ARC_1_2/temp5[45] ,
         \MC_ARK_ARC_1_2/temp5[43] , \MC_ARK_ARC_1_2/temp5[42] ,
         \MC_ARK_ARC_1_2/temp5[40] , \MC_ARK_ARC_1_2/temp5[39] ,
         \MC_ARK_ARC_1_2/temp5[38] , \MC_ARK_ARC_1_2/temp5[37] ,
         \MC_ARK_ARC_1_2/temp5[36] , \MC_ARK_ARC_1_2/temp5[35] ,
         \MC_ARK_ARC_1_2/temp5[34] , \MC_ARK_ARC_1_2/temp5[33] ,
         \MC_ARK_ARC_1_2/temp5[32] , \MC_ARK_ARC_1_2/temp5[31] ,
         \MC_ARK_ARC_1_2/temp5[30] , \MC_ARK_ARC_1_2/temp5[28] ,
         \MC_ARK_ARC_1_2/temp5[27] , \MC_ARK_ARC_1_2/temp5[26] ,
         \MC_ARK_ARC_1_2/temp5[25] , \MC_ARK_ARC_1_2/temp5[24] ,
         \MC_ARK_ARC_1_2/temp5[22] , \MC_ARK_ARC_1_2/temp5[21] ,
         \MC_ARK_ARC_1_2/temp5[20] , \MC_ARK_ARC_1_2/temp5[19] ,
         \MC_ARK_ARC_1_2/temp5[18] , \MC_ARK_ARC_1_2/temp5[16] ,
         \MC_ARK_ARC_1_2/temp5[13] , \MC_ARK_ARC_1_2/temp5[12] ,
         \MC_ARK_ARC_1_2/temp5[11] , \MC_ARK_ARC_1_2/temp5[10] ,
         \MC_ARK_ARC_1_2/temp5[9] , \MC_ARK_ARC_1_2/temp5[8] ,
         \MC_ARK_ARC_1_2/temp5[7] , \MC_ARK_ARC_1_2/temp5[6] ,
         \MC_ARK_ARC_1_2/temp5[5] , \MC_ARK_ARC_1_2/temp5[4] ,
         \MC_ARK_ARC_1_2/temp5[3] , \MC_ARK_ARC_1_2/temp5[2] ,
         \MC_ARK_ARC_1_2/temp5[1] , \MC_ARK_ARC_1_2/temp5[0] ,
         \MC_ARK_ARC_1_2/temp4[191] , \MC_ARK_ARC_1_2/temp4[190] ,
         \MC_ARK_ARC_1_2/temp4[189] , \MC_ARK_ARC_1_2/temp4[188] ,
         \MC_ARK_ARC_1_2/temp4[187] , \MC_ARK_ARC_1_2/temp4[186] ,
         \MC_ARK_ARC_1_2/temp4[185] , \MC_ARK_ARC_1_2/temp4[184] ,
         \MC_ARK_ARC_1_2/temp4[183] , \MC_ARK_ARC_1_2/temp4[182] ,
         \MC_ARK_ARC_1_2/temp4[181] , \MC_ARK_ARC_1_2/temp4[180] ,
         \MC_ARK_ARC_1_2/temp4[179] , \MC_ARK_ARC_1_2/temp4[178] ,
         \MC_ARK_ARC_1_2/temp4[177] , \MC_ARK_ARC_1_2/temp4[176] ,
         \MC_ARK_ARC_1_2/temp4[175] , \MC_ARK_ARC_1_2/temp4[174] ,
         \MC_ARK_ARC_1_2/temp4[173] , \MC_ARK_ARC_1_2/temp4[172] ,
         \MC_ARK_ARC_1_2/temp4[171] , \MC_ARK_ARC_1_2/temp4[170] ,
         \MC_ARK_ARC_1_2/temp4[169] , \MC_ARK_ARC_1_2/temp4[168] ,
         \MC_ARK_ARC_1_2/temp4[167] , \MC_ARK_ARC_1_2/temp4[166] ,
         \MC_ARK_ARC_1_2/temp4[165] , \MC_ARK_ARC_1_2/temp4[164] ,
         \MC_ARK_ARC_1_2/temp4[163] , \MC_ARK_ARC_1_2/temp4[162] ,
         \MC_ARK_ARC_1_2/temp4[161] , \MC_ARK_ARC_1_2/temp4[160] ,
         \MC_ARK_ARC_1_2/temp4[159] , \MC_ARK_ARC_1_2/temp4[158] ,
         \MC_ARK_ARC_1_2/temp4[157] , \MC_ARK_ARC_1_2/temp4[156] ,
         \MC_ARK_ARC_1_2/temp4[155] , \MC_ARK_ARC_1_2/temp4[154] ,
         \MC_ARK_ARC_1_2/temp4[153] , \MC_ARK_ARC_1_2/temp4[152] ,
         \MC_ARK_ARC_1_2/temp4[151] , \MC_ARK_ARC_1_2/temp4[150] ,
         \MC_ARK_ARC_1_2/temp4[149] , \MC_ARK_ARC_1_2/temp4[148] ,
         \MC_ARK_ARC_1_2/temp4[147] , \MC_ARK_ARC_1_2/temp4[146] ,
         \MC_ARK_ARC_1_2/temp4[145] , \MC_ARK_ARC_1_2/temp4[144] ,
         \MC_ARK_ARC_1_2/temp4[143] , \MC_ARK_ARC_1_2/temp4[142] ,
         \MC_ARK_ARC_1_2/temp4[141] , \MC_ARK_ARC_1_2/temp4[140] ,
         \MC_ARK_ARC_1_2/temp4[139] , \MC_ARK_ARC_1_2/temp4[138] ,
         \MC_ARK_ARC_1_2/temp4[137] , \MC_ARK_ARC_1_2/temp4[136] ,
         \MC_ARK_ARC_1_2/temp4[135] , \MC_ARK_ARC_1_2/temp4[134] ,
         \MC_ARK_ARC_1_2/temp4[133] , \MC_ARK_ARC_1_2/temp4[132] ,
         \MC_ARK_ARC_1_2/temp4[131] , \MC_ARK_ARC_1_2/temp4[130] ,
         \MC_ARK_ARC_1_2/temp4[129] , \MC_ARK_ARC_1_2/temp4[128] ,
         \MC_ARK_ARC_1_2/temp4[127] , \MC_ARK_ARC_1_2/temp4[126] ,
         \MC_ARK_ARC_1_2/temp4[125] , \MC_ARK_ARC_1_2/temp4[124] ,
         \MC_ARK_ARC_1_2/temp4[123] , \MC_ARK_ARC_1_2/temp4[122] ,
         \MC_ARK_ARC_1_2/temp4[121] , \MC_ARK_ARC_1_2/temp4[120] ,
         \MC_ARK_ARC_1_2/temp4[119] , \MC_ARK_ARC_1_2/temp4[118] ,
         \MC_ARK_ARC_1_2/temp4[117] , \MC_ARK_ARC_1_2/temp4[116] ,
         \MC_ARK_ARC_1_2/temp4[115] , \MC_ARK_ARC_1_2/temp4[114] ,
         \MC_ARK_ARC_1_2/temp4[113] , \MC_ARK_ARC_1_2/temp4[112] ,
         \MC_ARK_ARC_1_2/temp4[111] , \MC_ARK_ARC_1_2/temp4[110] ,
         \MC_ARK_ARC_1_2/temp4[109] , \MC_ARK_ARC_1_2/temp4[108] ,
         \MC_ARK_ARC_1_2/temp4[107] , \MC_ARK_ARC_1_2/temp4[106] ,
         \MC_ARK_ARC_1_2/temp4[105] , \MC_ARK_ARC_1_2/temp4[104] ,
         \MC_ARK_ARC_1_2/temp4[103] , \MC_ARK_ARC_1_2/temp4[102] ,
         \MC_ARK_ARC_1_2/temp4[101] , \MC_ARK_ARC_1_2/temp4[100] ,
         \MC_ARK_ARC_1_2/temp4[99] , \MC_ARK_ARC_1_2/temp4[98] ,
         \MC_ARK_ARC_1_2/temp4[97] , \MC_ARK_ARC_1_2/temp4[96] ,
         \MC_ARK_ARC_1_2/temp4[95] , \MC_ARK_ARC_1_2/temp4[94] ,
         \MC_ARK_ARC_1_2/temp4[93] , \MC_ARK_ARC_1_2/temp4[92] ,
         \MC_ARK_ARC_1_2/temp4[91] , \MC_ARK_ARC_1_2/temp4[90] ,
         \MC_ARK_ARC_1_2/temp4[89] , \MC_ARK_ARC_1_2/temp4[88] ,
         \MC_ARK_ARC_1_2/temp4[87] , \MC_ARK_ARC_1_2/temp4[86] ,
         \MC_ARK_ARC_1_2/temp4[85] , \MC_ARK_ARC_1_2/temp4[84] ,
         \MC_ARK_ARC_1_2/temp4[83] , \MC_ARK_ARC_1_2/temp4[82] ,
         \MC_ARK_ARC_1_2/temp4[81] , \MC_ARK_ARC_1_2/temp4[80] ,
         \MC_ARK_ARC_1_2/temp4[79] , \MC_ARK_ARC_1_2/temp4[78] ,
         \MC_ARK_ARC_1_2/temp4[77] , \MC_ARK_ARC_1_2/temp4[76] ,
         \MC_ARK_ARC_1_2/temp4[75] , \MC_ARK_ARC_1_2/temp4[74] ,
         \MC_ARK_ARC_1_2/temp4[73] , \MC_ARK_ARC_1_2/temp4[72] ,
         \MC_ARK_ARC_1_2/temp4[71] , \MC_ARK_ARC_1_2/temp4[70] ,
         \MC_ARK_ARC_1_2/temp4[69] , \MC_ARK_ARC_1_2/temp4[68] ,
         \MC_ARK_ARC_1_2/temp4[67] , \MC_ARK_ARC_1_2/temp4[66] ,
         \MC_ARK_ARC_1_2/temp4[65] , \MC_ARK_ARC_1_2/temp4[64] ,
         \MC_ARK_ARC_1_2/temp4[63] , \MC_ARK_ARC_1_2/temp4[62] ,
         \MC_ARK_ARC_1_2/temp4[61] , \MC_ARK_ARC_1_2/temp4[60] ,
         \MC_ARK_ARC_1_2/temp4[59] , \MC_ARK_ARC_1_2/temp4[58] ,
         \MC_ARK_ARC_1_2/temp4[57] , \MC_ARK_ARC_1_2/temp4[56] ,
         \MC_ARK_ARC_1_2/temp4[55] , \MC_ARK_ARC_1_2/temp4[54] ,
         \MC_ARK_ARC_1_2/temp4[53] , \MC_ARK_ARC_1_2/temp4[52] ,
         \MC_ARK_ARC_1_2/temp4[51] , \MC_ARK_ARC_1_2/temp4[50] ,
         \MC_ARK_ARC_1_2/temp4[49] , \MC_ARK_ARC_1_2/temp4[48] ,
         \MC_ARK_ARC_1_2/temp4[47] , \MC_ARK_ARC_1_2/temp4[46] ,
         \MC_ARK_ARC_1_2/temp4[45] , \MC_ARK_ARC_1_2/temp4[44] ,
         \MC_ARK_ARC_1_2/temp4[43] , \MC_ARK_ARC_1_2/temp4[42] ,
         \MC_ARK_ARC_1_2/temp4[41] , \MC_ARK_ARC_1_2/temp4[40] ,
         \MC_ARK_ARC_1_2/temp4[39] , \MC_ARK_ARC_1_2/temp4[38] ,
         \MC_ARK_ARC_1_2/temp4[37] , \MC_ARK_ARC_1_2/temp4[36] ,
         \MC_ARK_ARC_1_2/temp4[35] , \MC_ARK_ARC_1_2/temp4[34] ,
         \MC_ARK_ARC_1_2/temp4[33] , \MC_ARK_ARC_1_2/temp4[32] ,
         \MC_ARK_ARC_1_2/temp4[31] , \MC_ARK_ARC_1_2/temp4[30] ,
         \MC_ARK_ARC_1_2/temp4[29] , \MC_ARK_ARC_1_2/temp4[28] ,
         \MC_ARK_ARC_1_2/temp4[27] , \MC_ARK_ARC_1_2/temp4[26] ,
         \MC_ARK_ARC_1_2/temp4[25] , \MC_ARK_ARC_1_2/temp4[24] ,
         \MC_ARK_ARC_1_2/temp4[23] , \MC_ARK_ARC_1_2/temp4[22] ,
         \MC_ARK_ARC_1_2/temp4[21] , \MC_ARK_ARC_1_2/temp4[20] ,
         \MC_ARK_ARC_1_2/temp4[19] , \MC_ARK_ARC_1_2/temp4[18] ,
         \MC_ARK_ARC_1_2/temp4[17] , \MC_ARK_ARC_1_2/temp4[16] ,
         \MC_ARK_ARC_1_2/temp4[15] , \MC_ARK_ARC_1_2/temp4[14] ,
         \MC_ARK_ARC_1_2/temp4[13] , \MC_ARK_ARC_1_2/temp4[12] ,
         \MC_ARK_ARC_1_2/temp4[11] , \MC_ARK_ARC_1_2/temp4[10] ,
         \MC_ARK_ARC_1_2/temp4[9] , \MC_ARK_ARC_1_2/temp4[8] ,
         \MC_ARK_ARC_1_2/temp4[7] , \MC_ARK_ARC_1_2/temp4[6] ,
         \MC_ARK_ARC_1_2/temp4[5] , \MC_ARK_ARC_1_2/temp4[4] ,
         \MC_ARK_ARC_1_2/temp4[3] , \MC_ARK_ARC_1_2/temp4[2] ,
         \MC_ARK_ARC_1_2/temp4[1] , \MC_ARK_ARC_1_2/temp4[0] ,
         \MC_ARK_ARC_1_2/temp3[191] , \MC_ARK_ARC_1_2/temp3[190] ,
         \MC_ARK_ARC_1_2/temp3[189] , \MC_ARK_ARC_1_2/temp3[188] ,
         \MC_ARK_ARC_1_2/temp3[187] , \MC_ARK_ARC_1_2/temp3[186] ,
         \MC_ARK_ARC_1_2/temp3[185] , \MC_ARK_ARC_1_2/temp3[184] ,
         \MC_ARK_ARC_1_2/temp3[183] , \MC_ARK_ARC_1_2/temp3[182] ,
         \MC_ARK_ARC_1_2/temp3[181] , \MC_ARK_ARC_1_2/temp3[180] ,
         \MC_ARK_ARC_1_2/temp3[179] , \MC_ARK_ARC_1_2/temp3[178] ,
         \MC_ARK_ARC_1_2/temp3[177] , \MC_ARK_ARC_1_2/temp3[176] ,
         \MC_ARK_ARC_1_2/temp3[175] , \MC_ARK_ARC_1_2/temp3[174] ,
         \MC_ARK_ARC_1_2/temp3[173] , \MC_ARK_ARC_1_2/temp3[172] ,
         \MC_ARK_ARC_1_2/temp3[171] , \MC_ARK_ARC_1_2/temp3[170] ,
         \MC_ARK_ARC_1_2/temp3[169] , \MC_ARK_ARC_1_2/temp3[168] ,
         \MC_ARK_ARC_1_2/temp3[167] , \MC_ARK_ARC_1_2/temp3[166] ,
         \MC_ARK_ARC_1_2/temp3[165] , \MC_ARK_ARC_1_2/temp3[164] ,
         \MC_ARK_ARC_1_2/temp3[163] , \MC_ARK_ARC_1_2/temp3[162] ,
         \MC_ARK_ARC_1_2/temp3[161] , \MC_ARK_ARC_1_2/temp3[160] ,
         \MC_ARK_ARC_1_2/temp3[159] , \MC_ARK_ARC_1_2/temp3[158] ,
         \MC_ARK_ARC_1_2/temp3[157] , \MC_ARK_ARC_1_2/temp3[156] ,
         \MC_ARK_ARC_1_2/temp3[155] , \MC_ARK_ARC_1_2/temp3[154] ,
         \MC_ARK_ARC_1_2/temp3[153] , \MC_ARK_ARC_1_2/temp3[152] ,
         \MC_ARK_ARC_1_2/temp3[151] , \MC_ARK_ARC_1_2/temp3[150] ,
         \MC_ARK_ARC_1_2/temp3[149] , \MC_ARK_ARC_1_2/temp3[148] ,
         \MC_ARK_ARC_1_2/temp3[147] , \MC_ARK_ARC_1_2/temp3[146] ,
         \MC_ARK_ARC_1_2/temp3[145] , \MC_ARK_ARC_1_2/temp3[144] ,
         \MC_ARK_ARC_1_2/temp3[143] , \MC_ARK_ARC_1_2/temp3[142] ,
         \MC_ARK_ARC_1_2/temp3[141] , \MC_ARK_ARC_1_2/temp3[140] ,
         \MC_ARK_ARC_1_2/temp3[139] , \MC_ARK_ARC_1_2/temp3[138] ,
         \MC_ARK_ARC_1_2/temp3[137] , \MC_ARK_ARC_1_2/temp3[136] ,
         \MC_ARK_ARC_1_2/temp3[135] , \MC_ARK_ARC_1_2/temp3[134] ,
         \MC_ARK_ARC_1_2/temp3[133] , \MC_ARK_ARC_1_2/temp3[132] ,
         \MC_ARK_ARC_1_2/temp3[131] , \MC_ARK_ARC_1_2/temp3[130] ,
         \MC_ARK_ARC_1_2/temp3[129] , \MC_ARK_ARC_1_2/temp3[128] ,
         \MC_ARK_ARC_1_2/temp3[127] , \MC_ARK_ARC_1_2/temp3[126] ,
         \MC_ARK_ARC_1_2/temp3[125] , \MC_ARK_ARC_1_2/temp3[124] ,
         \MC_ARK_ARC_1_2/temp3[123] , \MC_ARK_ARC_1_2/temp3[122] ,
         \MC_ARK_ARC_1_2/temp3[121] , \MC_ARK_ARC_1_2/temp3[120] ,
         \MC_ARK_ARC_1_2/temp3[119] , \MC_ARK_ARC_1_2/temp3[118] ,
         \MC_ARK_ARC_1_2/temp3[117] , \MC_ARK_ARC_1_2/temp3[116] ,
         \MC_ARK_ARC_1_2/temp3[115] , \MC_ARK_ARC_1_2/temp3[114] ,
         \MC_ARK_ARC_1_2/temp3[113] , \MC_ARK_ARC_1_2/temp3[112] ,
         \MC_ARK_ARC_1_2/temp3[111] , \MC_ARK_ARC_1_2/temp3[110] ,
         \MC_ARK_ARC_1_2/temp3[109] , \MC_ARK_ARC_1_2/temp3[108] ,
         \MC_ARK_ARC_1_2/temp3[107] , \MC_ARK_ARC_1_2/temp3[106] ,
         \MC_ARK_ARC_1_2/temp3[105] , \MC_ARK_ARC_1_2/temp3[104] ,
         \MC_ARK_ARC_1_2/temp3[103] , \MC_ARK_ARC_1_2/temp3[102] ,
         \MC_ARK_ARC_1_2/temp3[101] , \MC_ARK_ARC_1_2/temp3[100] ,
         \MC_ARK_ARC_1_2/temp3[99] , \MC_ARK_ARC_1_2/temp3[98] ,
         \MC_ARK_ARC_1_2/temp3[97] , \MC_ARK_ARC_1_2/temp3[96] ,
         \MC_ARK_ARC_1_2/temp3[95] , \MC_ARK_ARC_1_2/temp3[94] ,
         \MC_ARK_ARC_1_2/temp3[93] , \MC_ARK_ARC_1_2/temp3[92] ,
         \MC_ARK_ARC_1_2/temp3[91] , \MC_ARK_ARC_1_2/temp3[90] ,
         \MC_ARK_ARC_1_2/temp3[89] , \MC_ARK_ARC_1_2/temp3[88] ,
         \MC_ARK_ARC_1_2/temp3[87] , \MC_ARK_ARC_1_2/temp3[86] ,
         \MC_ARK_ARC_1_2/temp3[85] , \MC_ARK_ARC_1_2/temp3[84] ,
         \MC_ARK_ARC_1_2/temp3[83] , \MC_ARK_ARC_1_2/temp3[82] ,
         \MC_ARK_ARC_1_2/temp3[81] , \MC_ARK_ARC_1_2/temp3[80] ,
         \MC_ARK_ARC_1_2/temp3[79] , \MC_ARK_ARC_1_2/temp3[78] ,
         \MC_ARK_ARC_1_2/temp3[77] , \MC_ARK_ARC_1_2/temp3[76] ,
         \MC_ARK_ARC_1_2/temp3[75] , \MC_ARK_ARC_1_2/temp3[74] ,
         \MC_ARK_ARC_1_2/temp3[73] , \MC_ARK_ARC_1_2/temp3[72] ,
         \MC_ARK_ARC_1_2/temp3[71] , \MC_ARK_ARC_1_2/temp3[70] ,
         \MC_ARK_ARC_1_2/temp3[69] , \MC_ARK_ARC_1_2/temp3[68] ,
         \MC_ARK_ARC_1_2/temp3[67] , \MC_ARK_ARC_1_2/temp3[66] ,
         \MC_ARK_ARC_1_2/temp3[65] , \MC_ARK_ARC_1_2/temp3[64] ,
         \MC_ARK_ARC_1_2/temp3[63] , \MC_ARK_ARC_1_2/temp3[62] ,
         \MC_ARK_ARC_1_2/temp3[61] , \MC_ARK_ARC_1_2/temp3[60] ,
         \MC_ARK_ARC_1_2/temp3[59] , \MC_ARK_ARC_1_2/temp3[58] ,
         \MC_ARK_ARC_1_2/temp3[57] , \MC_ARK_ARC_1_2/temp3[56] ,
         \MC_ARK_ARC_1_2/temp3[55] , \MC_ARK_ARC_1_2/temp3[54] ,
         \MC_ARK_ARC_1_2/temp3[53] , \MC_ARK_ARC_1_2/temp3[52] ,
         \MC_ARK_ARC_1_2/temp3[51] , \MC_ARK_ARC_1_2/temp3[50] ,
         \MC_ARK_ARC_1_2/temp3[49] , \MC_ARK_ARC_1_2/temp3[48] ,
         \MC_ARK_ARC_1_2/temp3[47] , \MC_ARK_ARC_1_2/temp3[46] ,
         \MC_ARK_ARC_1_2/temp3[45] , \MC_ARK_ARC_1_2/temp3[44] ,
         \MC_ARK_ARC_1_2/temp3[43] , \MC_ARK_ARC_1_2/temp3[42] ,
         \MC_ARK_ARC_1_2/temp3[41] , \MC_ARK_ARC_1_2/temp3[40] ,
         \MC_ARK_ARC_1_2/temp3[39] , \MC_ARK_ARC_1_2/temp3[38] ,
         \MC_ARK_ARC_1_2/temp3[37] , \MC_ARK_ARC_1_2/temp3[36] ,
         \MC_ARK_ARC_1_2/temp3[35] , \MC_ARK_ARC_1_2/temp3[34] ,
         \MC_ARK_ARC_1_2/temp3[33] , \MC_ARK_ARC_1_2/temp3[32] ,
         \MC_ARK_ARC_1_2/temp3[31] , \MC_ARK_ARC_1_2/temp3[30] ,
         \MC_ARK_ARC_1_2/temp3[29] , \MC_ARK_ARC_1_2/temp3[28] ,
         \MC_ARK_ARC_1_2/temp3[27] , \MC_ARK_ARC_1_2/temp3[26] ,
         \MC_ARK_ARC_1_2/temp3[25] , \MC_ARK_ARC_1_2/temp3[24] ,
         \MC_ARK_ARC_1_2/temp3[23] , \MC_ARK_ARC_1_2/temp3[22] ,
         \MC_ARK_ARC_1_2/temp3[21] , \MC_ARK_ARC_1_2/temp3[20] ,
         \MC_ARK_ARC_1_2/temp3[19] , \MC_ARK_ARC_1_2/temp3[18] ,
         \MC_ARK_ARC_1_2/temp3[17] , \MC_ARK_ARC_1_2/temp3[16] ,
         \MC_ARK_ARC_1_2/temp3[15] , \MC_ARK_ARC_1_2/temp3[14] ,
         \MC_ARK_ARC_1_2/temp3[13] , \MC_ARK_ARC_1_2/temp3[12] ,
         \MC_ARK_ARC_1_2/temp3[11] , \MC_ARK_ARC_1_2/temp3[10] ,
         \MC_ARK_ARC_1_2/temp3[9] , \MC_ARK_ARC_1_2/temp3[8] ,
         \MC_ARK_ARC_1_2/temp3[7] , \MC_ARK_ARC_1_2/temp3[6] ,
         \MC_ARK_ARC_1_2/temp3[5] , \MC_ARK_ARC_1_2/temp3[4] ,
         \MC_ARK_ARC_1_2/temp3[3] , \MC_ARK_ARC_1_2/temp3[2] ,
         \MC_ARK_ARC_1_2/temp3[1] , \MC_ARK_ARC_1_2/temp3[0] ,
         \MC_ARK_ARC_1_2/temp2[191] , \MC_ARK_ARC_1_2/temp2[190] ,
         \MC_ARK_ARC_1_2/temp2[189] , \MC_ARK_ARC_1_2/temp2[188] ,
         \MC_ARK_ARC_1_2/temp2[187] , \MC_ARK_ARC_1_2/temp2[186] ,
         \MC_ARK_ARC_1_2/temp2[185] , \MC_ARK_ARC_1_2/temp2[184] ,
         \MC_ARK_ARC_1_2/temp2[183] , \MC_ARK_ARC_1_2/temp2[182] ,
         \MC_ARK_ARC_1_2/temp2[181] , \MC_ARK_ARC_1_2/temp2[180] ,
         \MC_ARK_ARC_1_2/temp2[179] , \MC_ARK_ARC_1_2/temp2[178] ,
         \MC_ARK_ARC_1_2/temp2[177] , \MC_ARK_ARC_1_2/temp2[176] ,
         \MC_ARK_ARC_1_2/temp2[175] , \MC_ARK_ARC_1_2/temp2[174] ,
         \MC_ARK_ARC_1_2/temp2[173] , \MC_ARK_ARC_1_2/temp2[172] ,
         \MC_ARK_ARC_1_2/temp2[171] , \MC_ARK_ARC_1_2/temp2[170] ,
         \MC_ARK_ARC_1_2/temp2[169] , \MC_ARK_ARC_1_2/temp2[168] ,
         \MC_ARK_ARC_1_2/temp2[167] , \MC_ARK_ARC_1_2/temp2[166] ,
         \MC_ARK_ARC_1_2/temp2[165] , \MC_ARK_ARC_1_2/temp2[164] ,
         \MC_ARK_ARC_1_2/temp2[163] , \MC_ARK_ARC_1_2/temp2[162] ,
         \MC_ARK_ARC_1_2/temp2[161] , \MC_ARK_ARC_1_2/temp2[160] ,
         \MC_ARK_ARC_1_2/temp2[159] , \MC_ARK_ARC_1_2/temp2[158] ,
         \MC_ARK_ARC_1_2/temp2[157] , \MC_ARK_ARC_1_2/temp2[156] ,
         \MC_ARK_ARC_1_2/temp2[155] , \MC_ARK_ARC_1_2/temp2[154] ,
         \MC_ARK_ARC_1_2/temp2[153] , \MC_ARK_ARC_1_2/temp2[152] ,
         \MC_ARK_ARC_1_2/temp2[151] , \MC_ARK_ARC_1_2/temp2[150] ,
         \MC_ARK_ARC_1_2/temp2[149] , \MC_ARK_ARC_1_2/temp2[148] ,
         \MC_ARK_ARC_1_2/temp2[147] , \MC_ARK_ARC_1_2/temp2[146] ,
         \MC_ARK_ARC_1_2/temp2[145] , \MC_ARK_ARC_1_2/temp2[144] ,
         \MC_ARK_ARC_1_2/temp2[143] , \MC_ARK_ARC_1_2/temp2[142] ,
         \MC_ARK_ARC_1_2/temp2[141] , \MC_ARK_ARC_1_2/temp2[140] ,
         \MC_ARK_ARC_1_2/temp2[139] , \MC_ARK_ARC_1_2/temp2[138] ,
         \MC_ARK_ARC_1_2/temp2[137] , \MC_ARK_ARC_1_2/temp2[136] ,
         \MC_ARK_ARC_1_2/temp2[135] , \MC_ARK_ARC_1_2/temp2[134] ,
         \MC_ARK_ARC_1_2/temp2[133] , \MC_ARK_ARC_1_2/temp2[132] ,
         \MC_ARK_ARC_1_2/temp2[131] , \MC_ARK_ARC_1_2/temp2[130] ,
         \MC_ARK_ARC_1_2/temp2[129] , \MC_ARK_ARC_1_2/temp2[128] ,
         \MC_ARK_ARC_1_2/temp2[127] , \MC_ARK_ARC_1_2/temp2[126] ,
         \MC_ARK_ARC_1_2/temp2[125] , \MC_ARK_ARC_1_2/temp2[124] ,
         \MC_ARK_ARC_1_2/temp2[123] , \MC_ARK_ARC_1_2/temp2[122] ,
         \MC_ARK_ARC_1_2/temp2[121] , \MC_ARK_ARC_1_2/temp2[120] ,
         \MC_ARK_ARC_1_2/temp2[119] , \MC_ARK_ARC_1_2/temp2[118] ,
         \MC_ARK_ARC_1_2/temp2[117] , \MC_ARK_ARC_1_2/temp2[116] ,
         \MC_ARK_ARC_1_2/temp2[115] , \MC_ARK_ARC_1_2/temp2[114] ,
         \MC_ARK_ARC_1_2/temp2[113] , \MC_ARK_ARC_1_2/temp2[112] ,
         \MC_ARK_ARC_1_2/temp2[111] , \MC_ARK_ARC_1_2/temp2[110] ,
         \MC_ARK_ARC_1_2/temp2[109] , \MC_ARK_ARC_1_2/temp2[108] ,
         \MC_ARK_ARC_1_2/temp2[107] , \MC_ARK_ARC_1_2/temp2[106] ,
         \MC_ARK_ARC_1_2/temp2[105] , \MC_ARK_ARC_1_2/temp2[104] ,
         \MC_ARK_ARC_1_2/temp2[103] , \MC_ARK_ARC_1_2/temp2[102] ,
         \MC_ARK_ARC_1_2/temp2[101] , \MC_ARK_ARC_1_2/temp2[100] ,
         \MC_ARK_ARC_1_2/temp2[99] , \MC_ARK_ARC_1_2/temp2[98] ,
         \MC_ARK_ARC_1_2/temp2[97] , \MC_ARK_ARC_1_2/temp2[96] ,
         \MC_ARK_ARC_1_2/temp2[95] , \MC_ARK_ARC_1_2/temp2[94] ,
         \MC_ARK_ARC_1_2/temp2[93] , \MC_ARK_ARC_1_2/temp2[92] ,
         \MC_ARK_ARC_1_2/temp2[91] , \MC_ARK_ARC_1_2/temp2[90] ,
         \MC_ARK_ARC_1_2/temp2[89] , \MC_ARK_ARC_1_2/temp2[88] ,
         \MC_ARK_ARC_1_2/temp2[87] , \MC_ARK_ARC_1_2/temp2[86] ,
         \MC_ARK_ARC_1_2/temp2[85] , \MC_ARK_ARC_1_2/temp2[84] ,
         \MC_ARK_ARC_1_2/temp2[83] , \MC_ARK_ARC_1_2/temp2[82] ,
         \MC_ARK_ARC_1_2/temp2[81] , \MC_ARK_ARC_1_2/temp2[80] ,
         \MC_ARK_ARC_1_2/temp2[79] , \MC_ARK_ARC_1_2/temp2[78] ,
         \MC_ARK_ARC_1_2/temp2[77] , \MC_ARK_ARC_1_2/temp2[76] ,
         \MC_ARK_ARC_1_2/temp2[75] , \MC_ARK_ARC_1_2/temp2[74] ,
         \MC_ARK_ARC_1_2/temp2[73] , \MC_ARK_ARC_1_2/temp2[72] ,
         \MC_ARK_ARC_1_2/temp2[71] , \MC_ARK_ARC_1_2/temp2[70] ,
         \MC_ARK_ARC_1_2/temp2[69] , \MC_ARK_ARC_1_2/temp2[68] ,
         \MC_ARK_ARC_1_2/temp2[67] , \MC_ARK_ARC_1_2/temp2[66] ,
         \MC_ARK_ARC_1_2/temp2[65] , \MC_ARK_ARC_1_2/temp2[64] ,
         \MC_ARK_ARC_1_2/temp2[63] , \MC_ARK_ARC_1_2/temp2[62] ,
         \MC_ARK_ARC_1_2/temp2[61] , \MC_ARK_ARC_1_2/temp2[60] ,
         \MC_ARK_ARC_1_2/temp2[59] , \MC_ARK_ARC_1_2/temp2[58] ,
         \MC_ARK_ARC_1_2/temp2[57] , \MC_ARK_ARC_1_2/temp2[56] ,
         \MC_ARK_ARC_1_2/temp2[55] , \MC_ARK_ARC_1_2/temp2[54] ,
         \MC_ARK_ARC_1_2/temp2[53] , \MC_ARK_ARC_1_2/temp2[52] ,
         \MC_ARK_ARC_1_2/temp2[51] , \MC_ARK_ARC_1_2/temp2[50] ,
         \MC_ARK_ARC_1_2/temp2[49] , \MC_ARK_ARC_1_2/temp2[48] ,
         \MC_ARK_ARC_1_2/temp2[47] , \MC_ARK_ARC_1_2/temp2[46] ,
         \MC_ARK_ARC_1_2/temp2[45] , \MC_ARK_ARC_1_2/temp2[44] ,
         \MC_ARK_ARC_1_2/temp2[43] , \MC_ARK_ARC_1_2/temp2[42] ,
         \MC_ARK_ARC_1_2/temp2[41] , \MC_ARK_ARC_1_2/temp2[40] ,
         \MC_ARK_ARC_1_2/temp2[39] , \MC_ARK_ARC_1_2/temp2[38] ,
         \MC_ARK_ARC_1_2/temp2[37] , \MC_ARK_ARC_1_2/temp2[36] ,
         \MC_ARK_ARC_1_2/temp2[35] , \MC_ARK_ARC_1_2/temp2[34] ,
         \MC_ARK_ARC_1_2/temp2[33] , \MC_ARK_ARC_1_2/temp2[32] ,
         \MC_ARK_ARC_1_2/temp2[31] , \MC_ARK_ARC_1_2/temp2[30] ,
         \MC_ARK_ARC_1_2/temp2[29] , \MC_ARK_ARC_1_2/temp2[28] ,
         \MC_ARK_ARC_1_2/temp2[27] , \MC_ARK_ARC_1_2/temp2[26] ,
         \MC_ARK_ARC_1_2/temp2[25] , \MC_ARK_ARC_1_2/temp2[24] ,
         \MC_ARK_ARC_1_2/temp2[23] , \MC_ARK_ARC_1_2/temp2[22] ,
         \MC_ARK_ARC_1_2/temp2[21] , \MC_ARK_ARC_1_2/temp2[20] ,
         \MC_ARK_ARC_1_2/temp2[19] , \MC_ARK_ARC_1_2/temp2[18] ,
         \MC_ARK_ARC_1_2/temp2[17] , \MC_ARK_ARC_1_2/temp2[16] ,
         \MC_ARK_ARC_1_2/temp2[15] , \MC_ARK_ARC_1_2/temp2[14] ,
         \MC_ARK_ARC_1_2/temp2[13] , \MC_ARK_ARC_1_2/temp2[12] ,
         \MC_ARK_ARC_1_2/temp2[11] , \MC_ARK_ARC_1_2/temp2[10] ,
         \MC_ARK_ARC_1_2/temp2[9] , \MC_ARK_ARC_1_2/temp2[8] ,
         \MC_ARK_ARC_1_2/temp2[7] , \MC_ARK_ARC_1_2/temp2[6] ,
         \MC_ARK_ARC_1_2/temp2[5] , \MC_ARK_ARC_1_2/temp2[4] ,
         \MC_ARK_ARC_1_2/temp2[3] , \MC_ARK_ARC_1_2/temp2[2] ,
         \MC_ARK_ARC_1_2/temp2[1] , \MC_ARK_ARC_1_2/temp2[0] ,
         \MC_ARK_ARC_1_2/temp1[191] , \MC_ARK_ARC_1_2/temp1[190] ,
         \MC_ARK_ARC_1_2/temp1[189] , \MC_ARK_ARC_1_2/temp1[188] ,
         \MC_ARK_ARC_1_2/temp1[187] , \MC_ARK_ARC_1_2/temp1[186] ,
         \MC_ARK_ARC_1_2/temp1[185] , \MC_ARK_ARC_1_2/temp1[184] ,
         \MC_ARK_ARC_1_2/temp1[183] , \MC_ARK_ARC_1_2/temp1[182] ,
         \MC_ARK_ARC_1_2/temp1[181] , \MC_ARK_ARC_1_2/temp1[180] ,
         \MC_ARK_ARC_1_2/temp1[179] , \MC_ARK_ARC_1_2/temp1[178] ,
         \MC_ARK_ARC_1_2/temp1[177] , \MC_ARK_ARC_1_2/temp1[176] ,
         \MC_ARK_ARC_1_2/temp1[175] , \MC_ARK_ARC_1_2/temp1[174] ,
         \MC_ARK_ARC_1_2/temp1[173] , \MC_ARK_ARC_1_2/temp1[172] ,
         \MC_ARK_ARC_1_2/temp1[171] , \MC_ARK_ARC_1_2/temp1[170] ,
         \MC_ARK_ARC_1_2/temp1[169] , \MC_ARK_ARC_1_2/temp1[168] ,
         \MC_ARK_ARC_1_2/temp1[167] , \MC_ARK_ARC_1_2/temp1[166] ,
         \MC_ARK_ARC_1_2/temp1[165] , \MC_ARK_ARC_1_2/temp1[164] ,
         \MC_ARK_ARC_1_2/temp1[163] , \MC_ARK_ARC_1_2/temp1[162] ,
         \MC_ARK_ARC_1_2/temp1[161] , \MC_ARK_ARC_1_2/temp1[160] ,
         \MC_ARK_ARC_1_2/temp1[159] , \MC_ARK_ARC_1_2/temp1[158] ,
         \MC_ARK_ARC_1_2/temp1[157] , \MC_ARK_ARC_1_2/temp1[156] ,
         \MC_ARK_ARC_1_2/temp1[155] , \MC_ARK_ARC_1_2/temp1[154] ,
         \MC_ARK_ARC_1_2/temp1[153] , \MC_ARK_ARC_1_2/temp1[152] ,
         \MC_ARK_ARC_1_2/temp1[151] , \MC_ARK_ARC_1_2/temp1[150] ,
         \MC_ARK_ARC_1_2/temp1[149] , \MC_ARK_ARC_1_2/temp1[148] ,
         \MC_ARK_ARC_1_2/temp1[147] , \MC_ARK_ARC_1_2/temp1[146] ,
         \MC_ARK_ARC_1_2/temp1[145] , \MC_ARK_ARC_1_2/temp1[144] ,
         \MC_ARK_ARC_1_2/temp1[143] , \MC_ARK_ARC_1_2/temp1[142] ,
         \MC_ARK_ARC_1_2/temp1[141] , \MC_ARK_ARC_1_2/temp1[140] ,
         \MC_ARK_ARC_1_2/temp1[139] , \MC_ARK_ARC_1_2/temp1[138] ,
         \MC_ARK_ARC_1_2/temp1[137] , \MC_ARK_ARC_1_2/temp1[136] ,
         \MC_ARK_ARC_1_2/temp1[135] , \MC_ARK_ARC_1_2/temp1[134] ,
         \MC_ARK_ARC_1_2/temp1[133] , \MC_ARK_ARC_1_2/temp1[132] ,
         \MC_ARK_ARC_1_2/temp1[131] , \MC_ARK_ARC_1_2/temp1[130] ,
         \MC_ARK_ARC_1_2/temp1[129] , \MC_ARK_ARC_1_2/temp1[128] ,
         \MC_ARK_ARC_1_2/temp1[127] , \MC_ARK_ARC_1_2/temp1[126] ,
         \MC_ARK_ARC_1_2/temp1[125] , \MC_ARK_ARC_1_2/temp1[124] ,
         \MC_ARK_ARC_1_2/temp1[123] , \MC_ARK_ARC_1_2/temp1[122] ,
         \MC_ARK_ARC_1_2/temp1[121] , \MC_ARK_ARC_1_2/temp1[120] ,
         \MC_ARK_ARC_1_2/temp1[119] , \MC_ARK_ARC_1_2/temp1[118] ,
         \MC_ARK_ARC_1_2/temp1[117] , \MC_ARK_ARC_1_2/temp1[116] ,
         \MC_ARK_ARC_1_2/temp1[115] , \MC_ARK_ARC_1_2/temp1[114] ,
         \MC_ARK_ARC_1_2/temp1[113] , \MC_ARK_ARC_1_2/temp1[112] ,
         \MC_ARK_ARC_1_2/temp1[111] , \MC_ARK_ARC_1_2/temp1[110] ,
         \MC_ARK_ARC_1_2/temp1[109] , \MC_ARK_ARC_1_2/temp1[108] ,
         \MC_ARK_ARC_1_2/temp1[107] , \MC_ARK_ARC_1_2/temp1[106] ,
         \MC_ARK_ARC_1_2/temp1[105] , \MC_ARK_ARC_1_2/temp1[104] ,
         \MC_ARK_ARC_1_2/temp1[103] , \MC_ARK_ARC_1_2/temp1[102] ,
         \MC_ARK_ARC_1_2/temp1[101] , \MC_ARK_ARC_1_2/temp1[100] ,
         \MC_ARK_ARC_1_2/temp1[99] , \MC_ARK_ARC_1_2/temp1[98] ,
         \MC_ARK_ARC_1_2/temp1[97] , \MC_ARK_ARC_1_2/temp1[96] ,
         \MC_ARK_ARC_1_2/temp1[95] , \MC_ARK_ARC_1_2/temp1[94] ,
         \MC_ARK_ARC_1_2/temp1[93] , \MC_ARK_ARC_1_2/temp1[92] ,
         \MC_ARK_ARC_1_2/temp1[91] , \MC_ARK_ARC_1_2/temp1[90] ,
         \MC_ARK_ARC_1_2/temp1[89] , \MC_ARK_ARC_1_2/temp1[88] ,
         \MC_ARK_ARC_1_2/temp1[87] , \MC_ARK_ARC_1_2/temp1[86] ,
         \MC_ARK_ARC_1_2/temp1[85] , \MC_ARK_ARC_1_2/temp1[84] ,
         \MC_ARK_ARC_1_2/temp1[83] , \MC_ARK_ARC_1_2/temp1[82] ,
         \MC_ARK_ARC_1_2/temp1[81] , \MC_ARK_ARC_1_2/temp1[80] ,
         \MC_ARK_ARC_1_2/temp1[79] , \MC_ARK_ARC_1_2/temp1[78] ,
         \MC_ARK_ARC_1_2/temp1[77] , \MC_ARK_ARC_1_2/temp1[76] ,
         \MC_ARK_ARC_1_2/temp1[75] , \MC_ARK_ARC_1_2/temp1[74] ,
         \MC_ARK_ARC_1_2/temp1[73] , \MC_ARK_ARC_1_2/temp1[72] ,
         \MC_ARK_ARC_1_2/temp1[71] , \MC_ARK_ARC_1_2/temp1[70] ,
         \MC_ARK_ARC_1_2/temp1[69] , \MC_ARK_ARC_1_2/temp1[68] ,
         \MC_ARK_ARC_1_2/temp1[67] , \MC_ARK_ARC_1_2/temp1[66] ,
         \MC_ARK_ARC_1_2/temp1[65] , \MC_ARK_ARC_1_2/temp1[64] ,
         \MC_ARK_ARC_1_2/temp1[63] , \MC_ARK_ARC_1_2/temp1[62] ,
         \MC_ARK_ARC_1_2/temp1[61] , \MC_ARK_ARC_1_2/temp1[60] ,
         \MC_ARK_ARC_1_2/temp1[59] , \MC_ARK_ARC_1_2/temp1[58] ,
         \MC_ARK_ARC_1_2/temp1[57] , \MC_ARK_ARC_1_2/temp1[56] ,
         \MC_ARK_ARC_1_2/temp1[55] , \MC_ARK_ARC_1_2/temp1[54] ,
         \MC_ARK_ARC_1_2/temp1[53] , \MC_ARK_ARC_1_2/temp1[52] ,
         \MC_ARK_ARC_1_2/temp1[51] , \MC_ARK_ARC_1_2/temp1[50] ,
         \MC_ARK_ARC_1_2/temp1[49] , \MC_ARK_ARC_1_2/temp1[48] ,
         \MC_ARK_ARC_1_2/temp1[47] , \MC_ARK_ARC_1_2/temp1[46] ,
         \MC_ARK_ARC_1_2/temp1[45] , \MC_ARK_ARC_1_2/temp1[44] ,
         \MC_ARK_ARC_1_2/temp1[43] , \MC_ARK_ARC_1_2/temp1[42] ,
         \MC_ARK_ARC_1_2/temp1[41] , \MC_ARK_ARC_1_2/temp1[40] ,
         \MC_ARK_ARC_1_2/temp1[39] , \MC_ARK_ARC_1_2/temp1[38] ,
         \MC_ARK_ARC_1_2/temp1[37] , \MC_ARK_ARC_1_2/temp1[36] ,
         \MC_ARK_ARC_1_2/temp1[35] , \MC_ARK_ARC_1_2/temp1[34] ,
         \MC_ARK_ARC_1_2/temp1[33] , \MC_ARK_ARC_1_2/temp1[32] ,
         \MC_ARK_ARC_1_2/temp1[31] , \MC_ARK_ARC_1_2/temp1[30] ,
         \MC_ARK_ARC_1_2/temp1[29] , \MC_ARK_ARC_1_2/temp1[28] ,
         \MC_ARK_ARC_1_2/temp1[27] , \MC_ARK_ARC_1_2/temp1[26] ,
         \MC_ARK_ARC_1_2/temp1[25] , \MC_ARK_ARC_1_2/temp1[24] ,
         \MC_ARK_ARC_1_2/temp1[23] , \MC_ARK_ARC_1_2/temp1[22] ,
         \MC_ARK_ARC_1_2/temp1[21] , \MC_ARK_ARC_1_2/temp1[20] ,
         \MC_ARK_ARC_1_2/temp1[19] , \MC_ARK_ARC_1_2/temp1[18] ,
         \MC_ARK_ARC_1_2/temp1[17] , \MC_ARK_ARC_1_2/temp1[16] ,
         \MC_ARK_ARC_1_2/temp1[15] , \MC_ARK_ARC_1_2/temp1[14] ,
         \MC_ARK_ARC_1_2/temp1[13] , \MC_ARK_ARC_1_2/temp1[12] ,
         \MC_ARK_ARC_1_2/temp1[11] , \MC_ARK_ARC_1_2/temp1[10] ,
         \MC_ARK_ARC_1_2/temp1[9] , \MC_ARK_ARC_1_2/temp1[8] ,
         \MC_ARK_ARC_1_2/temp1[7] , \MC_ARK_ARC_1_2/temp1[6] ,
         \MC_ARK_ARC_1_2/temp1[5] , \MC_ARK_ARC_1_2/temp1[4] ,
         \MC_ARK_ARC_1_2/temp1[3] , \MC_ARK_ARC_1_2/temp1[2] ,
         \MC_ARK_ARC_1_2/temp1[1] , \MC_ARK_ARC_1_2/temp1[0] ,
         \MC_ARK_ARC_1_2/buf_keyinput[184] ,
         \MC_ARK_ARC_1_2/buf_keyinput[177] ,
         \MC_ARK_ARC_1_2/buf_keyinput[172] ,
         \MC_ARK_ARC_1_2/buf_keyinput[143] ,
         \MC_ARK_ARC_1_2/buf_keyinput[129] ,
         \MC_ARK_ARC_1_2/buf_keyinput[118] ,
         \MC_ARK_ARC_1_2/buf_keyinput[112] ,
         \MC_ARK_ARC_1_2/buf_keyinput[107] , \MC_ARK_ARC_1_2/buf_keyinput[94] ,
         \MC_ARK_ARC_1_2/buf_keyinput[87] , \MC_ARK_ARC_1_2/buf_keyinput[76] ,
         \MC_ARK_ARC_1_2/buf_keyinput[69] , \MC_ARK_ARC_1_2/buf_keyinput[45] ,
         \MC_ARK_ARC_1_2/buf_keyinput[33] ,
         \MC_ARK_ARC_1_2/buf_datainput[191] ,
         \MC_ARK_ARC_1_2/buf_datainput[190] ,
         \MC_ARK_ARC_1_2/buf_datainput[189] ,
         \MC_ARK_ARC_1_2/buf_datainput[188] ,
         \MC_ARK_ARC_1_2/buf_datainput[186] ,
         \MC_ARK_ARC_1_2/buf_datainput[185] ,
         \MC_ARK_ARC_1_2/buf_datainput[184] ,
         \MC_ARK_ARC_1_2/buf_datainput[183] ,
         \MC_ARK_ARC_1_2/buf_datainput[182] ,
         \MC_ARK_ARC_1_2/buf_datainput[181] ,
         \MC_ARK_ARC_1_2/buf_datainput[180] ,
         \MC_ARK_ARC_1_2/buf_datainput[178] ,
         \MC_ARK_ARC_1_2/buf_datainput[176] ,
         \MC_ARK_ARC_1_2/buf_datainput[175] ,
         \MC_ARK_ARC_1_2/buf_datainput[174] ,
         \MC_ARK_ARC_1_2/buf_datainput[173] ,
         \MC_ARK_ARC_1_2/buf_datainput[172] ,
         \MC_ARK_ARC_1_2/buf_datainput[169] ,
         \MC_ARK_ARC_1_2/buf_datainput[168] ,
         \MC_ARK_ARC_1_2/buf_datainput[167] ,
         \MC_ARK_ARC_1_2/buf_datainput[166] ,
         \MC_ARK_ARC_1_2/buf_datainput[165] ,
         \MC_ARK_ARC_1_2/buf_datainput[164] ,
         \MC_ARK_ARC_1_2/buf_datainput[163] ,
         \MC_ARK_ARC_1_2/buf_datainput[162] ,
         \MC_ARK_ARC_1_2/buf_datainput[161] ,
         \MC_ARK_ARC_1_2/buf_datainput[160] ,
         \MC_ARK_ARC_1_2/buf_datainput[158] ,
         \MC_ARK_ARC_1_2/buf_datainput[157] ,
         \MC_ARK_ARC_1_2/buf_datainput[156] ,
         \MC_ARK_ARC_1_2/buf_datainput[155] ,
         \MC_ARK_ARC_1_2/buf_datainput[154] ,
         \MC_ARK_ARC_1_2/buf_datainput[153] ,
         \MC_ARK_ARC_1_2/buf_datainput[152] ,
         \MC_ARK_ARC_1_2/buf_datainput[151] ,
         \MC_ARK_ARC_1_2/buf_datainput[150] ,
         \MC_ARK_ARC_1_2/buf_datainput[148] ,
         \MC_ARK_ARC_1_2/buf_datainput[146] ,
         \MC_ARK_ARC_1_2/buf_datainput[145] ,
         \MC_ARK_ARC_1_2/buf_datainput[144] ,
         \MC_ARK_ARC_1_2/buf_datainput[143] ,
         \MC_ARK_ARC_1_2/buf_datainput[142] ,
         \MC_ARK_ARC_1_2/buf_datainput[140] ,
         \MC_ARK_ARC_1_2/buf_datainput[139] ,
         \MC_ARK_ARC_1_2/buf_datainput[138] ,
         \MC_ARK_ARC_1_2/buf_datainput[137] ,
         \MC_ARK_ARC_1_2/buf_datainput[136] ,
         \MC_ARK_ARC_1_2/buf_datainput[134] ,
         \MC_ARK_ARC_1_2/buf_datainput[132] ,
         \MC_ARK_ARC_1_2/buf_datainput[131] ,
         \MC_ARK_ARC_1_2/buf_datainput[130] ,
         \MC_ARK_ARC_1_2/buf_datainput[129] ,
         \MC_ARK_ARC_1_2/buf_datainput[128] ,
         \MC_ARK_ARC_1_2/buf_datainput[127] ,
         \MC_ARK_ARC_1_2/buf_datainput[126] ,
         \MC_ARK_ARC_1_2/buf_datainput[125] ,
         \MC_ARK_ARC_1_2/buf_datainput[124] ,
         \MC_ARK_ARC_1_2/buf_datainput[122] ,
         \MC_ARK_ARC_1_2/buf_datainput[121] ,
         \MC_ARK_ARC_1_2/buf_datainput[120] ,
         \MC_ARK_ARC_1_2/buf_datainput[118] ,
         \MC_ARK_ARC_1_2/buf_datainput[116] ,
         \MC_ARK_ARC_1_2/buf_datainput[115] ,
         \MC_ARK_ARC_1_2/buf_datainput[114] ,
         \MC_ARK_ARC_1_2/buf_datainput[113] ,
         \MC_ARK_ARC_1_2/buf_datainput[112] ,
         \MC_ARK_ARC_1_2/buf_datainput[110] ,
         \MC_ARK_ARC_1_2/buf_datainput[109] ,
         \MC_ARK_ARC_1_2/buf_datainput[107] ,
         \MC_ARK_ARC_1_2/buf_datainput[106] ,
         \MC_ARK_ARC_1_2/buf_datainput[105] ,
         \MC_ARK_ARC_1_2/buf_datainput[104] ,
         \MC_ARK_ARC_1_2/buf_datainput[103] ,
         \MC_ARK_ARC_1_2/buf_datainput[102] ,
         \MC_ARK_ARC_1_2/buf_datainput[101] ,
         \MC_ARK_ARC_1_2/buf_datainput[100] ,
         \MC_ARK_ARC_1_2/buf_datainput[98] ,
         \MC_ARK_ARC_1_2/buf_datainput[97] ,
         \MC_ARK_ARC_1_2/buf_datainput[96] ,
         \MC_ARK_ARC_1_2/buf_datainput[95] ,
         \MC_ARK_ARC_1_2/buf_datainput[94] ,
         \MC_ARK_ARC_1_2/buf_datainput[92] ,
         \MC_ARK_ARC_1_2/buf_datainput[91] ,
         \MC_ARK_ARC_1_2/buf_datainput[90] ,
         \MC_ARK_ARC_1_2/buf_datainput[89] ,
         \MC_ARK_ARC_1_2/buf_datainput[88] ,
         \MC_ARK_ARC_1_2/buf_datainput[86] ,
         \MC_ARK_ARC_1_2/buf_datainput[85] ,
         \MC_ARK_ARC_1_2/buf_datainput[84] ,
         \MC_ARK_ARC_1_2/buf_datainput[83] ,
         \MC_ARK_ARC_1_2/buf_datainput[82] ,
         \MC_ARK_ARC_1_2/buf_datainput[81] ,
         \MC_ARK_ARC_1_2/buf_datainput[80] ,
         \MC_ARK_ARC_1_2/buf_datainput[79] ,
         \MC_ARK_ARC_1_2/buf_datainput[78] ,
         \MC_ARK_ARC_1_2/buf_datainput[77] ,
         \MC_ARK_ARC_1_2/buf_datainput[76] ,
         \MC_ARK_ARC_1_2/buf_datainput[75] ,
         \MC_ARK_ARC_1_2/buf_datainput[74] ,
         \MC_ARK_ARC_1_2/buf_datainput[73] ,
         \MC_ARK_ARC_1_2/buf_datainput[72] ,
         \MC_ARK_ARC_1_2/buf_datainput[71] ,
         \MC_ARK_ARC_1_2/buf_datainput[70] ,
         \MC_ARK_ARC_1_2/buf_datainput[68] ,
         \MC_ARK_ARC_1_2/buf_datainput[67] ,
         \MC_ARK_ARC_1_2/buf_datainput[66] ,
         \MC_ARK_ARC_1_2/buf_datainput[65] ,
         \MC_ARK_ARC_1_2/buf_datainput[64] ,
         \MC_ARK_ARC_1_2/buf_datainput[63] ,
         \MC_ARK_ARC_1_2/buf_datainput[62] ,
         \MC_ARK_ARC_1_2/buf_datainput[61] ,
         \MC_ARK_ARC_1_2/buf_datainput[60] ,
         \MC_ARK_ARC_1_2/buf_datainput[58] ,
         \MC_ARK_ARC_1_2/buf_datainput[57] ,
         \MC_ARK_ARC_1_2/buf_datainput[56] ,
         \MC_ARK_ARC_1_2/buf_datainput[55] ,
         \MC_ARK_ARC_1_2/buf_datainput[54] ,
         \MC_ARK_ARC_1_2/buf_datainput[53] ,
         \MC_ARK_ARC_1_2/buf_datainput[52] ,
         \MC_ARK_ARC_1_2/buf_datainput[50] ,
         \MC_ARK_ARC_1_2/buf_datainput[49] ,
         \MC_ARK_ARC_1_2/buf_datainput[48] ,
         \MC_ARK_ARC_1_2/buf_datainput[47] ,
         \MC_ARK_ARC_1_2/buf_datainput[46] ,
         \MC_ARK_ARC_1_2/buf_datainput[45] ,
         \MC_ARK_ARC_1_2/buf_datainput[44] ,
         \MC_ARK_ARC_1_2/buf_datainput[43] ,
         \MC_ARK_ARC_1_2/buf_datainput[42] ,
         \MC_ARK_ARC_1_2/buf_datainput[41] ,
         \MC_ARK_ARC_1_2/buf_datainput[40] ,
         \MC_ARK_ARC_1_2/buf_datainput[38] ,
         \MC_ARK_ARC_1_2/buf_datainput[37] ,
         \MC_ARK_ARC_1_2/buf_datainput[36] ,
         \MC_ARK_ARC_1_2/buf_datainput[35] ,
         \MC_ARK_ARC_1_2/buf_datainput[34] ,
         \MC_ARK_ARC_1_2/buf_datainput[33] ,
         \MC_ARK_ARC_1_2/buf_datainput[31] ,
         \MC_ARK_ARC_1_2/buf_datainput[30] ,
         \MC_ARK_ARC_1_2/buf_datainput[29] ,
         \MC_ARK_ARC_1_2/buf_datainput[27] ,
         \MC_ARK_ARC_1_2/buf_datainput[26] ,
         \MC_ARK_ARC_1_2/buf_datainput[25] ,
         \MC_ARK_ARC_1_2/buf_datainput[24] ,
         \MC_ARK_ARC_1_2/buf_datainput[23] ,
         \MC_ARK_ARC_1_2/buf_datainput[22] ,
         \MC_ARK_ARC_1_2/buf_datainput[20] ,
         \MC_ARK_ARC_1_2/buf_datainput[19] ,
         \MC_ARK_ARC_1_2/buf_datainput[18] ,
         \MC_ARK_ARC_1_2/buf_datainput[17] ,
         \MC_ARK_ARC_1_2/buf_datainput[16] ,
         \MC_ARK_ARC_1_2/buf_datainput[15] ,
         \MC_ARK_ARC_1_2/buf_datainput[14] ,
         \MC_ARK_ARC_1_2/buf_datainput[13] ,
         \MC_ARK_ARC_1_2/buf_datainput[12] ,
         \MC_ARK_ARC_1_2/buf_datainput[11] ,
         \MC_ARK_ARC_1_2/buf_datainput[10] , \MC_ARK_ARC_1_2/buf_datainput[9] ,
         \MC_ARK_ARC_1_2/buf_datainput[8] , \MC_ARK_ARC_1_2/buf_datainput[7] ,
         \MC_ARK_ARC_1_2/buf_datainput[6] , \MC_ARK_ARC_1_2/buf_datainput[5] ,
         \MC_ARK_ARC_1_2/buf_datainput[4] , \MC_ARK_ARC_1_2/buf_datainput[1] ,
         \MC_ARK_ARC_1_2/buf_datainput[0] , \MC_ARK_ARC_1_3/temp6[191] ,
         \MC_ARK_ARC_1_3/temp6[190] , \MC_ARK_ARC_1_3/temp6[189] ,
         \MC_ARK_ARC_1_3/temp6[188] , \MC_ARK_ARC_1_3/temp6[187] ,
         \MC_ARK_ARC_1_3/temp6[186] , \MC_ARK_ARC_1_3/temp6[185] ,
         \MC_ARK_ARC_1_3/temp6[184] , \MC_ARK_ARC_1_3/temp6[183] ,
         \MC_ARK_ARC_1_3/temp6[182] , \MC_ARK_ARC_1_3/temp6[181] ,
         \MC_ARK_ARC_1_3/temp6[180] , \MC_ARK_ARC_1_3/temp6[177] ,
         \MC_ARK_ARC_1_3/temp6[176] , \MC_ARK_ARC_1_3/temp6[175] ,
         \MC_ARK_ARC_1_3/temp6[174] , \MC_ARK_ARC_1_3/temp6[173] ,
         \MC_ARK_ARC_1_3/temp6[172] , \MC_ARK_ARC_1_3/temp6[171] ,
         \MC_ARK_ARC_1_3/temp6[170] , \MC_ARK_ARC_1_3/temp6[169] ,
         \MC_ARK_ARC_1_3/temp6[168] , \MC_ARK_ARC_1_3/temp6[166] ,
         \MC_ARK_ARC_1_3/temp6[165] , \MC_ARK_ARC_1_3/temp6[164] ,
         \MC_ARK_ARC_1_3/temp6[163] , \MC_ARK_ARC_1_3/temp6[162] ,
         \MC_ARK_ARC_1_3/temp6[161] , \MC_ARK_ARC_1_3/temp6[160] ,
         \MC_ARK_ARC_1_3/temp6[159] , \MC_ARK_ARC_1_3/temp6[158] ,
         \MC_ARK_ARC_1_3/temp6[157] , \MC_ARK_ARC_1_3/temp6[156] ,
         \MC_ARK_ARC_1_3/temp6[155] , \MC_ARK_ARC_1_3/temp6[154] ,
         \MC_ARK_ARC_1_3/temp6[153] , \MC_ARK_ARC_1_3/temp6[152] ,
         \MC_ARK_ARC_1_3/temp6[151] , \MC_ARK_ARC_1_3/temp6[150] ,
         \MC_ARK_ARC_1_3/temp6[149] , \MC_ARK_ARC_1_3/temp6[148] ,
         \MC_ARK_ARC_1_3/temp6[147] , \MC_ARK_ARC_1_3/temp6[145] ,
         \MC_ARK_ARC_1_3/temp6[144] , \MC_ARK_ARC_1_3/temp6[143] ,
         \MC_ARK_ARC_1_3/temp6[142] , \MC_ARK_ARC_1_3/temp6[141] ,
         \MC_ARK_ARC_1_3/temp6[140] , \MC_ARK_ARC_1_3/temp6[139] ,
         \MC_ARK_ARC_1_3/temp6[138] , \MC_ARK_ARC_1_3/temp6[137] ,
         \MC_ARK_ARC_1_3/temp6[136] , \MC_ARK_ARC_1_3/temp6[135] ,
         \MC_ARK_ARC_1_3/temp6[134] , \MC_ARK_ARC_1_3/temp6[133] ,
         \MC_ARK_ARC_1_3/temp6[132] , \MC_ARK_ARC_1_3/temp6[129] ,
         \MC_ARK_ARC_1_3/temp6[128] , \MC_ARK_ARC_1_3/temp6[127] ,
         \MC_ARK_ARC_1_3/temp6[126] , \MC_ARK_ARC_1_3/temp6[125] ,
         \MC_ARK_ARC_1_3/temp6[124] , \MC_ARK_ARC_1_3/temp6[123] ,
         \MC_ARK_ARC_1_3/temp6[122] , \MC_ARK_ARC_1_3/temp6[121] ,
         \MC_ARK_ARC_1_3/temp6[120] , \MC_ARK_ARC_1_3/temp6[119] ,
         \MC_ARK_ARC_1_3/temp6[118] , \MC_ARK_ARC_1_3/temp6[117] ,
         \MC_ARK_ARC_1_3/temp6[116] , \MC_ARK_ARC_1_3/temp6[115] ,
         \MC_ARK_ARC_1_3/temp6[114] , \MC_ARK_ARC_1_3/temp6[113] ,
         \MC_ARK_ARC_1_3/temp6[112] , \MC_ARK_ARC_1_3/temp6[111] ,
         \MC_ARK_ARC_1_3/temp6[110] , \MC_ARK_ARC_1_3/temp6[109] ,
         \MC_ARK_ARC_1_3/temp6[108] , \MC_ARK_ARC_1_3/temp6[107] ,
         \MC_ARK_ARC_1_3/temp6[106] , \MC_ARK_ARC_1_3/temp6[105] ,
         \MC_ARK_ARC_1_3/temp6[104] , \MC_ARK_ARC_1_3/temp6[103] ,
         \MC_ARK_ARC_1_3/temp6[102] , \MC_ARK_ARC_1_3/temp6[101] ,
         \MC_ARK_ARC_1_3/temp6[100] , \MC_ARK_ARC_1_3/temp6[99] ,
         \MC_ARK_ARC_1_3/temp6[98] , \MC_ARK_ARC_1_3/temp6[97] ,
         \MC_ARK_ARC_1_3/temp6[96] , \MC_ARK_ARC_1_3/temp6[95] ,
         \MC_ARK_ARC_1_3/temp6[94] , \MC_ARK_ARC_1_3/temp6[93] ,
         \MC_ARK_ARC_1_3/temp6[91] , \MC_ARK_ARC_1_3/temp6[90] ,
         \MC_ARK_ARC_1_3/temp6[89] , \MC_ARK_ARC_1_3/temp6[88] ,
         \MC_ARK_ARC_1_3/temp6[87] , \MC_ARK_ARC_1_3/temp6[86] ,
         \MC_ARK_ARC_1_3/temp6[85] , \MC_ARK_ARC_1_3/temp6[84] ,
         \MC_ARK_ARC_1_3/temp6[82] , \MC_ARK_ARC_1_3/temp6[81] ,
         \MC_ARK_ARC_1_3/temp6[80] , \MC_ARK_ARC_1_3/temp6[79] ,
         \MC_ARK_ARC_1_3/temp6[78] , \MC_ARK_ARC_1_3/temp6[76] ,
         \MC_ARK_ARC_1_3/temp6[75] , \MC_ARK_ARC_1_3/temp6[74] ,
         \MC_ARK_ARC_1_3/temp6[73] , \MC_ARK_ARC_1_3/temp6[72] ,
         \MC_ARK_ARC_1_3/temp6[71] , \MC_ARK_ARC_1_3/temp6[70] ,
         \MC_ARK_ARC_1_3/temp6[69] , \MC_ARK_ARC_1_3/temp6[68] ,
         \MC_ARK_ARC_1_3/temp6[67] , \MC_ARK_ARC_1_3/temp6[66] ,
         \MC_ARK_ARC_1_3/temp6[65] , \MC_ARK_ARC_1_3/temp6[64] ,
         \MC_ARK_ARC_1_3/temp6[63] , \MC_ARK_ARC_1_3/temp6[62] ,
         \MC_ARK_ARC_1_3/temp6[61] , \MC_ARK_ARC_1_3/temp6[60] ,
         \MC_ARK_ARC_1_3/temp6[58] , \MC_ARK_ARC_1_3/temp6[57] ,
         \MC_ARK_ARC_1_3/temp6[56] , \MC_ARK_ARC_1_3/temp6[55] ,
         \MC_ARK_ARC_1_3/temp6[54] , \MC_ARK_ARC_1_3/temp6[53] ,
         \MC_ARK_ARC_1_3/temp6[52] , \MC_ARK_ARC_1_3/temp6[51] ,
         \MC_ARK_ARC_1_3/temp6[50] , \MC_ARK_ARC_1_3/temp6[49] ,
         \MC_ARK_ARC_1_3/temp6[48] , \MC_ARK_ARC_1_3/temp6[47] ,
         \MC_ARK_ARC_1_3/temp6[46] , \MC_ARK_ARC_1_3/temp6[45] ,
         \MC_ARK_ARC_1_3/temp6[44] , \MC_ARK_ARC_1_3/temp6[43] ,
         \MC_ARK_ARC_1_3/temp6[42] , \MC_ARK_ARC_1_3/temp6[41] ,
         \MC_ARK_ARC_1_3/temp6[40] , \MC_ARK_ARC_1_3/temp6[39] ,
         \MC_ARK_ARC_1_3/temp6[38] , \MC_ARK_ARC_1_3/temp6[37] ,
         \MC_ARK_ARC_1_3/temp6[36] , \MC_ARK_ARC_1_3/temp6[34] ,
         \MC_ARK_ARC_1_3/temp6[33] , \MC_ARK_ARC_1_3/temp6[32] ,
         \MC_ARK_ARC_1_3/temp6[31] , \MC_ARK_ARC_1_3/temp6[30] ,
         \MC_ARK_ARC_1_3/temp6[29] , \MC_ARK_ARC_1_3/temp6[28] ,
         \MC_ARK_ARC_1_3/temp6[27] , \MC_ARK_ARC_1_3/temp6[26] ,
         \MC_ARK_ARC_1_3/temp6[25] , \MC_ARK_ARC_1_3/temp6[24] ,
         \MC_ARK_ARC_1_3/temp6[23] , \MC_ARK_ARC_1_3/temp6[22] ,
         \MC_ARK_ARC_1_3/temp6[21] , \MC_ARK_ARC_1_3/temp6[20] ,
         \MC_ARK_ARC_1_3/temp6[19] , \MC_ARK_ARC_1_3/temp6[18] ,
         \MC_ARK_ARC_1_3/temp6[17] , \MC_ARK_ARC_1_3/temp6[16] ,
         \MC_ARK_ARC_1_3/temp6[15] , \MC_ARK_ARC_1_3/temp6[14] ,
         \MC_ARK_ARC_1_3/temp6[13] , \MC_ARK_ARC_1_3/temp6[12] ,
         \MC_ARK_ARC_1_3/temp6[11] , \MC_ARK_ARC_1_3/temp6[10] ,
         \MC_ARK_ARC_1_3/temp6[9] , \MC_ARK_ARC_1_3/temp6[8] ,
         \MC_ARK_ARC_1_3/temp6[7] , \MC_ARK_ARC_1_3/temp6[6] ,
         \MC_ARK_ARC_1_3/temp6[4] , \MC_ARK_ARC_1_3/temp6[3] ,
         \MC_ARK_ARC_1_3/temp6[2] , \MC_ARK_ARC_1_3/temp6[1] ,
         \MC_ARK_ARC_1_3/temp6[0] , \MC_ARK_ARC_1_3/temp5[191] ,
         \MC_ARK_ARC_1_3/temp5[190] , \MC_ARK_ARC_1_3/temp5[189] ,
         \MC_ARK_ARC_1_3/temp5[188] , \MC_ARK_ARC_1_3/temp5[187] ,
         \MC_ARK_ARC_1_3/temp5[186] , \MC_ARK_ARC_1_3/temp5[185] ,
         \MC_ARK_ARC_1_3/temp5[184] , \MC_ARK_ARC_1_3/temp5[183] ,
         \MC_ARK_ARC_1_3/temp5[181] , \MC_ARK_ARC_1_3/temp5[180] ,
         \MC_ARK_ARC_1_3/temp5[179] , \MC_ARK_ARC_1_3/temp5[177] ,
         \MC_ARK_ARC_1_3/temp5[176] , \MC_ARK_ARC_1_3/temp5[175] ,
         \MC_ARK_ARC_1_3/temp5[174] , \MC_ARK_ARC_1_3/temp5[173] ,
         \MC_ARK_ARC_1_3/temp5[172] , \MC_ARK_ARC_1_3/temp5[171] ,
         \MC_ARK_ARC_1_3/temp5[170] , \MC_ARK_ARC_1_3/temp5[169] ,
         \MC_ARK_ARC_1_3/temp5[168] , \MC_ARK_ARC_1_3/temp5[166] ,
         \MC_ARK_ARC_1_3/temp5[165] , \MC_ARK_ARC_1_3/temp5[164] ,
         \MC_ARK_ARC_1_3/temp5[163] , \MC_ARK_ARC_1_3/temp5[162] ,
         \MC_ARK_ARC_1_3/temp5[161] , \MC_ARK_ARC_1_3/temp5[160] ,
         \MC_ARK_ARC_1_3/temp5[159] , \MC_ARK_ARC_1_3/temp5[158] ,
         \MC_ARK_ARC_1_3/temp5[157] , \MC_ARK_ARC_1_3/temp5[156] ,
         \MC_ARK_ARC_1_3/temp5[155] , \MC_ARK_ARC_1_3/temp5[154] ,
         \MC_ARK_ARC_1_3/temp5[153] , \MC_ARK_ARC_1_3/temp5[152] ,
         \MC_ARK_ARC_1_3/temp5[151] , \MC_ARK_ARC_1_3/temp5[150] ,
         \MC_ARK_ARC_1_3/temp5[149] , \MC_ARK_ARC_1_3/temp5[148] ,
         \MC_ARK_ARC_1_3/temp5[147] , \MC_ARK_ARC_1_3/temp5[145] ,
         \MC_ARK_ARC_1_3/temp5[144] , \MC_ARK_ARC_1_3/temp5[143] ,
         \MC_ARK_ARC_1_3/temp5[142] , \MC_ARK_ARC_1_3/temp5[141] ,
         \MC_ARK_ARC_1_3/temp5[140] , \MC_ARK_ARC_1_3/temp5[139] ,
         \MC_ARK_ARC_1_3/temp5[138] , \MC_ARK_ARC_1_3/temp5[137] ,
         \MC_ARK_ARC_1_3/temp5[136] , \MC_ARK_ARC_1_3/temp5[135] ,
         \MC_ARK_ARC_1_3/temp5[134] , \MC_ARK_ARC_1_3/temp5[133] ,
         \MC_ARK_ARC_1_3/temp5[132] , \MC_ARK_ARC_1_3/temp5[129] ,
         \MC_ARK_ARC_1_3/temp5[128] , \MC_ARK_ARC_1_3/temp5[127] ,
         \MC_ARK_ARC_1_3/temp5[126] , \MC_ARK_ARC_1_3/temp5[125] ,
         \MC_ARK_ARC_1_3/temp5[124] , \MC_ARK_ARC_1_3/temp5[122] ,
         \MC_ARK_ARC_1_3/temp5[120] , \MC_ARK_ARC_1_3/temp5[119] ,
         \MC_ARK_ARC_1_3/temp5[118] , \MC_ARK_ARC_1_3/temp5[117] ,
         \MC_ARK_ARC_1_3/temp5[116] , \MC_ARK_ARC_1_3/temp5[115] ,
         \MC_ARK_ARC_1_3/temp5[114] , \MC_ARK_ARC_1_3/temp5[113] ,
         \MC_ARK_ARC_1_3/temp5[112] , \MC_ARK_ARC_1_3/temp5[111] ,
         \MC_ARK_ARC_1_3/temp5[110] , \MC_ARK_ARC_1_3/temp5[109] ,
         \MC_ARK_ARC_1_3/temp5[108] , \MC_ARK_ARC_1_3/temp5[107] ,
         \MC_ARK_ARC_1_3/temp5[106] , \MC_ARK_ARC_1_3/temp5[105] ,
         \MC_ARK_ARC_1_3/temp5[104] , \MC_ARK_ARC_1_3/temp5[103] ,
         \MC_ARK_ARC_1_3/temp5[102] , \MC_ARK_ARC_1_3/temp5[101] ,
         \MC_ARK_ARC_1_3/temp5[100] , \MC_ARK_ARC_1_3/temp5[99] ,
         \MC_ARK_ARC_1_3/temp5[98] , \MC_ARK_ARC_1_3/temp5[97] ,
         \MC_ARK_ARC_1_3/temp5[96] , \MC_ARK_ARC_1_3/temp5[95] ,
         \MC_ARK_ARC_1_3/temp5[93] , \MC_ARK_ARC_1_3/temp5[92] ,
         \MC_ARK_ARC_1_3/temp5[91] , \MC_ARK_ARC_1_3/temp5[90] ,
         \MC_ARK_ARC_1_3/temp5[89] , \MC_ARK_ARC_1_3/temp5[88] ,
         \MC_ARK_ARC_1_3/temp5[87] , \MC_ARK_ARC_1_3/temp5[85] ,
         \MC_ARK_ARC_1_3/temp5[84] , \MC_ARK_ARC_1_3/temp5[81] ,
         \MC_ARK_ARC_1_3/temp5[80] , \MC_ARK_ARC_1_3/temp5[78] ,
         \MC_ARK_ARC_1_3/temp5[76] , \MC_ARK_ARC_1_3/temp5[75] ,
         \MC_ARK_ARC_1_3/temp5[74] , \MC_ARK_ARC_1_3/temp5[73] ,
         \MC_ARK_ARC_1_3/temp5[71] , \MC_ARK_ARC_1_3/temp5[70] ,
         \MC_ARK_ARC_1_3/temp5[69] , \MC_ARK_ARC_1_3/temp5[68] ,
         \MC_ARK_ARC_1_3/temp5[67] , \MC_ARK_ARC_1_3/temp5[66] ,
         \MC_ARK_ARC_1_3/temp5[65] , \MC_ARK_ARC_1_3/temp5[63] ,
         \MC_ARK_ARC_1_3/temp5[62] , \MC_ARK_ARC_1_3/temp5[61] ,
         \MC_ARK_ARC_1_3/temp5[60] , \MC_ARK_ARC_1_3/temp5[58] ,
         \MC_ARK_ARC_1_3/temp5[57] , \MC_ARK_ARC_1_3/temp5[56] ,
         \MC_ARK_ARC_1_3/temp5[55] , \MC_ARK_ARC_1_3/temp5[54] ,
         \MC_ARK_ARC_1_3/temp5[53] , \MC_ARK_ARC_1_3/temp5[52] ,
         \MC_ARK_ARC_1_3/temp5[51] , \MC_ARK_ARC_1_3/temp5[50] ,
         \MC_ARK_ARC_1_3/temp5[49] , \MC_ARK_ARC_1_3/temp5[48] ,
         \MC_ARK_ARC_1_3/temp5[47] , \MC_ARK_ARC_1_3/temp5[46] ,
         \MC_ARK_ARC_1_3/temp5[45] , \MC_ARK_ARC_1_3/temp5[44] ,
         \MC_ARK_ARC_1_3/temp5[42] , \MC_ARK_ARC_1_3/temp5[41] ,
         \MC_ARK_ARC_1_3/temp5[40] , \MC_ARK_ARC_1_3/temp5[39] ,
         \MC_ARK_ARC_1_3/temp5[38] , \MC_ARK_ARC_1_3/temp5[36] ,
         \MC_ARK_ARC_1_3/temp5[34] , \MC_ARK_ARC_1_3/temp5[33] ,
         \MC_ARK_ARC_1_3/temp5[32] , \MC_ARK_ARC_1_3/temp5[31] ,
         \MC_ARK_ARC_1_3/temp5[30] , \MC_ARK_ARC_1_3/temp5[29] ,
         \MC_ARK_ARC_1_3/temp5[28] , \MC_ARK_ARC_1_3/temp5[27] ,
         \MC_ARK_ARC_1_3/temp5[25] , \MC_ARK_ARC_1_3/temp5[24] ,
         \MC_ARK_ARC_1_3/temp5[23] , \MC_ARK_ARC_1_3/temp5[22] ,
         \MC_ARK_ARC_1_3/temp5[21] , \MC_ARK_ARC_1_3/temp5[20] ,
         \MC_ARK_ARC_1_3/temp5[19] , \MC_ARK_ARC_1_3/temp5[18] ,
         \MC_ARK_ARC_1_3/temp5[17] , \MC_ARK_ARC_1_3/temp5[16] ,
         \MC_ARK_ARC_1_3/temp5[15] , \MC_ARK_ARC_1_3/temp5[14] ,
         \MC_ARK_ARC_1_3/temp5[13] , \MC_ARK_ARC_1_3/temp5[12] ,
         \MC_ARK_ARC_1_3/temp5[11] , \MC_ARK_ARC_1_3/temp5[10] ,
         \MC_ARK_ARC_1_3/temp5[9] , \MC_ARK_ARC_1_3/temp5[8] ,
         \MC_ARK_ARC_1_3/temp5[7] , \MC_ARK_ARC_1_3/temp5[6] ,
         \MC_ARK_ARC_1_3/temp5[4] , \MC_ARK_ARC_1_3/temp5[3] ,
         \MC_ARK_ARC_1_3/temp5[2] , \MC_ARK_ARC_1_3/temp5[1] ,
         \MC_ARK_ARC_1_3/temp5[0] , \MC_ARK_ARC_1_3/temp4[191] ,
         \MC_ARK_ARC_1_3/temp4[190] , \MC_ARK_ARC_1_3/temp4[189] ,
         \MC_ARK_ARC_1_3/temp4[188] , \MC_ARK_ARC_1_3/temp4[187] ,
         \MC_ARK_ARC_1_3/temp4[186] , \MC_ARK_ARC_1_3/temp4[185] ,
         \MC_ARK_ARC_1_3/temp4[184] , \MC_ARK_ARC_1_3/temp4[183] ,
         \MC_ARK_ARC_1_3/temp4[182] , \MC_ARK_ARC_1_3/temp4[181] ,
         \MC_ARK_ARC_1_3/temp4[180] , \MC_ARK_ARC_1_3/temp4[179] ,
         \MC_ARK_ARC_1_3/temp4[178] , \MC_ARK_ARC_1_3/temp4[177] ,
         \MC_ARK_ARC_1_3/temp4[176] , \MC_ARK_ARC_1_3/temp4[175] ,
         \MC_ARK_ARC_1_3/temp4[174] , \MC_ARK_ARC_1_3/temp4[173] ,
         \MC_ARK_ARC_1_3/temp4[172] , \MC_ARK_ARC_1_3/temp4[171] ,
         \MC_ARK_ARC_1_3/temp4[170] , \MC_ARK_ARC_1_3/temp4[169] ,
         \MC_ARK_ARC_1_3/temp4[168] , \MC_ARK_ARC_1_3/temp4[167] ,
         \MC_ARK_ARC_1_3/temp4[166] , \MC_ARK_ARC_1_3/temp4[165] ,
         \MC_ARK_ARC_1_3/temp4[164] , \MC_ARK_ARC_1_3/temp4[163] ,
         \MC_ARK_ARC_1_3/temp4[162] , \MC_ARK_ARC_1_3/temp4[161] ,
         \MC_ARK_ARC_1_3/temp4[160] , \MC_ARK_ARC_1_3/temp4[159] ,
         \MC_ARK_ARC_1_3/temp4[158] , \MC_ARK_ARC_1_3/temp4[157] ,
         \MC_ARK_ARC_1_3/temp4[156] , \MC_ARK_ARC_1_3/temp4[155] ,
         \MC_ARK_ARC_1_3/temp4[154] , \MC_ARK_ARC_1_3/temp4[153] ,
         \MC_ARK_ARC_1_3/temp4[152] , \MC_ARK_ARC_1_3/temp4[151] ,
         \MC_ARK_ARC_1_3/temp4[150] , \MC_ARK_ARC_1_3/temp4[149] ,
         \MC_ARK_ARC_1_3/temp4[148] , \MC_ARK_ARC_1_3/temp4[147] ,
         \MC_ARK_ARC_1_3/temp4[146] , \MC_ARK_ARC_1_3/temp4[145] ,
         \MC_ARK_ARC_1_3/temp4[144] , \MC_ARK_ARC_1_3/temp4[143] ,
         \MC_ARK_ARC_1_3/temp4[142] , \MC_ARK_ARC_1_3/temp4[141] ,
         \MC_ARK_ARC_1_3/temp4[140] , \MC_ARK_ARC_1_3/temp4[139] ,
         \MC_ARK_ARC_1_3/temp4[138] , \MC_ARK_ARC_1_3/temp4[137] ,
         \MC_ARK_ARC_1_3/temp4[136] , \MC_ARK_ARC_1_3/temp4[135] ,
         \MC_ARK_ARC_1_3/temp4[134] , \MC_ARK_ARC_1_3/temp4[133] ,
         \MC_ARK_ARC_1_3/temp4[132] , \MC_ARK_ARC_1_3/temp4[131] ,
         \MC_ARK_ARC_1_3/temp4[130] , \MC_ARK_ARC_1_3/temp4[129] ,
         \MC_ARK_ARC_1_3/temp4[128] , \MC_ARK_ARC_1_3/temp4[127] ,
         \MC_ARK_ARC_1_3/temp4[126] , \MC_ARK_ARC_1_3/temp4[125] ,
         \MC_ARK_ARC_1_3/temp4[124] , \MC_ARK_ARC_1_3/temp4[123] ,
         \MC_ARK_ARC_1_3/temp4[122] , \MC_ARK_ARC_1_3/temp4[121] ,
         \MC_ARK_ARC_1_3/temp4[120] , \MC_ARK_ARC_1_3/temp4[119] ,
         \MC_ARK_ARC_1_3/temp4[118] , \MC_ARK_ARC_1_3/temp4[117] ,
         \MC_ARK_ARC_1_3/temp4[116] , \MC_ARK_ARC_1_3/temp4[115] ,
         \MC_ARK_ARC_1_3/temp4[114] , \MC_ARK_ARC_1_3/temp4[113] ,
         \MC_ARK_ARC_1_3/temp4[112] , \MC_ARK_ARC_1_3/temp4[111] ,
         \MC_ARK_ARC_1_3/temp4[110] , \MC_ARK_ARC_1_3/temp4[109] ,
         \MC_ARK_ARC_1_3/temp4[108] , \MC_ARK_ARC_1_3/temp4[107] ,
         \MC_ARK_ARC_1_3/temp4[106] , \MC_ARK_ARC_1_3/temp4[105] ,
         \MC_ARK_ARC_1_3/temp4[104] , \MC_ARK_ARC_1_3/temp4[103] ,
         \MC_ARK_ARC_1_3/temp4[102] , \MC_ARK_ARC_1_3/temp4[101] ,
         \MC_ARK_ARC_1_3/temp4[100] , \MC_ARK_ARC_1_3/temp4[99] ,
         \MC_ARK_ARC_1_3/temp4[98] , \MC_ARK_ARC_1_3/temp4[97] ,
         \MC_ARK_ARC_1_3/temp4[96] , \MC_ARK_ARC_1_3/temp4[95] ,
         \MC_ARK_ARC_1_3/temp4[94] , \MC_ARK_ARC_1_3/temp4[93] ,
         \MC_ARK_ARC_1_3/temp4[92] , \MC_ARK_ARC_1_3/temp4[91] ,
         \MC_ARK_ARC_1_3/temp4[90] , \MC_ARK_ARC_1_3/temp4[89] ,
         \MC_ARK_ARC_1_3/temp4[88] , \MC_ARK_ARC_1_3/temp4[87] ,
         \MC_ARK_ARC_1_3/temp4[86] , \MC_ARK_ARC_1_3/temp4[85] ,
         \MC_ARK_ARC_1_3/temp4[84] , \MC_ARK_ARC_1_3/temp4[83] ,
         \MC_ARK_ARC_1_3/temp4[82] , \MC_ARK_ARC_1_3/temp4[81] ,
         \MC_ARK_ARC_1_3/temp4[80] , \MC_ARK_ARC_1_3/temp4[79] ,
         \MC_ARK_ARC_1_3/temp4[78] , \MC_ARK_ARC_1_3/temp4[77] ,
         \MC_ARK_ARC_1_3/temp4[76] , \MC_ARK_ARC_1_3/temp4[75] ,
         \MC_ARK_ARC_1_3/temp4[74] , \MC_ARK_ARC_1_3/temp4[73] ,
         \MC_ARK_ARC_1_3/temp4[72] , \MC_ARK_ARC_1_3/temp4[71] ,
         \MC_ARK_ARC_1_3/temp4[70] , \MC_ARK_ARC_1_3/temp4[69] ,
         \MC_ARK_ARC_1_3/temp4[68] , \MC_ARK_ARC_1_3/temp4[67] ,
         \MC_ARK_ARC_1_3/temp4[66] , \MC_ARK_ARC_1_3/temp4[65] ,
         \MC_ARK_ARC_1_3/temp4[64] , \MC_ARK_ARC_1_3/temp4[63] ,
         \MC_ARK_ARC_1_3/temp4[62] , \MC_ARK_ARC_1_3/temp4[61] ,
         \MC_ARK_ARC_1_3/temp4[60] , \MC_ARK_ARC_1_3/temp4[59] ,
         \MC_ARK_ARC_1_3/temp4[58] , \MC_ARK_ARC_1_3/temp4[57] ,
         \MC_ARK_ARC_1_3/temp4[56] , \MC_ARK_ARC_1_3/temp4[55] ,
         \MC_ARK_ARC_1_3/temp4[54] , \MC_ARK_ARC_1_3/temp4[53] ,
         \MC_ARK_ARC_1_3/temp4[52] , \MC_ARK_ARC_1_3/temp4[51] ,
         \MC_ARK_ARC_1_3/temp4[50] , \MC_ARK_ARC_1_3/temp4[49] ,
         \MC_ARK_ARC_1_3/temp4[48] , \MC_ARK_ARC_1_3/temp4[47] ,
         \MC_ARK_ARC_1_3/temp4[46] , \MC_ARK_ARC_1_3/temp4[45] ,
         \MC_ARK_ARC_1_3/temp4[44] , \MC_ARK_ARC_1_3/temp4[43] ,
         \MC_ARK_ARC_1_3/temp4[42] , \MC_ARK_ARC_1_3/temp4[41] ,
         \MC_ARK_ARC_1_3/temp4[40] , \MC_ARK_ARC_1_3/temp4[39] ,
         \MC_ARK_ARC_1_3/temp4[38] , \MC_ARK_ARC_1_3/temp4[37] ,
         \MC_ARK_ARC_1_3/temp4[36] , \MC_ARK_ARC_1_3/temp4[35] ,
         \MC_ARK_ARC_1_3/temp4[34] , \MC_ARK_ARC_1_3/temp4[33] ,
         \MC_ARK_ARC_1_3/temp4[32] , \MC_ARK_ARC_1_3/temp4[31] ,
         \MC_ARK_ARC_1_3/temp4[30] , \MC_ARK_ARC_1_3/temp4[29] ,
         \MC_ARK_ARC_1_3/temp4[28] , \MC_ARK_ARC_1_3/temp4[27] ,
         \MC_ARK_ARC_1_3/temp4[26] , \MC_ARK_ARC_1_3/temp4[25] ,
         \MC_ARK_ARC_1_3/temp4[24] , \MC_ARK_ARC_1_3/temp4[23] ,
         \MC_ARK_ARC_1_3/temp4[22] , \MC_ARK_ARC_1_3/temp4[21] ,
         \MC_ARK_ARC_1_3/temp4[20] , \MC_ARK_ARC_1_3/temp4[19] ,
         \MC_ARK_ARC_1_3/temp4[18] , \MC_ARK_ARC_1_3/temp4[17] ,
         \MC_ARK_ARC_1_3/temp4[16] , \MC_ARK_ARC_1_3/temp4[15] ,
         \MC_ARK_ARC_1_3/temp4[14] , \MC_ARK_ARC_1_3/temp4[13] ,
         \MC_ARK_ARC_1_3/temp4[12] , \MC_ARK_ARC_1_3/temp4[11] ,
         \MC_ARK_ARC_1_3/temp4[10] , \MC_ARK_ARC_1_3/temp4[9] ,
         \MC_ARK_ARC_1_3/temp4[8] , \MC_ARK_ARC_1_3/temp4[7] ,
         \MC_ARK_ARC_1_3/temp4[6] , \MC_ARK_ARC_1_3/temp4[5] ,
         \MC_ARK_ARC_1_3/temp4[4] , \MC_ARK_ARC_1_3/temp4[3] ,
         \MC_ARK_ARC_1_3/temp4[2] , \MC_ARK_ARC_1_3/temp4[1] ,
         \MC_ARK_ARC_1_3/temp4[0] , \MC_ARK_ARC_1_3/temp3[191] ,
         \MC_ARK_ARC_1_3/temp3[190] , \MC_ARK_ARC_1_3/temp3[189] ,
         \MC_ARK_ARC_1_3/temp3[188] , \MC_ARK_ARC_1_3/temp3[187] ,
         \MC_ARK_ARC_1_3/temp3[186] , \MC_ARK_ARC_1_3/temp3[185] ,
         \MC_ARK_ARC_1_3/temp3[184] , \MC_ARK_ARC_1_3/temp3[183] ,
         \MC_ARK_ARC_1_3/temp3[182] , \MC_ARK_ARC_1_3/temp3[181] ,
         \MC_ARK_ARC_1_3/temp3[180] , \MC_ARK_ARC_1_3/temp3[179] ,
         \MC_ARK_ARC_1_3/temp3[178] , \MC_ARK_ARC_1_3/temp3[177] ,
         \MC_ARK_ARC_1_3/temp3[176] , \MC_ARK_ARC_1_3/temp3[175] ,
         \MC_ARK_ARC_1_3/temp3[174] , \MC_ARK_ARC_1_3/temp3[173] ,
         \MC_ARK_ARC_1_3/temp3[172] , \MC_ARK_ARC_1_3/temp3[171] ,
         \MC_ARK_ARC_1_3/temp3[170] , \MC_ARK_ARC_1_3/temp3[169] ,
         \MC_ARK_ARC_1_3/temp3[168] , \MC_ARK_ARC_1_3/temp3[167] ,
         \MC_ARK_ARC_1_3/temp3[166] , \MC_ARK_ARC_1_3/temp3[165] ,
         \MC_ARK_ARC_1_3/temp3[164] , \MC_ARK_ARC_1_3/temp3[163] ,
         \MC_ARK_ARC_1_3/temp3[162] , \MC_ARK_ARC_1_3/temp3[161] ,
         \MC_ARK_ARC_1_3/temp3[160] , \MC_ARK_ARC_1_3/temp3[159] ,
         \MC_ARK_ARC_1_3/temp3[158] , \MC_ARK_ARC_1_3/temp3[157] ,
         \MC_ARK_ARC_1_3/temp3[156] , \MC_ARK_ARC_1_3/temp3[155] ,
         \MC_ARK_ARC_1_3/temp3[154] , \MC_ARK_ARC_1_3/temp3[153] ,
         \MC_ARK_ARC_1_3/temp3[152] , \MC_ARK_ARC_1_3/temp3[151] ,
         \MC_ARK_ARC_1_3/temp3[150] , \MC_ARK_ARC_1_3/temp3[149] ,
         \MC_ARK_ARC_1_3/temp3[148] , \MC_ARK_ARC_1_3/temp3[147] ,
         \MC_ARK_ARC_1_3/temp3[146] , \MC_ARK_ARC_1_3/temp3[145] ,
         \MC_ARK_ARC_1_3/temp3[144] , \MC_ARK_ARC_1_3/temp3[143] ,
         \MC_ARK_ARC_1_3/temp3[142] , \MC_ARK_ARC_1_3/temp3[141] ,
         \MC_ARK_ARC_1_3/temp3[140] , \MC_ARK_ARC_1_3/temp3[139] ,
         \MC_ARK_ARC_1_3/temp3[138] , \MC_ARK_ARC_1_3/temp3[137] ,
         \MC_ARK_ARC_1_3/temp3[136] , \MC_ARK_ARC_1_3/temp3[135] ,
         \MC_ARK_ARC_1_3/temp3[134] , \MC_ARK_ARC_1_3/temp3[133] ,
         \MC_ARK_ARC_1_3/temp3[132] , \MC_ARK_ARC_1_3/temp3[131] ,
         \MC_ARK_ARC_1_3/temp3[130] , \MC_ARK_ARC_1_3/temp3[129] ,
         \MC_ARK_ARC_1_3/temp3[128] , \MC_ARK_ARC_1_3/temp3[127] ,
         \MC_ARK_ARC_1_3/temp3[126] , \MC_ARK_ARC_1_3/temp3[125] ,
         \MC_ARK_ARC_1_3/temp3[124] , \MC_ARK_ARC_1_3/temp3[123] ,
         \MC_ARK_ARC_1_3/temp3[122] , \MC_ARK_ARC_1_3/temp3[121] ,
         \MC_ARK_ARC_1_3/temp3[120] , \MC_ARK_ARC_1_3/temp3[119] ,
         \MC_ARK_ARC_1_3/temp3[118] , \MC_ARK_ARC_1_3/temp3[117] ,
         \MC_ARK_ARC_1_3/temp3[116] , \MC_ARK_ARC_1_3/temp3[115] ,
         \MC_ARK_ARC_1_3/temp3[114] , \MC_ARK_ARC_1_3/temp3[113] ,
         \MC_ARK_ARC_1_3/temp3[112] , \MC_ARK_ARC_1_3/temp3[111] ,
         \MC_ARK_ARC_1_3/temp3[110] , \MC_ARK_ARC_1_3/temp3[109] ,
         \MC_ARK_ARC_1_3/temp3[108] , \MC_ARK_ARC_1_3/temp3[107] ,
         \MC_ARK_ARC_1_3/temp3[106] , \MC_ARK_ARC_1_3/temp3[105] ,
         \MC_ARK_ARC_1_3/temp3[104] , \MC_ARK_ARC_1_3/temp3[103] ,
         \MC_ARK_ARC_1_3/temp3[102] , \MC_ARK_ARC_1_3/temp3[101] ,
         \MC_ARK_ARC_1_3/temp3[100] , \MC_ARK_ARC_1_3/temp3[99] ,
         \MC_ARK_ARC_1_3/temp3[98] , \MC_ARK_ARC_1_3/temp3[97] ,
         \MC_ARK_ARC_1_3/temp3[96] , \MC_ARK_ARC_1_3/temp3[95] ,
         \MC_ARK_ARC_1_3/temp3[94] , \MC_ARK_ARC_1_3/temp3[93] ,
         \MC_ARK_ARC_1_3/temp3[92] , \MC_ARK_ARC_1_3/temp3[91] ,
         \MC_ARK_ARC_1_3/temp3[90] , \MC_ARK_ARC_1_3/temp3[89] ,
         \MC_ARK_ARC_1_3/temp3[88] , \MC_ARK_ARC_1_3/temp3[87] ,
         \MC_ARK_ARC_1_3/temp3[86] , \MC_ARK_ARC_1_3/temp3[85] ,
         \MC_ARK_ARC_1_3/temp3[84] , \MC_ARK_ARC_1_3/temp3[83] ,
         \MC_ARK_ARC_1_3/temp3[82] , \MC_ARK_ARC_1_3/temp3[81] ,
         \MC_ARK_ARC_1_3/temp3[80] , \MC_ARK_ARC_1_3/temp3[79] ,
         \MC_ARK_ARC_1_3/temp3[78] , \MC_ARK_ARC_1_3/temp3[77] ,
         \MC_ARK_ARC_1_3/temp3[76] , \MC_ARK_ARC_1_3/temp3[75] ,
         \MC_ARK_ARC_1_3/temp3[74] , \MC_ARK_ARC_1_3/temp3[73] ,
         \MC_ARK_ARC_1_3/temp3[72] , \MC_ARK_ARC_1_3/temp3[71] ,
         \MC_ARK_ARC_1_3/temp3[70] , \MC_ARK_ARC_1_3/temp3[69] ,
         \MC_ARK_ARC_1_3/temp3[68] , \MC_ARK_ARC_1_3/temp3[67] ,
         \MC_ARK_ARC_1_3/temp3[66] , \MC_ARK_ARC_1_3/temp3[65] ,
         \MC_ARK_ARC_1_3/temp3[64] , \MC_ARK_ARC_1_3/temp3[63] ,
         \MC_ARK_ARC_1_3/temp3[62] , \MC_ARK_ARC_1_3/temp3[61] ,
         \MC_ARK_ARC_1_3/temp3[60] , \MC_ARK_ARC_1_3/temp3[59] ,
         \MC_ARK_ARC_1_3/temp3[58] , \MC_ARK_ARC_1_3/temp3[57] ,
         \MC_ARK_ARC_1_3/temp3[56] , \MC_ARK_ARC_1_3/temp3[55] ,
         \MC_ARK_ARC_1_3/temp3[54] , \MC_ARK_ARC_1_3/temp3[53] ,
         \MC_ARK_ARC_1_3/temp3[52] , \MC_ARK_ARC_1_3/temp3[51] ,
         \MC_ARK_ARC_1_3/temp3[50] , \MC_ARK_ARC_1_3/temp3[49] ,
         \MC_ARK_ARC_1_3/temp3[48] , \MC_ARK_ARC_1_3/temp3[47] ,
         \MC_ARK_ARC_1_3/temp3[46] , \MC_ARK_ARC_1_3/temp3[45] ,
         \MC_ARK_ARC_1_3/temp3[44] , \MC_ARK_ARC_1_3/temp3[43] ,
         \MC_ARK_ARC_1_3/temp3[42] , \MC_ARK_ARC_1_3/temp3[41] ,
         \MC_ARK_ARC_1_3/temp3[40] , \MC_ARK_ARC_1_3/temp3[39] ,
         \MC_ARK_ARC_1_3/temp3[38] , \MC_ARK_ARC_1_3/temp3[37] ,
         \MC_ARK_ARC_1_3/temp3[36] , \MC_ARK_ARC_1_3/temp3[35] ,
         \MC_ARK_ARC_1_3/temp3[34] , \MC_ARK_ARC_1_3/temp3[33] ,
         \MC_ARK_ARC_1_3/temp3[32] , \MC_ARK_ARC_1_3/temp3[31] ,
         \MC_ARK_ARC_1_3/temp3[30] , \MC_ARK_ARC_1_3/temp3[29] ,
         \MC_ARK_ARC_1_3/temp3[28] , \MC_ARK_ARC_1_3/temp3[27] ,
         \MC_ARK_ARC_1_3/temp3[26] , \MC_ARK_ARC_1_3/temp3[25] ,
         \MC_ARK_ARC_1_3/temp3[24] , \MC_ARK_ARC_1_3/temp3[23] ,
         \MC_ARK_ARC_1_3/temp3[22] , \MC_ARK_ARC_1_3/temp3[21] ,
         \MC_ARK_ARC_1_3/temp3[20] , \MC_ARK_ARC_1_3/temp3[19] ,
         \MC_ARK_ARC_1_3/temp3[18] , \MC_ARK_ARC_1_3/temp3[17] ,
         \MC_ARK_ARC_1_3/temp3[16] , \MC_ARK_ARC_1_3/temp3[15] ,
         \MC_ARK_ARC_1_3/temp3[14] , \MC_ARK_ARC_1_3/temp3[13] ,
         \MC_ARK_ARC_1_3/temp3[12] , \MC_ARK_ARC_1_3/temp3[11] ,
         \MC_ARK_ARC_1_3/temp3[10] , \MC_ARK_ARC_1_3/temp3[9] ,
         \MC_ARK_ARC_1_3/temp3[8] , \MC_ARK_ARC_1_3/temp3[7] ,
         \MC_ARK_ARC_1_3/temp3[6] , \MC_ARK_ARC_1_3/temp3[5] ,
         \MC_ARK_ARC_1_3/temp3[4] , \MC_ARK_ARC_1_3/temp3[3] ,
         \MC_ARK_ARC_1_3/temp3[2] , \MC_ARK_ARC_1_3/temp3[1] ,
         \MC_ARK_ARC_1_3/temp3[0] , \MC_ARK_ARC_1_3/temp2[191] ,
         \MC_ARK_ARC_1_3/temp2[190] , \MC_ARK_ARC_1_3/temp2[189] ,
         \MC_ARK_ARC_1_3/temp2[188] , \MC_ARK_ARC_1_3/temp2[187] ,
         \MC_ARK_ARC_1_3/temp2[186] , \MC_ARK_ARC_1_3/temp2[185] ,
         \MC_ARK_ARC_1_3/temp2[184] , \MC_ARK_ARC_1_3/temp2[183] ,
         \MC_ARK_ARC_1_3/temp2[182] , \MC_ARK_ARC_1_3/temp2[181] ,
         \MC_ARK_ARC_1_3/temp2[180] , \MC_ARK_ARC_1_3/temp2[179] ,
         \MC_ARK_ARC_1_3/temp2[178] , \MC_ARK_ARC_1_3/temp2[177] ,
         \MC_ARK_ARC_1_3/temp2[176] , \MC_ARK_ARC_1_3/temp2[175] ,
         \MC_ARK_ARC_1_3/temp2[174] , \MC_ARK_ARC_1_3/temp2[173] ,
         \MC_ARK_ARC_1_3/temp2[172] , \MC_ARK_ARC_1_3/temp2[171] ,
         \MC_ARK_ARC_1_3/temp2[170] , \MC_ARK_ARC_1_3/temp2[169] ,
         \MC_ARK_ARC_1_3/temp2[168] , \MC_ARK_ARC_1_3/temp2[167] ,
         \MC_ARK_ARC_1_3/temp2[166] , \MC_ARK_ARC_1_3/temp2[165] ,
         \MC_ARK_ARC_1_3/temp2[164] , \MC_ARK_ARC_1_3/temp2[163] ,
         \MC_ARK_ARC_1_3/temp2[162] , \MC_ARK_ARC_1_3/temp2[161] ,
         \MC_ARK_ARC_1_3/temp2[160] , \MC_ARK_ARC_1_3/temp2[159] ,
         \MC_ARK_ARC_1_3/temp2[158] , \MC_ARK_ARC_1_3/temp2[157] ,
         \MC_ARK_ARC_1_3/temp2[156] , \MC_ARK_ARC_1_3/temp2[155] ,
         \MC_ARK_ARC_1_3/temp2[154] , \MC_ARK_ARC_1_3/temp2[153] ,
         \MC_ARK_ARC_1_3/temp2[152] , \MC_ARK_ARC_1_3/temp2[151] ,
         \MC_ARK_ARC_1_3/temp2[150] , \MC_ARK_ARC_1_3/temp2[149] ,
         \MC_ARK_ARC_1_3/temp2[148] , \MC_ARK_ARC_1_3/temp2[147] ,
         \MC_ARK_ARC_1_3/temp2[146] , \MC_ARK_ARC_1_3/temp2[145] ,
         \MC_ARK_ARC_1_3/temp2[144] , \MC_ARK_ARC_1_3/temp2[143] ,
         \MC_ARK_ARC_1_3/temp2[142] , \MC_ARK_ARC_1_3/temp2[141] ,
         \MC_ARK_ARC_1_3/temp2[140] , \MC_ARK_ARC_1_3/temp2[139] ,
         \MC_ARK_ARC_1_3/temp2[138] , \MC_ARK_ARC_1_3/temp2[137] ,
         \MC_ARK_ARC_1_3/temp2[136] , \MC_ARK_ARC_1_3/temp2[135] ,
         \MC_ARK_ARC_1_3/temp2[134] , \MC_ARK_ARC_1_3/temp2[133] ,
         \MC_ARK_ARC_1_3/temp2[132] , \MC_ARK_ARC_1_3/temp2[131] ,
         \MC_ARK_ARC_1_3/temp2[130] , \MC_ARK_ARC_1_3/temp2[129] ,
         \MC_ARK_ARC_1_3/temp2[128] , \MC_ARK_ARC_1_3/temp2[127] ,
         \MC_ARK_ARC_1_3/temp2[126] , \MC_ARK_ARC_1_3/temp2[125] ,
         \MC_ARK_ARC_1_3/temp2[124] , \MC_ARK_ARC_1_3/temp2[123] ,
         \MC_ARK_ARC_1_3/temp2[122] , \MC_ARK_ARC_1_3/temp2[121] ,
         \MC_ARK_ARC_1_3/temp2[120] , \MC_ARK_ARC_1_3/temp2[119] ,
         \MC_ARK_ARC_1_3/temp2[118] , \MC_ARK_ARC_1_3/temp2[117] ,
         \MC_ARK_ARC_1_3/temp2[116] , \MC_ARK_ARC_1_3/temp2[115] ,
         \MC_ARK_ARC_1_3/temp2[114] , \MC_ARK_ARC_1_3/temp2[113] ,
         \MC_ARK_ARC_1_3/temp2[112] , \MC_ARK_ARC_1_3/temp2[111] ,
         \MC_ARK_ARC_1_3/temp2[110] , \MC_ARK_ARC_1_3/temp2[109] ,
         \MC_ARK_ARC_1_3/temp2[108] , \MC_ARK_ARC_1_3/temp2[107] ,
         \MC_ARK_ARC_1_3/temp2[106] , \MC_ARK_ARC_1_3/temp2[105] ,
         \MC_ARK_ARC_1_3/temp2[104] , \MC_ARK_ARC_1_3/temp2[103] ,
         \MC_ARK_ARC_1_3/temp2[102] , \MC_ARK_ARC_1_3/temp2[101] ,
         \MC_ARK_ARC_1_3/temp2[100] , \MC_ARK_ARC_1_3/temp2[99] ,
         \MC_ARK_ARC_1_3/temp2[98] , \MC_ARK_ARC_1_3/temp2[97] ,
         \MC_ARK_ARC_1_3/temp2[96] , \MC_ARK_ARC_1_3/temp2[95] ,
         \MC_ARK_ARC_1_3/temp2[94] , \MC_ARK_ARC_1_3/temp2[93] ,
         \MC_ARK_ARC_1_3/temp2[92] , \MC_ARK_ARC_1_3/temp2[91] ,
         \MC_ARK_ARC_1_3/temp2[90] , \MC_ARK_ARC_1_3/temp2[89] ,
         \MC_ARK_ARC_1_3/temp2[88] , \MC_ARK_ARC_1_3/temp2[87] ,
         \MC_ARK_ARC_1_3/temp2[86] , \MC_ARK_ARC_1_3/temp2[85] ,
         \MC_ARK_ARC_1_3/temp2[84] , \MC_ARK_ARC_1_3/temp2[83] ,
         \MC_ARK_ARC_1_3/temp2[82] , \MC_ARK_ARC_1_3/temp2[81] ,
         \MC_ARK_ARC_1_3/temp2[80] , \MC_ARK_ARC_1_3/temp2[79] ,
         \MC_ARK_ARC_1_3/temp2[78] , \MC_ARK_ARC_1_3/temp2[77] ,
         \MC_ARK_ARC_1_3/temp2[76] , \MC_ARK_ARC_1_3/temp2[75] ,
         \MC_ARK_ARC_1_3/temp2[74] , \MC_ARK_ARC_1_3/temp2[73] ,
         \MC_ARK_ARC_1_3/temp2[72] , \MC_ARK_ARC_1_3/temp2[71] ,
         \MC_ARK_ARC_1_3/temp2[70] , \MC_ARK_ARC_1_3/temp2[69] ,
         \MC_ARK_ARC_1_3/temp2[68] , \MC_ARK_ARC_1_3/temp2[67] ,
         \MC_ARK_ARC_1_3/temp2[66] , \MC_ARK_ARC_1_3/temp2[65] ,
         \MC_ARK_ARC_1_3/temp2[64] , \MC_ARK_ARC_1_3/temp2[63] ,
         \MC_ARK_ARC_1_3/temp2[62] , \MC_ARK_ARC_1_3/temp2[61] ,
         \MC_ARK_ARC_1_3/temp2[60] , \MC_ARK_ARC_1_3/temp2[59] ,
         \MC_ARK_ARC_1_3/temp2[58] , \MC_ARK_ARC_1_3/temp2[57] ,
         \MC_ARK_ARC_1_3/temp2[56] , \MC_ARK_ARC_1_3/temp2[55] ,
         \MC_ARK_ARC_1_3/temp2[54] , \MC_ARK_ARC_1_3/temp2[53] ,
         \MC_ARK_ARC_1_3/temp2[52] , \MC_ARK_ARC_1_3/temp2[51] ,
         \MC_ARK_ARC_1_3/temp2[50] , \MC_ARK_ARC_1_3/temp2[49] ,
         \MC_ARK_ARC_1_3/temp2[48] , \MC_ARK_ARC_1_3/temp2[47] ,
         \MC_ARK_ARC_1_3/temp2[46] , \MC_ARK_ARC_1_3/temp2[45] ,
         \MC_ARK_ARC_1_3/temp2[44] , \MC_ARK_ARC_1_3/temp2[43] ,
         \MC_ARK_ARC_1_3/temp2[42] , \MC_ARK_ARC_1_3/temp2[41] ,
         \MC_ARK_ARC_1_3/temp2[40] , \MC_ARK_ARC_1_3/temp2[39] ,
         \MC_ARK_ARC_1_3/temp2[38] , \MC_ARK_ARC_1_3/temp2[37] ,
         \MC_ARK_ARC_1_3/temp2[36] , \MC_ARK_ARC_1_3/temp2[35] ,
         \MC_ARK_ARC_1_3/temp2[34] , \MC_ARK_ARC_1_3/temp2[33] ,
         \MC_ARK_ARC_1_3/temp2[32] , \MC_ARK_ARC_1_3/temp2[31] ,
         \MC_ARK_ARC_1_3/temp2[30] , \MC_ARK_ARC_1_3/temp2[29] ,
         \MC_ARK_ARC_1_3/temp2[28] , \MC_ARK_ARC_1_3/temp2[27] ,
         \MC_ARK_ARC_1_3/temp2[26] , \MC_ARK_ARC_1_3/temp2[25] ,
         \MC_ARK_ARC_1_3/temp2[24] , \MC_ARK_ARC_1_3/temp2[23] ,
         \MC_ARK_ARC_1_3/temp2[22] , \MC_ARK_ARC_1_3/temp2[21] ,
         \MC_ARK_ARC_1_3/temp2[20] , \MC_ARK_ARC_1_3/temp2[19] ,
         \MC_ARK_ARC_1_3/temp2[18] , \MC_ARK_ARC_1_3/temp2[17] ,
         \MC_ARK_ARC_1_3/temp2[16] , \MC_ARK_ARC_1_3/temp2[15] ,
         \MC_ARK_ARC_1_3/temp2[14] , \MC_ARK_ARC_1_3/temp2[13] ,
         \MC_ARK_ARC_1_3/temp2[12] , \MC_ARK_ARC_1_3/temp2[11] ,
         \MC_ARK_ARC_1_3/temp2[10] , \MC_ARK_ARC_1_3/temp2[9] ,
         \MC_ARK_ARC_1_3/temp2[8] , \MC_ARK_ARC_1_3/temp2[7] ,
         \MC_ARK_ARC_1_3/temp2[6] , \MC_ARK_ARC_1_3/temp2[5] ,
         \MC_ARK_ARC_1_3/temp2[4] , \MC_ARK_ARC_1_3/temp2[3] ,
         \MC_ARK_ARC_1_3/temp2[2] , \MC_ARK_ARC_1_3/temp2[1] ,
         \MC_ARK_ARC_1_3/temp2[0] , \MC_ARK_ARC_1_3/temp1[191] ,
         \MC_ARK_ARC_1_3/temp1[190] , \MC_ARK_ARC_1_3/temp1[189] ,
         \MC_ARK_ARC_1_3/temp1[188] , \MC_ARK_ARC_1_3/temp1[187] ,
         \MC_ARK_ARC_1_3/temp1[186] , \MC_ARK_ARC_1_3/temp1[185] ,
         \MC_ARK_ARC_1_3/temp1[184] , \MC_ARK_ARC_1_3/temp1[183] ,
         \MC_ARK_ARC_1_3/temp1[182] , \MC_ARK_ARC_1_3/temp1[181] ,
         \MC_ARK_ARC_1_3/temp1[180] , \MC_ARK_ARC_1_3/temp1[179] ,
         \MC_ARK_ARC_1_3/temp1[178] , \MC_ARK_ARC_1_3/temp1[177] ,
         \MC_ARK_ARC_1_3/temp1[176] , \MC_ARK_ARC_1_3/temp1[175] ,
         \MC_ARK_ARC_1_3/temp1[174] , \MC_ARK_ARC_1_3/temp1[173] ,
         \MC_ARK_ARC_1_3/temp1[172] , \MC_ARK_ARC_1_3/temp1[171] ,
         \MC_ARK_ARC_1_3/temp1[170] , \MC_ARK_ARC_1_3/temp1[169] ,
         \MC_ARK_ARC_1_3/temp1[168] , \MC_ARK_ARC_1_3/temp1[167] ,
         \MC_ARK_ARC_1_3/temp1[166] , \MC_ARK_ARC_1_3/temp1[165] ,
         \MC_ARK_ARC_1_3/temp1[164] , \MC_ARK_ARC_1_3/temp1[163] ,
         \MC_ARK_ARC_1_3/temp1[162] , \MC_ARK_ARC_1_3/temp1[161] ,
         \MC_ARK_ARC_1_3/temp1[160] , \MC_ARK_ARC_1_3/temp1[159] ,
         \MC_ARK_ARC_1_3/temp1[158] , \MC_ARK_ARC_1_3/temp1[157] ,
         \MC_ARK_ARC_1_3/temp1[156] , \MC_ARK_ARC_1_3/temp1[155] ,
         \MC_ARK_ARC_1_3/temp1[154] , \MC_ARK_ARC_1_3/temp1[153] ,
         \MC_ARK_ARC_1_3/temp1[152] , \MC_ARK_ARC_1_3/temp1[151] ,
         \MC_ARK_ARC_1_3/temp1[150] , \MC_ARK_ARC_1_3/temp1[149] ,
         \MC_ARK_ARC_1_3/temp1[148] , \MC_ARK_ARC_1_3/temp1[147] ,
         \MC_ARK_ARC_1_3/temp1[146] , \MC_ARK_ARC_1_3/temp1[145] ,
         \MC_ARK_ARC_1_3/temp1[144] , \MC_ARK_ARC_1_3/temp1[143] ,
         \MC_ARK_ARC_1_3/temp1[142] , \MC_ARK_ARC_1_3/temp1[141] ,
         \MC_ARK_ARC_1_3/temp1[140] , \MC_ARK_ARC_1_3/temp1[139] ,
         \MC_ARK_ARC_1_3/temp1[138] , \MC_ARK_ARC_1_3/temp1[137] ,
         \MC_ARK_ARC_1_3/temp1[136] , \MC_ARK_ARC_1_3/temp1[135] ,
         \MC_ARK_ARC_1_3/temp1[134] , \MC_ARK_ARC_1_3/temp1[133] ,
         \MC_ARK_ARC_1_3/temp1[132] , \MC_ARK_ARC_1_3/temp1[131] ,
         \MC_ARK_ARC_1_3/temp1[130] , \MC_ARK_ARC_1_3/temp1[129] ,
         \MC_ARK_ARC_1_3/temp1[128] , \MC_ARK_ARC_1_3/temp1[127] ,
         \MC_ARK_ARC_1_3/temp1[126] , \MC_ARK_ARC_1_3/temp1[125] ,
         \MC_ARK_ARC_1_3/temp1[124] , \MC_ARK_ARC_1_3/temp1[123] ,
         \MC_ARK_ARC_1_3/temp1[122] , \MC_ARK_ARC_1_3/temp1[121] ,
         \MC_ARK_ARC_1_3/temp1[120] , \MC_ARK_ARC_1_3/temp1[119] ,
         \MC_ARK_ARC_1_3/temp1[118] , \MC_ARK_ARC_1_3/temp1[117] ,
         \MC_ARK_ARC_1_3/temp1[116] , \MC_ARK_ARC_1_3/temp1[115] ,
         \MC_ARK_ARC_1_3/temp1[114] , \MC_ARK_ARC_1_3/temp1[113] ,
         \MC_ARK_ARC_1_3/temp1[112] , \MC_ARK_ARC_1_3/temp1[111] ,
         \MC_ARK_ARC_1_3/temp1[110] , \MC_ARK_ARC_1_3/temp1[109] ,
         \MC_ARK_ARC_1_3/temp1[108] , \MC_ARK_ARC_1_3/temp1[107] ,
         \MC_ARK_ARC_1_3/temp1[106] , \MC_ARK_ARC_1_3/temp1[105] ,
         \MC_ARK_ARC_1_3/temp1[104] , \MC_ARK_ARC_1_3/temp1[103] ,
         \MC_ARK_ARC_1_3/temp1[102] , \MC_ARK_ARC_1_3/temp1[101] ,
         \MC_ARK_ARC_1_3/temp1[100] , \MC_ARK_ARC_1_3/temp1[99] ,
         \MC_ARK_ARC_1_3/temp1[98] , \MC_ARK_ARC_1_3/temp1[97] ,
         \MC_ARK_ARC_1_3/temp1[96] , \MC_ARK_ARC_1_3/temp1[95] ,
         \MC_ARK_ARC_1_3/temp1[94] , \MC_ARK_ARC_1_3/temp1[93] ,
         \MC_ARK_ARC_1_3/temp1[92] , \MC_ARK_ARC_1_3/temp1[91] ,
         \MC_ARK_ARC_1_3/temp1[90] , \MC_ARK_ARC_1_3/temp1[89] ,
         \MC_ARK_ARC_1_3/temp1[88] , \MC_ARK_ARC_1_3/temp1[87] ,
         \MC_ARK_ARC_1_3/temp1[86] , \MC_ARK_ARC_1_3/temp1[85] ,
         \MC_ARK_ARC_1_3/temp1[84] , \MC_ARK_ARC_1_3/temp1[83] ,
         \MC_ARK_ARC_1_3/temp1[82] , \MC_ARK_ARC_1_3/temp1[81] ,
         \MC_ARK_ARC_1_3/temp1[80] , \MC_ARK_ARC_1_3/temp1[79] ,
         \MC_ARK_ARC_1_3/temp1[78] , \MC_ARK_ARC_1_3/temp1[77] ,
         \MC_ARK_ARC_1_3/temp1[76] , \MC_ARK_ARC_1_3/temp1[75] ,
         \MC_ARK_ARC_1_3/temp1[74] , \MC_ARK_ARC_1_3/temp1[73] ,
         \MC_ARK_ARC_1_3/temp1[72] , \MC_ARK_ARC_1_3/temp1[71] ,
         \MC_ARK_ARC_1_3/temp1[70] , \MC_ARK_ARC_1_3/temp1[69] ,
         \MC_ARK_ARC_1_3/temp1[68] , \MC_ARK_ARC_1_3/temp1[67] ,
         \MC_ARK_ARC_1_3/temp1[66] , \MC_ARK_ARC_1_3/temp1[65] ,
         \MC_ARK_ARC_1_3/temp1[64] , \MC_ARK_ARC_1_3/temp1[63] ,
         \MC_ARK_ARC_1_3/temp1[62] , \MC_ARK_ARC_1_3/temp1[61] ,
         \MC_ARK_ARC_1_3/temp1[60] , \MC_ARK_ARC_1_3/temp1[59] ,
         \MC_ARK_ARC_1_3/temp1[58] , \MC_ARK_ARC_1_3/temp1[57] ,
         \MC_ARK_ARC_1_3/temp1[56] , \MC_ARK_ARC_1_3/temp1[55] ,
         \MC_ARK_ARC_1_3/temp1[54] , \MC_ARK_ARC_1_3/temp1[53] ,
         \MC_ARK_ARC_1_3/temp1[52] , \MC_ARK_ARC_1_3/temp1[51] ,
         \MC_ARK_ARC_1_3/temp1[50] , \MC_ARK_ARC_1_3/temp1[49] ,
         \MC_ARK_ARC_1_3/temp1[48] , \MC_ARK_ARC_1_3/temp1[47] ,
         \MC_ARK_ARC_1_3/temp1[46] , \MC_ARK_ARC_1_3/temp1[45] ,
         \MC_ARK_ARC_1_3/temp1[44] , \MC_ARK_ARC_1_3/temp1[43] ,
         \MC_ARK_ARC_1_3/temp1[42] , \MC_ARK_ARC_1_3/temp1[41] ,
         \MC_ARK_ARC_1_3/temp1[40] , \MC_ARK_ARC_1_3/temp1[39] ,
         \MC_ARK_ARC_1_3/temp1[38] , \MC_ARK_ARC_1_3/temp1[37] ,
         \MC_ARK_ARC_1_3/temp1[36] , \MC_ARK_ARC_1_3/temp1[35] ,
         \MC_ARK_ARC_1_3/temp1[34] , \MC_ARK_ARC_1_3/temp1[33] ,
         \MC_ARK_ARC_1_3/temp1[32] , \MC_ARK_ARC_1_3/temp1[31] ,
         \MC_ARK_ARC_1_3/temp1[30] , \MC_ARK_ARC_1_3/temp1[29] ,
         \MC_ARK_ARC_1_3/temp1[28] , \MC_ARK_ARC_1_3/temp1[27] ,
         \MC_ARK_ARC_1_3/temp1[26] , \MC_ARK_ARC_1_3/temp1[25] ,
         \MC_ARK_ARC_1_3/temp1[24] , \MC_ARK_ARC_1_3/temp1[23] ,
         \MC_ARK_ARC_1_3/temp1[22] , \MC_ARK_ARC_1_3/temp1[21] ,
         \MC_ARK_ARC_1_3/temp1[20] , \MC_ARK_ARC_1_3/temp1[19] ,
         \MC_ARK_ARC_1_3/temp1[18] , \MC_ARK_ARC_1_3/temp1[17] ,
         \MC_ARK_ARC_1_3/temp1[16] , \MC_ARK_ARC_1_3/temp1[15] ,
         \MC_ARK_ARC_1_3/temp1[14] , \MC_ARK_ARC_1_3/temp1[13] ,
         \MC_ARK_ARC_1_3/temp1[12] , \MC_ARK_ARC_1_3/temp1[11] ,
         \MC_ARK_ARC_1_3/temp1[10] , \MC_ARK_ARC_1_3/temp1[9] ,
         \MC_ARK_ARC_1_3/temp1[8] , \MC_ARK_ARC_1_3/temp1[7] ,
         \MC_ARK_ARC_1_3/temp1[6] , \MC_ARK_ARC_1_3/temp1[5] ,
         \MC_ARK_ARC_1_3/temp1[4] , \MC_ARK_ARC_1_3/temp1[3] ,
         \MC_ARK_ARC_1_3/temp1[2] , \MC_ARK_ARC_1_3/temp1[1] ,
         \MC_ARK_ARC_1_3/temp1[0] , \MC_ARK_ARC_1_3/buf_keyinput[179] ,
         \MC_ARK_ARC_1_3/buf_keyinput[173] ,
         \MC_ARK_ARC_1_3/buf_keyinput[172] ,
         \MC_ARK_ARC_1_3/buf_keyinput[166] ,
         \MC_ARK_ARC_1_3/buf_keyinput[154] ,
         \MC_ARK_ARC_1_3/buf_keyinput[142] ,
         \MC_ARK_ARC_1_3/buf_keyinput[137] , \MC_ARK_ARC_1_3/buf_keyinput[89] ,
         \MC_ARK_ARC_1_3/buf_keyinput[70] , \MC_ARK_ARC_1_3/buf_keyinput[44] ,
         \MC_ARK_ARC_1_3/buf_datainput[191] ,
         \MC_ARK_ARC_1_3/buf_datainput[185] ,
         \MC_ARK_ARC_1_3/buf_datainput[183] ,
         \MC_ARK_ARC_1_3/buf_datainput[182] ,
         \MC_ARK_ARC_1_3/buf_datainput[179] ,
         \MC_ARK_ARC_1_3/buf_datainput[178] ,
         \MC_ARK_ARC_1_3/buf_datainput[176] ,
         \MC_ARK_ARC_1_3/buf_datainput[174] ,
         \MC_ARK_ARC_1_3/buf_datainput[173] ,
         \MC_ARK_ARC_1_3/buf_datainput[172] ,
         \MC_ARK_ARC_1_3/buf_datainput[167] ,
         \MC_ARK_ARC_1_3/buf_datainput[166] ,
         \MC_ARK_ARC_1_3/buf_datainput[161] ,
         \MC_ARK_ARC_1_3/buf_datainput[155] ,
         \MC_ARK_ARC_1_3/buf_datainput[154] ,
         \MC_ARK_ARC_1_3/buf_datainput[146] ,
         \MC_ARK_ARC_1_3/buf_datainput[144] ,
         \MC_ARK_ARC_1_3/buf_datainput[143] ,
         \MC_ARK_ARC_1_3/buf_datainput[142] ,
         \MC_ARK_ARC_1_3/buf_datainput[141] ,
         \MC_ARK_ARC_1_3/buf_datainput[137] ,
         \MC_ARK_ARC_1_3/buf_datainput[136] ,
         \MC_ARK_ARC_1_3/buf_datainput[132] ,
         \MC_ARK_ARC_1_3/buf_datainput[131] ,
         \MC_ARK_ARC_1_3/buf_datainput[128] ,
         \MC_ARK_ARC_1_3/buf_datainput[125] ,
         \MC_ARK_ARC_1_3/buf_datainput[124] ,
         \MC_ARK_ARC_1_3/buf_datainput[122] ,
         \MC_ARK_ARC_1_3/buf_datainput[119] ,
         \MC_ARK_ARC_1_3/buf_datainput[117] ,
         \MC_ARK_ARC_1_3/buf_datainput[116] ,
         \MC_ARK_ARC_1_3/buf_datainput[114] ,
         \MC_ARK_ARC_1_3/buf_datainput[112] ,
         \MC_ARK_ARC_1_3/buf_datainput[111] ,
         \MC_ARK_ARC_1_3/buf_datainput[110] ,
         \MC_ARK_ARC_1_3/buf_datainput[107] ,
         \MC_ARK_ARC_1_3/buf_datainput[106] ,
         \MC_ARK_ARC_1_3/buf_datainput[104] ,
         \MC_ARK_ARC_1_3/buf_datainput[102] ,
         \MC_ARK_ARC_1_3/buf_datainput[101] ,
         \MC_ARK_ARC_1_3/buf_datainput[100] ,
         \MC_ARK_ARC_1_3/buf_datainput[95] ,
         \MC_ARK_ARC_1_3/buf_datainput[91] ,
         \MC_ARK_ARC_1_3/buf_datainput[89] ,
         \MC_ARK_ARC_1_3/buf_datainput[88] ,
         \MC_ARK_ARC_1_3/buf_datainput[83] ,
         \MC_ARK_ARC_1_3/buf_datainput[77] ,
         \MC_ARK_ARC_1_3/buf_datainput[76] ,
         \MC_ARK_ARC_1_3/buf_datainput[74] ,
         \MC_ARK_ARC_1_3/buf_datainput[71] ,
         \MC_ARK_ARC_1_3/buf_datainput[70] ,
         \MC_ARK_ARC_1_3/buf_datainput[68] ,
         \MC_ARK_ARC_1_3/buf_datainput[65] ,
         \MC_ARK_ARC_1_3/buf_datainput[64] ,
         \MC_ARK_ARC_1_3/buf_datainput[62] ,
         \MC_ARK_ARC_1_3/buf_datainput[59] ,
         \MC_ARK_ARC_1_3/buf_datainput[53] ,
         \MC_ARK_ARC_1_3/buf_datainput[52] ,
         \MC_ARK_ARC_1_3/buf_datainput[47] ,
         \MC_ARK_ARC_1_3/buf_datainput[42] ,
         \MC_ARK_ARC_1_3/buf_datainput[40] ,
         \MC_ARK_ARC_1_3/buf_datainput[35] ,
         \MC_ARK_ARC_1_3/buf_datainput[34] ,
         \MC_ARK_ARC_1_3/buf_datainput[32] ,
         \MC_ARK_ARC_1_3/buf_datainput[29] ,
         \MC_ARK_ARC_1_3/buf_datainput[26] ,
         \MC_ARK_ARC_1_3/buf_datainput[23] ,
         \MC_ARK_ARC_1_3/buf_datainput[22] ,
         \MC_ARK_ARC_1_3/buf_datainput[21] ,
         \MC_ARK_ARC_1_3/buf_datainput[20] ,
         \MC_ARK_ARC_1_3/buf_datainput[17] ,
         \MC_ARK_ARC_1_3/buf_datainput[16] ,
         \MC_ARK_ARC_1_3/buf_datainput[14] ,
         \MC_ARK_ARC_1_3/buf_datainput[12] ,
         \MC_ARK_ARC_1_3/buf_datainput[11] ,
         \MC_ARK_ARC_1_3/buf_datainput[10] , \MC_ARK_ARC_1_3/buf_datainput[5] ,
         \MC_ARK_ARC_1_3/buf_datainput[4] , \MC_ARK_ARC_1_3/buf_datainput[2] ,
         \SB1_0_0/i3[0] , \SB1_0_0/i1_7 , \SB1_0_0/i1[9] , \SB1_0_0/i0_0 ,
         \SB1_0_0/i0_3 , \SB1_0_0/i0_4 , \SB1_0_0/i0[10] , \SB1_0_0/i0[9] ,
         \SB1_0_0/i0[8] , \SB1_0_0/i0[7] , \SB1_0_0/i0[6] , \SB1_0_1/i3[0] ,
         \SB1_0_1/i1_5 , \SB1_0_1/i1_7 , \SB1_0_1/i1[9] , \SB1_0_1/i0_0 ,
         \SB1_0_1/i0_3 , \SB1_0_1/i0_4 , \SB1_0_1/i0[10] , \SB1_0_1/i0[9] ,
         \SB1_0_1/i0[8] , \SB1_0_1/i0[7] , \SB1_0_1/i0[6] , \SB1_0_2/i3[0] ,
         \SB1_0_2/i1_5 , \SB1_0_2/i1_7 , \SB1_0_2/i1[9] , \SB1_0_2/i0_0 ,
         \SB1_0_2/i0_3 , \SB1_0_2/i0_4 , \SB1_0_2/i0[10] , \SB1_0_2/i0[9] ,
         \SB1_0_2/i0[8] , \SB1_0_2/i0[7] , \SB1_0_2/i0[6] , \SB1_0_3/i3[0] ,
         \SB1_0_3/i1_5 , \SB1_0_3/i1_7 , \SB1_0_3/i1[9] , \SB1_0_3/i0_0 ,
         \SB1_0_3/i0_3 , \SB1_0_3/i0_4 , \SB1_0_3/i0[10] , \SB1_0_3/i0[9] ,
         \SB1_0_3/i0[8] , \SB1_0_3/i0[7] , \SB1_0_3/i0[6] , \SB1_0_4/i3[0] ,
         \SB1_0_4/i1_5 , \SB1_0_4/i1_7 , \SB1_0_4/i1[9] , \SB1_0_4/i0_0 ,
         \SB1_0_4/i0_3 , \SB1_0_4/i0_4 , \SB1_0_4/i0[10] , \SB1_0_4/i0[9] ,
         \SB1_0_4/i0[8] , \SB1_0_4/i0[7] , \SB1_0_4/i0[6] , \SB1_0_5/i3[0] ,
         \SB1_0_5/i1_5 , \SB1_0_5/i1_7 , \SB1_0_5/i1[9] , \SB1_0_5/i0_0 ,
         \SB1_0_5/i0_3 , \SB1_0_5/i0_4 , \SB1_0_5/i0[10] , \SB1_0_5/i0[9] ,
         \SB1_0_5/i0[8] , \SB1_0_5/i0[7] , \SB1_0_5/i0[6] , \SB1_0_6/i3[0] ,
         \SB1_0_6/i1_5 , \SB1_0_6/i1_7 , \SB1_0_6/i1[9] , \SB1_0_6/i0_0 ,
         \SB1_0_6/i0_3 , \SB1_0_6/i0_4 , \SB1_0_6/i0[10] , \SB1_0_6/i0[9] ,
         \SB1_0_6/i0[8] , \SB1_0_6/i0[7] , \SB1_0_6/i0[6] , \SB1_0_7/i3[0] ,
         \SB1_0_7/i1_5 , \SB1_0_7/i1_7 , \SB1_0_7/i1[9] , \SB1_0_7/i0_0 ,
         \SB1_0_7/i0_3 , \SB1_0_7/i0_4 , \SB1_0_7/i0[10] , \SB1_0_7/i0[9] ,
         \SB1_0_7/i0[8] , \SB1_0_7/i0[7] , \SB1_0_7/i0[6] , \SB1_0_8/i3[0] ,
         \SB1_0_8/i1_5 , \SB1_0_8/i1_7 , \SB1_0_8/i1[9] , \SB1_0_8/i0_0 ,
         \SB1_0_8/i0_3 , \SB1_0_8/i0_4 , \SB1_0_8/i0[10] , \SB1_0_8/i0[9] ,
         \SB1_0_8/i0[8] , \SB1_0_8/i0[7] , \SB1_0_8/i0[6] , \SB1_0_9/i3[0] ,
         \SB1_0_9/i1_5 , \SB1_0_9/i1_7 , \SB1_0_9/i1[9] , \SB1_0_9/i0_0 ,
         \SB1_0_9/i0_3 , \SB1_0_9/i0_4 , \SB1_0_9/i0[10] , \SB1_0_9/i0[9] ,
         \SB1_0_9/i0[8] , \SB1_0_9/i0[7] , \SB1_0_9/i0[6] , \SB1_0_10/i3[0] ,
         \SB1_0_10/i1_5 , \SB1_0_10/i1_7 , \SB1_0_10/i1[9] , \SB1_0_10/i0_0 ,
         \SB1_0_10/i0_3 , \SB1_0_10/i0_4 , \SB1_0_10/i0[10] , \SB1_0_10/i0[9] ,
         \SB1_0_10/i0[8] , \SB1_0_10/i0[7] , \SB1_0_10/i0[6] ,
         \SB1_0_11/i3[0] , \SB1_0_11/i1_5 , \SB1_0_11/i1_7 , \SB1_0_11/i1[9] ,
         \SB1_0_11/i0_0 , \SB1_0_11/i0_3 , \SB1_0_11/i0_4 , \SB1_0_11/i0[10] ,
         \SB1_0_11/i0[9] , \SB1_0_11/i0[8] , \SB1_0_11/i0[7] ,
         \SB1_0_11/i0[6] , \SB1_0_12/i3[0] , \SB1_0_12/i1_7 , \SB1_0_12/i1[9] ,
         \SB1_0_12/i0_0 , \SB1_0_12/i0_3 , \SB1_0_12/i0_4 , \SB1_0_12/i0[10] ,
         \SB1_0_12/i0[9] , \SB1_0_12/i0[8] , \SB1_0_12/i0[7] ,
         \SB1_0_12/i0[6] , \SB1_0_13/i3[0] , \SB1_0_13/i1_5 , \SB1_0_13/i1_7 ,
         \SB1_0_13/i1[9] , \SB1_0_13/i0_0 , \SB1_0_13/i0_3 , \SB1_0_13/i0_4 ,
         \SB1_0_13/i0[10] , \SB1_0_13/i0[9] , \SB1_0_13/i0[8] ,
         \SB1_0_13/i0[7] , \SB1_0_13/i0[6] , \SB1_0_14/i3[0] , \SB1_0_14/i1_5 ,
         \SB1_0_14/i1_7 , \SB1_0_14/i1[9] , \SB1_0_14/i0_0 , \SB1_0_14/i0_3 ,
         \SB1_0_14/i0_4 , \SB1_0_14/i0[10] , \SB1_0_14/i0[9] ,
         \SB1_0_14/i0[8] , \SB1_0_14/i0[7] , \SB1_0_14/i0[6] ,
         \SB1_0_15/i3[0] , \SB1_0_15/i1_5 , \SB1_0_15/i1_7 , \SB1_0_15/i1[9] ,
         \SB1_0_15/i0_0 , \SB1_0_15/i0_3 , \SB1_0_15/i0_4 , \SB1_0_15/i0[10] ,
         \SB1_0_15/i0[9] , \SB1_0_15/i0[8] , \SB1_0_15/i0[7] ,
         \SB1_0_15/i0[6] , \SB1_0_16/i3[0] , \SB1_0_16/i1_5 , \SB1_0_16/i1_7 ,
         \SB1_0_16/i1[9] , \SB1_0_16/i0_0 , \SB1_0_16/i0_3 , \SB1_0_16/i0_4 ,
         \SB1_0_16/i0[10] , \SB1_0_16/i0[9] , \SB1_0_16/i0[8] ,
         \SB1_0_16/i0[7] , \SB1_0_16/i0[6] , \SB1_0_17/i3[0] , \SB1_0_17/i1_5 ,
         \SB1_0_17/i1_7 , \SB1_0_17/i1[9] , \SB1_0_17/i0_0 , \SB1_0_17/i0_3 ,
         \SB1_0_17/i0_4 , \SB1_0_17/i0[10] , \SB1_0_17/i0[9] ,
         \SB1_0_17/i0[8] , \SB1_0_17/i0[7] , \SB1_0_17/i0[6] ,
         \SB1_0_18/i3[0] , \SB1_0_18/i1_5 , \SB1_0_18/i1_7 , \SB1_0_18/i1[9] ,
         \SB1_0_18/i0_0 , \SB1_0_18/i0_3 , \SB1_0_18/i0_4 , \SB1_0_18/i0[10] ,
         \SB1_0_18/i0[9] , \SB1_0_18/i0[8] , \SB1_0_18/i0[7] ,
         \SB1_0_18/i0[6] , \SB1_0_19/i3[0] , \SB1_0_19/i1_5 , \SB1_0_19/i1_7 ,
         \SB1_0_19/i1[9] , \SB1_0_19/i0_0 , \SB1_0_19/i0_3 , \SB1_0_19/i0_4 ,
         \SB1_0_19/i0[10] , \SB1_0_19/i0[9] , \SB1_0_19/i0[8] ,
         \SB1_0_19/i0[7] , \SB1_0_19/i0[6] , \SB1_0_20/i3[0] , \SB1_0_20/i1_5 ,
         \SB1_0_20/i1_7 , \SB1_0_20/i1[9] , \SB1_0_20/i0_0 , \SB1_0_20/i0_3 ,
         \SB1_0_20/i0_4 , \SB1_0_20/i0[10] , \SB1_0_20/i0[9] ,
         \SB1_0_20/i0[8] , \SB1_0_20/i0[7] , \SB1_0_20/i0[6] ,
         \SB1_0_21/i3[0] , \SB1_0_21/i1_5 , \SB1_0_21/i1_7 , \SB1_0_21/i1[9] ,
         \SB1_0_21/i0_0 , \SB1_0_21/i0_3 , \SB1_0_21/i0_4 , \SB1_0_21/i0[10] ,
         \SB1_0_21/i0[9] , \SB1_0_21/i0[8] , \SB1_0_21/i0[7] ,
         \SB1_0_21/i0[6] , \SB1_0_22/i3[0] , \SB1_0_22/i1_5 , \SB1_0_22/i1_7 ,
         \SB1_0_22/i1[9] , \SB1_0_22/i0_0 , \SB1_0_22/i0_3 , \SB1_0_22/i0_4 ,
         \SB1_0_22/i0[10] , \SB1_0_22/i0[9] , \SB1_0_22/i0[8] ,
         \SB1_0_22/i0[7] , \SB1_0_22/i0[6] , \SB1_0_23/i3[0] , \SB1_0_23/i1_5 ,
         \SB1_0_23/i1_7 , \SB1_0_23/i1[9] , \SB1_0_23/i0_0 , \SB1_0_23/i0_3 ,
         \SB1_0_23/i0_4 , \SB1_0_23/i0[10] , \SB1_0_23/i0[9] ,
         \SB1_0_23/i0[8] , \SB1_0_23/i0[7] , \SB1_0_23/i0[6] ,
         \SB1_0_24/i3[0] , \SB1_0_24/i1_5 , \SB1_0_24/i1_7 , \SB1_0_24/i1[9] ,
         \SB1_0_24/i0_0 , \SB1_0_24/i0_3 , \SB1_0_24/i0_4 , \SB1_0_24/i0[10] ,
         \SB1_0_24/i0[9] , \SB1_0_24/i0[8] , \SB1_0_24/i0[7] ,
         \SB1_0_24/i0[6] , \SB1_0_25/i3[0] , \SB1_0_25/i1_5 , \SB1_0_25/i1_7 ,
         \SB1_0_25/i1[9] , \SB1_0_25/i0_0 , \SB1_0_25/i0_3 , \SB1_0_25/i0_4 ,
         \SB1_0_25/i0[10] , \SB1_0_25/i0[9] , \SB1_0_25/i0[8] ,
         \SB1_0_25/i0[7] , \SB1_0_25/i0[6] , \SB1_0_26/i3[0] , \SB1_0_26/i1_5 ,
         \SB1_0_26/i1_7 , \SB1_0_26/i1[9] , \SB1_0_26/i0_0 , \SB1_0_26/i0_3 ,
         \SB1_0_26/i0_4 , \SB1_0_26/i0[10] , \SB1_0_26/i0[9] ,
         \SB1_0_26/i0[8] , \SB1_0_26/i0[7] , \SB1_0_26/i0[6] ,
         \SB1_0_27/i3[0] , \SB1_0_27/i1_5 , \SB1_0_27/i1_7 , \SB1_0_27/i1[9] ,
         \SB1_0_27/i0_0 , \SB1_0_27/i0_3 , \SB1_0_27/i0_4 , \SB1_0_27/i0[10] ,
         \SB1_0_27/i0[9] , \SB1_0_27/i0[8] , \SB1_0_27/i0[7] ,
         \SB1_0_27/i0[6] , \SB1_0_28/i3[0] , \SB1_0_28/i1_5 , \SB1_0_28/i1_7 ,
         \SB1_0_28/i1[9] , \SB1_0_28/i0_0 , \SB1_0_28/i0_3 , \SB1_0_28/i0_4 ,
         \SB1_0_28/i0[10] , \SB1_0_28/i0[9] , \SB1_0_28/i0[8] ,
         \SB1_0_28/i0[7] , \SB1_0_28/i0[6] , \SB1_0_29/i3[0] , \SB1_0_29/i1_5 ,
         \SB1_0_29/i1_7 , \SB1_0_29/i1[9] , \SB1_0_29/i0_0 , \SB1_0_29/i0_3 ,
         \SB1_0_29/i0_4 , \SB1_0_29/i0[10] , \SB1_0_29/i0[9] ,
         \SB1_0_29/i0[8] , \SB1_0_29/i0[7] , \SB1_0_29/i0[6] ,
         \SB1_0_30/i3[0] , \SB1_0_30/i1_5 , \SB1_0_30/i1_7 , \SB1_0_30/i1[9] ,
         \SB1_0_30/i0_0 , \SB1_0_30/i0_3 , \SB1_0_30/i0_4 , \SB1_0_30/i0[10] ,
         \SB1_0_30/i0[9] , \SB1_0_30/i0[8] , \SB1_0_30/i0[7] ,
         \SB1_0_30/i0[6] , \SB1_0_31/i3[0] , \SB1_0_31/i1_5 , \SB1_0_31/i1_7 ,
         \SB1_0_31/i1[9] , \SB1_0_31/i0_0 , \SB1_0_31/i0_3 , \SB1_0_31/i0_4 ,
         \SB1_0_31/i0[10] , \SB1_0_31/i0[9] , \SB1_0_31/i0[8] ,
         \SB1_0_31/i0[7] , \SB1_0_31/i0[6] , \SB1_1_0/i3[0] , \SB1_1_0/i1_5 ,
         \SB1_1_0/i1_7 , \SB1_1_0/i1[9] , \SB1_1_0/i0_0 , \SB1_1_0/i0_3 ,
         \SB1_1_0/i0_4 , \SB1_1_0/i0[10] , \SB1_1_0/i0[9] , \SB1_1_0/i0[8] ,
         \SB1_1_0/i0[7] , \SB1_1_0/i0[6] , \SB1_1_1/i3[0] , \SB1_1_1/i1_5 ,
         \SB1_1_1/i1_7 , \SB1_1_1/i1[9] , \SB1_1_1/i0_0 , \SB1_1_1/i0_3 ,
         \SB1_1_1/i0_4 , \SB1_1_1/i0[10] , \SB1_1_1/i0[9] , \SB1_1_1/i0[8] ,
         \SB1_1_1/i0[7] , \SB1_1_1/i0[6] , \SB1_1_2/i3[0] , \SB1_1_2/i1_5 ,
         \SB1_1_2/i1_7 , \SB1_1_2/i1[9] , \SB1_1_2/i0_0 , \SB1_1_2/i0_3 ,
         \SB1_1_2/i0_4 , \SB1_1_2/i0[10] , \SB1_1_2/i0[9] , \SB1_1_2/i0[8] ,
         \SB1_1_2/i0[7] , \SB1_1_2/i0[6] , \SB1_1_3/i3[0] , \SB1_1_3/i1_5 ,
         \SB1_1_3/i1_7 , \SB1_1_3/i1[9] , \SB1_1_3/i0_0 , \SB1_1_3/i0_3 ,
         \SB1_1_3/i0_4 , \SB1_1_3/i0[10] , \SB1_1_3/i0[9] , \SB1_1_3/i0[8] ,
         \SB1_1_3/i0[7] , \SB1_1_3/i0[6] , \SB1_1_4/i3[0] , \SB1_1_4/i1_5 ,
         \SB1_1_4/i1_7 , \SB1_1_4/i1[9] , \SB1_1_4/i0_0 , \SB1_1_4/i0_3 ,
         \SB1_1_4/i0_4 , \SB1_1_4/i0[10] , \SB1_1_4/i0[9] , \SB1_1_4/i0[8] ,
         \SB1_1_4/i0[7] , \SB1_1_4/i0[6] , \SB1_1_5/i3[0] , \SB1_1_5/i1_5 ,
         \SB1_1_5/i1_7 , \SB1_1_5/i1[9] , \SB1_1_5/i0_0 , \SB1_1_5/i0_3 ,
         \SB1_1_5/i0_4 , \SB1_1_5/i0[10] , \SB1_1_5/i0[9] , \SB1_1_5/i0[8] ,
         \SB1_1_5/i0[7] , \SB1_1_5/i0[6] , \SB1_1_6/i3[0] , \SB1_1_6/i1_5 ,
         \SB1_1_6/i1_7 , \SB1_1_6/i1[9] , \SB1_1_6/i0_0 , \SB1_1_6/i0_3 ,
         \SB1_1_6/i0_4 , \SB1_1_6/i0[10] , \SB1_1_6/i0[9] , \SB1_1_6/i0[8] ,
         \SB1_1_6/i0[7] , \SB1_1_6/i0[6] , \SB1_1_7/i3[0] , \SB1_1_7/i1_5 ,
         \SB1_1_7/i1_7 , \SB1_1_7/i1[9] , \SB1_1_7/i0_0 , \SB1_1_7/i0_3 ,
         \SB1_1_7/i0_4 , \SB1_1_7/i0[10] , \SB1_1_7/i0[9] , \SB1_1_7/i0[8] ,
         \SB1_1_7/i0[7] , \SB1_1_7/i0[6] , \SB1_1_8/i3[0] , \SB1_1_8/i1_5 ,
         \SB1_1_8/i1_7 , \SB1_1_8/i1[9] , \SB1_1_8/i0_0 , \SB1_1_8/i0_3 ,
         \SB1_1_8/i0_4 , \SB1_1_8/i0[10] , \SB1_1_8/i0[9] , \SB1_1_8/i0[8] ,
         \SB1_1_8/i0[7] , \SB1_1_8/i0[6] , \SB1_1_9/i3[0] , \SB1_1_9/i1_5 ,
         \SB1_1_9/i1_7 , \SB1_1_9/i1[9] , \SB1_1_9/i0_0 , \SB1_1_9/i0_3 ,
         \SB1_1_9/i0_4 , \SB1_1_9/i0[10] , \SB1_1_9/i0[9] , \SB1_1_9/i0[8] ,
         \SB1_1_9/i0[7] , \SB1_1_9/i0[6] , \SB1_1_10/i3[0] , \SB1_1_10/i1_5 ,
         \SB1_1_10/i1_7 , \SB1_1_10/i1[9] , \SB1_1_10/i0_0 , \SB1_1_10/i0_3 ,
         \SB1_1_10/i0_4 , \SB1_1_10/i0[10] , \SB1_1_10/i0[9] ,
         \SB1_1_10/i0[8] , \SB1_1_10/i0[7] , \SB1_1_10/i0[6] ,
         \SB1_1_11/i3[0] , \SB1_1_11/i1_5 , \SB1_1_11/i1_7 , \SB1_1_11/i1[9] ,
         \SB1_1_11/i0_0 , \SB1_1_11/i0_3 , \SB1_1_11/i0_4 , \SB1_1_11/i0[10] ,
         \SB1_1_11/i0[9] , \SB1_1_11/i0[8] , \SB1_1_11/i0[7] ,
         \SB1_1_11/i0[6] , \SB1_1_12/i3[0] , \SB1_1_12/i1_5 , \SB1_1_12/i1_7 ,
         \SB1_1_12/i1[9] , \SB1_1_12/i0_0 , \SB1_1_12/i0_3 , \SB1_1_12/i0_4 ,
         \SB1_1_12/i0[10] , \SB1_1_12/i0[9] , \SB1_1_12/i0[8] ,
         \SB1_1_12/i0[7] , \SB1_1_12/i0[6] , \SB1_1_13/i3[0] , \SB1_1_13/i1_5 ,
         \SB1_1_13/i1_7 , \SB1_1_13/i1[9] , \SB1_1_13/i0_0 , \SB1_1_13/i0_3 ,
         \SB1_1_13/i0_4 , \SB1_1_13/i0[10] , \SB1_1_13/i0[9] ,
         \SB1_1_13/i0[8] , \SB1_1_13/i0[7] , \SB1_1_13/i0[6] ,
         \SB1_1_14/i3[0] , \SB1_1_14/i1_5 , \SB1_1_14/i1_7 , \SB1_1_14/i1[9] ,
         \SB1_1_14/i0_0 , \SB1_1_14/i0_3 , \SB1_1_14/i0_4 , \SB1_1_14/i0[10] ,
         \SB1_1_14/i0[9] , \SB1_1_14/i0[8] , \SB1_1_14/i0[7] ,
         \SB1_1_14/i0[6] , \SB1_1_15/i3[0] , \SB1_1_15/i1_5 , \SB1_1_15/i1_7 ,
         \SB1_1_15/i1[9] , \SB1_1_15/i0_0 , \SB1_1_15/i0_3 , \SB1_1_15/i0_4 ,
         \SB1_1_15/i0[10] , \SB1_1_15/i0[9] , \SB1_1_15/i0[8] ,
         \SB1_1_15/i0[7] , \SB1_1_15/i0[6] , \SB1_1_16/i3[0] , \SB1_1_16/i1_5 ,
         \SB1_1_16/i1_7 , \SB1_1_16/i1[9] , \SB1_1_16/i0_0 , \SB1_1_16/i0_3 ,
         \SB1_1_16/i0_4 , \SB1_1_16/i0[10] , \SB1_1_16/i0[9] ,
         \SB1_1_16/i0[8] , \SB1_1_16/i0[7] , \SB1_1_16/i0[6] ,
         \SB1_1_17/i3[0] , \SB1_1_17/i1_5 , \SB1_1_17/i1_7 , \SB1_1_17/i1[9] ,
         \SB1_1_17/i0_0 , \SB1_1_17/i0_3 , \SB1_1_17/i0_4 , \SB1_1_17/i0[10] ,
         \SB1_1_17/i0[9] , \SB1_1_17/i0[8] , \SB1_1_17/i0[7] ,
         \SB1_1_17/i0[6] , \SB1_1_18/i3[0] , \SB1_1_18/i1_5 , \SB1_1_18/i1_7 ,
         \SB1_1_18/i1[9] , \SB1_1_18/i0_0 , \SB1_1_18/i0_3 , \SB1_1_18/i0_4 ,
         \SB1_1_18/i0[10] , \SB1_1_18/i0[9] , \SB1_1_18/i0[8] ,
         \SB1_1_18/i0[7] , \SB1_1_18/i0[6] , \SB1_1_19/i3[0] , \SB1_1_19/i1_5 ,
         \SB1_1_19/i1_7 , \SB1_1_19/i1[9] , \SB1_1_19/i0_0 , \SB1_1_19/i0_3 ,
         \SB1_1_19/i0_4 , \SB1_1_19/i0[10] , \SB1_1_19/i0[9] ,
         \SB1_1_19/i0[8] , \SB1_1_19/i0[7] , \SB1_1_19/i0[6] ,
         \SB1_1_20/i3[0] , \SB1_1_20/i1_5 , \SB1_1_20/i1_7 , \SB1_1_20/i1[9] ,
         \SB1_1_20/i0_0 , \SB1_1_20/i0_3 , \SB1_1_20/i0_4 , \SB1_1_20/i0[10] ,
         \SB1_1_20/i0[9] , \SB1_1_20/i0[8] , \SB1_1_20/i0[7] ,
         \SB1_1_20/i0[6] , \SB1_1_21/i3[0] , \SB1_1_21/i1_5 , \SB1_1_21/i1_7 ,
         \SB1_1_21/i1[9] , \SB1_1_21/i0_0 , \SB1_1_21/i0_3 , \SB1_1_21/i0_4 ,
         \SB1_1_21/i0[10] , \SB1_1_21/i0[9] , \SB1_1_21/i0[8] ,
         \SB1_1_21/i0[7] , \SB1_1_21/i0[6] , \SB1_1_22/i3[0] , \SB1_1_22/i1_5 ,
         \SB1_1_22/i1_7 , \SB1_1_22/i1[9] , \SB1_1_22/i0_0 , \SB1_1_22/i0_3 ,
         \SB1_1_22/i0_4 , \SB1_1_22/i0[10] , \SB1_1_22/i0[9] ,
         \SB1_1_22/i0[8] , \SB1_1_22/i0[7] , \SB1_1_22/i0[6] ,
         \SB1_1_23/i3[0] , \SB1_1_23/i1_5 , \SB1_1_23/i1_7 , \SB1_1_23/i1[9] ,
         \SB1_1_23/i0_0 , \SB1_1_23/i0_3 , \SB1_1_23/i0_4 , \SB1_1_23/i0[10] ,
         \SB1_1_23/i0[9] , \SB1_1_23/i0[8] , \SB1_1_23/i0[7] ,
         \SB1_1_23/i0[6] , \SB1_1_24/i3[0] , \SB1_1_24/i1_5 , \SB1_1_24/i1_7 ,
         \SB1_1_24/i1[9] , \SB1_1_24/i0_0 , \SB1_1_24/i0_3 , \SB1_1_24/i0_4 ,
         \SB1_1_24/i0[10] , \SB1_1_24/i0[9] , \SB1_1_24/i0[8] ,
         \SB1_1_24/i0[7] , \SB1_1_24/i0[6] , \SB1_1_25/i3[0] , \SB1_1_25/i1_5 ,
         \SB1_1_25/i1_7 , \SB1_1_25/i1[9] , \SB1_1_25/i0_0 , \SB1_1_25/i0_3 ,
         \SB1_1_25/i0_4 , \SB1_1_25/i0[10] , \SB1_1_25/i0[9] ,
         \SB1_1_25/i0[8] , \SB1_1_25/i0[7] , \SB1_1_25/i0[6] ,
         \SB1_1_26/i3[0] , \SB1_1_26/i1_5 , \SB1_1_26/i1_7 , \SB1_1_26/i1[9] ,
         \SB1_1_26/i0_0 , \SB1_1_26/i0_3 , \SB1_1_26/i0_4 , \SB1_1_26/i0[10] ,
         \SB1_1_26/i0[9] , \SB1_1_26/i0[8] , \SB1_1_26/i0[7] ,
         \SB1_1_26/i0[6] , \SB1_1_27/i3[0] , \SB1_1_27/i1_5 , \SB1_1_27/i1_7 ,
         \SB1_1_27/i1[9] , \SB1_1_27/i0_0 , \SB1_1_27/i0_3 , \SB1_1_27/i0_4 ,
         \SB1_1_27/i0[10] , \SB1_1_27/i0[9] , \SB1_1_27/i0[8] ,
         \SB1_1_27/i0[7] , \SB1_1_27/i0[6] , \SB1_1_28/i3[0] , \SB1_1_28/i1_5 ,
         \SB1_1_28/i1_7 , \SB1_1_28/i1[9] , \SB1_1_28/i0_0 , \SB1_1_28/i0_3 ,
         \SB1_1_28/i0_4 , \SB1_1_28/i0[10] , \SB1_1_28/i0[9] ,
         \SB1_1_28/i0[8] , \SB1_1_28/i0[7] , \SB1_1_28/i0[6] ,
         \SB1_1_29/i3[0] , \SB1_1_29/i1_5 , \SB1_1_29/i1_7 , \SB1_1_29/i1[9] ,
         \SB1_1_29/i0_0 , \SB1_1_29/i0_3 , \SB1_1_29/i0_4 , \SB1_1_29/i0[10] ,
         \SB1_1_29/i0[9] , \SB1_1_29/i0[8] , \SB1_1_29/i0[7] ,
         \SB1_1_29/i0[6] , \SB1_1_30/i3[0] , \SB1_1_30/i1_5 , \SB1_1_30/i1_7 ,
         \SB1_1_30/i1[9] , \SB1_1_30/i0_0 , \SB1_1_30/i0_3 , \SB1_1_30/i0_4 ,
         \SB1_1_30/i0[10] , \SB1_1_30/i0[9] , \SB1_1_30/i0[8] ,
         \SB1_1_30/i0[7] , \SB1_1_30/i0[6] , \SB1_1_31/i3[0] , \SB1_1_31/i1_5 ,
         \SB1_1_31/i1_7 , \SB1_1_31/i1[9] , \SB1_1_31/i0_0 , \SB1_1_31/i0_3 ,
         \SB1_1_31/i0_4 , \SB1_1_31/i0[10] , \SB1_1_31/i0[9] ,
         \SB1_1_31/i0[8] , \SB1_1_31/i0[7] , \SB1_1_31/i0[6] , \SB1_2_0/i3[0] ,
         \SB1_2_0/i1_5 , \SB1_2_0/i1_7 , \SB1_2_0/i1[9] , \SB1_2_0/i0_0 ,
         \SB1_2_0/i0_3 , \SB1_2_0/i0_4 , \SB1_2_0/i0[10] , \SB1_2_0/i0[9] ,
         \SB1_2_0/i0[8] , \SB1_2_0/i0[7] , \SB1_2_0/i0[6] , \SB1_2_1/i3[0] ,
         \SB1_2_1/i1_5 , \SB1_2_1/i1_7 , \SB1_2_1/i1[9] , \SB1_2_1/i0_0 ,
         \SB1_2_1/i0_3 , \SB1_2_1/i0_4 , \SB1_2_1/i0[10] , \SB1_2_1/i0[9] ,
         \SB1_2_1/i0[8] , \SB1_2_1/i0[7] , \SB1_2_1/i0[6] , \SB1_2_2/i3[0] ,
         \SB1_2_2/i1_5 , \SB1_2_2/i1_7 , \SB1_2_2/i1[9] , \SB1_2_2/i0_0 ,
         \SB1_2_2/i0_3 , \SB1_2_2/i0_4 , \SB1_2_2/i0[10] , \SB1_2_2/i0[9] ,
         \SB1_2_2/i0[8] , \SB1_2_2/i0[7] , \SB1_2_2/i0[6] , \SB1_2_3/i3[0] ,
         \SB1_2_3/i1_5 , \SB1_2_3/i1_7 , \SB1_2_3/i1[9] , \SB1_2_3/i0_0 ,
         \SB1_2_3/i0_3 , \SB1_2_3/i0_4 , \SB1_2_3/i0[10] , \SB1_2_3/i0[9] ,
         \SB1_2_3/i0[8] , \SB1_2_3/i0[7] , \SB1_2_3/i0[6] , \SB1_2_4/i3[0] ,
         \SB1_2_4/i1_5 , \SB1_2_4/i1_7 , \SB1_2_4/i1[9] , \SB1_2_4/i0_0 ,
         \SB1_2_4/i0_3 , \SB1_2_4/i0_4 , \SB1_2_4/i0[10] , \SB1_2_4/i0[9] ,
         \SB1_2_4/i0[8] , \SB1_2_4/i0[7] , \SB1_2_4/i0[6] , \SB1_2_5/i3[0] ,
         \SB1_2_5/i1_5 , \SB1_2_5/i1_7 , \SB1_2_5/i1[9] , \SB1_2_5/i0_0 ,
         \SB1_2_5/i0_3 , \SB1_2_5/i0_4 , \SB1_2_5/i0[10] , \SB1_2_5/i0[9] ,
         \SB1_2_5/i0[8] , \SB1_2_5/i0[7] , \SB1_2_5/i0[6] , \SB1_2_6/i3[0] ,
         \SB1_2_6/i1_5 , \SB1_2_6/i1_7 , \SB1_2_6/i1[9] , \SB1_2_6/i0_0 ,
         \SB1_2_6/i0_3 , \SB1_2_6/i0_4 , \SB1_2_6/i0[10] , \SB1_2_6/i0[9] ,
         \SB1_2_6/i0[8] , \SB1_2_6/i0[7] , \SB1_2_6/i0[6] , \SB1_2_7/i3[0] ,
         \SB1_2_7/i1_5 , \SB1_2_7/i1_7 , \SB1_2_7/i1[9] , \SB1_2_7/i0_0 ,
         \SB1_2_7/i0_3 , \SB1_2_7/i0_4 , \SB1_2_7/i0[10] , \SB1_2_7/i0[9] ,
         \SB1_2_7/i0[8] , \SB1_2_7/i0[7] , \SB1_2_7/i0[6] , \SB1_2_8/i3[0] ,
         \SB1_2_8/i1_5 , \SB1_2_8/i1_7 , \SB1_2_8/i1[9] , \SB1_2_8/i0_0 ,
         \SB1_2_8/i0_3 , \SB1_2_8/i0_4 , \SB1_2_8/i0[10] , \SB1_2_8/i0[9] ,
         \SB1_2_8/i0[8] , \SB1_2_8/i0[7] , \SB1_2_8/i0[6] , \SB1_2_9/i3[0] ,
         \SB1_2_9/i1_5 , \SB1_2_9/i1_7 , \SB1_2_9/i1[9] , \SB1_2_9/i0_0 ,
         \SB1_2_9/i0_4 , \SB1_2_9/i0[10] , \SB1_2_9/i0[9] , \SB1_2_9/i0[8] ,
         \SB1_2_9/i0[7] , \SB1_2_9/i0[6] , \SB1_2_10/i3[0] , \SB1_2_10/i1_5 ,
         \SB1_2_10/i1_7 , \SB1_2_10/i1[9] , \SB1_2_10/i0_0 , \SB1_2_10/i0_3 ,
         \SB1_2_10/i0_4 , \SB1_2_10/i0[10] , \SB1_2_10/i0[9] ,
         \SB1_2_10/i0[8] , \SB1_2_10/i0[7] , \SB1_2_10/i0[6] ,
         \SB1_2_11/i3[0] , \SB1_2_11/i1_5 , \SB1_2_11/i1_7 , \SB1_2_11/i1[9] ,
         \SB1_2_11/i0_0 , \SB1_2_11/i0_3 , \SB1_2_11/i0_4 , \SB1_2_11/i0[10] ,
         \SB1_2_11/i0[9] , \SB1_2_11/i0[8] , \SB1_2_11/i0[7] ,
         \SB1_2_11/i0[6] , \SB1_2_12/i3[0] , \SB1_2_12/i1_5 , \SB1_2_12/i1_7 ,
         \SB1_2_12/i1[9] , \SB1_2_12/i0_0 , \SB1_2_12/i0_3 , \SB1_2_12/i0_4 ,
         \SB1_2_12/i0[10] , \SB1_2_12/i0[9] , \SB1_2_12/i0[8] ,
         \SB1_2_12/i0[7] , \SB1_2_12/i0[6] , \SB1_2_13/i3[0] , \SB1_2_13/i1_5 ,
         \SB1_2_13/i1_7 , \SB1_2_13/i1[9] , \SB1_2_13/i0_0 , \SB1_2_13/i0_3 ,
         \SB1_2_13/i0_4 , \SB1_2_13/i0[10] , \SB1_2_13/i0[9] ,
         \SB1_2_13/i0[8] , \SB1_2_13/i0[7] , \SB1_2_13/i0[6] ,
         \SB1_2_14/i3[0] , \SB1_2_14/i1_5 , \SB1_2_14/i1_7 , \SB1_2_14/i1[9] ,
         \SB1_2_14/i0_0 , \SB1_2_14/i0_3 , \SB1_2_14/i0_4 , \SB1_2_14/i0[10] ,
         \SB1_2_14/i0[9] , \SB1_2_14/i0[8] , \SB1_2_14/i0[7] ,
         \SB1_2_14/i0[6] , \SB1_2_15/i3[0] , \SB1_2_15/i1_5 , \SB1_2_15/i1_7 ,
         \SB1_2_15/i1[9] , \SB1_2_15/i0_0 , \SB1_2_15/i0_3 , \SB1_2_15/i0_4 ,
         \SB1_2_15/i0[10] , \SB1_2_15/i0[9] , \SB1_2_15/i0[8] ,
         \SB1_2_15/i0[7] , \SB1_2_15/i0[6] , \SB1_2_16/i3[0] , \SB1_2_16/i1_5 ,
         \SB1_2_16/i1_7 , \SB1_2_16/i1[9] , \SB1_2_16/i0_0 , \SB1_2_16/i0_3 ,
         \SB1_2_16/i0_4 , \SB1_2_16/i0[10] , \SB1_2_16/i0[9] ,
         \SB1_2_16/i0[8] , \SB1_2_16/i0[7] , \SB1_2_16/i0[6] ,
         \SB1_2_17/i3[0] , \SB1_2_17/i1_5 , \SB1_2_17/i1_7 , \SB1_2_17/i1[9] ,
         \SB1_2_17/i0_0 , \SB1_2_17/i0_3 , \SB1_2_17/i0_4 , \SB1_2_17/i0[10] ,
         \SB1_2_17/i0[9] , \SB1_2_17/i0[8] , \SB1_2_17/i0[7] ,
         \SB1_2_17/i0[6] , \SB1_2_18/i3[0] , \SB1_2_18/i1_5 , \SB1_2_18/i1_7 ,
         \SB1_2_18/i1[9] , \SB1_2_18/i0_0 , \SB1_2_18/i0_3 , \SB1_2_18/i0_4 ,
         \SB1_2_18/i0[10] , \SB1_2_18/i0[9] , \SB1_2_18/i0[8] ,
         \SB1_2_18/i0[7] , \SB1_2_18/i0[6] , \SB1_2_19/i3[0] , \SB1_2_19/i1_5 ,
         \SB1_2_19/i1_7 , \SB1_2_19/i1[9] , \SB1_2_19/i0_0 , \SB1_2_19/i0_3 ,
         \SB1_2_19/i0_4 , \SB1_2_19/i0[10] , \SB1_2_19/i0[9] ,
         \SB1_2_19/i0[8] , \SB1_2_19/i0[7] , \SB1_2_19/i0[6] ,
         \SB1_2_20/i3[0] , \SB1_2_20/i1_5 , \SB1_2_20/i1_7 , \SB1_2_20/i1[9] ,
         \SB1_2_20/i0_0 , \SB1_2_20/i0_3 , \SB1_2_20/i0_4 , \SB1_2_20/i0[10] ,
         \SB1_2_20/i0[9] , \SB1_2_20/i0[8] , \SB1_2_20/i0[7] ,
         \SB1_2_20/i0[6] , \SB1_2_21/i3[0] , \SB1_2_21/i1_5 , \SB1_2_21/i1_7 ,
         \SB1_2_21/i1[9] , \SB1_2_21/i0_0 , \SB1_2_21/i0_3 , \SB1_2_21/i0_4 ,
         \SB1_2_21/i0[10] , \SB1_2_21/i0[9] , \SB1_2_21/i0[8] ,
         \SB1_2_21/i0[7] , \SB1_2_21/i0[6] , \SB1_2_22/i3[0] , \SB1_2_22/i1_5 ,
         \SB1_2_22/i1_7 , \SB1_2_22/i1[9] , \SB1_2_22/i0_0 , \SB1_2_22/i0_3 ,
         \SB1_2_22/i0_4 , \SB1_2_22/i0[10] , \SB1_2_22/i0[9] ,
         \SB1_2_22/i0[8] , \SB1_2_22/i0[7] , \SB1_2_22/i0[6] ,
         \SB1_2_23/i3[0] , \SB1_2_23/i1_5 , \SB1_2_23/i1_7 , \SB1_2_23/i1[9] ,
         \SB1_2_23/i0_0 , \SB1_2_23/i0_3 , \SB1_2_23/i0_4 , \SB1_2_23/i0[10] ,
         \SB1_2_23/i0[9] , \SB1_2_23/i0[8] , \SB1_2_23/i0[7] ,
         \SB1_2_23/i0[6] , \SB1_2_24/i3[0] , \SB1_2_24/i1_5 , \SB1_2_24/i1_7 ,
         \SB1_2_24/i1[9] , \SB1_2_24/i0_0 , \SB1_2_24/i0_3 , \SB1_2_24/i0_4 ,
         \SB1_2_24/i0[10] , \SB1_2_24/i0[9] , \SB1_2_24/i0[8] ,
         \SB1_2_24/i0[7] , \SB1_2_24/i0[6] , \SB1_2_25/i3[0] , \SB1_2_25/i1_5 ,
         \SB1_2_25/i1_7 , \SB1_2_25/i1[9] , \SB1_2_25/i0_0 , \SB1_2_25/i0_3 ,
         \SB1_2_25/i0_4 , \SB1_2_25/i0[10] , \SB1_2_25/i0[9] ,
         \SB1_2_25/i0[8] , \SB1_2_25/i0[7] , \SB1_2_25/i0[6] ,
         \SB1_2_26/i3[0] , \SB1_2_26/i1_5 , \SB1_2_26/i1_7 , \SB1_2_26/i1[9] ,
         \SB1_2_26/i0_0 , \SB1_2_26/i0_3 , \SB1_2_26/i0_4 , \SB1_2_26/i0[10] ,
         \SB1_2_26/i0[9] , \SB1_2_26/i0[8] , \SB1_2_26/i0[7] ,
         \SB1_2_26/i0[6] , \SB1_2_27/i3[0] , \SB1_2_27/i1_5 , \SB1_2_27/i1_7 ,
         \SB1_2_27/i1[9] , \SB1_2_27/i0_0 , \SB1_2_27/i0_3 , \SB1_2_27/i0_4 ,
         \SB1_2_27/i0[10] , \SB1_2_27/i0[9] , \SB1_2_27/i0[8] ,
         \SB1_2_27/i0[7] , \SB1_2_27/i0[6] , \SB1_2_28/i3[0] , \SB1_2_28/i1_5 ,
         \SB1_2_28/i1_7 , \SB1_2_28/i1[9] , \SB1_2_28/i0_0 , \SB1_2_28/i0_3 ,
         \SB1_2_28/i0_4 , \SB1_2_28/i0[10] , \SB1_2_28/i0[9] ,
         \SB1_2_28/i0[8] , \SB1_2_28/i0[7] , \SB1_2_28/i0[6] ,
         \SB1_2_29/i3[0] , \SB1_2_29/i1_5 , \SB1_2_29/i1_7 , \SB1_2_29/i1[9] ,
         \SB1_2_29/i0_0 , \SB1_2_29/i0_3 , \SB1_2_29/i0_4 , \SB1_2_29/i0[10] ,
         \SB1_2_29/i0[9] , \SB1_2_29/i0[8] , \SB1_2_29/i0[7] ,
         \SB1_2_29/i0[6] , \SB1_2_30/i3[0] , \SB1_2_30/i1_5 , \SB1_2_30/i1_7 ,
         \SB1_2_30/i1[9] , \SB1_2_30/i0_0 , \SB1_2_30/i0_3 , \SB1_2_30/i0_4 ,
         \SB1_2_30/i0[10] , \SB1_2_30/i0[9] , \SB1_2_30/i0[8] ,
         \SB1_2_30/i0[7] , \SB1_2_30/i0[6] , \SB1_2_31/i3[0] , \SB1_2_31/i1_5 ,
         \SB1_2_31/i1_7 , \SB1_2_31/i1[9] , \SB1_2_31/i0_0 , \SB1_2_31/i0_3 ,
         \SB1_2_31/i0_4 , \SB1_2_31/i0[10] , \SB1_2_31/i0[9] ,
         \SB1_2_31/i0[8] , \SB1_2_31/i0[7] , \SB1_2_31/i0[6] , \SB1_3_0/i3[0] ,
         \SB1_3_0/i1_5 , \SB1_3_0/i1_7 , \SB1_3_0/i1[9] , \SB1_3_0/i0_0 ,
         \SB1_3_0/i0_4 , \SB1_3_0/i0[10] , \SB1_3_0/i0[9] , \SB1_3_0/i0[8] ,
         \SB1_3_0/i0[7] , \SB1_3_0/i0[6] , \SB1_3_1/i3[0] , \SB1_3_1/i1_5 ,
         \SB1_3_1/i1_7 , \SB1_3_1/i1[9] , \SB1_3_1/i0_0 , \SB1_3_1/i0_3 ,
         \SB1_3_1/i0_4 , \SB1_3_1/i0[10] , \SB1_3_1/i0[9] , \SB1_3_1/i0[8] ,
         \SB1_3_1/i0[7] , \SB1_3_1/i0[6] , \SB1_3_2/i3[0] , \SB1_3_2/i1_5 ,
         \SB1_3_2/i1_7 , \SB1_3_2/i1[9] , \SB1_3_2/i0_0 , \SB1_3_2/i0_3 ,
         \SB1_3_2/i0_4 , \SB1_3_2/i0[10] , \SB1_3_2/i0[9] , \SB1_3_2/i0[8] ,
         \SB1_3_2/i0[7] , \SB1_3_2/i0[6] , \SB1_3_3/i3[0] , \SB1_3_3/i1_5 ,
         \SB1_3_3/i1_7 , \SB1_3_3/i1[9] , \SB1_3_3/i0_0 , \SB1_3_3/i0_3 ,
         \SB1_3_3/i0_4 , \SB1_3_3/i0[10] , \SB1_3_3/i0[9] , \SB1_3_3/i0[8] ,
         \SB1_3_3/i0[7] , \SB1_3_3/i0[6] , \SB1_3_4/i3[0] , \SB1_3_4/i1_5 ,
         \SB1_3_4/i1_7 , \SB1_3_4/i1[9] , \SB1_3_4/i0_0 , \SB1_3_4/i0_3 ,
         \SB1_3_4/i0_4 , \SB1_3_4/i0[10] , \SB1_3_4/i0[9] , \SB1_3_4/i0[8] ,
         \SB1_3_4/i0[7] , \SB1_3_4/i0[6] , \SB1_3_5/i3[0] , \SB1_3_5/i1_5 ,
         \SB1_3_5/i1_7 , \SB1_3_5/i1[9] , \SB1_3_5/i0_0 , \SB1_3_5/i0_3 ,
         \SB1_3_5/i0_4 , \SB1_3_5/i0[10] , \SB1_3_5/i0[9] , \SB1_3_5/i0[8] ,
         \SB1_3_5/i0[7] , \SB1_3_5/i0[6] , \SB1_3_6/i3[0] , \SB1_3_6/i1_5 ,
         \SB1_3_6/i1_7 , \SB1_3_6/i1[9] , \SB1_3_6/i0_0 , \SB1_3_6/i0_3 ,
         \SB1_3_6/i0_4 , \SB1_3_6/i0[10] , \SB1_3_6/i0[9] , \SB1_3_6/i0[8] ,
         \SB1_3_6/i0[7] , \SB1_3_6/i0[6] , \SB1_3_7/i3[0] , \SB1_3_7/i1_5 ,
         \SB1_3_7/i1_7 , \SB1_3_7/i1[9] , \SB1_3_7/i0_0 , \SB1_3_7/i0_3 ,
         \SB1_3_7/i0_4 , \SB1_3_7/i0[10] , \SB1_3_7/i0[9] , \SB1_3_7/i0[8] ,
         \SB1_3_7/i0[7] , \SB1_3_7/i0[6] , \SB1_3_8/i3[0] , \SB1_3_8/i1_5 ,
         \SB1_3_8/i1_7 , \SB1_3_8/i1[9] , \SB1_3_8/i0_0 , \SB1_3_8/i0_3 ,
         \SB1_3_8/i0_4 , \SB1_3_8/i0[10] , \SB1_3_8/i0[9] , \SB1_3_8/i0[8] ,
         \SB1_3_8/i0[7] , \SB1_3_8/i0[6] , \SB1_3_9/i3[0] , \SB1_3_9/i1_5 ,
         \SB1_3_9/i1_7 , \SB1_3_9/i1[9] , \SB1_3_9/i0_0 , \SB1_3_9/i0_3 ,
         \SB1_3_9/i0_4 , \SB1_3_9/i0[10] , \SB1_3_9/i0[9] , \SB1_3_9/i0[8] ,
         \SB1_3_9/i0[7] , \SB1_3_9/i0[6] , \SB1_3_10/i3[0] , \SB1_3_10/i1_5 ,
         \SB1_3_10/i1_7 , \SB1_3_10/i1[9] , \SB1_3_10/i0_0 , \SB1_3_10/i0_3 ,
         \SB1_3_10/i0_4 , \SB1_3_10/i0[10] , \SB1_3_10/i0[9] ,
         \SB1_3_10/i0[8] , \SB1_3_10/i0[7] , \SB1_3_10/i0[6] ,
         \SB1_3_11/i3[0] , \SB1_3_11/i1_5 , \SB1_3_11/i1_7 , \SB1_3_11/i1[9] ,
         \SB1_3_11/i0_0 , \SB1_3_11/i0_3 , \SB1_3_11/i0_4 , \SB1_3_11/i0[10] ,
         \SB1_3_11/i0[9] , \SB1_3_11/i0[8] , \SB1_3_11/i0[7] ,
         \SB1_3_11/i0[6] , \SB1_3_12/i3[0] , \SB1_3_12/i1_5 , \SB1_3_12/i1_7 ,
         \SB1_3_12/i1[9] , \SB1_3_12/i0_0 , \SB1_3_12/i0_3 , \SB1_3_12/i0_4 ,
         \SB1_3_12/i0[10] , \SB1_3_12/i0[9] , \SB1_3_12/i0[8] ,
         \SB1_3_12/i0[7] , \SB1_3_12/i0[6] , \SB1_3_13/i3[0] , \SB1_3_13/i1_5 ,
         \SB1_3_13/i1_7 , \SB1_3_13/i1[9] , \SB1_3_13/i0_0 , \SB1_3_13/i0_3 ,
         \SB1_3_13/i0_4 , \SB1_3_13/i0[10] , \SB1_3_13/i0[9] ,
         \SB1_3_13/i0[8] , \SB1_3_13/i0[7] , \SB1_3_13/i0[6] ,
         \SB1_3_14/i3[0] , \SB1_3_14/i1_5 , \SB1_3_14/i1_7 , \SB1_3_14/i1[9] ,
         \SB1_3_14/i0_0 , \SB1_3_14/i0_3 , \SB1_3_14/i0_4 , \SB1_3_14/i0[10] ,
         \SB1_3_14/i0[9] , \SB1_3_14/i0[8] , \SB1_3_14/i0[7] ,
         \SB1_3_14/i0[6] , \SB1_3_15/i3[0] , \SB1_3_15/i1_5 , \SB1_3_15/i1_7 ,
         \SB1_3_15/i1[9] , \SB1_3_15/i0_0 , \SB1_3_15/i0_3 , \SB1_3_15/i0_4 ,
         \SB1_3_15/i0[10] , \SB1_3_15/i0[9] , \SB1_3_15/i0[8] ,
         \SB1_3_15/i0[7] , \SB1_3_15/i0[6] , \SB1_3_16/i3[0] , \SB1_3_16/i1_5 ,
         \SB1_3_16/i1_7 , \SB1_3_16/i1[9] , \SB1_3_16/i0_0 , \SB1_3_16/i0_3 ,
         \SB1_3_16/i0_4 , \SB1_3_16/i0[10] , \SB1_3_16/i0[9] ,
         \SB1_3_16/i0[8] , \SB1_3_16/i0[7] , \SB1_3_16/i0[6] ,
         \SB1_3_17/i3[0] , \SB1_3_17/i1_5 , \SB1_3_17/i1_7 , \SB1_3_17/i1[9] ,
         \SB1_3_17/i0_0 , \SB1_3_17/i0_3 , \SB1_3_17/i0_4 , \SB1_3_17/i0[10] ,
         \SB1_3_17/i0[9] , \SB1_3_17/i0[8] , \SB1_3_17/i0[7] ,
         \SB1_3_17/i0[6] , \SB1_3_18/i3[0] , \SB1_3_18/i1_5 , \SB1_3_18/i1_7 ,
         \SB1_3_18/i1[9] , \SB1_3_18/i0_0 , \SB1_3_18/i0_3 , \SB1_3_18/i0_4 ,
         \SB1_3_18/i0[10] , \SB1_3_18/i0[9] , \SB1_3_18/i0[8] ,
         \SB1_3_18/i0[7] , \SB1_3_18/i0[6] , \SB1_3_19/i3[0] , \SB1_3_19/i1_5 ,
         \SB1_3_19/i1_7 , \SB1_3_19/i1[9] , \SB1_3_19/i0_0 , \SB1_3_19/i0_3 ,
         \SB1_3_19/i0_4 , \SB1_3_19/i0[10] , \SB1_3_19/i0[9] ,
         \SB1_3_19/i0[8] , \SB1_3_19/i0[7] , \SB1_3_19/i0[6] ,
         \SB1_3_20/i3[0] , \SB1_3_20/i1_5 , \SB1_3_20/i1_7 , \SB1_3_20/i1[9] ,
         \SB1_3_20/i0_0 , \SB1_3_20/i0_3 , \SB1_3_20/i0_4 , \SB1_3_20/i0[10] ,
         \SB1_3_20/i0[9] , \SB1_3_20/i0[8] , \SB1_3_20/i0[7] ,
         \SB1_3_20/i0[6] , \SB1_3_21/i3[0] , \SB1_3_21/i1_5 , \SB1_3_21/i1_7 ,
         \SB1_3_21/i1[9] , \SB1_3_21/i0_0 , \SB1_3_21/i0_3 , \SB1_3_21/i0_4 ,
         \SB1_3_21/i0[10] , \SB1_3_21/i0[9] , \SB1_3_21/i0[8] ,
         \SB1_3_21/i0[7] , \SB1_3_21/i0[6] , \SB1_3_22/i3[0] , \SB1_3_22/i1_5 ,
         \SB1_3_22/i1_7 , \SB1_3_22/i1[9] , \SB1_3_22/i0_0 , \SB1_3_22/i0_3 ,
         \SB1_3_22/i0_4 , \SB1_3_22/i0[10] , \SB1_3_22/i0[9] ,
         \SB1_3_22/i0[8] , \SB1_3_22/i0[7] , \SB1_3_22/i0[6] ,
         \SB1_3_23/i3[0] , \SB1_3_23/i1_5 , \SB1_3_23/i1_7 , \SB1_3_23/i1[9] ,
         \SB1_3_23/i0_0 , \SB1_3_23/i0_3 , \SB1_3_23/i0_4 , \SB1_3_23/i0[10] ,
         \SB1_3_23/i0[9] , \SB1_3_23/i0[8] , \SB1_3_23/i0[7] ,
         \SB1_3_23/i0[6] , \SB1_3_24/i3[0] , \SB1_3_24/i1_5 , \SB1_3_24/i1_7 ,
         \SB1_3_24/i1[9] , \SB1_3_24/i0_0 , \SB1_3_24/i0_3 , \SB1_3_24/i0_4 ,
         \SB1_3_24/i0[10] , \SB1_3_24/i0[9] , \SB1_3_24/i0[8] ,
         \SB1_3_24/i0[7] , \SB1_3_24/i0[6] , \SB1_3_25/i3[0] , \SB1_3_25/i1_5 ,
         \SB1_3_25/i1_7 , \SB1_3_25/i1[9] , \SB1_3_25/i0_0 , \SB1_3_25/i0_3 ,
         \SB1_3_25/i0_4 , \SB1_3_25/i0[10] , \SB1_3_25/i0[9] ,
         \SB1_3_25/i0[8] , \SB1_3_25/i0[7] , \SB1_3_25/i0[6] ,
         \SB1_3_26/i3[0] , \SB1_3_26/i1_5 , \SB1_3_26/i1_7 , \SB1_3_26/i1[9] ,
         \SB1_3_26/i0_0 , \SB1_3_26/i0_3 , \SB1_3_26/i0_4 , \SB1_3_26/i0[10] ,
         \SB1_3_26/i0[9] , \SB1_3_26/i0[8] , \SB1_3_26/i0[7] ,
         \SB1_3_26/i0[6] , \SB1_3_27/i3[0] , \SB1_3_27/i1_5 , \SB1_3_27/i1_7 ,
         \SB1_3_27/i1[9] , \SB1_3_27/i0_0 , \SB1_3_27/i0_3 , \SB1_3_27/i0_4 ,
         \SB1_3_27/i0[10] , \SB1_3_27/i0[9] , \SB1_3_27/i0[8] ,
         \SB1_3_27/i0[7] , \SB1_3_27/i0[6] , \SB1_3_28/i3[0] , \SB1_3_28/i1_5 ,
         \SB1_3_28/i1_7 , \SB1_3_28/i1[9] , \SB1_3_28/i0_0 , \SB1_3_28/i0_3 ,
         \SB1_3_28/i0_4 , \SB1_3_28/i0[10] , \SB1_3_28/i0[9] ,
         \SB1_3_28/i0[8] , \SB1_3_28/i0[7] , \SB1_3_28/i0[6] ,
         \SB1_3_29/i3[0] , \SB1_3_29/i1_5 , \SB1_3_29/i1_7 , \SB1_3_29/i1[9] ,
         \SB1_3_29/i0_0 , \SB1_3_29/i0_3 , \SB1_3_29/i0_4 , \SB1_3_29/i0[10] ,
         \SB1_3_29/i0[9] , \SB1_3_29/i0[8] , \SB1_3_29/i0[7] ,
         \SB1_3_29/i0[6] , \SB1_3_30/i3[0] , \SB1_3_30/i1_5 , \SB1_3_30/i1_7 ,
         \SB1_3_30/i1[9] , \SB1_3_30/i0_0 , \SB1_3_30/i0_3 , \SB1_3_30/i0_4 ,
         \SB1_3_30/i0[10] , \SB1_3_30/i0[9] , \SB1_3_30/i0[8] ,
         \SB1_3_30/i0[7] , \SB1_3_30/i0[6] , \SB1_3_31/i3[0] , \SB1_3_31/i1_5 ,
         \SB1_3_31/i1_7 , \SB1_3_31/i1[9] , \SB1_3_31/i0_0 , \SB1_3_31/i0_3 ,
         \SB1_3_31/i0_4 , \SB1_3_31/i0[10] , \SB1_3_31/i0[9] ,
         \SB1_3_31/i0[8] , \SB1_3_31/i0[7] , \SB1_3_31/i0[6] , \SB3_0/i3[0] ,
         \SB3_0/i1_5 , \SB3_0/i1_7 , \SB3_0/i1[9] , \SB3_0/i0_0 , \SB3_0/i0_3 ,
         \SB3_0/i0_4 , \SB3_0/i0[10] , \SB3_0/i0[9] , \SB3_0/i0[8] ,
         \SB3_0/i0[7] , \SB3_0/i0[6] , \SB3_1/i3[0] , \SB3_1/i1_5 ,
         \SB3_1/i1_7 , \SB3_1/i1[9] , \SB3_1/i0_0 , \SB3_1/i0_3 , \SB3_1/i0_4 ,
         \SB3_1/i0[10] , \SB3_1/i0[9] , \SB3_1/i0[8] , \SB3_1/i0[7] ,
         \SB3_1/i0[6] , \SB3_2/i3[0] , \SB3_2/i1_5 , \SB3_2/i1_7 ,
         \SB3_2/i1[9] , \SB3_2/i0_0 , \SB3_2/i0_3 , \SB3_2/i0_4 ,
         \SB3_2/i0[10] , \SB3_2/i0[9] , \SB3_2/i0[8] , \SB3_2/i0[7] ,
         \SB3_2/i0[6] , \SB3_3/i3[0] , \SB3_3/i1_5 , \SB3_3/i1_7 ,
         \SB3_3/i1[9] , \SB3_3/i0_0 , \SB3_3/i0_3 , \SB3_3/i0_4 ,
         \SB3_3/i0[10] , \SB3_3/i0[9] , \SB3_3/i0[8] , \SB3_3/i0[7] ,
         \SB3_3/i0[6] , \SB3_4/i3[0] , \SB3_4/i1_5 , \SB3_4/i1_7 ,
         \SB3_4/i1[9] , \SB3_4/i0_0 , \SB3_4/i0_3 , \SB3_4/i0_4 ,
         \SB3_4/i0[10] , \SB3_4/i0[9] , \SB3_4/i0[8] , \SB3_4/i0[7] ,
         \SB3_4/i0[6] , \SB3_5/i3[0] , \SB3_5/i1_5 , \SB3_5/i1_7 ,
         \SB3_5/i1[9] , \SB3_5/i0_0 , \SB3_5/i0_3 , \SB3_5/i0_4 ,
         \SB3_5/i0[10] , \SB3_5/i0[9] , \SB3_5/i0[8] , \SB3_5/i0[7] ,
         \SB3_5/i0[6] , \SB3_6/i3[0] , \SB3_6/i1_5 , \SB3_6/i1_7 ,
         \SB3_6/i1[9] , \SB3_6/i0_0 , \SB3_6/i0_3 , \SB3_6/i0_4 ,
         \SB3_6/i0[10] , \SB3_6/i0[9] , \SB3_6/i0[8] , \SB3_6/i0[7] ,
         \SB3_6/i0[6] , \SB3_7/i3[0] , \SB3_7/i1_5 , \SB3_7/i1_7 ,
         \SB3_7/i1[9] , \SB3_7/i0_0 , \SB3_7/i0_3 , \SB3_7/i0_4 ,
         \SB3_7/i0[10] , \SB3_7/i0[9] , \SB3_7/i0[7] , \SB3_7/i0[6] ,
         \SB3_8/i3[0] , \SB3_8/i1_5 , \SB3_8/i1_7 , \SB3_8/i1[9] ,
         \SB3_8/i0_0 , \SB3_8/i0_3 , \SB3_8/i0_4 , \SB3_8/i0[10] ,
         \SB3_8/i0[9] , \SB3_8/i0[8] , \SB3_8/i0[7] , \SB3_8/i0[6] ,
         \SB3_9/i3[0] , \SB3_9/i1_5 , \SB3_9/i1_7 , \SB3_9/i1[9] ,
         \SB3_9/i0_0 , \SB3_9/i0_3 , \SB3_9/i0_4 , \SB3_9/i0[10] ,
         \SB3_9/i0[9] , \SB3_9/i0[8] , \SB3_9/i0[7] , \SB3_9/i0[6] ,
         \SB3_10/i3[0] , \SB3_10/i1_5 , \SB3_10/i1_7 , \SB3_10/i1[9] ,
         \SB3_10/i0_0 , \SB3_10/i0_3 , \SB3_10/i0_4 , \SB3_10/i0[10] ,
         \SB3_10/i0[9] , \SB3_10/i0[8] , \SB3_10/i0[7] , \SB3_10/i0[6] ,
         \SB3_11/i3[0] , \SB3_11/i1_5 , \SB3_11/i1_7 , \SB3_11/i1[9] ,
         \SB3_11/i0_0 , \SB3_11/i0_3 , \SB3_11/i0_4 , \SB3_11/i0[10] ,
         \SB3_11/i0[9] , \SB3_11/i0[8] , \SB3_11/i0[7] , \SB3_11/i0[6] ,
         \SB3_12/i3[0] , \SB3_12/i1_5 , \SB3_12/i1_7 , \SB3_12/i1[9] ,
         \SB3_12/i0_0 , \SB3_12/i0_3 , \SB3_12/i0_4 , \SB3_12/i0[10] ,
         \SB3_12/i0[9] , \SB3_12/i0[8] , \SB3_12/i0[7] , \SB3_12/i0[6] ,
         \SB3_13/i3[0] , \SB3_13/i1_5 , \SB3_13/i1_7 , \SB3_13/i1[9] ,
         \SB3_13/i0_0 , \SB3_13/i0_3 , \SB3_13/i0_4 , \SB3_13/i0[10] ,
         \SB3_13/i0[9] , \SB3_13/i0[8] , \SB3_13/i0[7] , \SB3_13/i0[6] ,
         \SB3_14/i3[0] , \SB3_14/i1_5 , \SB3_14/i1_7 , \SB3_14/i1[9] ,
         \SB3_14/i0_0 , \SB3_14/i0_3 , \SB3_14/i0_4 , \SB3_14/i0[10] ,
         \SB3_14/i0[9] , \SB3_14/i0[8] , \SB3_14/i0[7] , \SB3_14/i0[6] ,
         \SB3_15/i3[0] , \SB3_15/i1_5 , \SB3_15/i1_7 , \SB3_15/i1[9] ,
         \SB3_15/i0_0 , \SB3_15/i0_3 , \SB3_15/i0_4 , \SB3_15/i0[10] ,
         \SB3_15/i0[9] , \SB3_15/i0[8] , \SB3_15/i0[7] , \SB3_15/i0[6] ,
         \SB3_16/i3[0] , \SB3_16/i1_5 , \SB3_16/i1_7 , \SB3_16/i1[9] ,
         \SB3_16/i0_0 , \SB3_16/i0_3 , \SB3_16/i0_4 , \SB3_16/i0[10] ,
         \SB3_16/i0[9] , \SB3_16/i0[8] , \SB3_16/i0[7] , \SB3_16/i0[6] ,
         \SB3_17/i3[0] , \SB3_17/i1_5 , \SB3_17/i1_7 , \SB3_17/i1[9] ,
         \SB3_17/i0_0 , \SB3_17/i0_3 , \SB3_17/i0_4 , \SB3_17/i0[10] ,
         \SB3_17/i0[9] , \SB3_17/i0[8] , \SB3_17/i0[7] , \SB3_17/i0[6] ,
         \SB3_18/i3[0] , \SB3_18/i1_5 , \SB3_18/i1_7 , \SB3_18/i1[9] ,
         \SB3_18/i0_0 , \SB3_18/i0_3 , \SB3_18/i0_4 , \SB3_18/i0[10] ,
         \SB3_18/i0[9] , \SB3_18/i0[8] , \SB3_18/i0[7] , \SB3_18/i0[6] ,
         \SB3_19/i3[0] , \SB3_19/i1_5 , \SB3_19/i1_7 , \SB3_19/i1[9] ,
         \SB3_19/i0_0 , \SB3_19/i0_3 , \SB3_19/i0_4 , \SB3_19/i0[10] ,
         \SB3_19/i0[9] , \SB3_19/i0[8] , \SB3_19/i0[7] , \SB3_19/i0[6] ,
         \SB3_20/i3[0] , \SB3_20/i1_5 , \SB3_20/i1_7 , \SB3_20/i1[9] ,
         \SB3_20/i0_0 , \SB3_20/i0_3 , \SB3_20/i0_4 , \SB3_20/i0[10] ,
         \SB3_20/i0[9] , \SB3_20/i0[8] , \SB3_20/i0[7] , \SB3_20/i0[6] ,
         \SB3_21/i3[0] , \SB3_21/i1_5 , \SB3_21/i1_7 , \SB3_21/i1[9] ,
         \SB3_21/i0_0 , \SB3_21/i0_3 , \SB3_21/i0_4 , \SB3_21/i0[10] ,
         \SB3_21/i0[9] , \SB3_21/i0[8] , \SB3_21/i0[7] , \SB3_21/i0[6] ,
         \SB3_22/i3[0] , \SB3_22/i1_5 , \SB3_22/i1_7 , \SB3_22/i1[9] ,
         \SB3_22/i0_0 , \SB3_22/i0_3 , \SB3_22/i0_4 , \SB3_22/i0[10] ,
         \SB3_22/i0[9] , \SB3_22/i0[8] , \SB3_22/i0[7] , \SB3_22/i0[6] ,
         \SB3_23/i3[0] , \SB3_23/i1_5 , \SB3_23/i1_7 , \SB3_23/i1[9] ,
         \SB3_23/i0_0 , \SB3_23/i0_3 , \SB3_23/i0_4 , \SB3_23/i0[10] ,
         \SB3_23/i0[9] , \SB3_23/i0[8] , \SB3_23/i0[7] , \SB3_23/i0[6] ,
         \SB3_24/i3[0] , \SB3_24/i1_5 , \SB3_24/i1_7 , \SB3_24/i1[9] ,
         \SB3_24/i0_0 , \SB3_24/i0_3 , \SB3_24/i0_4 , \SB3_24/i0[10] ,
         \SB3_24/i0[9] , \SB3_24/i0[8] , \SB3_24/i0[7] , \SB3_24/i0[6] ,
         \SB3_25/i3[0] , \SB3_25/i1_5 , \SB3_25/i1_7 , \SB3_25/i1[9] ,
         \SB3_25/i0_0 , \SB3_25/i0_3 , \SB3_25/i0_4 , \SB3_25/i0[10] ,
         \SB3_25/i0[9] , \SB3_25/i0[8] , \SB3_25/i0[7] , \SB3_25/i0[6] ,
         \SB3_26/i3[0] , \SB3_26/i1_5 , \SB3_26/i1_7 , \SB3_26/i1[9] ,
         \SB3_26/i0_0 , \SB3_26/i0_3 , \SB3_26/i0_4 , \SB3_26/i0[10] ,
         \SB3_26/i0[9] , \SB3_26/i0[8] , \SB3_26/i0[7] , \SB3_26/i0[6] ,
         \SB3_27/i3[0] , \SB3_27/i1_5 , \SB3_27/i1_7 , \SB3_27/i1[9] ,
         \SB3_27/i0_0 , \SB3_27/i0_3 , \SB3_27/i0_4 , \SB3_27/i0[10] ,
         \SB3_27/i0[9] , \SB3_27/i0[8] , \SB3_27/i0[7] , \SB3_27/i0[6] ,
         \SB3_28/i3[0] , \SB3_28/i1_5 , \SB3_28/i1_7 , \SB3_28/i1[9] ,
         \SB3_28/i0_0 , \SB3_28/i0_3 , \SB3_28/i0_4 , \SB3_28/i0[10] ,
         \SB3_28/i0[9] , \SB3_28/i0[8] , \SB3_28/i0[7] , \SB3_28/i0[6] ,
         \SB3_29/i3[0] , \SB3_29/i1_5 , \SB3_29/i1_7 , \SB3_29/i1[9] ,
         \SB3_29/i0_0 , \SB3_29/i0_3 , \SB3_29/i0_4 , \SB3_29/i0[10] ,
         \SB3_29/i0[9] , \SB3_29/i0[8] , \SB3_29/i0[7] , \SB3_29/i0[6] ,
         \SB3_30/i3[0] , \SB3_30/i1_5 , \SB3_30/i1_7 , \SB3_30/i1[9] ,
         \SB3_30/i0_0 , \SB3_30/i0_3 , \SB3_30/i0_4 , \SB3_30/i0[10] ,
         \SB3_30/i0[9] , \SB3_30/i0[8] , \SB3_30/i0[7] , \SB3_30/i0[6] ,
         \SB3_31/i3[0] , \SB3_31/i1_5 , \SB3_31/i1_7 , \SB3_31/i1[9] ,
         \SB3_31/i0_0 , \SB3_31/i0_3 , \SB3_31/i0_4 , \SB3_31/i0[10] ,
         \SB3_31/i0[9] , \SB3_31/i0[8] , \SB3_31/i0[7] , \SB3_31/i0[6] ,
         \SB2_0_0/i3[0] , \SB2_0_0/i1_5 , \SB2_0_0/i1_7 , \SB2_0_0/i1[9] ,
         \SB2_0_0/i0_0 , \SB2_0_0/i0_3 , \SB2_0_0/i0_4 , \SB2_0_0/i0[10] ,
         \SB2_0_0/i0[9] , \SB2_0_0/i0[8] , \SB2_0_0/i0[7] , \SB2_0_0/i0[6] ,
         \SB2_0_1/i3[0] , \SB2_0_1/i1_5 , \SB2_0_1/i1_7 , \SB2_0_1/i1[9] ,
         \SB2_0_1/i0_0 , \SB2_0_1/i0_3 , \SB2_0_1/i0_4 , \SB2_0_1/i0[10] ,
         \SB2_0_1/i0[9] , \SB2_0_1/i0[8] , \SB2_0_1/i0[7] , \SB2_0_1/i0[6] ,
         \SB2_0_2/i3[0] , \SB2_0_2/i1_5 , \SB2_0_2/i1_7 , \SB2_0_2/i1[9] ,
         \SB2_0_2/i0_0 , \SB2_0_2/i0_3 , \SB2_0_2/i0_4 , \SB2_0_2/i0[10] ,
         \SB2_0_2/i0[9] , \SB2_0_2/i0[8] , \SB2_0_2/i0[7] , \SB2_0_2/i0[6] ,
         \SB2_0_3/i3[0] , \SB2_0_3/i1_5 , \SB2_0_3/i1_7 , \SB2_0_3/i1[9] ,
         \SB2_0_3/i0_0 , \SB2_0_3/i0_3 , \SB2_0_3/i0_4 , \SB2_0_3/i0[10] ,
         \SB2_0_3/i0[9] , \SB2_0_3/i0[8] , \SB2_0_3/i0[7] , \SB2_0_3/i0[6] ,
         \SB2_0_4/i3[0] , \SB2_0_4/i1_5 , \SB2_0_4/i1_7 , \SB2_0_4/i1[9] ,
         \SB2_0_4/i0_0 , \SB2_0_4/i0_3 , \SB2_0_4/i0_4 , \SB2_0_4/i0[10] ,
         \SB2_0_4/i0[9] , \SB2_0_4/i0[8] , \SB2_0_4/i0[7] , \SB2_0_4/i0[6] ,
         \SB2_0_5/i3[0] , \SB2_0_5/i1_5 , \SB2_0_5/i1_7 , \SB2_0_5/i1[9] ,
         \SB2_0_5/i0_0 , \SB2_0_5/i0_3 , \SB2_0_5/i0_4 , \SB2_0_5/i0[10] ,
         \SB2_0_5/i0[9] , \SB2_0_5/i0[8] , \SB2_0_5/i0[7] , \SB2_0_5/i0[6] ,
         \SB2_0_6/i3[0] , \SB2_0_6/i1_5 , \SB2_0_6/i1_7 , \SB2_0_6/i1[9] ,
         \SB2_0_6/i0_0 , \SB2_0_6/i0_3 , \SB2_0_6/i0_4 , \SB2_0_6/i0[10] ,
         \SB2_0_6/i0[9] , \SB2_0_6/i0[8] , \SB2_0_6/i0[7] , \SB2_0_6/i0[6] ,
         \SB2_0_7/i3[0] , \SB2_0_7/i1_5 , \SB2_0_7/i1_7 , \SB2_0_7/i1[9] ,
         \SB2_0_7/i0_0 , \SB2_0_7/i0_3 , \SB2_0_7/i0_4 , \SB2_0_7/i0[10] ,
         \SB2_0_7/i0[9] , \SB2_0_7/i0[8] , \SB2_0_7/i0[7] , \SB2_0_7/i0[6] ,
         \SB2_0_8/i3[0] , \SB2_0_8/i1_5 , \SB2_0_8/i1_7 , \SB2_0_8/i1[9] ,
         \SB2_0_8/i0_0 , \SB2_0_8/i0_3 , \SB2_0_8/i0_4 , \SB2_0_8/i0[10] ,
         \SB2_0_8/i0[9] , \SB2_0_8/i0[8] , \SB2_0_8/i0[7] , \SB2_0_8/i0[6] ,
         \SB2_0_9/i3[0] , \SB2_0_9/i1_5 , \SB2_0_9/i1_7 , \SB2_0_9/i1[9] ,
         \SB2_0_9/i0_0 , \SB2_0_9/i0_3 , \SB2_0_9/i0_4 , \SB2_0_9/i0[10] ,
         \SB2_0_9/i0[9] , \SB2_0_9/i0[8] , \SB2_0_9/i0[7] , \SB2_0_9/i0[6] ,
         \SB2_0_10/i3[0] , \SB2_0_10/i1_5 , \SB2_0_10/i1_7 , \SB2_0_10/i1[9] ,
         \SB2_0_10/i0_0 , \SB2_0_10/i0_3 , \SB2_0_10/i0_4 , \SB2_0_10/i0[10] ,
         \SB2_0_10/i0[9] , \SB2_0_10/i0[8] , \SB2_0_10/i0[7] ,
         \SB2_0_10/i0[6] , \SB2_0_11/i3[0] , \SB2_0_11/i1_5 , \SB2_0_11/i1_7 ,
         \SB2_0_11/i1[9] , \SB2_0_11/i0_0 , \SB2_0_11/i0_3 , \SB2_0_11/i0_4 ,
         \SB2_0_11/i0[10] , \SB2_0_11/i0[9] , \SB2_0_11/i0[8] ,
         \SB2_0_11/i0[7] , \SB2_0_11/i0[6] , \SB2_0_12/i3[0] , \SB2_0_12/i1_5 ,
         \SB2_0_12/i1_7 , \SB2_0_12/i1[9] , \SB2_0_12/i0_0 , \SB2_0_12/i0_3 ,
         \SB2_0_12/i0_4 , \SB2_0_12/i0[10] , \SB2_0_12/i0[9] ,
         \SB2_0_12/i0[8] , \SB2_0_12/i0[7] , \SB2_0_12/i0[6] ,
         \SB2_0_13/i3[0] , \SB2_0_13/i1_5 , \SB2_0_13/i1_7 , \SB2_0_13/i1[9] ,
         \SB2_0_13/i0_0 , \SB2_0_13/i0_3 , \SB2_0_13/i0_4 , \SB2_0_13/i0[10] ,
         \SB2_0_13/i0[9] , \SB2_0_13/i0[8] , \SB2_0_13/i0[7] ,
         \SB2_0_13/i0[6] , \SB2_0_14/i3[0] , \SB2_0_14/i1_5 , \SB2_0_14/i1_7 ,
         \SB2_0_14/i1[9] , \SB2_0_14/i0_0 , \SB2_0_14/i0_3 , \SB2_0_14/i0_4 ,
         \SB2_0_14/i0[10] , \SB2_0_14/i0[9] , \SB2_0_14/i0[8] ,
         \SB2_0_14/i0[7] , \SB2_0_14/i0[6] , \SB2_0_15/i3[0] , \SB2_0_15/i1_5 ,
         \SB2_0_15/i1_7 , \SB2_0_15/i1[9] , \SB2_0_15/i0_0 , \SB2_0_15/i0_3 ,
         \SB2_0_15/i0_4 , \SB2_0_15/i0[10] , \SB2_0_15/i0[9] ,
         \SB2_0_15/i0[8] , \SB2_0_15/i0[7] , \SB2_0_15/i0[6] ,
         \SB2_0_16/i3[0] , \SB2_0_16/i1_5 , \SB2_0_16/i1_7 , \SB2_0_16/i1[9] ,
         \SB2_0_16/i0_0 , \SB2_0_16/i0_3 , \SB2_0_16/i0_4 , \SB2_0_16/i0[10] ,
         \SB2_0_16/i0[9] , \SB2_0_16/i0[8] , \SB2_0_16/i0[7] ,
         \SB2_0_16/i0[6] , \SB2_0_17/i3[0] , \SB2_0_17/i1_5 , \SB2_0_17/i1_7 ,
         \SB2_0_17/i1[9] , \SB2_0_17/i0_0 , \SB2_0_17/i0_3 , \SB2_0_17/i0_4 ,
         \SB2_0_17/i0[10] , \SB2_0_17/i0[9] , \SB2_0_17/i0[8] ,
         \SB2_0_17/i0[7] , \SB2_0_17/i0[6] , \SB2_0_18/i3[0] , \SB2_0_18/i1_5 ,
         \SB2_0_18/i1_7 , \SB2_0_18/i1[9] , \SB2_0_18/i0_0 , \SB2_0_18/i0_3 ,
         \SB2_0_18/i0_4 , \SB2_0_18/i0[10] , \SB2_0_18/i0[9] ,
         \SB2_0_18/i0[8] , \SB2_0_18/i0[7] , \SB2_0_18/i0[6] ,
         \SB2_0_19/i3[0] , \SB2_0_19/i1_5 , \SB2_0_19/i1_7 , \SB2_0_19/i1[9] ,
         \SB2_0_19/i0_0 , \SB2_0_19/i0_3 , \SB2_0_19/i0_4 , \SB2_0_19/i0[10] ,
         \SB2_0_19/i0[9] , \SB2_0_19/i0[8] , \SB2_0_19/i0[7] ,
         \SB2_0_19/i0[6] , \SB2_0_20/i3[0] , \SB2_0_20/i1_5 , \SB2_0_20/i1_7 ,
         \SB2_0_20/i1[9] , \SB2_0_20/i0_0 , \SB2_0_20/i0_3 , \SB2_0_20/i0_4 ,
         \SB2_0_20/i0[10] , \SB2_0_20/i0[9] , \SB2_0_20/i0[8] ,
         \SB2_0_20/i0[7] , \SB2_0_20/i0[6] , \SB2_0_21/i3[0] , \SB2_0_21/i1_5 ,
         \SB2_0_21/i1_7 , \SB2_0_21/i1[9] , \SB2_0_21/i0_0 , \SB2_0_21/i0_3 ,
         \SB2_0_21/i0_4 , \SB2_0_21/i0[10] , \SB2_0_21/i0[9] ,
         \SB2_0_21/i0[8] , \SB2_0_21/i0[7] , \SB2_0_21/i0[6] ,
         \SB2_0_22/i3[0] , \SB2_0_22/i1_5 , \SB2_0_22/i1_7 , \SB2_0_22/i1[9] ,
         \SB2_0_22/i0_0 , \SB2_0_22/i0_3 , \SB2_0_22/i0_4 , \SB2_0_22/i0[10] ,
         \SB2_0_22/i0[9] , \SB2_0_22/i0[8] , \SB2_0_22/i0[7] ,
         \SB2_0_22/i0[6] , \SB2_0_23/i3[0] , \SB2_0_23/i1_5 , \SB2_0_23/i1_7 ,
         \SB2_0_23/i1[9] , \SB2_0_23/i0_0 , \SB2_0_23/i0_3 , \SB2_0_23/i0_4 ,
         \SB2_0_23/i0[10] , \SB2_0_23/i0[9] , \SB2_0_23/i0[8] ,
         \SB2_0_23/i0[7] , \SB2_0_23/i0[6] , \SB2_0_24/i3[0] , \SB2_0_24/i1_5 ,
         \SB2_0_24/i1_7 , \SB2_0_24/i1[9] , \SB2_0_24/i0_0 , \SB2_0_24/i0_3 ,
         \SB2_0_24/i0_4 , \SB2_0_24/i0[10] , \SB2_0_24/i0[9] ,
         \SB2_0_24/i0[8] , \SB2_0_24/i0[7] , \SB2_0_24/i0[6] ,
         \SB2_0_25/i3[0] , \SB2_0_25/i1_5 , \SB2_0_25/i1_7 , \SB2_0_25/i1[9] ,
         \SB2_0_25/i0_0 , \SB2_0_25/i0_3 , \SB2_0_25/i0_4 , \SB2_0_25/i0[10] ,
         \SB2_0_25/i0[9] , \SB2_0_25/i0[8] , \SB2_0_25/i0[7] ,
         \SB2_0_25/i0[6] , \SB2_0_26/i3[0] , \SB2_0_26/i1_5 , \SB2_0_26/i1_7 ,
         \SB2_0_26/i1[9] , \SB2_0_26/i0_0 , \SB2_0_26/i0_3 , \SB2_0_26/i0_4 ,
         \SB2_0_26/i0[10] , \SB2_0_26/i0[8] , \SB2_0_26/i0[7] ,
         \SB2_0_26/i0[6] , \SB2_0_27/i3[0] , \SB2_0_27/i1_5 , \SB2_0_27/i1_7 ,
         \SB2_0_27/i1[9] , \SB2_0_27/i0_0 , \SB2_0_27/i0_3 , \SB2_0_27/i0_4 ,
         \SB2_0_27/i0[10] , \SB2_0_27/i0[9] , \SB2_0_27/i0[8] ,
         \SB2_0_27/i0[7] , \SB2_0_27/i0[6] , \SB2_0_28/i3[0] , \SB2_0_28/i1_5 ,
         \SB2_0_28/i1_7 , \SB2_0_28/i1[9] , \SB2_0_28/i0_0 , \SB2_0_28/i0_3 ,
         \SB2_0_28/i0_4 , \SB2_0_28/i0[10] , \SB2_0_28/i0[9] ,
         \SB2_0_28/i0[8] , \SB2_0_28/i0[7] , \SB2_0_28/i0[6] ,
         \SB2_0_29/i3[0] , \SB2_0_29/i1_5 , \SB2_0_29/i1_7 , \SB2_0_29/i1[9] ,
         \SB2_0_29/i0_0 , \SB2_0_29/i0_3 , \SB2_0_29/i0_4 , \SB2_0_29/i0[10] ,
         \SB2_0_29/i0[9] , \SB2_0_29/i0[8] , \SB2_0_29/i0[7] ,
         \SB2_0_29/i0[6] , \SB2_0_30/i3[0] , \SB2_0_30/i1_5 , \SB2_0_30/i1_7 ,
         \SB2_0_30/i1[9] , \SB2_0_30/i0_0 , \SB2_0_30/i0_3 , \SB2_0_30/i0_4 ,
         \SB2_0_30/i0[10] , \SB2_0_30/i0[9] , \SB2_0_30/i0[8] ,
         \SB2_0_30/i0[7] , \SB2_0_30/i0[6] , \SB2_0_31/i3[0] , \SB2_0_31/i1_5 ,
         \SB2_0_31/i1_7 , \SB2_0_31/i1[9] , \SB2_0_31/i0_0 , \SB2_0_31/i0_3 ,
         \SB2_0_31/i0_4 , \SB2_0_31/i0[10] , \SB2_0_31/i0[9] ,
         \SB2_0_31/i0[8] , \SB2_0_31/i0[7] , \SB2_0_31/i0[6] , \SB2_1_0/i3[0] ,
         \SB2_1_0/i1_5 , \SB2_1_0/i1_7 , \SB2_1_0/i1[9] , \SB2_1_0/i0_0 ,
         \SB2_1_0/i0_3 , \SB2_1_0/i0_4 , \SB2_1_0/i0[10] , \SB2_1_0/i0[9] ,
         \SB2_1_0/i0[8] , \SB2_1_0/i0[7] , \SB2_1_0/i0[6] , \SB2_1_1/i3[0] ,
         \SB2_1_1/i1_5 , \SB2_1_1/i1_7 , \SB2_1_1/i1[9] , \SB2_1_1/i0_0 ,
         \SB2_1_1/i0_3 , \SB2_1_1/i0_4 , \SB2_1_1/i0[10] , \SB2_1_1/i0[9] ,
         \SB2_1_1/i0[8] , \SB2_1_1/i0[7] , \SB2_1_1/i0[6] , \SB2_1_2/i3[0] ,
         \SB2_1_2/i1_5 , \SB2_1_2/i1_7 , \SB2_1_2/i1[9] , \SB2_1_2/i0_0 ,
         \SB2_1_2/i0_3 , \SB2_1_2/i0_4 , \SB2_1_2/i0[10] , \SB2_1_2/i0[9] ,
         \SB2_1_2/i0[8] , \SB2_1_2/i0[7] , \SB2_1_2/i0[6] , \SB2_1_3/i3[0] ,
         \SB2_1_3/i1_5 , \SB2_1_3/i1_7 , \SB2_1_3/i1[9] , \SB2_1_3/i0_0 ,
         \SB2_1_3/i0_3 , \SB2_1_3/i0_4 , \SB2_1_3/i0[10] , \SB2_1_3/i0[9] ,
         \SB2_1_3/i0[8] , \SB2_1_3/i0[7] , \SB2_1_3/i0[6] , \SB2_1_4/i3[0] ,
         \SB2_1_4/i1_5 , \SB2_1_4/i1_7 , \SB2_1_4/i1[9] , \SB2_1_4/i0_0 ,
         \SB2_1_4/i0_3 , \SB2_1_4/i0_4 , \SB2_1_4/i0[10] , \SB2_1_4/i0[9] ,
         \SB2_1_4/i0[8] , \SB2_1_4/i0[7] , \SB2_1_4/i0[6] , \SB2_1_5/i3[0] ,
         \SB2_1_5/i1_5 , \SB2_1_5/i1_7 , \SB2_1_5/i1[9] , \SB2_1_5/i0_0 ,
         \SB2_1_5/i0_3 , \SB2_1_5/i0_4 , \SB2_1_5/i0[10] , \SB2_1_5/i0[9] ,
         \SB2_1_5/i0[8] , \SB2_1_5/i0[7] , \SB2_1_5/i0[6] , \SB2_1_6/i3[0] ,
         \SB2_1_6/i1_5 , \SB2_1_6/i1_7 , \SB2_1_6/i1[9] , \SB2_1_6/i0_0 ,
         \SB2_1_6/i0_3 , \SB2_1_6/i0_4 , \SB2_1_6/i0[10] , \SB2_1_6/i0[9] ,
         \SB2_1_6/i0[8] , \SB2_1_6/i0[7] , \SB2_1_6/i0[6] , \SB2_1_7/i3[0] ,
         \SB2_1_7/i1_5 , \SB2_1_7/i1_7 , \SB2_1_7/i1[9] , \SB2_1_7/i0_0 ,
         \SB2_1_7/i0_3 , \SB2_1_7/i0_4 , \SB2_1_7/i0[10] , \SB2_1_7/i0[9] ,
         \SB2_1_7/i0[8] , \SB2_1_7/i0[7] , \SB2_1_7/i0[6] , \SB2_1_8/i3[0] ,
         \SB2_1_8/i1_5 , \SB2_1_8/i1_7 , \SB2_1_8/i1[9] , \SB2_1_8/i0_0 ,
         \SB2_1_8/i0_3 , \SB2_1_8/i0_4 , \SB2_1_8/i0[10] , \SB2_1_8/i0[9] ,
         \SB2_1_8/i0[8] , \SB2_1_8/i0[7] , \SB2_1_8/i0[6] , \SB2_1_9/i3[0] ,
         \SB2_1_9/i1_5 , \SB2_1_9/i1_7 , \SB2_1_9/i1[9] , \SB2_1_9/i0_0 ,
         \SB2_1_9/i0_3 , \SB2_1_9/i0_4 , \SB2_1_9/i0[10] , \SB2_1_9/i0[9] ,
         \SB2_1_9/i0[8] , \SB2_1_9/i0[7] , \SB2_1_9/i0[6] , \SB2_1_10/i3[0] ,
         \SB2_1_10/i1_5 , \SB2_1_10/i1_7 , \SB2_1_10/i1[9] , \SB2_1_10/i0_0 ,
         \SB2_1_10/i0_3 , \SB2_1_10/i0_4 , \SB2_1_10/i0[10] , \SB2_1_10/i0[9] ,
         \SB2_1_10/i0[8] , \SB2_1_10/i0[7] , \SB2_1_10/i0[6] ,
         \SB2_1_11/i3[0] , \SB2_1_11/i1_5 , \SB2_1_11/i1_7 , \SB2_1_11/i1[9] ,
         \SB2_1_11/i0_0 , \SB2_1_11/i0_3 , \SB2_1_11/i0_4 , \SB2_1_11/i0[10] ,
         \SB2_1_11/i0[9] , \SB2_1_11/i0[8] , \SB2_1_11/i0[7] ,
         \SB2_1_11/i0[6] , \SB2_1_12/i3[0] , \SB2_1_12/i1_5 , \SB2_1_12/i1_7 ,
         \SB2_1_12/i1[9] , \SB2_1_12/i0_0 , \SB2_1_12/i0_3 , \SB2_1_12/i0_4 ,
         \SB2_1_12/i0[10] , \SB2_1_12/i0[9] , \SB2_1_12/i0[8] ,
         \SB2_1_12/i0[7] , \SB2_1_12/i0[6] , \SB2_1_13/i3[0] , \SB2_1_13/i1_5 ,
         \SB2_1_13/i1_7 , \SB2_1_13/i1[9] , \SB2_1_13/i0_0 , \SB2_1_13/i0_3 ,
         \SB2_1_13/i0_4 , \SB2_1_13/i0[10] , \SB2_1_13/i0[9] ,
         \SB2_1_13/i0[8] , \SB2_1_13/i0[7] , \SB2_1_13/i0[6] ,
         \SB2_1_14/i3[0] , \SB2_1_14/i1_5 , \SB2_1_14/i1_7 , \SB2_1_14/i1[9] ,
         \SB2_1_14/i0_0 , \SB2_1_14/i0_3 , \SB2_1_14/i0_4 , \SB2_1_14/i0[10] ,
         \SB2_1_14/i0[9] , \SB2_1_14/i0[8] , \SB2_1_14/i0[7] ,
         \SB2_1_14/i0[6] , \SB2_1_15/i3[0] , \SB2_1_15/i1_5 , \SB2_1_15/i1_7 ,
         \SB2_1_15/i1[9] , \SB2_1_15/i0_0 , \SB2_1_15/i0_3 , \SB2_1_15/i0_4 ,
         \SB2_1_15/i0[10] , \SB2_1_15/i0[9] , \SB2_1_15/i0[8] ,
         \SB2_1_15/i0[7] , \SB2_1_15/i0[6] , \SB2_1_16/i3[0] , \SB2_1_16/i1_5 ,
         \SB2_1_16/i1_7 , \SB2_1_16/i1[9] , \SB2_1_16/i0_0 , \SB2_1_16/i0_3 ,
         \SB2_1_16/i0_4 , \SB2_1_16/i0[10] , \SB2_1_16/i0[9] ,
         \SB2_1_16/i0[8] , \SB2_1_16/i0[7] , \SB2_1_16/i0[6] ,
         \SB2_1_17/i3[0] , \SB2_1_17/i1_5 , \SB2_1_17/i1_7 , \SB2_1_17/i1[9] ,
         \SB2_1_17/i0_0 , \SB2_1_17/i0_3 , \SB2_1_17/i0_4 , \SB2_1_17/i0[10] ,
         \SB2_1_17/i0[9] , \SB2_1_17/i0[8] , \SB2_1_17/i0[7] ,
         \SB2_1_17/i0[6] , \SB2_1_18/i3[0] , \SB2_1_18/i1_5 , \SB2_1_18/i1_7 ,
         \SB2_1_18/i1[9] , \SB2_1_18/i0_0 , \SB2_1_18/i0_3 , \SB2_1_18/i0_4 ,
         \SB2_1_18/i0[10] , \SB2_1_18/i0[9] , \SB2_1_18/i0[8] ,
         \SB2_1_18/i0[7] , \SB2_1_18/i0[6] , \SB2_1_19/i3[0] , \SB2_1_19/i1_5 ,
         \SB2_1_19/i1_7 , \SB2_1_19/i1[9] , \SB2_1_19/i0_0 , \SB2_1_19/i0_3 ,
         \SB2_1_19/i0_4 , \SB2_1_19/i0[10] , \SB2_1_19/i0[9] ,
         \SB2_1_19/i0[8] , \SB2_1_19/i0[7] , \SB2_1_19/i0[6] ,
         \SB2_1_20/i3[0] , \SB2_1_20/i1_5 , \SB2_1_20/i1_7 , \SB2_1_20/i1[9] ,
         \SB2_1_20/i0_0 , \SB2_1_20/i0_3 , \SB2_1_20/i0_4 , \SB2_1_20/i0[10] ,
         \SB2_1_20/i0[9] , \SB2_1_20/i0[8] , \SB2_1_20/i0[7] ,
         \SB2_1_20/i0[6] , \SB2_1_21/i3[0] , \SB2_1_21/i1_5 , \SB2_1_21/i1_7 ,
         \SB2_1_21/i1[9] , \SB2_1_21/i0_0 , \SB2_1_21/i0_3 , \SB2_1_21/i0_4 ,
         \SB2_1_21/i0[10] , \SB2_1_21/i0[9] , \SB2_1_21/i0[8] ,
         \SB2_1_21/i0[7] , \SB2_1_21/i0[6] , \SB2_1_22/i3[0] , \SB2_1_22/i1_5 ,
         \SB2_1_22/i1_7 , \SB2_1_22/i1[9] , \SB2_1_22/i0_0 , \SB2_1_22/i0_3 ,
         \SB2_1_22/i0_4 , \SB2_1_22/i0[10] , \SB2_1_22/i0[9] ,
         \SB2_1_22/i0[8] , \SB2_1_22/i0[7] , \SB2_1_22/i0[6] ,
         \SB2_1_23/i3[0] , \SB2_1_23/i1_5 , \SB2_1_23/i1_7 , \SB2_1_23/i1[9] ,
         \SB2_1_23/i0_0 , \SB2_1_23/i0_3 , \SB2_1_23/i0_4 , \SB2_1_23/i0[10] ,
         \SB2_1_23/i0[9] , \SB2_1_23/i0[8] , \SB2_1_23/i0[7] ,
         \SB2_1_23/i0[6] , \SB2_1_24/i3[0] , \SB2_1_24/i1_5 , \SB2_1_24/i1_7 ,
         \SB2_1_24/i1[9] , \SB2_1_24/i0_0 , \SB2_1_24/i0_3 , \SB2_1_24/i0_4 ,
         \SB2_1_24/i0[10] , \SB2_1_24/i0[9] , \SB2_1_24/i0[8] ,
         \SB2_1_24/i0[7] , \SB2_1_24/i0[6] , \SB2_1_25/i3[0] , \SB2_1_25/i1_5 ,
         \SB2_1_25/i1_7 , \SB2_1_25/i1[9] , \SB2_1_25/i0_0 , \SB2_1_25/i0_3 ,
         \SB2_1_25/i0_4 , \SB2_1_25/i0[10] , \SB2_1_25/i0[9] ,
         \SB2_1_25/i0[8] , \SB2_1_25/i0[7] , \SB2_1_25/i0[6] ,
         \SB2_1_26/i3[0] , \SB2_1_26/i1_5 , \SB2_1_26/i1_7 , \SB2_1_26/i1[9] ,
         \SB2_1_26/i0_0 , \SB2_1_26/i0_3 , \SB2_1_26/i0_4 , \SB2_1_26/i0[10] ,
         \SB2_1_26/i0[9] , \SB2_1_26/i0[8] , \SB2_1_26/i0[7] ,
         \SB2_1_26/i0[6] , \SB2_1_27/i3[0] , \SB2_1_27/i1_5 , \SB2_1_27/i1_7 ,
         \SB2_1_27/i1[9] , \SB2_1_27/i0_0 , \SB2_1_27/i0_3 , \SB2_1_27/i0_4 ,
         \SB2_1_27/i0[10] , \SB2_1_27/i0[9] , \SB2_1_27/i0[8] ,
         \SB2_1_27/i0[7] , \SB2_1_27/i0[6] , \SB2_1_28/i3[0] , \SB2_1_28/i1_5 ,
         \SB2_1_28/i1_7 , \SB2_1_28/i1[9] , \SB2_1_28/i0_0 , \SB2_1_28/i0_3 ,
         \SB2_1_28/i0_4 , \SB2_1_28/i0[10] , \SB2_1_28/i0[9] ,
         \SB2_1_28/i0[8] , \SB2_1_28/i0[7] , \SB2_1_28/i0[6] ,
         \SB2_1_29/i3[0] , \SB2_1_29/i1_5 , \SB2_1_29/i1_7 , \SB2_1_29/i1[9] ,
         \SB2_1_29/i0_0 , \SB2_1_29/i0_3 , \SB2_1_29/i0_4 , \SB2_1_29/i0[10] ,
         \SB2_1_29/i0[9] , \SB2_1_29/i0[8] , \SB2_1_29/i0[7] ,
         \SB2_1_29/i0[6] , \SB2_1_30/i3[0] , \SB2_1_30/i1_5 , \SB2_1_30/i1_7 ,
         \SB2_1_30/i1[9] , \SB2_1_30/i0_0 , \SB2_1_30/i0_3 , \SB2_1_30/i0_4 ,
         \SB2_1_30/i0[10] , \SB2_1_30/i0[9] , \SB2_1_30/i0[8] ,
         \SB2_1_30/i0[7] , \SB2_1_30/i0[6] , \SB2_1_31/i3[0] , \SB2_1_31/i1_5 ,
         \SB2_1_31/i1_7 , \SB2_1_31/i1[9] , \SB2_1_31/i0_0 , \SB2_1_31/i0_3 ,
         \SB2_1_31/i0_4 , \SB2_1_31/i0[10] , \SB2_1_31/i0[9] ,
         \SB2_1_31/i0[8] , \SB2_1_31/i0[7] , \SB2_1_31/i0[6] , \SB2_2_0/i3[0] ,
         \SB2_2_0/i1_5 , \SB2_2_0/i1_7 , \SB2_2_0/i1[9] , \SB2_2_0/i0_0 ,
         \SB2_2_0/i0_3 , \SB2_2_0/i0_4 , \SB2_2_0/i0[10] , \SB2_2_0/i0[9] ,
         \SB2_2_0/i0[8] , \SB2_2_0/i0[7] , \SB2_2_0/i0[6] , \SB2_2_1/i3[0] ,
         \SB2_2_1/i1_5 , \SB2_2_1/i1_7 , \SB2_2_1/i1[9] , \SB2_2_1/i0_0 ,
         \SB2_2_1/i0_3 , \SB2_2_1/i0_4 , \SB2_2_1/i0[10] , \SB2_2_1/i0[9] ,
         \SB2_2_1/i0[8] , \SB2_2_1/i0[7] , \SB2_2_1/i0[6] , \SB2_2_2/i3[0] ,
         \SB2_2_2/i1_5 , \SB2_2_2/i1_7 , \SB2_2_2/i1[9] , \SB2_2_2/i0_0 ,
         \SB2_2_2/i0_3 , \SB2_2_2/i0_4 , \SB2_2_2/i0[10] , \SB2_2_2/i0[9] ,
         \SB2_2_2/i0[8] , \SB2_2_2/i0[7] , \SB2_2_2/i0[6] , \SB2_2_3/i3[0] ,
         \SB2_2_3/i1_5 , \SB2_2_3/i1_7 , \SB2_2_3/i1[9] , \SB2_2_3/i0_0 ,
         \SB2_2_3/i0_3 , \SB2_2_3/i0_4 , \SB2_2_3/i0[10] , \SB2_2_3/i0[9] ,
         \SB2_2_3/i0[8] , \SB2_2_3/i0[7] , \SB2_2_3/i0[6] , \SB2_2_4/i3[0] ,
         \SB2_2_4/i1_5 , \SB2_2_4/i1_7 , \SB2_2_4/i1[9] , \SB2_2_4/i0_0 ,
         \SB2_2_4/i0_3 , \SB2_2_4/i0_4 , \SB2_2_4/i0[10] , \SB2_2_4/i0[9] ,
         \SB2_2_4/i0[8] , \SB2_2_4/i0[7] , \SB2_2_4/i0[6] , \SB2_2_5/i3[0] ,
         \SB2_2_5/i1_5 , \SB2_2_5/i1_7 , \SB2_2_5/i1[9] , \SB2_2_5/i0_0 ,
         \SB2_2_5/i0_3 , \SB2_2_5/i0_4 , \SB2_2_5/i0[10] , \SB2_2_5/i0[9] ,
         \SB2_2_5/i0[8] , \SB2_2_5/i0[7] , \SB2_2_5/i0[6] , \SB2_2_6/i3[0] ,
         \SB2_2_6/i1_5 , \SB2_2_6/i1_7 , \SB2_2_6/i1[9] , \SB2_2_6/i0_0 ,
         \SB2_2_6/i0_3 , \SB2_2_6/i0_4 , \SB2_2_6/i0[10] , \SB2_2_6/i0[9] ,
         \SB2_2_6/i0[8] , \SB2_2_6/i0[7] , \SB2_2_6/i0[6] , \SB2_2_7/i3[0] ,
         \SB2_2_7/i1_5 , \SB2_2_7/i1_7 , \SB2_2_7/i1[9] , \SB2_2_7/i0_0 ,
         \SB2_2_7/i0_3 , \SB2_2_7/i0_4 , \SB2_2_7/i0[10] , \SB2_2_7/i0[9] ,
         \SB2_2_7/i0[8] , \SB2_2_7/i0[7] , \SB2_2_7/i0[6] , \SB2_2_8/i3[0] ,
         \SB2_2_8/i1_5 , \SB2_2_8/i1_7 , \SB2_2_8/i1[9] , \SB2_2_8/i0_0 ,
         \SB2_2_8/i0_3 , \SB2_2_8/i0_4 , \SB2_2_8/i0[10] , \SB2_2_8/i0[9] ,
         \SB2_2_8/i0[8] , \SB2_2_8/i0[7] , \SB2_2_8/i0[6] , \SB2_2_9/i3[0] ,
         \SB2_2_9/i1_5 , \SB2_2_9/i1_7 , \SB2_2_9/i1[9] , \SB2_2_9/i0_0 ,
         \SB2_2_9/i0_3 , \SB2_2_9/i0_4 , \SB2_2_9/i0[10] , \SB2_2_9/i0[9] ,
         \SB2_2_9/i0[8] , \SB2_2_9/i0[7] , \SB2_2_9/i0[6] , \SB2_2_10/i3[0] ,
         \SB2_2_10/i1_5 , \SB2_2_10/i1_7 , \SB2_2_10/i1[9] , \SB2_2_10/i0_0 ,
         \SB2_2_10/i0_3 , \SB2_2_10/i0_4 , \SB2_2_10/i0[10] , \SB2_2_10/i0[9] ,
         \SB2_2_10/i0[8] , \SB2_2_10/i0[7] , \SB2_2_10/i0[6] ,
         \SB2_2_11/i3[0] , \SB2_2_11/i1_5 , \SB2_2_11/i1_7 , \SB2_2_11/i1[9] ,
         \SB2_2_11/i0_0 , \SB2_2_11/i0_3 , \SB2_2_11/i0_4 , \SB2_2_11/i0[10] ,
         \SB2_2_11/i0[9] , \SB2_2_11/i0[8] , \SB2_2_11/i0[7] ,
         \SB2_2_11/i0[6] , \SB2_2_12/i3[0] , \SB2_2_12/i1_5 , \SB2_2_12/i1_7 ,
         \SB2_2_12/i1[9] , \SB2_2_12/i0_0 , \SB2_2_12/i0_3 , \SB2_2_12/i0_4 ,
         \SB2_2_12/i0[10] , \SB2_2_12/i0[9] , \SB2_2_12/i0[8] ,
         \SB2_2_12/i0[7] , \SB2_2_12/i0[6] , \SB2_2_13/i3[0] , \SB2_2_13/i1_5 ,
         \SB2_2_13/i1_7 , \SB2_2_13/i1[9] , \SB2_2_13/i0_0 , \SB2_2_13/i0_3 ,
         \SB2_2_13/i0_4 , \SB2_2_13/i0[10] , \SB2_2_13/i0[9] ,
         \SB2_2_13/i0[8] , \SB2_2_13/i0[7] , \SB2_2_13/i0[6] ,
         \SB2_2_14/i3[0] , \SB2_2_14/i1_5 , \SB2_2_14/i1_7 , \SB2_2_14/i1[9] ,
         \SB2_2_14/i0_0 , \SB2_2_14/i0_3 , \SB2_2_14/i0_4 , \SB2_2_14/i0[10] ,
         \SB2_2_14/i0[9] , \SB2_2_14/i0[8] , \SB2_2_14/i0[7] ,
         \SB2_2_14/i0[6] , \SB2_2_15/i3[0] , \SB2_2_15/i1_5 , \SB2_2_15/i1_7 ,
         \SB2_2_15/i1[9] , \SB2_2_15/i0_0 , \SB2_2_15/i0_3 , \SB2_2_15/i0_4 ,
         \SB2_2_15/i0[10] , \SB2_2_15/i0[9] , \SB2_2_15/i0[8] ,
         \SB2_2_15/i0[7] , \SB2_2_15/i0[6] , \SB2_2_16/i3[0] , \SB2_2_16/i1_5 ,
         \SB2_2_16/i1_7 , \SB2_2_16/i1[9] , \SB2_2_16/i0_0 , \SB2_2_16/i0_3 ,
         \SB2_2_16/i0_4 , \SB2_2_16/i0[10] , \SB2_2_16/i0[9] ,
         \SB2_2_16/i0[8] , \SB2_2_16/i0[7] , \SB2_2_16/i0[6] ,
         \SB2_2_17/i3[0] , \SB2_2_17/i1_5 , \SB2_2_17/i1_7 , \SB2_2_17/i1[9] ,
         \SB2_2_17/i0_0 , \SB2_2_17/i0_3 , \SB2_2_17/i0_4 , \SB2_2_17/i0[10] ,
         \SB2_2_17/i0[9] , \SB2_2_17/i0[8] , \SB2_2_17/i0[7] ,
         \SB2_2_17/i0[6] , \SB2_2_18/i3[0] , \SB2_2_18/i1_5 , \SB2_2_18/i1_7 ,
         \SB2_2_18/i1[9] , \SB2_2_18/i0_0 , \SB2_2_18/i0_3 , \SB2_2_18/i0_4 ,
         \SB2_2_18/i0[10] , \SB2_2_18/i0[9] , \SB2_2_18/i0[8] ,
         \SB2_2_18/i0[7] , \SB2_2_18/i0[6] , \SB2_2_19/i3[0] , \SB2_2_19/i1_5 ,
         \SB2_2_19/i1_7 , \SB2_2_19/i1[9] , \SB2_2_19/i0_0 , \SB2_2_19/i0_3 ,
         \SB2_2_19/i0_4 , \SB2_2_19/i0[10] , \SB2_2_19/i0[9] ,
         \SB2_2_19/i0[8] , \SB2_2_19/i0[7] , \SB2_2_19/i0[6] ,
         \SB2_2_20/i3[0] , \SB2_2_20/i1_5 , \SB2_2_20/i1_7 , \SB2_2_20/i1[9] ,
         \SB2_2_20/i0_0 , \SB2_2_20/i0_3 , \SB2_2_20/i0_4 , \SB2_2_20/i0[10] ,
         \SB2_2_20/i0[9] , \SB2_2_20/i0[8] , \SB2_2_20/i0[7] ,
         \SB2_2_20/i0[6] , \SB2_2_21/i3[0] , \SB2_2_21/i1_5 , \SB2_2_21/i1_7 ,
         \SB2_2_21/i1[9] , \SB2_2_21/i0_0 , \SB2_2_21/i0_3 , \SB2_2_21/i0_4 ,
         \SB2_2_21/i0[10] , \SB2_2_21/i0[9] , \SB2_2_21/i0[8] ,
         \SB2_2_21/i0[7] , \SB2_2_21/i0[6] , \SB2_2_22/i3[0] , \SB2_2_22/i1_5 ,
         \SB2_2_22/i1_7 , \SB2_2_22/i1[9] , \SB2_2_22/i0_0 , \SB2_2_22/i0_3 ,
         \SB2_2_22/i0_4 , \SB2_2_22/i0[10] , \SB2_2_22/i0[9] ,
         \SB2_2_22/i0[8] , \SB2_2_22/i0[7] , \SB2_2_22/i0[6] ,
         \SB2_2_23/i3[0] , \SB2_2_23/i1_5 , \SB2_2_23/i1_7 , \SB2_2_23/i1[9] ,
         \SB2_2_23/i0_0 , \SB2_2_23/i0_3 , \SB2_2_23/i0_4 , \SB2_2_23/i0[10] ,
         \SB2_2_23/i0[9] , \SB2_2_23/i0[8] , \SB2_2_23/i0[7] ,
         \SB2_2_23/i0[6] , \SB2_2_24/i3[0] , \SB2_2_24/i1_5 , \SB2_2_24/i1_7 ,
         \SB2_2_24/i1[9] , \SB2_2_24/i0_0 , \SB2_2_24/i0_3 , \SB2_2_24/i0_4 ,
         \SB2_2_24/i0[10] , \SB2_2_24/i0[9] , \SB2_2_24/i0[8] ,
         \SB2_2_24/i0[7] , \SB2_2_24/i0[6] , \SB2_2_25/i3[0] , \SB2_2_25/i1_5 ,
         \SB2_2_25/i1_7 , \SB2_2_25/i1[9] , \SB2_2_25/i0_0 , \SB2_2_25/i0_3 ,
         \SB2_2_25/i0_4 , \SB2_2_25/i0[10] , \SB2_2_25/i0[9] ,
         \SB2_2_25/i0[8] , \SB2_2_25/i0[7] , \SB2_2_25/i0[6] ,
         \SB2_2_26/i3[0] , \SB2_2_26/i1_5 , \SB2_2_26/i1_7 , \SB2_2_26/i1[9] ,
         \SB2_2_26/i0_0 , \SB2_2_26/i0_3 , \SB2_2_26/i0_4 , \SB2_2_26/i0[10] ,
         \SB2_2_26/i0[9] , \SB2_2_26/i0[8] , \SB2_2_26/i0[7] ,
         \SB2_2_26/i0[6] , \SB2_2_27/i3[0] , \SB2_2_27/i1_5 , \SB2_2_27/i1_7 ,
         \SB2_2_27/i1[9] , \SB2_2_27/i0_0 , \SB2_2_27/i0_3 , \SB2_2_27/i0_4 ,
         \SB2_2_27/i0[10] , \SB2_2_27/i0[9] , \SB2_2_27/i0[8] ,
         \SB2_2_27/i0[7] , \SB2_2_27/i0[6] , \SB2_2_28/i3[0] , \SB2_2_28/i1_5 ,
         \SB2_2_28/i1_7 , \SB2_2_28/i1[9] , \SB2_2_28/i0_0 , \SB2_2_28/i0_3 ,
         \SB2_2_28/i0_4 , \SB2_2_28/i0[10] , \SB2_2_28/i0[9] ,
         \SB2_2_28/i0[8] , \SB2_2_28/i0[7] , \SB2_2_28/i0[6] ,
         \SB2_2_29/i3[0] , \SB2_2_29/i1_5 , \SB2_2_29/i1_7 , \SB2_2_29/i1[9] ,
         \SB2_2_29/i0_0 , \SB2_2_29/i0_3 , \SB2_2_29/i0_4 , \SB2_2_29/i0[10] ,
         \SB2_2_29/i0[9] , \SB2_2_29/i0[8] , \SB2_2_29/i0[7] ,
         \SB2_2_29/i0[6] , \SB2_2_30/i3[0] , \SB2_2_30/i1_5 , \SB2_2_30/i1_7 ,
         \SB2_2_30/i0_0 , \SB2_2_30/i0_3 , \SB2_2_30/i0_4 , \SB2_2_30/i0[10] ,
         \SB2_2_30/i0[9] , \SB2_2_30/i0[8] , \SB2_2_30/i0[7] ,
         \SB2_2_30/i0[6] , \SB2_2_31/i3[0] , \SB2_2_31/i1_5 , \SB2_2_31/i1_7 ,
         \SB2_2_31/i1[9] , \SB2_2_31/i0_0 , \SB2_2_31/i0_3 , \SB2_2_31/i0_4 ,
         \SB2_2_31/i0[10] , \SB2_2_31/i0[9] , \SB2_2_31/i0[8] ,
         \SB2_2_31/i0[7] , \SB2_2_31/i0[6] , \SB2_3_0/i3[0] , \SB2_3_0/i1_5 ,
         \SB2_3_0/i1_7 , \SB2_3_0/i1[9] , \SB2_3_0/i0_0 , \SB2_3_0/i0_3 ,
         \SB2_3_0/i0_4 , \SB2_3_0/i0[10] , \SB2_3_0/i0[9] , \SB2_3_0/i0[8] ,
         \SB2_3_0/i0[7] , \SB2_3_0/i0[6] , \SB2_3_1/i3[0] , \SB2_3_1/i1_5 ,
         \SB2_3_1/i1_7 , \SB2_3_1/i1[9] , \SB2_3_1/i0_0 , \SB2_3_1/i0_3 ,
         \SB2_3_1/i0_4 , \SB2_3_1/i0[10] , \SB2_3_1/i0[9] , \SB2_3_1/i0[8] ,
         \SB2_3_1/i0[7] , \SB2_3_2/i3[0] , \SB2_3_2/i1_5 , \SB2_3_2/i1_7 ,
         \SB2_3_2/i1[9] , \SB2_3_2/i0_0 , \SB2_3_2/i0_3 , \SB2_3_2/i0_4 ,
         \SB2_3_2/i0[10] , \SB2_3_2/i0[9] , \SB2_3_2/i0[8] , \SB2_3_2/i0[7] ,
         \SB2_3_2/i0[6] , \SB2_3_3/i3[0] , \SB2_3_3/i1_5 , \SB2_3_3/i1_7 ,
         \SB2_3_3/i1[9] , \SB2_3_3/i0_0 , \SB2_3_3/i0_3 , \SB2_3_3/i0_4 ,
         \SB2_3_3/i0[10] , \SB2_3_3/i0[9] , \SB2_3_3/i0[8] , \SB2_3_3/i0[7] ,
         \SB2_3_3/i0[6] , \SB2_3_4/i3[0] , \SB2_3_4/i1_5 , \SB2_3_4/i1_7 ,
         \SB2_3_4/i1[9] , \SB2_3_4/i0_0 , \SB2_3_4/i0_3 , \SB2_3_4/i0_4 ,
         \SB2_3_4/i0[10] , \SB2_3_4/i0[8] , \SB2_3_4/i0[7] , \SB2_3_4/i0[6] ,
         \SB2_3_5/i3[0] , \SB2_3_5/i1_5 , \SB2_3_5/i1_7 , \SB2_3_5/i1[9] ,
         \SB2_3_5/i0_0 , \SB2_3_5/i0_3 , \SB2_3_5/i0_4 , \SB2_3_5/i0[10] ,
         \SB2_3_5/i0[8] , \SB2_3_5/i0[7] , \SB2_3_5/i0[6] , \SB2_3_6/i3[0] ,
         \SB2_3_6/i1_5 , \SB2_3_6/i1_7 , \SB2_3_6/i1[9] , \SB2_3_6/i0_0 ,
         \SB2_3_6/i0_3 , \SB2_3_6/i0[10] , \SB2_3_6/i0[9] , \SB2_3_6/i0[8] ,
         \SB2_3_6/i0[7] , \SB2_3_7/i3[0] , \SB2_3_7/i1_5 , \SB2_3_7/i1_7 ,
         \SB2_3_7/i1[9] , \SB2_3_7/i0_0 , \SB2_3_7/i0_3 , \SB2_3_7/i0_4 ,
         \SB2_3_7/i0[10] , \SB2_3_7/i0[9] , \SB2_3_7/i0[8] , \SB2_3_7/i0[7] ,
         \SB2_3_7/i0[6] , \SB2_3_8/i3[0] , \SB2_3_8/i1_5 , \SB2_3_8/i1_7 ,
         \SB2_3_8/i1[9] , \SB2_3_8/i0_0 , \SB2_3_8/i0_3 , \SB2_3_8/i0_4 ,
         \SB2_3_8/i0[10] , \SB2_3_8/i0[8] , \SB2_3_8/i0[7] , \SB2_3_8/i0[6] ,
         \SB2_3_9/i3[0] , \SB2_3_9/i1_5 , \SB2_3_9/i1_7 , \SB2_3_9/i1[9] ,
         \SB2_3_9/i0_0 , \SB2_3_9/i0_3 , \SB2_3_9/i0_4 , \SB2_3_9/i0[10] ,
         \SB2_3_9/i0[8] , \SB2_3_9/i0[7] , \SB2_3_9/i0[6] , \SB2_3_10/i3[0] ,
         \SB2_3_10/i1_5 , \SB2_3_10/i1_7 , \SB2_3_10/i1[9] , \SB2_3_10/i0_0 ,
         \SB2_3_10/i0_3 , \SB2_3_10/i0_4 , \SB2_3_10/i0[10] , \SB2_3_10/i0[9] ,
         \SB2_3_10/i0[8] , \SB2_3_10/i0[7] , \SB2_3_10/i0[6] ,
         \SB2_3_11/i3[0] , \SB2_3_11/i1_5 , \SB2_3_11/i1_7 , \SB2_3_11/i1[9] ,
         \SB2_3_11/i0_0 , \SB2_3_11/i0_3 , \SB2_3_11/i0[10] , \SB2_3_11/i0[9] ,
         \SB2_3_11/i0[8] , \SB2_3_11/i0[7] , \SB2_3_11/i0[6] ,
         \SB2_3_12/i3[0] , \SB2_3_12/i1_5 , \SB2_3_12/i1_7 , \SB2_3_12/i1[9] ,
         \SB2_3_12/i0_0 , \SB2_3_12/i0_3 , \SB2_3_12/i0_4 , \SB2_3_12/i0[10] ,
         \SB2_3_12/i0[9] , \SB2_3_12/i0[8] , \SB2_3_12/i0[7] ,
         \SB2_3_12/i0[6] , \SB2_3_13/i3[0] , \SB2_3_13/i1_5 , \SB2_3_13/i1_7 ,
         \SB2_3_13/i1[9] , \SB2_3_13/i0_0 , \SB2_3_13/i0_3 , \SB2_3_13/i0_4 ,
         \SB2_3_13/i0[10] , \SB2_3_13/i0[8] , \SB2_3_13/i0[7] ,
         \SB2_3_13/i0[6] , \SB2_3_14/i3[0] , \SB2_3_14/i1_5 , \SB2_3_14/i1_7 ,
         \SB2_3_14/i1[9] , \SB2_3_14/i0_0 , \SB2_3_14/i0_3 , \SB2_3_14/i0[10] ,
         \SB2_3_14/i0[9] , \SB2_3_14/i0[8] , \SB2_3_14/i0[7] ,
         \SB2_3_14/i0[6] , \SB2_3_15/i3[0] , \SB2_3_15/i1_5 , \SB2_3_15/i1[9] ,
         \SB2_3_15/i0_0 , \SB2_3_15/i0_3 , \SB2_3_15/i0_4 , \SB2_3_15/i0[10] ,
         \SB2_3_15/i0[9] , \SB2_3_15/i0[8] , \SB2_3_15/i0[7] ,
         \SB2_3_16/i3[0] , \SB2_3_16/i1_5 , \SB2_3_16/i1_7 , \SB2_3_16/i1[9] ,
         \SB2_3_16/i0_0 , \SB2_3_16/i0_3 , \SB2_3_16/i0[10] , \SB2_3_16/i0[8] ,
         \SB2_3_16/i0[6] , \SB2_3_17/i3[0] , \SB2_3_17/i1_5 , \SB2_3_17/i1_7 ,
         \SB2_3_17/i1[9] , \SB2_3_17/i0_0 , \SB2_3_17/i0_3 , \SB2_3_17/i0_4 ,
         \SB2_3_17/i0[10] , \SB2_3_17/i0[9] , \SB2_3_17/i0[8] ,
         \SB2_3_17/i0[7] , \SB2_3_17/i0[6] , \SB2_3_18/i3[0] , \SB2_3_18/i1_5 ,
         \SB2_3_18/i1_7 , \SB2_3_18/i1[9] , \SB2_3_18/i0_0 , \SB2_3_18/i0_3 ,
         \SB2_3_18/i0_4 , \SB2_3_18/i0[10] , \SB2_3_18/i0[9] ,
         \SB2_3_18/i0[8] , \SB2_3_18/i0[7] , \SB2_3_18/i0[6] ,
         \SB2_3_19/i3[0] , \SB2_3_19/i1_5 , \SB2_3_19/i1_7 , \SB2_3_19/i1[9] ,
         \SB2_3_19/i0_0 , \SB2_3_19/i0_3 , \SB2_3_19/i0_4 , \SB2_3_19/i0[10] ,
         \SB2_3_19/i0[8] , \SB2_3_19/i0[7] , \SB2_3_19/i0[6] ,
         \SB2_3_20/i3[0] , \SB2_3_20/i1_5 , \SB2_3_20/i1_7 , \SB2_3_20/i1[9] ,
         \SB2_3_20/i0_0 , \SB2_3_20/i0_3 , \SB2_3_20/i0_4 , \SB2_3_20/i0[10] ,
         \SB2_3_20/i0[9] , \SB2_3_20/i0[8] , \SB2_3_20/i0[7] ,
         \SB2_3_20/i0[6] , \SB2_3_21/i3[0] , \SB2_3_21/i1_5 , \SB2_3_21/i1_7 ,
         \SB2_3_21/i1[9] , \SB2_3_21/i0_0 , \SB2_3_21/i0_3 , \SB2_3_21/i0[10] ,
         \SB2_3_21/i0[9] , \SB2_3_21/i0[8] , \SB2_3_21/i0[7] ,
         \SB2_3_21/i0[6] , \SB2_3_22/i3[0] , \SB2_3_22/i1_5 , \SB2_3_22/i1_7 ,
         \SB2_3_22/i1[9] , \SB2_3_22/i0_0 , \SB2_3_22/i0_3 , \SB2_3_22/i0_4 ,
         \SB2_3_22/i0[10] , \SB2_3_22/i0[9] , \SB2_3_22/i0[8] ,
         \SB2_3_22/i0[7] , \SB2_3_22/i0[6] , \SB2_3_23/i3[0] , \SB2_3_23/i1_5 ,
         \SB2_3_23/i1_7 , \SB2_3_23/i1[9] , \SB2_3_23/i0_0 , \SB2_3_23/i0_3 ,
         \SB2_3_23/i0_4 , \SB2_3_23/i0[10] , \SB2_3_23/i0[9] ,
         \SB2_3_23/i0[8] , \SB2_3_23/i0[7] , \SB2_3_23/i0[6] ,
         \SB2_3_24/i3[0] , \SB2_3_24/i1_5 , \SB2_3_24/i1_7 , \SB2_3_24/i1[9] ,
         \SB2_3_24/i0_0 , \SB2_3_24/i0_3 , \SB2_3_24/i0_4 , \SB2_3_24/i0[10] ,
         \SB2_3_24/i0[9] , \SB2_3_24/i0[8] , \SB2_3_24/i0[7] ,
         \SB2_3_24/i0[6] , \SB2_3_25/i3[0] , \SB2_3_25/i1_5 , \SB2_3_25/i1_7 ,
         \SB2_3_25/i1[9] , \SB2_3_25/i0_0 , \SB2_3_25/i0_3 , \SB2_3_25/i0_4 ,
         \SB2_3_25/i0[10] , \SB2_3_25/i0[9] , \SB2_3_25/i0[8] ,
         \SB2_3_25/i0[7] , \SB2_3_25/i0[6] , \SB2_3_26/i3[0] , \SB2_3_26/i1_5 ,
         \SB2_3_26/i1_7 , \SB2_3_26/i1[9] , \SB2_3_26/i0_0 , \SB2_3_26/i0_3 ,
         \SB2_3_26/i0_4 , \SB2_3_26/i0[10] , \SB2_3_26/i0[9] ,
         \SB2_3_26/i0[8] , \SB2_3_26/i0[7] , \SB2_3_26/i0[6] ,
         \SB2_3_27/i3[0] , \SB2_3_27/i1_7 , \SB2_3_27/i1[9] , \SB2_3_27/i0_0 ,
         \SB2_3_27/i0_3 , \SB2_3_27/i0_4 , \SB2_3_27/i0[10] , \SB2_3_27/i0[9] ,
         \SB2_3_27/i0[8] , \SB2_3_27/i0[7] , \SB2_3_27/i0[6] ,
         \SB2_3_28/i3[0] , \SB2_3_28/i1_5 , \SB2_3_28/i1_7 , \SB2_3_28/i1[9] ,
         \SB2_3_28/i0_0 , \SB2_3_28/i0_3 , \SB2_3_28/i0_4 , \SB2_3_28/i0[10] ,
         \SB2_3_28/i0[9] , \SB2_3_28/i0[8] , \SB2_3_28/i0[7] ,
         \SB2_3_28/i0[6] , \SB2_3_29/i3[0] , \SB2_3_29/i1_5 , \SB2_3_29/i1_7 ,
         \SB2_3_29/i1[9] , \SB2_3_29/i0_0 , \SB2_3_29/i0_3 , \SB2_3_29/i0_4 ,
         \SB2_3_29/i0[10] , \SB2_3_29/i0[9] , \SB2_3_29/i0[8] ,
         \SB2_3_29/i0[7] , \SB2_3_30/i3[0] , \SB2_3_30/i1_5 , \SB2_3_30/i1_7 ,
         \SB2_3_30/i1[9] , \SB2_3_30/i0_0 , \SB2_3_30/i0_3 , \SB2_3_30/i0_4 ,
         \SB2_3_30/i0[10] , \SB2_3_30/i0[9] , \SB2_3_30/i0[8] ,
         \SB2_3_30/i0[7] , \SB2_3_30/i0[6] , \SB2_3_31/i3[0] , \SB2_3_31/i1_5 ,
         \SB2_3_31/i1_7 , \SB2_3_31/i1[9] , \SB2_3_31/i0_0 , \SB2_3_31/i0_3 ,
         \SB2_3_31/i0[10] , \SB2_3_31/i0[9] , \SB2_3_31/i0[8] ,
         \SB2_3_31/i0[6] , \SB4_0/i3[0] , \SB4_0/i1_5 , \SB4_0/i1_7 ,
         \SB4_0/i1[9] , \SB4_0/i0_0 , \SB4_0/i0_3 , \SB4_0/i0_4 ,
         \SB4_0/i0[10] , \SB4_0/i0[9] , \SB4_0/i0[8] , \SB4_0/i0[7] ,
         \SB4_0/i0[6] , \SB4_1/i3[0] , \SB4_1/i1_5 , \SB4_1/i1_7 ,
         \SB4_1/i1[9] , \SB4_1/i0_0 , \SB4_1/i0_3 , \SB4_1/i0_4 ,
         \SB4_1/i0[10] , \SB4_1/i0[9] , \SB4_1/i0[8] , \SB4_1/i0[7] ,
         \SB4_1/i0[6] , \SB4_2/i1_5 , \SB4_2/i1_7 , \SB4_2/i1[9] ,
         \SB4_2/i0_0 , \SB4_2/i0_3 , \SB4_2/i0_4 , \SB4_2/i0[10] ,
         \SB4_2/i0[8] , \SB4_2/i0[7] , \SB4_2/i0[6] , \SB4_3/i3[0] ,
         \SB4_3/i1_5 , \SB4_3/i1_7 , \SB4_3/i1[9] , \SB4_3/i0_0 , \SB4_3/i0_3 ,
         \SB4_3/i0_4 , \SB4_3/i0[10] , \SB4_3/i0[9] , \SB4_3/i0[8] ,
         \SB4_3/i0[7] , \SB4_3/i0[6] , \SB4_4/i3[0] , \SB4_4/i1_5 ,
         \SB4_4/i1_7 , \SB4_4/i1[9] , \SB4_4/i0_0 , \SB4_4/i0_3 , \SB4_4/i0_4 ,
         \SB4_4/i0[10] , \SB4_4/i0[9] , \SB4_4/i0[8] , \SB4_4/i0[7] ,
         \SB4_4/i0[6] , \SB4_5/i3[0] , \SB4_5/i1_5 , \SB4_5/i1_7 ,
         \SB4_5/i1[9] , \SB4_5/i0_0 , \SB4_5/i0_3 , \SB4_5/i0[10] ,
         \SB4_5/i0[9] , \SB4_5/i0[8] , \SB4_6/i3[0] , \SB4_6/i1_5 ,
         \SB4_6/i1_7 , \SB4_6/i1[9] , \SB4_6/i0_0 , \SB4_6/i0_3 , \SB4_6/i0_4 ,
         \SB4_6/i0[10] , \SB4_6/i0[9] , \SB4_6/i0[8] , \SB4_6/i0[7] ,
         \SB4_6/i0[6] , \SB4_7/i3[0] , \SB4_7/i1_5 , \SB4_7/i1_7 ,
         \SB4_7/i1[9] , \SB4_7/i0_0 , \SB4_7/i0_3 , \SB4_7/i0_4 ,
         \SB4_7/i0[10] , \SB4_7/i0[9] , \SB4_7/i0[8] , \SB4_7/i0[7] ,
         \SB4_7/i0[6] , \SB4_8/i3[0] , \SB4_8/i1_5 , \SB4_8/i1_7 ,
         \SB4_8/i1[9] , \SB4_8/i0_0 , \SB4_8/i0_3 , \SB4_8/i0[10] ,
         \SB4_8/i0[9] , \SB4_8/i0[8] , \SB4_8/i0[6] , \SB4_9/i3[0] ,
         \SB4_9/i1_5 , \SB4_9/i1_7 , \SB4_9/i1[9] , \SB4_9/i0_0 , \SB4_9/i0_3 ,
         \SB4_9/i0[10] , \SB4_9/i0[9] , \SB4_9/i0[8] , \SB4_9/i0[6] ,
         \SB4_10/i3[0] , \SB4_10/i1_5 , \SB4_10/i1_7 , \SB4_10/i1[9] ,
         \SB4_10/i0_0 , \SB4_10/i0_3 , \SB4_10/i0_4 , \SB4_10/i0[10] ,
         \SB4_10/i0[9] , \SB4_10/i0[8] , \SB4_10/i0[7] , \SB4_10/i0[6] ,
         \SB4_11/i3[0] , \SB4_11/i1_5 , \SB4_11/i1_7 , \SB4_11/i1[9] ,
         \SB4_11/i0_0 , \SB4_11/i0_3 , \SB4_11/i0[10] , \SB4_11/i0[9] ,
         \SB4_11/i0[8] , \SB4_11/i0[6] , \SB4_12/i3[0] , \SB4_12/i1_5 ,
         \SB4_12/i1_7 , \SB4_12/i1[9] , \SB4_12/i0_0 , \SB4_12/i0_3 ,
         \SB4_12/i0_4 , \SB4_12/i0[10] , \SB4_12/i0[9] , \SB4_12/i0[8] ,
         \SB4_12/i0[7] , \SB4_12/i0[6] , \SB4_13/i3[0] , \SB4_13/i1_5 ,
         \SB4_13/i1_7 , \SB4_13/i1[9] , \SB4_13/i0_0 , \SB4_13/i0_3 ,
         \SB4_13/i0_4 , \SB4_13/i0[10] , \SB4_13/i0[9] , \SB4_13/i0[8] ,
         \SB4_13/i0[7] , \SB4_13/i0[6] , \SB4_14/i3[0] , \SB4_14/i1_5 ,
         \SB4_14/i1_7 , \SB4_14/i1[9] , \SB4_14/i0_0 , \SB4_14/i0_3 ,
         \SB4_14/i0[10] , \SB4_14/i0[9] , \SB4_14/i0[8] , \SB4_15/i3[0] ,
         \SB4_15/i1_5 , \SB4_15/i1_7 , \SB4_15/i1[9] , \SB4_15/i0_0 ,
         \SB4_15/i0_3 , \SB4_15/i0_4 , \SB4_15/i0[10] , \SB4_15/i0[9] ,
         \SB4_15/i0[8] , \SB4_15/i0[7] , \SB4_15/i0[6] , \SB4_16/i3[0] ,
         \SB4_16/i1_5 , \SB4_16/i1_7 , \SB4_16/i1[9] , \SB4_16/i0_0 ,
         \SB4_16/i0_3 , \SB4_16/i0_4 , \SB4_16/i0[10] , \SB4_16/i0[9] ,
         \SB4_16/i0[8] , \SB4_16/i0[7] , \SB4_16/i0[6] , \SB4_17/i3[0] ,
         \SB4_17/i1_5 , \SB4_17/i1_7 , \SB4_17/i1[9] , \SB4_17/i0_0 ,
         \SB4_17/i0_3 , \SB4_17/i0_4 , \SB4_17/i0[10] , \SB4_17/i0[9] ,
         \SB4_17/i0[8] , \SB4_17/i0[7] , \SB4_17/i0[6] , \SB4_18/i3[0] ,
         \SB4_18/i1_5 , \SB4_18/i1_7 , \SB4_18/i0_0 , \SB4_18/i0_3 ,
         \SB4_18/i0_4 , \SB4_18/i0[10] , \SB4_18/i0[9] , \SB4_18/i0[8] ,
         \SB4_18/i0[7] , \SB4_18/i0[6] , \SB4_19/i3[0] , \SB4_19/i1_5 ,
         \SB4_19/i1_7 , \SB4_19/i1[9] , \SB4_19/i0_0 , \SB4_19/i0_3 ,
         \SB4_19/i0_4 , \SB4_19/i0[10] , \SB4_19/i0[9] , \SB4_19/i0[8] ,
         \SB4_19/i0[7] , \SB4_19/i0[6] , \SB4_20/i3[0] , \SB4_20/i1_5 ,
         \SB4_20/i1_7 , \SB4_20/i1[9] , \SB4_20/i0_0 , \SB4_20/i0_3 ,
         \SB4_20/i0[10] , \SB4_20/i0[9] , \SB4_20/i0[8] , \SB4_20/i0[6] ,
         \SB4_21/i3[0] , \SB4_21/i1_5 , \SB4_21/i1_7 , \SB4_21/i1[9] ,
         \SB4_21/i0_0 , \SB4_21/i0_3 , \SB4_21/i0_4 , \SB4_21/i0[10] ,
         \SB4_21/i0[9] , \SB4_21/i0[8] , \SB4_21/i0[7] , \SB4_21/i0[6] ,
         \SB4_22/i1_5 , \SB4_22/i1_7 , \SB4_22/i1[9] , \SB4_22/i0_0 ,
         \SB4_22/i0_3 , \SB4_22/i0_4 , \SB4_22/i0[10] , \SB4_22/i0[8] ,
         \SB4_22/i0[7] , \SB4_22/i0[6] , \SB4_23/i3[0] , \SB4_23/i1_5 ,
         \SB4_23/i1_7 , \SB4_23/i1[9] , \SB4_23/i0_0 , \SB4_23/i0_4 ,
         \SB4_23/i0[10] , \SB4_23/i0[9] , \SB4_23/i0[8] , \SB4_23/i0[7] ,
         \SB4_23/i0[6] , \SB4_24/i3[0] , \SB4_24/i1_5 , \SB4_24/i1_7 ,
         \SB4_24/i1[9] , \SB4_24/i0_0 , \SB4_24/i0_3 , \SB4_24/i0_4 ,
         \SB4_24/i0[10] , \SB4_24/i0[9] , \SB4_24/i0[8] , \SB4_24/i0[7] ,
         \SB4_24/i0[6] , \SB4_25/i3[0] , \SB4_25/i1_5 , \SB4_25/i1_7 ,
         \SB4_25/i1[9] , \SB4_25/i0_0 , \SB4_25/i0_3 , \SB4_25/i0_4 ,
         \SB4_25/i0[10] , \SB4_25/i0[9] , \SB4_25/i0[8] , \SB4_25/i0[6] ,
         \SB4_26/i3[0] , \SB4_26/i1_5 , \SB4_26/i1_7 , \SB4_26/i1[9] ,
         \SB4_26/i0_0 , \SB4_26/i0_3 , \SB4_26/i0_4 , \SB4_26/i0[10] ,
         \SB4_26/i0[9] , \SB4_26/i0[8] , \SB4_26/i0[7] , \SB4_26/i0[6] ,
         \SB4_27/i3[0] , \SB4_27/i1_5 , \SB4_27/i1_7 , \SB4_27/i1[9] ,
         \SB4_27/i0_0 , \SB4_27/i0[10] , \SB4_27/i0[9] , \SB4_27/i0[8] ,
         \SB4_27/i0[6] , \SB4_28/i3[0] , \SB4_28/i1_5 , \SB4_28/i1_7 ,
         \SB4_28/i1[9] , \SB4_28/i0_0 , \SB4_28/i0_3 , \SB4_28/i0_4 ,
         \SB4_28/i0[10] , \SB4_28/i0[9] , \SB4_28/i0[8] , \SB4_28/i0[7] ,
         \SB4_28/i0[6] , \SB4_29/i1_5 , \SB4_29/i1[9] , \SB4_29/i0_0 ,
         \SB4_29/i0_3 , \SB4_29/i0[10] , \SB4_29/i0[8] , \SB4_30/i3[0] ,
         \SB4_30/i1_5 , \SB4_30/i1_7 , \SB4_30/i1[9] , \SB4_30/i0_0 ,
         \SB4_30/i0_3 , \SB4_30/i0_4 , \SB4_30/i0[10] , \SB4_30/i0[9] ,
         \SB4_30/i0[8] , \SB4_30/i0[7] , \SB4_30/i0[6] , \SB4_31/i3[0] ,
         \SB4_31/i1_7 , \SB4_31/i1[9] , \SB4_31/i0_0 , \SB4_31/i0_4 ,
         \SB4_31/i0[10] , \SB4_31/i0[9] , \SB4_31/i0[8] , \SB4_31/i0[7] ,
         \SB4_31/i0[6] , \SB1_0_0/Component_Function_2/NAND4_in[3] ,
         \SB1_0_0/Component_Function_2/NAND4_in[2] ,
         \SB1_0_0/Component_Function_2/NAND4_in[1] ,
         \SB1_0_0/Component_Function_2/NAND4_in[0] ,
         \SB1_0_0/Component_Function_3/NAND4_in[3] ,
         \SB1_0_0/Component_Function_3/NAND4_in[2] ,
         \SB1_0_0/Component_Function_3/NAND4_in[1] ,
         \SB1_0_0/Component_Function_3/NAND4_in[0] ,
         \SB1_0_0/Component_Function_4/NAND4_in[3] ,
         \SB1_0_0/Component_Function_4/NAND4_in[2] ,
         \SB1_0_0/Component_Function_4/NAND4_in[1] ,
         \SB1_0_0/Component_Function_4/NAND4_in[0] ,
         \SB1_0_1/Component_Function_2/NAND4_in[2] ,
         \SB1_0_1/Component_Function_2/NAND4_in[1] ,
         \SB1_0_1/Component_Function_2/NAND4_in[0] ,
         \SB1_0_1/Component_Function_3/NAND4_in[3] ,
         \SB1_0_1/Component_Function_3/NAND4_in[2] ,
         \SB1_0_1/Component_Function_3/NAND4_in[1] ,
         \SB1_0_1/Component_Function_3/NAND4_in[0] ,
         \SB1_0_1/Component_Function_4/NAND4_in[3] ,
         \SB1_0_1/Component_Function_4/NAND4_in[2] ,
         \SB1_0_1/Component_Function_4/NAND4_in[1] ,
         \SB1_0_1/Component_Function_4/NAND4_in[0] ,
         \SB1_0_2/Component_Function_2/NAND4_in[3] ,
         \SB1_0_2/Component_Function_2/NAND4_in[2] ,
         \SB1_0_2/Component_Function_2/NAND4_in[1] ,
         \SB1_0_2/Component_Function_2/NAND4_in[0] ,
         \SB1_0_2/Component_Function_3/NAND4_in[3] ,
         \SB1_0_2/Component_Function_3/NAND4_in[2] ,
         \SB1_0_2/Component_Function_3/NAND4_in[1] ,
         \SB1_0_2/Component_Function_3/NAND4_in[0] ,
         \SB1_0_2/Component_Function_4/NAND4_in[3] ,
         \SB1_0_2/Component_Function_4/NAND4_in[2] ,
         \SB1_0_2/Component_Function_4/NAND4_in[1] ,
         \SB1_0_2/Component_Function_4/NAND4_in[0] ,
         \SB1_0_3/Component_Function_2/NAND4_in[3] ,
         \SB1_0_3/Component_Function_2/NAND4_in[2] ,
         \SB1_0_3/Component_Function_2/NAND4_in[1] ,
         \SB1_0_3/Component_Function_2/NAND4_in[0] ,
         \SB1_0_3/Component_Function_3/NAND4_in[3] ,
         \SB1_0_3/Component_Function_3/NAND4_in[2] ,
         \SB1_0_3/Component_Function_3/NAND4_in[1] ,
         \SB1_0_3/Component_Function_3/NAND4_in[0] ,
         \SB1_0_3/Component_Function_4/NAND4_in[3] ,
         \SB1_0_3/Component_Function_4/NAND4_in[2] ,
         \SB1_0_3/Component_Function_4/NAND4_in[1] ,
         \SB1_0_3/Component_Function_4/NAND4_in[0] ,
         \SB1_0_4/Component_Function_2/NAND4_in[3] ,
         \SB1_0_4/Component_Function_2/NAND4_in[2] ,
         \SB1_0_4/Component_Function_2/NAND4_in[1] ,
         \SB1_0_4/Component_Function_2/NAND4_in[0] ,
         \SB1_0_4/Component_Function_3/NAND4_in[3] ,
         \SB1_0_4/Component_Function_3/NAND4_in[2] ,
         \SB1_0_4/Component_Function_3/NAND4_in[1] ,
         \SB1_0_4/Component_Function_3/NAND4_in[0] ,
         \SB1_0_4/Component_Function_4/NAND4_in[3] ,
         \SB1_0_4/Component_Function_4/NAND4_in[2] ,
         \SB1_0_4/Component_Function_4/NAND4_in[1] ,
         \SB1_0_4/Component_Function_4/NAND4_in[0] ,
         \SB1_0_5/Component_Function_2/NAND4_in[3] ,
         \SB1_0_5/Component_Function_2/NAND4_in[2] ,
         \SB1_0_5/Component_Function_2/NAND4_in[1] ,
         \SB1_0_5/Component_Function_2/NAND4_in[0] ,
         \SB1_0_5/Component_Function_3/NAND4_in[3] ,
         \SB1_0_5/Component_Function_3/NAND4_in[2] ,
         \SB1_0_5/Component_Function_3/NAND4_in[1] ,
         \SB1_0_5/Component_Function_3/NAND4_in[0] ,
         \SB1_0_5/Component_Function_4/NAND4_in[3] ,
         \SB1_0_5/Component_Function_4/NAND4_in[2] ,
         \SB1_0_5/Component_Function_4/NAND4_in[1] ,
         \SB1_0_5/Component_Function_4/NAND4_in[0] ,
         \SB1_0_6/Component_Function_2/NAND4_in[3] ,
         \SB1_0_6/Component_Function_2/NAND4_in[2] ,
         \SB1_0_6/Component_Function_2/NAND4_in[1] ,
         \SB1_0_6/Component_Function_2/NAND4_in[0] ,
         \SB1_0_6/Component_Function_3/NAND4_in[3] ,
         \SB1_0_6/Component_Function_3/NAND4_in[2] ,
         \SB1_0_6/Component_Function_3/NAND4_in[1] ,
         \SB1_0_6/Component_Function_3/NAND4_in[0] ,
         \SB1_0_6/Component_Function_4/NAND4_in[3] ,
         \SB1_0_6/Component_Function_4/NAND4_in[2] ,
         \SB1_0_6/Component_Function_4/NAND4_in[1] ,
         \SB1_0_6/Component_Function_4/NAND4_in[0] ,
         \SB1_0_7/Component_Function_2/NAND4_in[3] ,
         \SB1_0_7/Component_Function_2/NAND4_in[2] ,
         \SB1_0_7/Component_Function_2/NAND4_in[1] ,
         \SB1_0_7/Component_Function_2/NAND4_in[0] ,
         \SB1_0_7/Component_Function_3/NAND4_in[3] ,
         \SB1_0_7/Component_Function_3/NAND4_in[2] ,
         \SB1_0_7/Component_Function_3/NAND4_in[1] ,
         \SB1_0_7/Component_Function_3/NAND4_in[0] ,
         \SB1_0_7/Component_Function_4/NAND4_in[3] ,
         \SB1_0_7/Component_Function_4/NAND4_in[2] ,
         \SB1_0_7/Component_Function_4/NAND4_in[1] ,
         \SB1_0_7/Component_Function_4/NAND4_in[0] ,
         \SB1_0_8/Component_Function_2/NAND4_in[2] ,
         \SB1_0_8/Component_Function_2/NAND4_in[1] ,
         \SB1_0_8/Component_Function_2/NAND4_in[0] ,
         \SB1_0_8/Component_Function_3/NAND4_in[3] ,
         \SB1_0_8/Component_Function_3/NAND4_in[1] ,
         \SB1_0_8/Component_Function_3/NAND4_in[0] ,
         \SB1_0_8/Component_Function_4/NAND4_in[3] ,
         \SB1_0_8/Component_Function_4/NAND4_in[2] ,
         \SB1_0_8/Component_Function_4/NAND4_in[0] ,
         \SB1_0_9/Component_Function_2/NAND4_in[3] ,
         \SB1_0_9/Component_Function_2/NAND4_in[2] ,
         \SB1_0_9/Component_Function_2/NAND4_in[1] ,
         \SB1_0_9/Component_Function_2/NAND4_in[0] ,
         \SB1_0_9/Component_Function_3/NAND4_in[3] ,
         \SB1_0_9/Component_Function_3/NAND4_in[2] ,
         \SB1_0_9/Component_Function_3/NAND4_in[1] ,
         \SB1_0_9/Component_Function_3/NAND4_in[0] ,
         \SB1_0_9/Component_Function_4/NAND4_in[3] ,
         \SB1_0_9/Component_Function_4/NAND4_in[2] ,
         \SB1_0_9/Component_Function_4/NAND4_in[1] ,
         \SB1_0_9/Component_Function_4/NAND4_in[0] ,
         \SB1_0_10/Component_Function_2/NAND4_in[3] ,
         \SB1_0_10/Component_Function_2/NAND4_in[2] ,
         \SB1_0_10/Component_Function_2/NAND4_in[1] ,
         \SB1_0_10/Component_Function_2/NAND4_in[0] ,
         \SB1_0_10/Component_Function_3/NAND4_in[3] ,
         \SB1_0_10/Component_Function_3/NAND4_in[2] ,
         \SB1_0_10/Component_Function_3/NAND4_in[1] ,
         \SB1_0_10/Component_Function_3/NAND4_in[0] ,
         \SB1_0_10/Component_Function_4/NAND4_in[3] ,
         \SB1_0_10/Component_Function_4/NAND4_in[2] ,
         \SB1_0_10/Component_Function_4/NAND4_in[1] ,
         \SB1_0_10/Component_Function_4/NAND4_in[0] ,
         \SB1_0_11/Component_Function_2/NAND4_in[3] ,
         \SB1_0_11/Component_Function_2/NAND4_in[2] ,
         \SB1_0_11/Component_Function_2/NAND4_in[1] ,
         \SB1_0_11/Component_Function_2/NAND4_in[0] ,
         \SB1_0_11/Component_Function_3/NAND4_in[3] ,
         \SB1_0_11/Component_Function_3/NAND4_in[2] ,
         \SB1_0_11/Component_Function_3/NAND4_in[1] ,
         \SB1_0_11/Component_Function_3/NAND4_in[0] ,
         \SB1_0_11/Component_Function_4/NAND4_in[3] ,
         \SB1_0_11/Component_Function_4/NAND4_in[2] ,
         \SB1_0_11/Component_Function_4/NAND4_in[1] ,
         \SB1_0_11/Component_Function_4/NAND4_in[0] ,
         \SB1_0_12/Component_Function_2/NAND4_in[3] ,
         \SB1_0_12/Component_Function_2/NAND4_in[2] ,
         \SB1_0_12/Component_Function_2/NAND4_in[1] ,
         \SB1_0_12/Component_Function_2/NAND4_in[0] ,
         \SB1_0_12/Component_Function_3/NAND4_in[3] ,
         \SB1_0_12/Component_Function_3/NAND4_in[2] ,
         \SB1_0_12/Component_Function_3/NAND4_in[1] ,
         \SB1_0_12/Component_Function_3/NAND4_in[0] ,
         \SB1_0_12/Component_Function_4/NAND4_in[3] ,
         \SB1_0_12/Component_Function_4/NAND4_in[2] ,
         \SB1_0_12/Component_Function_4/NAND4_in[1] ,
         \SB1_0_12/Component_Function_4/NAND4_in[0] ,
         \SB1_0_13/Component_Function_2/NAND4_in[2] ,
         \SB1_0_13/Component_Function_2/NAND4_in[1] ,
         \SB1_0_13/Component_Function_2/NAND4_in[0] ,
         \SB1_0_13/Component_Function_3/NAND4_in[3] ,
         \SB1_0_13/Component_Function_3/NAND4_in[2] ,
         \SB1_0_13/Component_Function_3/NAND4_in[1] ,
         \SB1_0_13/Component_Function_3/NAND4_in[0] ,
         \SB1_0_13/Component_Function_4/NAND4_in[3] ,
         \SB1_0_13/Component_Function_4/NAND4_in[2] ,
         \SB1_0_13/Component_Function_4/NAND4_in[1] ,
         \SB1_0_13/Component_Function_4/NAND4_in[0] ,
         \SB1_0_14/Component_Function_2/NAND4_in[3] ,
         \SB1_0_14/Component_Function_2/NAND4_in[2] ,
         \SB1_0_14/Component_Function_2/NAND4_in[1] ,
         \SB1_0_14/Component_Function_2/NAND4_in[0] ,
         \SB1_0_14/Component_Function_3/NAND4_in[3] ,
         \SB1_0_14/Component_Function_3/NAND4_in[2] ,
         \SB1_0_14/Component_Function_3/NAND4_in[1] ,
         \SB1_0_14/Component_Function_3/NAND4_in[0] ,
         \SB1_0_14/Component_Function_4/NAND4_in[3] ,
         \SB1_0_14/Component_Function_4/NAND4_in[2] ,
         \SB1_0_14/Component_Function_4/NAND4_in[1] ,
         \SB1_0_14/Component_Function_4/NAND4_in[0] ,
         \SB1_0_15/Component_Function_2/NAND4_in[3] ,
         \SB1_0_15/Component_Function_2/NAND4_in[2] ,
         \SB1_0_15/Component_Function_2/NAND4_in[1] ,
         \SB1_0_15/Component_Function_2/NAND4_in[0] ,
         \SB1_0_15/Component_Function_3/NAND4_in[3] ,
         \SB1_0_15/Component_Function_3/NAND4_in[2] ,
         \SB1_0_15/Component_Function_3/NAND4_in[1] ,
         \SB1_0_15/Component_Function_3/NAND4_in[0] ,
         \SB1_0_15/Component_Function_4/NAND4_in[3] ,
         \SB1_0_15/Component_Function_4/NAND4_in[2] ,
         \SB1_0_15/Component_Function_4/NAND4_in[1] ,
         \SB1_0_15/Component_Function_4/NAND4_in[0] ,
         \SB1_0_16/Component_Function_2/NAND4_in[3] ,
         \SB1_0_16/Component_Function_2/NAND4_in[2] ,
         \SB1_0_16/Component_Function_2/NAND4_in[1] ,
         \SB1_0_16/Component_Function_2/NAND4_in[0] ,
         \SB1_0_16/Component_Function_3/NAND4_in[3] ,
         \SB1_0_16/Component_Function_3/NAND4_in[2] ,
         \SB1_0_16/Component_Function_3/NAND4_in[1] ,
         \SB1_0_16/Component_Function_3/NAND4_in[0] ,
         \SB1_0_16/Component_Function_4/NAND4_in[3] ,
         \SB1_0_16/Component_Function_4/NAND4_in[2] ,
         \SB1_0_16/Component_Function_4/NAND4_in[1] ,
         \SB1_0_16/Component_Function_4/NAND4_in[0] ,
         \SB1_0_17/Component_Function_2/NAND4_in[3] ,
         \SB1_0_17/Component_Function_2/NAND4_in[2] ,
         \SB1_0_17/Component_Function_2/NAND4_in[1] ,
         \SB1_0_17/Component_Function_2/NAND4_in[0] ,
         \SB1_0_17/Component_Function_3/NAND4_in[3] ,
         \SB1_0_17/Component_Function_3/NAND4_in[2] ,
         \SB1_0_17/Component_Function_3/NAND4_in[1] ,
         \SB1_0_17/Component_Function_3/NAND4_in[0] ,
         \SB1_0_17/Component_Function_4/NAND4_in[3] ,
         \SB1_0_17/Component_Function_4/NAND4_in[2] ,
         \SB1_0_17/Component_Function_4/NAND4_in[1] ,
         \SB1_0_17/Component_Function_4/NAND4_in[0] ,
         \SB1_0_18/Component_Function_2/NAND4_in[3] ,
         \SB1_0_18/Component_Function_2/NAND4_in[2] ,
         \SB1_0_18/Component_Function_2/NAND4_in[1] ,
         \SB1_0_18/Component_Function_2/NAND4_in[0] ,
         \SB1_0_18/Component_Function_3/NAND4_in[3] ,
         \SB1_0_18/Component_Function_3/NAND4_in[2] ,
         \SB1_0_18/Component_Function_3/NAND4_in[1] ,
         \SB1_0_18/Component_Function_3/NAND4_in[0] ,
         \SB1_0_18/Component_Function_4/NAND4_in[2] ,
         \SB1_0_18/Component_Function_4/NAND4_in[1] ,
         \SB1_0_19/Component_Function_2/NAND4_in[3] ,
         \SB1_0_19/Component_Function_2/NAND4_in[2] ,
         \SB1_0_19/Component_Function_2/NAND4_in[1] ,
         \SB1_0_19/Component_Function_2/NAND4_in[0] ,
         \SB1_0_19/Component_Function_3/NAND4_in[3] ,
         \SB1_0_19/Component_Function_3/NAND4_in[1] ,
         \SB1_0_19/Component_Function_3/NAND4_in[0] ,
         \SB1_0_19/Component_Function_4/NAND4_in[3] ,
         \SB1_0_19/Component_Function_4/NAND4_in[2] ,
         \SB1_0_19/Component_Function_4/NAND4_in[1] ,
         \SB1_0_19/Component_Function_4/NAND4_in[0] ,
         \SB1_0_20/Component_Function_2/NAND4_in[3] ,
         \SB1_0_20/Component_Function_2/NAND4_in[2] ,
         \SB1_0_20/Component_Function_2/NAND4_in[1] ,
         \SB1_0_20/Component_Function_2/NAND4_in[0] ,
         \SB1_0_20/Component_Function_3/NAND4_in[3] ,
         \SB1_0_20/Component_Function_3/NAND4_in[2] ,
         \SB1_0_20/Component_Function_3/NAND4_in[1] ,
         \SB1_0_20/Component_Function_3/NAND4_in[0] ,
         \SB1_0_20/Component_Function_4/NAND4_in[3] ,
         \SB1_0_20/Component_Function_4/NAND4_in[2] ,
         \SB1_0_20/Component_Function_4/NAND4_in[1] ,
         \SB1_0_20/Component_Function_4/NAND4_in[0] ,
         \SB1_0_21/Component_Function_2/NAND4_in[3] ,
         \SB1_0_21/Component_Function_2/NAND4_in[2] ,
         \SB1_0_21/Component_Function_2/NAND4_in[1] ,
         \SB1_0_21/Component_Function_2/NAND4_in[0] ,
         \SB1_0_21/Component_Function_3/NAND4_in[3] ,
         \SB1_0_21/Component_Function_3/NAND4_in[2] ,
         \SB1_0_21/Component_Function_3/NAND4_in[1] ,
         \SB1_0_21/Component_Function_3/NAND4_in[0] ,
         \SB1_0_21/Component_Function_4/NAND4_in[3] ,
         \SB1_0_21/Component_Function_4/NAND4_in[2] ,
         \SB1_0_21/Component_Function_4/NAND4_in[1] ,
         \SB1_0_21/Component_Function_4/NAND4_in[0] ,
         \SB1_0_22/Component_Function_2/NAND4_in[3] ,
         \SB1_0_22/Component_Function_2/NAND4_in[2] ,
         \SB1_0_22/Component_Function_2/NAND4_in[1] ,
         \SB1_0_22/Component_Function_2/NAND4_in[0] ,
         \SB1_0_22/Component_Function_3/NAND4_in[3] ,
         \SB1_0_22/Component_Function_3/NAND4_in[2] ,
         \SB1_0_22/Component_Function_3/NAND4_in[1] ,
         \SB1_0_22/Component_Function_3/NAND4_in[0] ,
         \SB1_0_22/Component_Function_4/NAND4_in[3] ,
         \SB1_0_22/Component_Function_4/NAND4_in[2] ,
         \SB1_0_22/Component_Function_4/NAND4_in[1] ,
         \SB1_0_22/Component_Function_4/NAND4_in[0] ,
         \SB1_0_23/Component_Function_2/NAND4_in[3] ,
         \SB1_0_23/Component_Function_2/NAND4_in[2] ,
         \SB1_0_23/Component_Function_2/NAND4_in[1] ,
         \SB1_0_23/Component_Function_2/NAND4_in[0] ,
         \SB1_0_23/Component_Function_3/NAND4_in[3] ,
         \SB1_0_23/Component_Function_3/NAND4_in[2] ,
         \SB1_0_23/Component_Function_3/NAND4_in[1] ,
         \SB1_0_23/Component_Function_3/NAND4_in[0] ,
         \SB1_0_23/Component_Function_4/NAND4_in[2] ,
         \SB1_0_23/Component_Function_4/NAND4_in[1] ,
         \SB1_0_23/Component_Function_4/NAND4_in[0] ,
         \SB1_0_24/Component_Function_2/NAND4_in[3] ,
         \SB1_0_24/Component_Function_2/NAND4_in[2] ,
         \SB1_0_24/Component_Function_2/NAND4_in[1] ,
         \SB1_0_24/Component_Function_2/NAND4_in[0] ,
         \SB1_0_24/Component_Function_3/NAND4_in[3] ,
         \SB1_0_24/Component_Function_3/NAND4_in[2] ,
         \SB1_0_24/Component_Function_3/NAND4_in[1] ,
         \SB1_0_24/Component_Function_3/NAND4_in[0] ,
         \SB1_0_24/Component_Function_4/NAND4_in[3] ,
         \SB1_0_24/Component_Function_4/NAND4_in[2] ,
         \SB1_0_24/Component_Function_4/NAND4_in[1] ,
         \SB1_0_24/Component_Function_4/NAND4_in[0] ,
         \SB1_0_25/Component_Function_2/NAND4_in[3] ,
         \SB1_0_25/Component_Function_2/NAND4_in[2] ,
         \SB1_0_25/Component_Function_2/NAND4_in[1] ,
         \SB1_0_25/Component_Function_2/NAND4_in[0] ,
         \SB1_0_25/Component_Function_3/NAND4_in[3] ,
         \SB1_0_25/Component_Function_3/NAND4_in[2] ,
         \SB1_0_25/Component_Function_3/NAND4_in[1] ,
         \SB1_0_25/Component_Function_3/NAND4_in[0] ,
         \SB1_0_25/Component_Function_4/NAND4_in[3] ,
         \SB1_0_25/Component_Function_4/NAND4_in[2] ,
         \SB1_0_25/Component_Function_4/NAND4_in[1] ,
         \SB1_0_25/Component_Function_4/NAND4_in[0] ,
         \SB1_0_26/Component_Function_2/NAND4_in[3] ,
         \SB1_0_26/Component_Function_2/NAND4_in[2] ,
         \SB1_0_26/Component_Function_2/NAND4_in[1] ,
         \SB1_0_26/Component_Function_2/NAND4_in[0] ,
         \SB1_0_26/Component_Function_3/NAND4_in[3] ,
         \SB1_0_26/Component_Function_3/NAND4_in[2] ,
         \SB1_0_26/Component_Function_3/NAND4_in[1] ,
         \SB1_0_26/Component_Function_3/NAND4_in[0] ,
         \SB1_0_26/Component_Function_4/NAND4_in[3] ,
         \SB1_0_26/Component_Function_4/NAND4_in[2] ,
         \SB1_0_26/Component_Function_4/NAND4_in[1] ,
         \SB1_0_26/Component_Function_4/NAND4_in[0] ,
         \SB1_0_27/Component_Function_2/NAND4_in[3] ,
         \SB1_0_27/Component_Function_2/NAND4_in[2] ,
         \SB1_0_27/Component_Function_2/NAND4_in[1] ,
         \SB1_0_27/Component_Function_2/NAND4_in[0] ,
         \SB1_0_27/Component_Function_3/NAND4_in[3] ,
         \SB1_0_27/Component_Function_3/NAND4_in[2] ,
         \SB1_0_27/Component_Function_3/NAND4_in[1] ,
         \SB1_0_27/Component_Function_3/NAND4_in[0] ,
         \SB1_0_27/Component_Function_4/NAND4_in[3] ,
         \SB1_0_27/Component_Function_4/NAND4_in[2] ,
         \SB1_0_27/Component_Function_4/NAND4_in[1] ,
         \SB1_0_27/Component_Function_4/NAND4_in[0] ,
         \SB1_0_28/Component_Function_2/NAND4_in[3] ,
         \SB1_0_28/Component_Function_2/NAND4_in[2] ,
         \SB1_0_28/Component_Function_2/NAND4_in[1] ,
         \SB1_0_28/Component_Function_2/NAND4_in[0] ,
         \SB1_0_28/Component_Function_3/NAND4_in[3] ,
         \SB1_0_28/Component_Function_3/NAND4_in[2] ,
         \SB1_0_28/Component_Function_3/NAND4_in[1] ,
         \SB1_0_28/Component_Function_3/NAND4_in[0] ,
         \SB1_0_28/Component_Function_4/NAND4_in[3] ,
         \SB1_0_28/Component_Function_4/NAND4_in[2] ,
         \SB1_0_28/Component_Function_4/NAND4_in[1] ,
         \SB1_0_28/Component_Function_4/NAND4_in[0] ,
         \SB1_0_29/Component_Function_2/NAND4_in[3] ,
         \SB1_0_29/Component_Function_2/NAND4_in[2] ,
         \SB1_0_29/Component_Function_2/NAND4_in[1] ,
         \SB1_0_29/Component_Function_2/NAND4_in[0] ,
         \SB1_0_29/Component_Function_3/NAND4_in[3] ,
         \SB1_0_29/Component_Function_3/NAND4_in[2] ,
         \SB1_0_29/Component_Function_3/NAND4_in[1] ,
         \SB1_0_29/Component_Function_3/NAND4_in[0] ,
         \SB1_0_29/Component_Function_4/NAND4_in[3] ,
         \SB1_0_29/Component_Function_4/NAND4_in[2] ,
         \SB1_0_29/Component_Function_4/NAND4_in[1] ,
         \SB1_0_29/Component_Function_4/NAND4_in[0] ,
         \SB1_0_30/Component_Function_2/NAND4_in[3] ,
         \SB1_0_30/Component_Function_2/NAND4_in[2] ,
         \SB1_0_30/Component_Function_2/NAND4_in[1] ,
         \SB1_0_30/Component_Function_2/NAND4_in[0] ,
         \SB1_0_30/Component_Function_3/NAND4_in[1] ,
         \SB1_0_30/Component_Function_3/NAND4_in[0] ,
         \SB1_0_30/Component_Function_4/NAND4_in[3] ,
         \SB1_0_30/Component_Function_4/NAND4_in[2] ,
         \SB1_0_30/Component_Function_4/NAND4_in[1] ,
         \SB1_0_30/Component_Function_4/NAND4_in[0] ,
         \SB1_0_31/Component_Function_2/NAND4_in[2] ,
         \SB1_0_31/Component_Function_2/NAND4_in[1] ,
         \SB1_0_31/Component_Function_2/NAND4_in[0] ,
         \SB1_0_31/Component_Function_3/NAND4_in[3] ,
         \SB1_0_31/Component_Function_3/NAND4_in[2] ,
         \SB1_0_31/Component_Function_3/NAND4_in[1] ,
         \SB1_0_31/Component_Function_3/NAND4_in[0] ,
         \SB1_0_31/Component_Function_4/NAND4_in[3] ,
         \SB1_0_31/Component_Function_4/NAND4_in[2] ,
         \SB1_0_31/Component_Function_4/NAND4_in[1] ,
         \SB1_0_31/Component_Function_4/NAND4_in[0] ,
         \SB2_0_0/Component_Function_2/NAND4_in[1] ,
         \SB2_0_0/Component_Function_2/NAND4_in[0] ,
         \SB2_0_0/Component_Function_3/NAND4_in[2] ,
         \SB2_0_0/Component_Function_3/NAND4_in[0] ,
         \SB2_0_0/Component_Function_4/NAND4_in[2] ,
         \SB2_0_0/Component_Function_4/NAND4_in[1] ,
         \SB2_0_0/Component_Function_4/NAND4_in[0] ,
         \SB2_0_1/Component_Function_2/NAND4_in[2] ,
         \SB2_0_1/Component_Function_2/NAND4_in[1] ,
         \SB2_0_1/Component_Function_2/NAND4_in[0] ,
         \SB2_0_1/Component_Function_3/NAND4_in[2] ,
         \SB2_0_1/Component_Function_3/NAND4_in[1] ,
         \SB2_0_1/Component_Function_3/NAND4_in[0] ,
         \SB2_0_1/Component_Function_4/NAND4_in[2] ,
         \SB2_0_1/Component_Function_4/NAND4_in[1] ,
         \SB2_0_1/Component_Function_4/NAND4_in[0] ,
         \SB2_0_2/Component_Function_2/NAND4_in[3] ,
         \SB2_0_2/Component_Function_2/NAND4_in[2] ,
         \SB2_0_2/Component_Function_2/NAND4_in[1] ,
         \SB2_0_2/Component_Function_2/NAND4_in[0] ,
         \SB2_0_2/Component_Function_3/NAND4_in[3] ,
         \SB2_0_2/Component_Function_3/NAND4_in[2] ,
         \SB2_0_2/Component_Function_3/NAND4_in[1] ,
         \SB2_0_2/Component_Function_3/NAND4_in[0] ,
         \SB2_0_2/Component_Function_4/NAND4_in[3] ,
         \SB2_0_2/Component_Function_4/NAND4_in[2] ,
         \SB2_0_2/Component_Function_4/NAND4_in[1] ,
         \SB2_0_2/Component_Function_4/NAND4_in[0] ,
         \SB2_0_3/Component_Function_2/NAND4_in[2] ,
         \SB2_0_3/Component_Function_2/NAND4_in[1] ,
         \SB2_0_3/Component_Function_2/NAND4_in[0] ,
         \SB2_0_3/Component_Function_3/NAND4_in[3] ,
         \SB2_0_3/Component_Function_3/NAND4_in[2] ,
         \SB2_0_3/Component_Function_3/NAND4_in[1] ,
         \SB2_0_3/Component_Function_3/NAND4_in[0] ,
         \SB2_0_3/Component_Function_4/NAND4_in[3] ,
         \SB2_0_3/Component_Function_4/NAND4_in[2] ,
         \SB2_0_3/Component_Function_4/NAND4_in[1] ,
         \SB2_0_3/Component_Function_4/NAND4_in[0] ,
         \SB2_0_4/Component_Function_2/NAND4_in[3] ,
         \SB2_0_4/Component_Function_2/NAND4_in[2] ,
         \SB2_0_4/Component_Function_2/NAND4_in[1] ,
         \SB2_0_4/Component_Function_2/NAND4_in[0] ,
         \SB2_0_4/Component_Function_3/NAND4_in[1] ,
         \SB2_0_4/Component_Function_4/NAND4_in[2] ,
         \SB2_0_4/Component_Function_4/NAND4_in[1] ,
         \SB2_0_4/Component_Function_4/NAND4_in[0] ,
         \SB2_0_5/Component_Function_2/NAND4_in[3] ,
         \SB2_0_5/Component_Function_2/NAND4_in[2] ,
         \SB2_0_5/Component_Function_2/NAND4_in[1] ,
         \SB2_0_5/Component_Function_2/NAND4_in[0] ,
         \SB2_0_5/Component_Function_3/NAND4_in[2] ,
         \SB2_0_5/Component_Function_3/NAND4_in[0] ,
         \SB2_0_5/Component_Function_4/NAND4_in[3] ,
         \SB2_0_5/Component_Function_4/NAND4_in[2] ,
         \SB2_0_5/Component_Function_4/NAND4_in[1] ,
         \SB2_0_5/Component_Function_4/NAND4_in[0] ,
         \SB2_0_6/Component_Function_2/NAND4_in[3] ,
         \SB2_0_6/Component_Function_2/NAND4_in[2] ,
         \SB2_0_6/Component_Function_2/NAND4_in[1] ,
         \SB2_0_6/Component_Function_2/NAND4_in[0] ,
         \SB2_0_6/Component_Function_3/NAND4_in[3] ,
         \SB2_0_6/Component_Function_3/NAND4_in[2] ,
         \SB2_0_6/Component_Function_3/NAND4_in[1] ,
         \SB2_0_6/Component_Function_3/NAND4_in[0] ,
         \SB2_0_6/Component_Function_4/NAND4_in[2] ,
         \SB2_0_6/Component_Function_4/NAND4_in[1] ,
         \SB2_0_6/Component_Function_4/NAND4_in[0] ,
         \SB2_0_7/Component_Function_2/NAND4_in[2] ,
         \SB2_0_7/Component_Function_2/NAND4_in[1] ,
         \SB2_0_7/Component_Function_2/NAND4_in[0] ,
         \SB2_0_7/Component_Function_3/NAND4_in[2] ,
         \SB2_0_7/Component_Function_3/NAND4_in[1] ,
         \SB2_0_7/Component_Function_3/NAND4_in[0] ,
         \SB2_0_7/Component_Function_4/NAND4_in[1] ,
         \SB2_0_7/Component_Function_4/NAND4_in[0] ,
         \SB2_0_8/Component_Function_2/NAND4_in[3] ,
         \SB2_0_8/Component_Function_2/NAND4_in[2] ,
         \SB2_0_8/Component_Function_2/NAND4_in[1] ,
         \SB2_0_8/Component_Function_2/NAND4_in[0] ,
         \SB2_0_8/Component_Function_3/NAND4_in[2] ,
         \SB2_0_8/Component_Function_3/NAND4_in[1] ,
         \SB2_0_8/Component_Function_3/NAND4_in[0] ,
         \SB2_0_8/Component_Function_4/NAND4_in[3] ,
         \SB2_0_8/Component_Function_4/NAND4_in[1] ,
         \SB2_0_8/Component_Function_4/NAND4_in[0] ,
         \SB2_0_9/Component_Function_2/NAND4_in[2] ,
         \SB2_0_9/Component_Function_2/NAND4_in[1] ,
         \SB2_0_9/Component_Function_2/NAND4_in[0] ,
         \SB2_0_9/Component_Function_3/NAND4_in[3] ,
         \SB2_0_9/Component_Function_3/NAND4_in[2] ,
         \SB2_0_9/Component_Function_3/NAND4_in[1] ,
         \SB2_0_9/Component_Function_3/NAND4_in[0] ,
         \SB2_0_9/Component_Function_4/NAND4_in[2] ,
         \SB2_0_9/Component_Function_4/NAND4_in[1] ,
         \SB2_0_9/Component_Function_4/NAND4_in[0] ,
         \SB2_0_10/Component_Function_2/NAND4_in[3] ,
         \SB2_0_10/Component_Function_2/NAND4_in[1] ,
         \SB2_0_10/Component_Function_2/NAND4_in[0] ,
         \SB2_0_10/Component_Function_3/NAND4_in[2] ,
         \SB2_0_10/Component_Function_3/NAND4_in[1] ,
         \SB2_0_10/Component_Function_3/NAND4_in[0] ,
         \SB2_0_10/Component_Function_4/NAND4_in[3] ,
         \SB2_0_10/Component_Function_4/NAND4_in[2] ,
         \SB2_0_10/Component_Function_4/NAND4_in[1] ,
         \SB2_0_10/Component_Function_4/NAND4_in[0] ,
         \SB2_0_11/Component_Function_2/NAND4_in[3] ,
         \SB2_0_11/Component_Function_2/NAND4_in[2] ,
         \SB2_0_11/Component_Function_2/NAND4_in[1] ,
         \SB2_0_11/Component_Function_2/NAND4_in[0] ,
         \SB2_0_11/Component_Function_3/NAND4_in[3] ,
         \SB2_0_11/Component_Function_3/NAND4_in[2] ,
         \SB2_0_11/Component_Function_3/NAND4_in[1] ,
         \SB2_0_11/Component_Function_3/NAND4_in[0] ,
         \SB2_0_11/Component_Function_4/NAND4_in[2] ,
         \SB2_0_11/Component_Function_4/NAND4_in[1] ,
         \SB2_0_11/Component_Function_4/NAND4_in[0] ,
         \SB2_0_12/Component_Function_2/NAND4_in[3] ,
         \SB2_0_12/Component_Function_2/NAND4_in[2] ,
         \SB2_0_12/Component_Function_2/NAND4_in[1] ,
         \SB2_0_12/Component_Function_2/NAND4_in[0] ,
         \SB2_0_12/Component_Function_3/NAND4_in[2] ,
         \SB2_0_12/Component_Function_3/NAND4_in[1] ,
         \SB2_0_12/Component_Function_3/NAND4_in[0] ,
         \SB2_0_12/Component_Function_4/NAND4_in[3] ,
         \SB2_0_12/Component_Function_4/NAND4_in[2] ,
         \SB2_0_12/Component_Function_4/NAND4_in[1] ,
         \SB2_0_12/Component_Function_4/NAND4_in[0] ,
         \SB2_0_13/Component_Function_2/NAND4_in[2] ,
         \SB2_0_13/Component_Function_2/NAND4_in[1] ,
         \SB2_0_13/Component_Function_2/NAND4_in[0] ,
         \SB2_0_13/Component_Function_3/NAND4_in[3] ,
         \SB2_0_13/Component_Function_3/NAND4_in[2] ,
         \SB2_0_13/Component_Function_3/NAND4_in[1] ,
         \SB2_0_13/Component_Function_3/NAND4_in[0] ,
         \SB2_0_13/Component_Function_4/NAND4_in[3] ,
         \SB2_0_13/Component_Function_4/NAND4_in[2] ,
         \SB2_0_13/Component_Function_4/NAND4_in[1] ,
         \SB2_0_13/Component_Function_4/NAND4_in[0] ,
         \SB2_0_14/Component_Function_2/NAND4_in[2] ,
         \SB2_0_14/Component_Function_2/NAND4_in[1] ,
         \SB2_0_14/Component_Function_2/NAND4_in[0] ,
         \SB2_0_14/Component_Function_3/NAND4_in[3] ,
         \SB2_0_14/Component_Function_3/NAND4_in[2] ,
         \SB2_0_14/Component_Function_3/NAND4_in[0] ,
         \SB2_0_14/Component_Function_4/NAND4_in[3] ,
         \SB2_0_14/Component_Function_4/NAND4_in[2] ,
         \SB2_0_14/Component_Function_4/NAND4_in[1] ,
         \SB2_0_14/Component_Function_4/NAND4_in[0] ,
         \SB2_0_15/Component_Function_2/NAND4_in[3] ,
         \SB2_0_15/Component_Function_2/NAND4_in[2] ,
         \SB2_0_15/Component_Function_2/NAND4_in[1] ,
         \SB2_0_15/Component_Function_2/NAND4_in[0] ,
         \SB2_0_15/Component_Function_3/NAND4_in[3] ,
         \SB2_0_15/Component_Function_3/NAND4_in[2] ,
         \SB2_0_15/Component_Function_3/NAND4_in[1] ,
         \SB2_0_15/Component_Function_3/NAND4_in[0] ,
         \SB2_0_15/Component_Function_4/NAND4_in[3] ,
         \SB2_0_15/Component_Function_4/NAND4_in[2] ,
         \SB2_0_15/Component_Function_4/NAND4_in[1] ,
         \SB2_0_15/Component_Function_4/NAND4_in[0] ,
         \SB2_0_16/Component_Function_2/NAND4_in[3] ,
         \SB2_0_16/Component_Function_2/NAND4_in[2] ,
         \SB2_0_16/Component_Function_2/NAND4_in[0] ,
         \SB2_0_16/Component_Function_3/NAND4_in[3] ,
         \SB2_0_16/Component_Function_3/NAND4_in[2] ,
         \SB2_0_16/Component_Function_3/NAND4_in[1] ,
         \SB2_0_16/Component_Function_3/NAND4_in[0] ,
         \SB2_0_16/Component_Function_4/NAND4_in[3] ,
         \SB2_0_16/Component_Function_4/NAND4_in[1] ,
         \SB2_0_16/Component_Function_4/NAND4_in[0] ,
         \SB2_0_17/Component_Function_2/NAND4_in[3] ,
         \SB2_0_17/Component_Function_2/NAND4_in[1] ,
         \SB2_0_17/Component_Function_2/NAND4_in[0] ,
         \SB2_0_17/Component_Function_3/NAND4_in[3] ,
         \SB2_0_17/Component_Function_3/NAND4_in[2] ,
         \SB2_0_17/Component_Function_3/NAND4_in[1] ,
         \SB2_0_17/Component_Function_3/NAND4_in[0] ,
         \SB2_0_17/Component_Function_4/NAND4_in[3] ,
         \SB2_0_17/Component_Function_4/NAND4_in[2] ,
         \SB2_0_17/Component_Function_4/NAND4_in[1] ,
         \SB2_0_17/Component_Function_4/NAND4_in[0] ,
         \SB2_0_18/Component_Function_2/NAND4_in[2] ,
         \SB2_0_18/Component_Function_2/NAND4_in[1] ,
         \SB2_0_18/Component_Function_2/NAND4_in[0] ,
         \SB2_0_18/Component_Function_3/NAND4_in[2] ,
         \SB2_0_18/Component_Function_3/NAND4_in[1] ,
         \SB2_0_18/Component_Function_3/NAND4_in[0] ,
         \SB2_0_18/Component_Function_4/NAND4_in[3] ,
         \SB2_0_18/Component_Function_4/NAND4_in[2] ,
         \SB2_0_18/Component_Function_4/NAND4_in[1] ,
         \SB2_0_18/Component_Function_4/NAND4_in[0] ,
         \SB2_0_19/Component_Function_2/NAND4_in[2] ,
         \SB2_0_19/Component_Function_2/NAND4_in[1] ,
         \SB2_0_19/Component_Function_2/NAND4_in[0] ,
         \SB2_0_19/Component_Function_3/NAND4_in[3] ,
         \SB2_0_19/Component_Function_3/NAND4_in[2] ,
         \SB2_0_19/Component_Function_3/NAND4_in[1] ,
         \SB2_0_19/Component_Function_3/NAND4_in[0] ,
         \SB2_0_19/Component_Function_4/NAND4_in[3] ,
         \SB2_0_19/Component_Function_4/NAND4_in[2] ,
         \SB2_0_19/Component_Function_4/NAND4_in[1] ,
         \SB2_0_19/Component_Function_4/NAND4_in[0] ,
         \SB2_0_20/Component_Function_2/NAND4_in[2] ,
         \SB2_0_20/Component_Function_2/NAND4_in[1] ,
         \SB2_0_20/Component_Function_3/NAND4_in[3] ,
         \SB2_0_20/Component_Function_3/NAND4_in[2] ,
         \SB2_0_20/Component_Function_3/NAND4_in[1] ,
         \SB2_0_20/Component_Function_3/NAND4_in[0] ,
         \SB2_0_20/Component_Function_4/NAND4_in[3] ,
         \SB2_0_20/Component_Function_4/NAND4_in[2] ,
         \SB2_0_20/Component_Function_4/NAND4_in[1] ,
         \SB2_0_20/Component_Function_4/NAND4_in[0] ,
         \SB2_0_21/Component_Function_2/NAND4_in[2] ,
         \SB2_0_21/Component_Function_2/NAND4_in[1] ,
         \SB2_0_21/Component_Function_2/NAND4_in[0] ,
         \SB2_0_21/Component_Function_3/NAND4_in[3] ,
         \SB2_0_21/Component_Function_3/NAND4_in[2] ,
         \SB2_0_21/Component_Function_3/NAND4_in[1] ,
         \SB2_0_21/Component_Function_3/NAND4_in[0] ,
         \SB2_0_21/Component_Function_4/NAND4_in[1] ,
         \SB2_0_21/Component_Function_4/NAND4_in[0] ,
         \SB2_0_22/Component_Function_2/NAND4_in[2] ,
         \SB2_0_22/Component_Function_2/NAND4_in[1] ,
         \SB2_0_22/Component_Function_2/NAND4_in[0] ,
         \SB2_0_22/Component_Function_3/NAND4_in[3] ,
         \SB2_0_22/Component_Function_3/NAND4_in[2] ,
         \SB2_0_22/Component_Function_3/NAND4_in[1] ,
         \SB2_0_22/Component_Function_3/NAND4_in[0] ,
         \SB2_0_22/Component_Function_4/NAND4_in[2] ,
         \SB2_0_22/Component_Function_4/NAND4_in[1] ,
         \SB2_0_22/Component_Function_4/NAND4_in[0] ,
         \SB2_0_23/Component_Function_2/NAND4_in[2] ,
         \SB2_0_23/Component_Function_2/NAND4_in[1] ,
         \SB2_0_23/Component_Function_2/NAND4_in[0] ,
         \SB2_0_23/Component_Function_3/NAND4_in[2] ,
         \SB2_0_23/Component_Function_4/NAND4_in[3] ,
         \SB2_0_23/Component_Function_4/NAND4_in[1] ,
         \SB2_0_23/Component_Function_4/NAND4_in[0] ,
         \SB2_0_24/Component_Function_2/NAND4_in[2] ,
         \SB2_0_24/Component_Function_2/NAND4_in[1] ,
         \SB2_0_24/Component_Function_2/NAND4_in[0] ,
         \SB2_0_24/Component_Function_3/NAND4_in[3] ,
         \SB2_0_24/Component_Function_3/NAND4_in[2] ,
         \SB2_0_24/Component_Function_3/NAND4_in[1] ,
         \SB2_0_24/Component_Function_3/NAND4_in[0] ,
         \SB2_0_24/Component_Function_4/NAND4_in[2] ,
         \SB2_0_24/Component_Function_4/NAND4_in[1] ,
         \SB2_0_24/Component_Function_4/NAND4_in[0] ,
         \SB2_0_25/Component_Function_2/NAND4_in[3] ,
         \SB2_0_25/Component_Function_2/NAND4_in[2] ,
         \SB2_0_25/Component_Function_2/NAND4_in[1] ,
         \SB2_0_25/Component_Function_2/NAND4_in[0] ,
         \SB2_0_25/Component_Function_3/NAND4_in[3] ,
         \SB2_0_25/Component_Function_3/NAND4_in[2] ,
         \SB2_0_25/Component_Function_3/NAND4_in[1] ,
         \SB2_0_25/Component_Function_3/NAND4_in[0] ,
         \SB2_0_25/Component_Function_4/NAND4_in[3] ,
         \SB2_0_25/Component_Function_4/NAND4_in[1] ,
         \SB2_0_25/Component_Function_4/NAND4_in[0] ,
         \SB2_0_26/Component_Function_2/NAND4_in[3] ,
         \SB2_0_26/Component_Function_2/NAND4_in[2] ,
         \SB2_0_26/Component_Function_2/NAND4_in[1] ,
         \SB2_0_26/Component_Function_2/NAND4_in[0] ,
         \SB2_0_26/Component_Function_3/NAND4_in[3] ,
         \SB2_0_26/Component_Function_3/NAND4_in[1] ,
         \SB2_0_26/Component_Function_3/NAND4_in[0] ,
         \SB2_0_26/Component_Function_4/NAND4_in[3] ,
         \SB2_0_26/Component_Function_4/NAND4_in[1] ,
         \SB2_0_26/Component_Function_4/NAND4_in[0] ,
         \SB2_0_27/Component_Function_2/NAND4_in[3] ,
         \SB2_0_27/Component_Function_2/NAND4_in[2] ,
         \SB2_0_27/Component_Function_2/NAND4_in[1] ,
         \SB2_0_27/Component_Function_2/NAND4_in[0] ,
         \SB2_0_27/Component_Function_3/NAND4_in[2] ,
         \SB2_0_27/Component_Function_3/NAND4_in[1] ,
         \SB2_0_27/Component_Function_3/NAND4_in[0] ,
         \SB2_0_27/Component_Function_4/NAND4_in[3] ,
         \SB2_0_27/Component_Function_4/NAND4_in[1] ,
         \SB2_0_27/Component_Function_4/NAND4_in[0] ,
         \SB2_0_28/Component_Function_2/NAND4_in[2] ,
         \SB2_0_28/Component_Function_2/NAND4_in[1] ,
         \SB2_0_28/Component_Function_2/NAND4_in[0] ,
         \SB2_0_28/Component_Function_3/NAND4_in[2] ,
         \SB2_0_28/Component_Function_3/NAND4_in[1] ,
         \SB2_0_28/Component_Function_3/NAND4_in[0] ,
         \SB2_0_28/Component_Function_4/NAND4_in[3] ,
         \SB2_0_28/Component_Function_4/NAND4_in[2] ,
         \SB2_0_28/Component_Function_4/NAND4_in[1] ,
         \SB2_0_28/Component_Function_4/NAND4_in[0] ,
         \SB2_0_29/Component_Function_2/NAND4_in[2] ,
         \SB2_0_29/Component_Function_2/NAND4_in[1] ,
         \SB2_0_29/Component_Function_2/NAND4_in[0] ,
         \SB2_0_29/Component_Function_3/NAND4_in[3] ,
         \SB2_0_29/Component_Function_3/NAND4_in[2] ,
         \SB2_0_29/Component_Function_3/NAND4_in[1] ,
         \SB2_0_29/Component_Function_3/NAND4_in[0] ,
         \SB2_0_29/Component_Function_4/NAND4_in[3] ,
         \SB2_0_29/Component_Function_4/NAND4_in[2] ,
         \SB2_0_29/Component_Function_4/NAND4_in[1] ,
         \SB2_0_29/Component_Function_4/NAND4_in[0] ,
         \SB2_0_30/Component_Function_2/NAND4_in[2] ,
         \SB2_0_30/Component_Function_2/NAND4_in[1] ,
         \SB2_0_30/Component_Function_2/NAND4_in[0] ,
         \SB2_0_30/Component_Function_3/NAND4_in[3] ,
         \SB2_0_30/Component_Function_3/NAND4_in[2] ,
         \SB2_0_30/Component_Function_3/NAND4_in[1] ,
         \SB2_0_30/Component_Function_3/NAND4_in[0] ,
         \SB2_0_30/Component_Function_4/NAND4_in[2] ,
         \SB2_0_30/Component_Function_4/NAND4_in[1] ,
         \SB2_0_30/Component_Function_4/NAND4_in[0] ,
         \SB2_0_31/Component_Function_2/NAND4_in[3] ,
         \SB2_0_31/Component_Function_2/NAND4_in[2] ,
         \SB2_0_31/Component_Function_2/NAND4_in[1] ,
         \SB2_0_31/Component_Function_2/NAND4_in[0] ,
         \SB2_0_31/Component_Function_3/NAND4_in[3] ,
         \SB2_0_31/Component_Function_3/NAND4_in[2] ,
         \SB2_0_31/Component_Function_3/NAND4_in[1] ,
         \SB2_0_31/Component_Function_3/NAND4_in[0] ,
         \SB2_0_31/Component_Function_4/NAND4_in[3] ,
         \SB2_0_31/Component_Function_4/NAND4_in[1] ,
         \SB2_0_31/Component_Function_4/NAND4_in[0] ,
         \SB1_1_0/Component_Function_2/NAND4_in[3] ,
         \SB1_1_0/Component_Function_2/NAND4_in[2] ,
         \SB1_1_0/Component_Function_2/NAND4_in[1] ,
         \SB1_1_0/Component_Function_2/NAND4_in[0] ,
         \SB1_1_0/Component_Function_3/NAND4_in[3] ,
         \SB1_1_0/Component_Function_3/NAND4_in[2] ,
         \SB1_1_0/Component_Function_3/NAND4_in[1] ,
         \SB1_1_0/Component_Function_3/NAND4_in[0] ,
         \SB1_1_0/Component_Function_4/NAND4_in[3] ,
         \SB1_1_0/Component_Function_4/NAND4_in[2] ,
         \SB1_1_0/Component_Function_4/NAND4_in[1] ,
         \SB1_1_0/Component_Function_4/NAND4_in[0] ,
         \SB1_1_1/Component_Function_2/NAND4_in[2] ,
         \SB1_1_1/Component_Function_2/NAND4_in[1] ,
         \SB1_1_1/Component_Function_2/NAND4_in[0] ,
         \SB1_1_1/Component_Function_3/NAND4_in[3] ,
         \SB1_1_1/Component_Function_3/NAND4_in[2] ,
         \SB1_1_1/Component_Function_3/NAND4_in[1] ,
         \SB1_1_1/Component_Function_3/NAND4_in[0] ,
         \SB1_1_1/Component_Function_4/NAND4_in[3] ,
         \SB1_1_1/Component_Function_4/NAND4_in[2] ,
         \SB1_1_1/Component_Function_4/NAND4_in[1] ,
         \SB1_1_1/Component_Function_4/NAND4_in[0] ,
         \SB1_1_2/Component_Function_2/NAND4_in[3] ,
         \SB1_1_2/Component_Function_2/NAND4_in[2] ,
         \SB1_1_2/Component_Function_2/NAND4_in[1] ,
         \SB1_1_2/Component_Function_2/NAND4_in[0] ,
         \SB1_1_2/Component_Function_3/NAND4_in[3] ,
         \SB1_1_2/Component_Function_3/NAND4_in[2] ,
         \SB1_1_2/Component_Function_3/NAND4_in[1] ,
         \SB1_1_2/Component_Function_3/NAND4_in[0] ,
         \SB1_1_2/Component_Function_4/NAND4_in[3] ,
         \SB1_1_2/Component_Function_4/NAND4_in[1] ,
         \SB1_1_2/Component_Function_4/NAND4_in[0] ,
         \SB1_1_3/Component_Function_2/NAND4_in[2] ,
         \SB1_1_3/Component_Function_2/NAND4_in[1] ,
         \SB1_1_3/Component_Function_2/NAND4_in[0] ,
         \SB1_1_3/Component_Function_3/NAND4_in[3] ,
         \SB1_1_3/Component_Function_3/NAND4_in[2] ,
         \SB1_1_3/Component_Function_3/NAND4_in[1] ,
         \SB1_1_3/Component_Function_3/NAND4_in[0] ,
         \SB1_1_3/Component_Function_4/NAND4_in[3] ,
         \SB1_1_3/Component_Function_4/NAND4_in[2] ,
         \SB1_1_3/Component_Function_4/NAND4_in[1] ,
         \SB1_1_3/Component_Function_4/NAND4_in[0] ,
         \SB1_1_4/Component_Function_2/NAND4_in[2] ,
         \SB1_1_4/Component_Function_2/NAND4_in[1] ,
         \SB1_1_4/Component_Function_2/NAND4_in[0] ,
         \SB1_1_4/Component_Function_3/NAND4_in[3] ,
         \SB1_1_4/Component_Function_3/NAND4_in[2] ,
         \SB1_1_4/Component_Function_3/NAND4_in[1] ,
         \SB1_1_4/Component_Function_3/NAND4_in[0] ,
         \SB1_1_4/Component_Function_4/NAND4_in[3] ,
         \SB1_1_4/Component_Function_4/NAND4_in[1] ,
         \SB1_1_4/Component_Function_4/NAND4_in[0] ,
         \SB1_1_5/Component_Function_2/NAND4_in[3] ,
         \SB1_1_5/Component_Function_2/NAND4_in[2] ,
         \SB1_1_5/Component_Function_2/NAND4_in[1] ,
         \SB1_1_5/Component_Function_2/NAND4_in[0] ,
         \SB1_1_5/Component_Function_3/NAND4_in[3] ,
         \SB1_1_5/Component_Function_3/NAND4_in[2] ,
         \SB1_1_5/Component_Function_3/NAND4_in[1] ,
         \SB1_1_5/Component_Function_3/NAND4_in[0] ,
         \SB1_1_5/Component_Function_4/NAND4_in[3] ,
         \SB1_1_5/Component_Function_4/NAND4_in[2] ,
         \SB1_1_5/Component_Function_4/NAND4_in[1] ,
         \SB1_1_5/Component_Function_4/NAND4_in[0] ,
         \SB1_1_6/Component_Function_2/NAND4_in[2] ,
         \SB1_1_6/Component_Function_2/NAND4_in[1] ,
         \SB1_1_6/Component_Function_2/NAND4_in[0] ,
         \SB1_1_6/Component_Function_3/NAND4_in[3] ,
         \SB1_1_6/Component_Function_3/NAND4_in[2] ,
         \SB1_1_6/Component_Function_3/NAND4_in[1] ,
         \SB1_1_6/Component_Function_3/NAND4_in[0] ,
         \SB1_1_6/Component_Function_4/NAND4_in[3] ,
         \SB1_1_6/Component_Function_4/NAND4_in[2] ,
         \SB1_1_6/Component_Function_4/NAND4_in[1] ,
         \SB1_1_6/Component_Function_4/NAND4_in[0] ,
         \SB1_1_7/Component_Function_2/NAND4_in[2] ,
         \SB1_1_7/Component_Function_2/NAND4_in[1] ,
         \SB1_1_7/Component_Function_2/NAND4_in[0] ,
         \SB1_1_7/Component_Function_3/NAND4_in[3] ,
         \SB1_1_7/Component_Function_3/NAND4_in[1] ,
         \SB1_1_7/Component_Function_3/NAND4_in[0] ,
         \SB1_1_7/Component_Function_4/NAND4_in[3] ,
         \SB1_1_7/Component_Function_4/NAND4_in[1] ,
         \SB1_1_7/Component_Function_4/NAND4_in[0] ,
         \SB1_1_8/Component_Function_2/NAND4_in[3] ,
         \SB1_1_8/Component_Function_2/NAND4_in[2] ,
         \SB1_1_8/Component_Function_2/NAND4_in[1] ,
         \SB1_1_8/Component_Function_2/NAND4_in[0] ,
         \SB1_1_8/Component_Function_3/NAND4_in[2] ,
         \SB1_1_8/Component_Function_3/NAND4_in[1] ,
         \SB1_1_8/Component_Function_3/NAND4_in[0] ,
         \SB1_1_8/Component_Function_4/NAND4_in[3] ,
         \SB1_1_8/Component_Function_4/NAND4_in[2] ,
         \SB1_1_8/Component_Function_4/NAND4_in[1] ,
         \SB1_1_8/Component_Function_4/NAND4_in[0] ,
         \SB1_1_9/Component_Function_2/NAND4_in[3] ,
         \SB1_1_9/Component_Function_2/NAND4_in[2] ,
         \SB1_1_9/Component_Function_2/NAND4_in[1] ,
         \SB1_1_9/Component_Function_2/NAND4_in[0] ,
         \SB1_1_9/Component_Function_3/NAND4_in[3] ,
         \SB1_1_9/Component_Function_3/NAND4_in[2] ,
         \SB1_1_9/Component_Function_3/NAND4_in[1] ,
         \SB1_1_9/Component_Function_3/NAND4_in[0] ,
         \SB1_1_9/Component_Function_4/NAND4_in[3] ,
         \SB1_1_9/Component_Function_4/NAND4_in[2] ,
         \SB1_1_9/Component_Function_4/NAND4_in[1] ,
         \SB1_1_9/Component_Function_4/NAND4_in[0] ,
         \SB1_1_10/Component_Function_2/NAND4_in[2] ,
         \SB1_1_10/Component_Function_2/NAND4_in[1] ,
         \SB1_1_10/Component_Function_2/NAND4_in[0] ,
         \SB1_1_10/Component_Function_3/NAND4_in[3] ,
         \SB1_1_10/Component_Function_3/NAND4_in[2] ,
         \SB1_1_10/Component_Function_3/NAND4_in[1] ,
         \SB1_1_10/Component_Function_3/NAND4_in[0] ,
         \SB1_1_10/Component_Function_4/NAND4_in[3] ,
         \SB1_1_10/Component_Function_4/NAND4_in[2] ,
         \SB1_1_10/Component_Function_4/NAND4_in[1] ,
         \SB1_1_10/Component_Function_4/NAND4_in[0] ,
         \SB1_1_11/Component_Function_2/NAND4_in[2] ,
         \SB1_1_11/Component_Function_2/NAND4_in[1] ,
         \SB1_1_11/Component_Function_2/NAND4_in[0] ,
         \SB1_1_11/Component_Function_3/NAND4_in[3] ,
         \SB1_1_11/Component_Function_3/NAND4_in[2] ,
         \SB1_1_11/Component_Function_3/NAND4_in[1] ,
         \SB1_1_11/Component_Function_3/NAND4_in[0] ,
         \SB1_1_11/Component_Function_4/NAND4_in[3] ,
         \SB1_1_11/Component_Function_4/NAND4_in[2] ,
         \SB1_1_11/Component_Function_4/NAND4_in[1] ,
         \SB1_1_11/Component_Function_4/NAND4_in[0] ,
         \SB1_1_12/Component_Function_2/NAND4_in[2] ,
         \SB1_1_12/Component_Function_2/NAND4_in[1] ,
         \SB1_1_12/Component_Function_2/NAND4_in[0] ,
         \SB1_1_12/Component_Function_3/NAND4_in[3] ,
         \SB1_1_12/Component_Function_3/NAND4_in[2] ,
         \SB1_1_12/Component_Function_3/NAND4_in[1] ,
         \SB1_1_12/Component_Function_3/NAND4_in[0] ,
         \SB1_1_12/Component_Function_4/NAND4_in[3] ,
         \SB1_1_12/Component_Function_4/NAND4_in[1] ,
         \SB1_1_12/Component_Function_4/NAND4_in[0] ,
         \SB1_1_13/Component_Function_2/NAND4_in[2] ,
         \SB1_1_13/Component_Function_2/NAND4_in[1] ,
         \SB1_1_13/Component_Function_2/NAND4_in[0] ,
         \SB1_1_13/Component_Function_3/NAND4_in[3] ,
         \SB1_1_13/Component_Function_3/NAND4_in[2] ,
         \SB1_1_13/Component_Function_3/NAND4_in[1] ,
         \SB1_1_13/Component_Function_3/NAND4_in[0] ,
         \SB1_1_13/Component_Function_4/NAND4_in[3] ,
         \SB1_1_13/Component_Function_4/NAND4_in[2] ,
         \SB1_1_13/Component_Function_4/NAND4_in[1] ,
         \SB1_1_13/Component_Function_4/NAND4_in[0] ,
         \SB1_1_14/Component_Function_2/NAND4_in[3] ,
         \SB1_1_14/Component_Function_2/NAND4_in[2] ,
         \SB1_1_14/Component_Function_2/NAND4_in[1] ,
         \SB1_1_14/Component_Function_2/NAND4_in[0] ,
         \SB1_1_14/Component_Function_3/NAND4_in[3] ,
         \SB1_1_14/Component_Function_3/NAND4_in[2] ,
         \SB1_1_14/Component_Function_3/NAND4_in[1] ,
         \SB1_1_14/Component_Function_3/NAND4_in[0] ,
         \SB1_1_14/Component_Function_4/NAND4_in[3] ,
         \SB1_1_14/Component_Function_4/NAND4_in[2] ,
         \SB1_1_14/Component_Function_4/NAND4_in[1] ,
         \SB1_1_14/Component_Function_4/NAND4_in[0] ,
         \SB1_1_15/Component_Function_2/NAND4_in[3] ,
         \SB1_1_15/Component_Function_2/NAND4_in[2] ,
         \SB1_1_15/Component_Function_2/NAND4_in[1] ,
         \SB1_1_15/Component_Function_2/NAND4_in[0] ,
         \SB1_1_15/Component_Function_3/NAND4_in[3] ,
         \SB1_1_15/Component_Function_3/NAND4_in[2] ,
         \SB1_1_15/Component_Function_3/NAND4_in[1] ,
         \SB1_1_15/Component_Function_3/NAND4_in[0] ,
         \SB1_1_15/Component_Function_4/NAND4_in[3] ,
         \SB1_1_15/Component_Function_4/NAND4_in[2] ,
         \SB1_1_15/Component_Function_4/NAND4_in[1] ,
         \SB1_1_15/Component_Function_4/NAND4_in[0] ,
         \SB1_1_16/Component_Function_2/NAND4_in[3] ,
         \SB1_1_16/Component_Function_2/NAND4_in[2] ,
         \SB1_1_16/Component_Function_2/NAND4_in[1] ,
         \SB1_1_16/Component_Function_2/NAND4_in[0] ,
         \SB1_1_16/Component_Function_3/NAND4_in[3] ,
         \SB1_1_16/Component_Function_3/NAND4_in[2] ,
         \SB1_1_16/Component_Function_3/NAND4_in[1] ,
         \SB1_1_16/Component_Function_3/NAND4_in[0] ,
         \SB1_1_16/Component_Function_4/NAND4_in[2] ,
         \SB1_1_16/Component_Function_4/NAND4_in[1] ,
         \SB1_1_16/Component_Function_4/NAND4_in[0] ,
         \SB1_1_17/Component_Function_2/NAND4_in[2] ,
         \SB1_1_17/Component_Function_2/NAND4_in[1] ,
         \SB1_1_17/Component_Function_2/NAND4_in[0] ,
         \SB1_1_17/Component_Function_3/NAND4_in[3] ,
         \SB1_1_17/Component_Function_3/NAND4_in[2] ,
         \SB1_1_17/Component_Function_3/NAND4_in[1] ,
         \SB1_1_17/Component_Function_3/NAND4_in[0] ,
         \SB1_1_17/Component_Function_4/NAND4_in[3] ,
         \SB1_1_17/Component_Function_4/NAND4_in[2] ,
         \SB1_1_17/Component_Function_4/NAND4_in[1] ,
         \SB1_1_17/Component_Function_4/NAND4_in[0] ,
         \SB1_1_18/Component_Function_2/NAND4_in[3] ,
         \SB1_1_18/Component_Function_2/NAND4_in[2] ,
         \SB1_1_18/Component_Function_2/NAND4_in[1] ,
         \SB1_1_18/Component_Function_2/NAND4_in[0] ,
         \SB1_1_18/Component_Function_3/NAND4_in[3] ,
         \SB1_1_18/Component_Function_3/NAND4_in[2] ,
         \SB1_1_18/Component_Function_3/NAND4_in[1] ,
         \SB1_1_18/Component_Function_3/NAND4_in[0] ,
         \SB1_1_18/Component_Function_4/NAND4_in[3] ,
         \SB1_1_18/Component_Function_4/NAND4_in[2] ,
         \SB1_1_18/Component_Function_4/NAND4_in[1] ,
         \SB1_1_18/Component_Function_4/NAND4_in[0] ,
         \SB1_1_19/Component_Function_2/NAND4_in[3] ,
         \SB1_1_19/Component_Function_2/NAND4_in[2] ,
         \SB1_1_19/Component_Function_2/NAND4_in[1] ,
         \SB1_1_19/Component_Function_2/NAND4_in[0] ,
         \SB1_1_19/Component_Function_3/NAND4_in[3] ,
         \SB1_1_19/Component_Function_3/NAND4_in[2] ,
         \SB1_1_19/Component_Function_3/NAND4_in[1] ,
         \SB1_1_19/Component_Function_3/NAND4_in[0] ,
         \SB1_1_19/Component_Function_4/NAND4_in[3] ,
         \SB1_1_19/Component_Function_4/NAND4_in[2] ,
         \SB1_1_19/Component_Function_4/NAND4_in[1] ,
         \SB1_1_19/Component_Function_4/NAND4_in[0] ,
         \SB1_1_20/Component_Function_2/NAND4_in[3] ,
         \SB1_1_20/Component_Function_2/NAND4_in[2] ,
         \SB1_1_20/Component_Function_2/NAND4_in[1] ,
         \SB1_1_20/Component_Function_2/NAND4_in[0] ,
         \SB1_1_20/Component_Function_3/NAND4_in[2] ,
         \SB1_1_20/Component_Function_3/NAND4_in[1] ,
         \SB1_1_20/Component_Function_3/NAND4_in[0] ,
         \SB1_1_20/Component_Function_4/NAND4_in[3] ,
         \SB1_1_20/Component_Function_4/NAND4_in[2] ,
         \SB1_1_20/Component_Function_4/NAND4_in[1] ,
         \SB1_1_20/Component_Function_4/NAND4_in[0] ,
         \SB1_1_21/Component_Function_2/NAND4_in[3] ,
         \SB1_1_21/Component_Function_2/NAND4_in[2] ,
         \SB1_1_21/Component_Function_2/NAND4_in[1] ,
         \SB1_1_21/Component_Function_2/NAND4_in[0] ,
         \SB1_1_21/Component_Function_3/NAND4_in[3] ,
         \SB1_1_21/Component_Function_3/NAND4_in[2] ,
         \SB1_1_21/Component_Function_3/NAND4_in[1] ,
         \SB1_1_21/Component_Function_3/NAND4_in[0] ,
         \SB1_1_21/Component_Function_4/NAND4_in[3] ,
         \SB1_1_21/Component_Function_4/NAND4_in[2] ,
         \SB1_1_21/Component_Function_4/NAND4_in[1] ,
         \SB1_1_21/Component_Function_4/NAND4_in[0] ,
         \SB1_1_22/Component_Function_2/NAND4_in[2] ,
         \SB1_1_22/Component_Function_2/NAND4_in[1] ,
         \SB1_1_22/Component_Function_2/NAND4_in[0] ,
         \SB1_1_22/Component_Function_3/NAND4_in[3] ,
         \SB1_1_22/Component_Function_3/NAND4_in[2] ,
         \SB1_1_22/Component_Function_3/NAND4_in[1] ,
         \SB1_1_22/Component_Function_3/NAND4_in[0] ,
         \SB1_1_22/Component_Function_4/NAND4_in[3] ,
         \SB1_1_22/Component_Function_4/NAND4_in[2] ,
         \SB1_1_22/Component_Function_4/NAND4_in[1] ,
         \SB1_1_22/Component_Function_4/NAND4_in[0] ,
         \SB1_1_23/Component_Function_2/NAND4_in[3] ,
         \SB1_1_23/Component_Function_2/NAND4_in[2] ,
         \SB1_1_23/Component_Function_2/NAND4_in[1] ,
         \SB1_1_23/Component_Function_2/NAND4_in[0] ,
         \SB1_1_23/Component_Function_3/NAND4_in[3] ,
         \SB1_1_23/Component_Function_3/NAND4_in[2] ,
         \SB1_1_23/Component_Function_3/NAND4_in[1] ,
         \SB1_1_23/Component_Function_3/NAND4_in[0] ,
         \SB1_1_23/Component_Function_4/NAND4_in[3] ,
         \SB1_1_23/Component_Function_4/NAND4_in[2] ,
         \SB1_1_23/Component_Function_4/NAND4_in[1] ,
         \SB1_1_23/Component_Function_4/NAND4_in[0] ,
         \SB1_1_24/Component_Function_2/NAND4_in[2] ,
         \SB1_1_24/Component_Function_2/NAND4_in[1] ,
         \SB1_1_24/Component_Function_2/NAND4_in[0] ,
         \SB1_1_24/Component_Function_3/NAND4_in[3] ,
         \SB1_1_24/Component_Function_3/NAND4_in[2] ,
         \SB1_1_24/Component_Function_3/NAND4_in[1] ,
         \SB1_1_24/Component_Function_3/NAND4_in[0] ,
         \SB1_1_24/Component_Function_4/NAND4_in[3] ,
         \SB1_1_24/Component_Function_4/NAND4_in[2] ,
         \SB1_1_24/Component_Function_4/NAND4_in[1] ,
         \SB1_1_24/Component_Function_4/NAND4_in[0] ,
         \SB1_1_25/Component_Function_2/NAND4_in[2] ,
         \SB1_1_25/Component_Function_2/NAND4_in[1] ,
         \SB1_1_25/Component_Function_2/NAND4_in[0] ,
         \SB1_1_25/Component_Function_3/NAND4_in[3] ,
         \SB1_1_25/Component_Function_3/NAND4_in[2] ,
         \SB1_1_25/Component_Function_3/NAND4_in[1] ,
         \SB1_1_25/Component_Function_3/NAND4_in[0] ,
         \SB1_1_25/Component_Function_4/NAND4_in[3] ,
         \SB1_1_25/Component_Function_4/NAND4_in[2] ,
         \SB1_1_25/Component_Function_4/NAND4_in[1] ,
         \SB1_1_25/Component_Function_4/NAND4_in[0] ,
         \SB1_1_26/Component_Function_2/NAND4_in[3] ,
         \SB1_1_26/Component_Function_2/NAND4_in[2] ,
         \SB1_1_26/Component_Function_2/NAND4_in[1] ,
         \SB1_1_26/Component_Function_2/NAND4_in[0] ,
         \SB1_1_26/Component_Function_3/NAND4_in[3] ,
         \SB1_1_26/Component_Function_3/NAND4_in[2] ,
         \SB1_1_26/Component_Function_3/NAND4_in[1] ,
         \SB1_1_26/Component_Function_3/NAND4_in[0] ,
         \SB1_1_26/Component_Function_4/NAND4_in[3] ,
         \SB1_1_26/Component_Function_4/NAND4_in[2] ,
         \SB1_1_26/Component_Function_4/NAND4_in[1] ,
         \SB1_1_26/Component_Function_4/NAND4_in[0] ,
         \SB1_1_27/Component_Function_2/NAND4_in[2] ,
         \SB1_1_27/Component_Function_2/NAND4_in[1] ,
         \SB1_1_27/Component_Function_2/NAND4_in[0] ,
         \SB1_1_27/Component_Function_3/NAND4_in[3] ,
         \SB1_1_27/Component_Function_3/NAND4_in[2] ,
         \SB1_1_27/Component_Function_3/NAND4_in[1] ,
         \SB1_1_27/Component_Function_3/NAND4_in[0] ,
         \SB1_1_27/Component_Function_4/NAND4_in[3] ,
         \SB1_1_27/Component_Function_4/NAND4_in[2] ,
         \SB1_1_27/Component_Function_4/NAND4_in[1] ,
         \SB1_1_27/Component_Function_4/NAND4_in[0] ,
         \SB1_1_28/Component_Function_2/NAND4_in[2] ,
         \SB1_1_28/Component_Function_2/NAND4_in[1] ,
         \SB1_1_28/Component_Function_2/NAND4_in[0] ,
         \SB1_1_28/Component_Function_3/NAND4_in[3] ,
         \SB1_1_28/Component_Function_3/NAND4_in[2] ,
         \SB1_1_28/Component_Function_3/NAND4_in[1] ,
         \SB1_1_28/Component_Function_3/NAND4_in[0] ,
         \SB1_1_28/Component_Function_4/NAND4_in[3] ,
         \SB1_1_28/Component_Function_4/NAND4_in[1] ,
         \SB1_1_28/Component_Function_4/NAND4_in[0] ,
         \SB1_1_29/Component_Function_2/NAND4_in[3] ,
         \SB1_1_29/Component_Function_2/NAND4_in[2] ,
         \SB1_1_29/Component_Function_2/NAND4_in[1] ,
         \SB1_1_29/Component_Function_2/NAND4_in[0] ,
         \SB1_1_29/Component_Function_3/NAND4_in[3] ,
         \SB1_1_29/Component_Function_3/NAND4_in[2] ,
         \SB1_1_29/Component_Function_3/NAND4_in[1] ,
         \SB1_1_29/Component_Function_3/NAND4_in[0] ,
         \SB1_1_29/Component_Function_4/NAND4_in[3] ,
         \SB1_1_29/Component_Function_4/NAND4_in[2] ,
         \SB1_1_29/Component_Function_4/NAND4_in[1] ,
         \SB1_1_29/Component_Function_4/NAND4_in[0] ,
         \SB1_1_30/Component_Function_2/NAND4_in[2] ,
         \SB1_1_30/Component_Function_2/NAND4_in[1] ,
         \SB1_1_30/Component_Function_2/NAND4_in[0] ,
         \SB1_1_30/Component_Function_3/NAND4_in[3] ,
         \SB1_1_30/Component_Function_3/NAND4_in[2] ,
         \SB1_1_30/Component_Function_3/NAND4_in[1] ,
         \SB1_1_30/Component_Function_3/NAND4_in[0] ,
         \SB1_1_30/Component_Function_4/NAND4_in[3] ,
         \SB1_1_30/Component_Function_4/NAND4_in[2] ,
         \SB1_1_30/Component_Function_4/NAND4_in[1] ,
         \SB1_1_30/Component_Function_4/NAND4_in[0] ,
         \SB1_1_31/Component_Function_2/NAND4_in[3] ,
         \SB1_1_31/Component_Function_2/NAND4_in[2] ,
         \SB1_1_31/Component_Function_2/NAND4_in[1] ,
         \SB1_1_31/Component_Function_2/NAND4_in[0] ,
         \SB1_1_31/Component_Function_3/NAND4_in[3] ,
         \SB1_1_31/Component_Function_3/NAND4_in[2] ,
         \SB1_1_31/Component_Function_3/NAND4_in[1] ,
         \SB1_1_31/Component_Function_3/NAND4_in[0] ,
         \SB1_1_31/Component_Function_4/NAND4_in[2] ,
         \SB1_1_31/Component_Function_4/NAND4_in[1] ,
         \SB1_1_31/Component_Function_4/NAND4_in[0] ,
         \SB2_1_0/Component_Function_2/NAND4_in[2] ,
         \SB2_1_0/Component_Function_2/NAND4_in[1] ,
         \SB2_1_0/Component_Function_2/NAND4_in[0] ,
         \SB2_1_0/Component_Function_3/NAND4_in[2] ,
         \SB2_1_0/Component_Function_3/NAND4_in[1] ,
         \SB2_1_0/Component_Function_3/NAND4_in[0] ,
         \SB2_1_0/Component_Function_4/NAND4_in[3] ,
         \SB2_1_0/Component_Function_4/NAND4_in[2] ,
         \SB2_1_0/Component_Function_4/NAND4_in[1] ,
         \SB2_1_0/Component_Function_4/NAND4_in[0] ,
         \SB2_1_1/Component_Function_2/NAND4_in[3] ,
         \SB2_1_1/Component_Function_2/NAND4_in[1] ,
         \SB2_1_1/Component_Function_2/NAND4_in[0] ,
         \SB2_1_1/Component_Function_3/NAND4_in[3] ,
         \SB2_1_1/Component_Function_3/NAND4_in[2] ,
         \SB2_1_1/Component_Function_3/NAND4_in[1] ,
         \SB2_1_1/Component_Function_3/NAND4_in[0] ,
         \SB2_1_1/Component_Function_4/NAND4_in[3] ,
         \SB2_1_1/Component_Function_4/NAND4_in[2] ,
         \SB2_1_1/Component_Function_4/NAND4_in[1] ,
         \SB2_1_1/Component_Function_4/NAND4_in[0] ,
         \SB2_1_2/Component_Function_2/NAND4_in[2] ,
         \SB2_1_2/Component_Function_2/NAND4_in[1] ,
         \SB2_1_2/Component_Function_2/NAND4_in[0] ,
         \SB2_1_2/Component_Function_3/NAND4_in[2] ,
         \SB2_1_2/Component_Function_3/NAND4_in[1] ,
         \SB2_1_2/Component_Function_3/NAND4_in[0] ,
         \SB2_1_2/Component_Function_4/NAND4_in[3] ,
         \SB2_1_2/Component_Function_4/NAND4_in[2] ,
         \SB2_1_2/Component_Function_4/NAND4_in[1] ,
         \SB2_1_2/Component_Function_4/NAND4_in[0] ,
         \SB2_1_3/Component_Function_2/NAND4_in[2] ,
         \SB2_1_3/Component_Function_2/NAND4_in[1] ,
         \SB2_1_3/Component_Function_2/NAND4_in[0] ,
         \SB2_1_3/Component_Function_3/NAND4_in[3] ,
         \SB2_1_3/Component_Function_3/NAND4_in[2] ,
         \SB2_1_3/Component_Function_3/NAND4_in[1] ,
         \SB2_1_3/Component_Function_3/NAND4_in[0] ,
         \SB2_1_3/Component_Function_4/NAND4_in[2] ,
         \SB2_1_3/Component_Function_4/NAND4_in[1] ,
         \SB2_1_3/Component_Function_4/NAND4_in[0] ,
         \SB2_1_4/Component_Function_2/NAND4_in[3] ,
         \SB2_1_4/Component_Function_2/NAND4_in[2] ,
         \SB2_1_4/Component_Function_2/NAND4_in[1] ,
         \SB2_1_4/Component_Function_2/NAND4_in[0] ,
         \SB2_1_4/Component_Function_3/NAND4_in[3] ,
         \SB2_1_4/Component_Function_3/NAND4_in[2] ,
         \SB2_1_4/Component_Function_3/NAND4_in[1] ,
         \SB2_1_4/Component_Function_3/NAND4_in[0] ,
         \SB2_1_4/Component_Function_4/NAND4_in[3] ,
         \SB2_1_4/Component_Function_4/NAND4_in[2] ,
         \SB2_1_4/Component_Function_4/NAND4_in[1] ,
         \SB2_1_4/Component_Function_4/NAND4_in[0] ,
         \SB2_1_5/Component_Function_2/NAND4_in[3] ,
         \SB2_1_5/Component_Function_2/NAND4_in[2] ,
         \SB2_1_5/Component_Function_2/NAND4_in[1] ,
         \SB2_1_5/Component_Function_2/NAND4_in[0] ,
         \SB2_1_5/Component_Function_3/NAND4_in[3] ,
         \SB2_1_5/Component_Function_3/NAND4_in[2] ,
         \SB2_1_5/Component_Function_3/NAND4_in[1] ,
         \SB2_1_5/Component_Function_3/NAND4_in[0] ,
         \SB2_1_5/Component_Function_4/NAND4_in[3] ,
         \SB2_1_5/Component_Function_4/NAND4_in[1] ,
         \SB2_1_5/Component_Function_4/NAND4_in[0] ,
         \SB2_1_6/Component_Function_2/NAND4_in[2] ,
         \SB2_1_6/Component_Function_2/NAND4_in[1] ,
         \SB2_1_6/Component_Function_2/NAND4_in[0] ,
         \SB2_1_6/Component_Function_3/NAND4_in[3] ,
         \SB2_1_6/Component_Function_3/NAND4_in[1] ,
         \SB2_1_6/Component_Function_3/NAND4_in[0] ,
         \SB2_1_6/Component_Function_4/NAND4_in[3] ,
         \SB2_1_6/Component_Function_4/NAND4_in[1] ,
         \SB2_1_6/Component_Function_4/NAND4_in[0] ,
         \SB2_1_7/Component_Function_2/NAND4_in[2] ,
         \SB2_1_7/Component_Function_2/NAND4_in[1] ,
         \SB2_1_7/Component_Function_2/NAND4_in[0] ,
         \SB2_1_7/Component_Function_3/NAND4_in[3] ,
         \SB2_1_7/Component_Function_3/NAND4_in[2] ,
         \SB2_1_7/Component_Function_3/NAND4_in[1] ,
         \SB2_1_7/Component_Function_3/NAND4_in[0] ,
         \SB2_1_7/Component_Function_4/NAND4_in[3] ,
         \SB2_1_7/Component_Function_4/NAND4_in[2] ,
         \SB2_1_7/Component_Function_4/NAND4_in[1] ,
         \SB2_1_7/Component_Function_4/NAND4_in[0] ,
         \SB2_1_8/Component_Function_2/NAND4_in[2] ,
         \SB2_1_8/Component_Function_2/NAND4_in[1] ,
         \SB2_1_8/Component_Function_2/NAND4_in[0] ,
         \SB2_1_8/Component_Function_3/NAND4_in[2] ,
         \SB2_1_8/Component_Function_3/NAND4_in[1] ,
         \SB2_1_8/Component_Function_3/NAND4_in[0] ,
         \SB2_1_8/Component_Function_4/NAND4_in[3] ,
         \SB2_1_8/Component_Function_4/NAND4_in[2] ,
         \SB2_1_8/Component_Function_4/NAND4_in[1] ,
         \SB2_1_8/Component_Function_4/NAND4_in[0] ,
         \SB2_1_9/Component_Function_2/NAND4_in[2] ,
         \SB2_1_9/Component_Function_2/NAND4_in[1] ,
         \SB2_1_9/Component_Function_2/NAND4_in[0] ,
         \SB2_1_9/Component_Function_3/NAND4_in[3] ,
         \SB2_1_9/Component_Function_3/NAND4_in[2] ,
         \SB2_1_9/Component_Function_3/NAND4_in[1] ,
         \SB2_1_9/Component_Function_3/NAND4_in[0] ,
         \SB2_1_9/Component_Function_4/NAND4_in[3] ,
         \SB2_1_9/Component_Function_4/NAND4_in[2] ,
         \SB2_1_9/Component_Function_4/NAND4_in[1] ,
         \SB2_1_9/Component_Function_4/NAND4_in[0] ,
         \SB2_1_10/Component_Function_2/NAND4_in[3] ,
         \SB2_1_10/Component_Function_2/NAND4_in[1] ,
         \SB2_1_10/Component_Function_3/NAND4_in[2] ,
         \SB2_1_10/Component_Function_3/NAND4_in[1] ,
         \SB2_1_10/Component_Function_3/NAND4_in[0] ,
         \SB2_1_10/Component_Function_4/NAND4_in[3] ,
         \SB2_1_10/Component_Function_4/NAND4_in[2] ,
         \SB2_1_10/Component_Function_4/NAND4_in[1] ,
         \SB2_1_10/Component_Function_4/NAND4_in[0] ,
         \SB2_1_11/Component_Function_2/NAND4_in[2] ,
         \SB2_1_11/Component_Function_2/NAND4_in[1] ,
         \SB2_1_11/Component_Function_2/NAND4_in[0] ,
         \SB2_1_11/Component_Function_3/NAND4_in[3] ,
         \SB2_1_11/Component_Function_3/NAND4_in[2] ,
         \SB2_1_11/Component_Function_3/NAND4_in[1] ,
         \SB2_1_11/Component_Function_3/NAND4_in[0] ,
         \SB2_1_11/Component_Function_4/NAND4_in[2] ,
         \SB2_1_11/Component_Function_4/NAND4_in[1] ,
         \SB2_1_11/Component_Function_4/NAND4_in[0] ,
         \SB2_1_12/Component_Function_2/NAND4_in[3] ,
         \SB2_1_12/Component_Function_2/NAND4_in[1] ,
         \SB2_1_12/Component_Function_2/NAND4_in[0] ,
         \SB2_1_12/Component_Function_3/NAND4_in[3] ,
         \SB2_1_12/Component_Function_3/NAND4_in[2] ,
         \SB2_1_12/Component_Function_3/NAND4_in[1] ,
         \SB2_1_12/Component_Function_3/NAND4_in[0] ,
         \SB2_1_12/Component_Function_4/NAND4_in[3] ,
         \SB2_1_12/Component_Function_4/NAND4_in[2] ,
         \SB2_1_12/Component_Function_4/NAND4_in[1] ,
         \SB2_1_12/Component_Function_4/NAND4_in[0] ,
         \SB2_1_13/Component_Function_2/NAND4_in[3] ,
         \SB2_1_13/Component_Function_2/NAND4_in[2] ,
         \SB2_1_13/Component_Function_2/NAND4_in[1] ,
         \SB2_1_13/Component_Function_2/NAND4_in[0] ,
         \SB2_1_13/Component_Function_3/NAND4_in[2] ,
         \SB2_1_13/Component_Function_3/NAND4_in[1] ,
         \SB2_1_13/Component_Function_3/NAND4_in[0] ,
         \SB2_1_13/Component_Function_4/NAND4_in[3] ,
         \SB2_1_13/Component_Function_4/NAND4_in[2] ,
         \SB2_1_13/Component_Function_4/NAND4_in[1] ,
         \SB2_1_13/Component_Function_4/NAND4_in[0] ,
         \SB2_1_14/Component_Function_2/NAND4_in[2] ,
         \SB2_1_14/Component_Function_2/NAND4_in[1] ,
         \SB2_1_14/Component_Function_2/NAND4_in[0] ,
         \SB2_1_14/Component_Function_3/NAND4_in[3] ,
         \SB2_1_14/Component_Function_3/NAND4_in[2] ,
         \SB2_1_14/Component_Function_3/NAND4_in[1] ,
         \SB2_1_14/Component_Function_3/NAND4_in[0] ,
         \SB2_1_14/Component_Function_4/NAND4_in[2] ,
         \SB2_1_14/Component_Function_4/NAND4_in[1] ,
         \SB2_1_14/Component_Function_4/NAND4_in[0] ,
         \SB2_1_15/Component_Function_2/NAND4_in[3] ,
         \SB2_1_15/Component_Function_2/NAND4_in[1] ,
         \SB2_1_15/Component_Function_2/NAND4_in[0] ,
         \SB2_1_15/Component_Function_3/NAND4_in[3] ,
         \SB2_1_15/Component_Function_3/NAND4_in[2] ,
         \SB2_1_15/Component_Function_3/NAND4_in[1] ,
         \SB2_1_15/Component_Function_3/NAND4_in[0] ,
         \SB2_1_15/Component_Function_4/NAND4_in[2] ,
         \SB2_1_15/Component_Function_4/NAND4_in[1] ,
         \SB2_1_15/Component_Function_4/NAND4_in[0] ,
         \SB2_1_16/Component_Function_2/NAND4_in[3] ,
         \SB2_1_16/Component_Function_2/NAND4_in[1] ,
         \SB2_1_16/Component_Function_2/NAND4_in[0] ,
         \SB2_1_16/Component_Function_3/NAND4_in[2] ,
         \SB2_1_16/Component_Function_3/NAND4_in[1] ,
         \SB2_1_16/Component_Function_3/NAND4_in[0] ,
         \SB2_1_16/Component_Function_4/NAND4_in[3] ,
         \SB2_1_16/Component_Function_4/NAND4_in[2] ,
         \SB2_1_16/Component_Function_4/NAND4_in[1] ,
         \SB2_1_16/Component_Function_4/NAND4_in[0] ,
         \SB2_1_17/Component_Function_2/NAND4_in[2] ,
         \SB2_1_17/Component_Function_2/NAND4_in[1] ,
         \SB2_1_17/Component_Function_2/NAND4_in[0] ,
         \SB2_1_17/Component_Function_3/NAND4_in[2] ,
         \SB2_1_17/Component_Function_3/NAND4_in[0] ,
         \SB2_1_17/Component_Function_4/NAND4_in[3] ,
         \SB2_1_17/Component_Function_4/NAND4_in[2] ,
         \SB2_1_17/Component_Function_4/NAND4_in[1] ,
         \SB2_1_17/Component_Function_4/NAND4_in[0] ,
         \SB2_1_18/Component_Function_2/NAND4_in[2] ,
         \SB2_1_18/Component_Function_2/NAND4_in[1] ,
         \SB2_1_18/Component_Function_2/NAND4_in[0] ,
         \SB2_1_18/Component_Function_3/NAND4_in[3] ,
         \SB2_1_18/Component_Function_3/NAND4_in[2] ,
         \SB2_1_18/Component_Function_3/NAND4_in[1] ,
         \SB2_1_18/Component_Function_3/NAND4_in[0] ,
         \SB2_1_18/Component_Function_4/NAND4_in[3] ,
         \SB2_1_18/Component_Function_4/NAND4_in[2] ,
         \SB2_1_18/Component_Function_4/NAND4_in[1] ,
         \SB2_1_18/Component_Function_4/NAND4_in[0] ,
         \SB2_1_19/Component_Function_2/NAND4_in[2] ,
         \SB2_1_19/Component_Function_2/NAND4_in[1] ,
         \SB2_1_19/Component_Function_2/NAND4_in[0] ,
         \SB2_1_19/Component_Function_3/NAND4_in[2] ,
         \SB2_1_19/Component_Function_3/NAND4_in[1] ,
         \SB2_1_19/Component_Function_3/NAND4_in[0] ,
         \SB2_1_19/Component_Function_4/NAND4_in[3] ,
         \SB2_1_19/Component_Function_4/NAND4_in[1] ,
         \SB2_1_19/Component_Function_4/NAND4_in[0] ,
         \SB2_1_20/Component_Function_2/NAND4_in[2] ,
         \SB2_1_20/Component_Function_2/NAND4_in[1] ,
         \SB2_1_20/Component_Function_2/NAND4_in[0] ,
         \SB2_1_20/Component_Function_3/NAND4_in[2] ,
         \SB2_1_20/Component_Function_3/NAND4_in[1] ,
         \SB2_1_20/Component_Function_3/NAND4_in[0] ,
         \SB2_1_20/Component_Function_4/NAND4_in[2] ,
         \SB2_1_20/Component_Function_4/NAND4_in[1] ,
         \SB2_1_20/Component_Function_4/NAND4_in[0] ,
         \SB2_1_21/Component_Function_2/NAND4_in[3] ,
         \SB2_1_21/Component_Function_2/NAND4_in[1] ,
         \SB2_1_21/Component_Function_2/NAND4_in[0] ,
         \SB2_1_21/Component_Function_3/NAND4_in[3] ,
         \SB2_1_21/Component_Function_3/NAND4_in[1] ,
         \SB2_1_21/Component_Function_3/NAND4_in[0] ,
         \SB2_1_21/Component_Function_4/NAND4_in[3] ,
         \SB2_1_21/Component_Function_4/NAND4_in[2] ,
         \SB2_1_21/Component_Function_4/NAND4_in[1] ,
         \SB2_1_21/Component_Function_4/NAND4_in[0] ,
         \SB2_1_22/Component_Function_2/NAND4_in[2] ,
         \SB2_1_22/Component_Function_2/NAND4_in[1] ,
         \SB2_1_22/Component_Function_2/NAND4_in[0] ,
         \SB2_1_22/Component_Function_3/NAND4_in[2] ,
         \SB2_1_22/Component_Function_3/NAND4_in[0] ,
         \SB2_1_22/Component_Function_4/NAND4_in[3] ,
         \SB2_1_22/Component_Function_4/NAND4_in[1] ,
         \SB2_1_22/Component_Function_4/NAND4_in[0] ,
         \SB2_1_23/Component_Function_2/NAND4_in[3] ,
         \SB2_1_23/Component_Function_2/NAND4_in[1] ,
         \SB2_1_23/Component_Function_2/NAND4_in[0] ,
         \SB2_1_23/Component_Function_3/NAND4_in[3] ,
         \SB2_1_23/Component_Function_3/NAND4_in[2] ,
         \SB2_1_23/Component_Function_3/NAND4_in[1] ,
         \SB2_1_23/Component_Function_3/NAND4_in[0] ,
         \SB2_1_23/Component_Function_4/NAND4_in[3] ,
         \SB2_1_23/Component_Function_4/NAND4_in[2] ,
         \SB2_1_23/Component_Function_4/NAND4_in[1] ,
         \SB2_1_23/Component_Function_4/NAND4_in[0] ,
         \SB2_1_24/Component_Function_2/NAND4_in[2] ,
         \SB2_1_24/Component_Function_2/NAND4_in[1] ,
         \SB2_1_24/Component_Function_2/NAND4_in[0] ,
         \SB2_1_24/Component_Function_3/NAND4_in[3] ,
         \SB2_1_24/Component_Function_3/NAND4_in[2] ,
         \SB2_1_24/Component_Function_3/NAND4_in[1] ,
         \SB2_1_24/Component_Function_3/NAND4_in[0] ,
         \SB2_1_24/Component_Function_4/NAND4_in[3] ,
         \SB2_1_24/Component_Function_4/NAND4_in[2] ,
         \SB2_1_24/Component_Function_4/NAND4_in[1] ,
         \SB2_1_24/Component_Function_4/NAND4_in[0] ,
         \SB2_1_25/Component_Function_2/NAND4_in[3] ,
         \SB2_1_25/Component_Function_2/NAND4_in[2] ,
         \SB2_1_25/Component_Function_2/NAND4_in[1] ,
         \SB2_1_25/Component_Function_2/NAND4_in[0] ,
         \SB2_1_25/Component_Function_3/NAND4_in[2] ,
         \SB2_1_25/Component_Function_3/NAND4_in[1] ,
         \SB2_1_25/Component_Function_3/NAND4_in[0] ,
         \SB2_1_25/Component_Function_4/NAND4_in[3] ,
         \SB2_1_25/Component_Function_4/NAND4_in[2] ,
         \SB2_1_25/Component_Function_4/NAND4_in[1] ,
         \SB2_1_25/Component_Function_4/NAND4_in[0] ,
         \SB2_1_26/Component_Function_2/NAND4_in[3] ,
         \SB2_1_26/Component_Function_2/NAND4_in[2] ,
         \SB2_1_26/Component_Function_2/NAND4_in[1] ,
         \SB2_1_26/Component_Function_3/NAND4_in[2] ,
         \SB2_1_26/Component_Function_3/NAND4_in[1] ,
         \SB2_1_26/Component_Function_3/NAND4_in[0] ,
         \SB2_1_26/Component_Function_4/NAND4_in[3] ,
         \SB2_1_26/Component_Function_4/NAND4_in[2] ,
         \SB2_1_26/Component_Function_4/NAND4_in[1] ,
         \SB2_1_26/Component_Function_4/NAND4_in[0] ,
         \SB2_1_27/Component_Function_2/NAND4_in[3] ,
         \SB2_1_27/Component_Function_2/NAND4_in[2] ,
         \SB2_1_27/Component_Function_2/NAND4_in[1] ,
         \SB2_1_27/Component_Function_2/NAND4_in[0] ,
         \SB2_1_27/Component_Function_3/NAND4_in[3] ,
         \SB2_1_27/Component_Function_3/NAND4_in[2] ,
         \SB2_1_27/Component_Function_3/NAND4_in[1] ,
         \SB2_1_27/Component_Function_3/NAND4_in[0] ,
         \SB2_1_27/Component_Function_4/NAND4_in[3] ,
         \SB2_1_27/Component_Function_4/NAND4_in[1] ,
         \SB2_1_27/Component_Function_4/NAND4_in[0] ,
         \SB2_1_28/Component_Function_2/NAND4_in[3] ,
         \SB2_1_28/Component_Function_2/NAND4_in[1] ,
         \SB2_1_28/Component_Function_2/NAND4_in[0] ,
         \SB2_1_28/Component_Function_3/NAND4_in[3] ,
         \SB2_1_28/Component_Function_3/NAND4_in[2] ,
         \SB2_1_28/Component_Function_3/NAND4_in[1] ,
         \SB2_1_28/Component_Function_3/NAND4_in[0] ,
         \SB2_1_28/Component_Function_4/NAND4_in[3] ,
         \SB2_1_28/Component_Function_4/NAND4_in[1] ,
         \SB2_1_28/Component_Function_4/NAND4_in[0] ,
         \SB2_1_29/Component_Function_2/NAND4_in[2] ,
         \SB2_1_29/Component_Function_2/NAND4_in[1] ,
         \SB2_1_29/Component_Function_2/NAND4_in[0] ,
         \SB2_1_29/Component_Function_3/NAND4_in[2] ,
         \SB2_1_29/Component_Function_3/NAND4_in[0] ,
         \SB2_1_29/Component_Function_4/NAND4_in[2] ,
         \SB2_1_29/Component_Function_4/NAND4_in[1] ,
         \SB2_1_29/Component_Function_4/NAND4_in[0] ,
         \SB2_1_30/Component_Function_2/NAND4_in[2] ,
         \SB2_1_30/Component_Function_2/NAND4_in[1] ,
         \SB2_1_30/Component_Function_2/NAND4_in[0] ,
         \SB2_1_30/Component_Function_3/NAND4_in[3] ,
         \SB2_1_30/Component_Function_3/NAND4_in[2] ,
         \SB2_1_30/Component_Function_3/NAND4_in[1] ,
         \SB2_1_30/Component_Function_3/NAND4_in[0] ,
         \SB2_1_30/Component_Function_4/NAND4_in[3] ,
         \SB2_1_30/Component_Function_4/NAND4_in[1] ,
         \SB2_1_30/Component_Function_4/NAND4_in[0] ,
         \SB2_1_31/Component_Function_2/NAND4_in[3] ,
         \SB2_1_31/Component_Function_2/NAND4_in[2] ,
         \SB2_1_31/Component_Function_2/NAND4_in[1] ,
         \SB2_1_31/Component_Function_2/NAND4_in[0] ,
         \SB2_1_31/Component_Function_3/NAND4_in[3] ,
         \SB2_1_31/Component_Function_3/NAND4_in[2] ,
         \SB2_1_31/Component_Function_3/NAND4_in[1] ,
         \SB2_1_31/Component_Function_3/NAND4_in[0] ,
         \SB2_1_31/Component_Function_4/NAND4_in[3] ,
         \SB2_1_31/Component_Function_4/NAND4_in[1] ,
         \SB2_1_31/Component_Function_4/NAND4_in[0] ,
         \SB1_2_0/Component_Function_2/NAND4_in[2] ,
         \SB1_2_0/Component_Function_2/NAND4_in[1] ,
         \SB1_2_0/Component_Function_2/NAND4_in[0] ,
         \SB1_2_0/Component_Function_3/NAND4_in[3] ,
         \SB1_2_0/Component_Function_3/NAND4_in[2] ,
         \SB1_2_0/Component_Function_3/NAND4_in[1] ,
         \SB1_2_0/Component_Function_3/NAND4_in[0] ,
         \SB1_2_0/Component_Function_4/NAND4_in[3] ,
         \SB1_2_0/Component_Function_4/NAND4_in[2] ,
         \SB1_2_0/Component_Function_4/NAND4_in[1] ,
         \SB1_2_0/Component_Function_4/NAND4_in[0] ,
         \SB1_2_1/Component_Function_2/NAND4_in[2] ,
         \SB1_2_1/Component_Function_2/NAND4_in[1] ,
         \SB1_2_1/Component_Function_2/NAND4_in[0] ,
         \SB1_2_1/Component_Function_3/NAND4_in[2] ,
         \SB1_2_1/Component_Function_3/NAND4_in[1] ,
         \SB1_2_1/Component_Function_3/NAND4_in[0] ,
         \SB1_2_1/Component_Function_4/NAND4_in[3] ,
         \SB1_2_1/Component_Function_4/NAND4_in[2] ,
         \SB1_2_1/Component_Function_4/NAND4_in[1] ,
         \SB1_2_1/Component_Function_4/NAND4_in[0] ,
         \SB1_2_2/Component_Function_2/NAND4_in[3] ,
         \SB1_2_2/Component_Function_2/NAND4_in[2] ,
         \SB1_2_2/Component_Function_2/NAND4_in[1] ,
         \SB1_2_2/Component_Function_2/NAND4_in[0] ,
         \SB1_2_2/Component_Function_3/NAND4_in[3] ,
         \SB1_2_2/Component_Function_3/NAND4_in[2] ,
         \SB1_2_2/Component_Function_3/NAND4_in[1] ,
         \SB1_2_2/Component_Function_3/NAND4_in[0] ,
         \SB1_2_2/Component_Function_4/NAND4_in[3] ,
         \SB1_2_2/Component_Function_4/NAND4_in[2] ,
         \SB1_2_2/Component_Function_4/NAND4_in[1] ,
         \SB1_2_2/Component_Function_4/NAND4_in[0] ,
         \SB1_2_3/Component_Function_2/NAND4_in[2] ,
         \SB1_2_3/Component_Function_2/NAND4_in[1] ,
         \SB1_2_3/Component_Function_2/NAND4_in[0] ,
         \SB1_2_3/Component_Function_3/NAND4_in[3] ,
         \SB1_2_3/Component_Function_3/NAND4_in[2] ,
         \SB1_2_3/Component_Function_3/NAND4_in[1] ,
         \SB1_2_3/Component_Function_3/NAND4_in[0] ,
         \SB1_2_3/Component_Function_4/NAND4_in[3] ,
         \SB1_2_3/Component_Function_4/NAND4_in[2] ,
         \SB1_2_3/Component_Function_4/NAND4_in[1] ,
         \SB1_2_3/Component_Function_4/NAND4_in[0] ,
         \SB1_2_4/Component_Function_2/NAND4_in[3] ,
         \SB1_2_4/Component_Function_2/NAND4_in[2] ,
         \SB1_2_4/Component_Function_2/NAND4_in[1] ,
         \SB1_2_4/Component_Function_2/NAND4_in[0] ,
         \SB1_2_4/Component_Function_3/NAND4_in[3] ,
         \SB1_2_4/Component_Function_3/NAND4_in[2] ,
         \SB1_2_4/Component_Function_3/NAND4_in[1] ,
         \SB1_2_4/Component_Function_3/NAND4_in[0] ,
         \SB1_2_4/Component_Function_4/NAND4_in[3] ,
         \SB1_2_4/Component_Function_4/NAND4_in[2] ,
         \SB1_2_4/Component_Function_4/NAND4_in[1] ,
         \SB1_2_4/Component_Function_4/NAND4_in[0] ,
         \SB1_2_5/Component_Function_2/NAND4_in[2] ,
         \SB1_2_5/Component_Function_2/NAND4_in[1] ,
         \SB1_2_5/Component_Function_2/NAND4_in[0] ,
         \SB1_2_5/Component_Function_3/NAND4_in[3] ,
         \SB1_2_5/Component_Function_3/NAND4_in[2] ,
         \SB1_2_5/Component_Function_3/NAND4_in[1] ,
         \SB1_2_5/Component_Function_3/NAND4_in[0] ,
         \SB1_2_5/Component_Function_4/NAND4_in[3] ,
         \SB1_2_5/Component_Function_4/NAND4_in[2] ,
         \SB1_2_5/Component_Function_4/NAND4_in[1] ,
         \SB1_2_5/Component_Function_4/NAND4_in[0] ,
         \SB1_2_6/Component_Function_2/NAND4_in[2] ,
         \SB1_2_6/Component_Function_2/NAND4_in[1] ,
         \SB1_2_6/Component_Function_2/NAND4_in[0] ,
         \SB1_2_6/Component_Function_3/NAND4_in[3] ,
         \SB1_2_6/Component_Function_3/NAND4_in[2] ,
         \SB1_2_6/Component_Function_3/NAND4_in[1] ,
         \SB1_2_6/Component_Function_3/NAND4_in[0] ,
         \SB1_2_6/Component_Function_4/NAND4_in[3] ,
         \SB1_2_6/Component_Function_4/NAND4_in[2] ,
         \SB1_2_6/Component_Function_4/NAND4_in[1] ,
         \SB1_2_6/Component_Function_4/NAND4_in[0] ,
         \SB1_2_7/Component_Function_2/NAND4_in[2] ,
         \SB1_2_7/Component_Function_2/NAND4_in[1] ,
         \SB1_2_7/Component_Function_2/NAND4_in[0] ,
         \SB1_2_7/Component_Function_3/NAND4_in[3] ,
         \SB1_2_7/Component_Function_3/NAND4_in[2] ,
         \SB1_2_7/Component_Function_3/NAND4_in[1] ,
         \SB1_2_7/Component_Function_3/NAND4_in[0] ,
         \SB1_2_7/Component_Function_4/NAND4_in[3] ,
         \SB1_2_7/Component_Function_4/NAND4_in[2] ,
         \SB1_2_7/Component_Function_4/NAND4_in[1] ,
         \SB1_2_7/Component_Function_4/NAND4_in[0] ,
         \SB1_2_8/Component_Function_2/NAND4_in[3] ,
         \SB1_2_8/Component_Function_2/NAND4_in[2] ,
         \SB1_2_8/Component_Function_2/NAND4_in[1] ,
         \SB1_2_8/Component_Function_2/NAND4_in[0] ,
         \SB1_2_8/Component_Function_3/NAND4_in[3] ,
         \SB1_2_8/Component_Function_3/NAND4_in[2] ,
         \SB1_2_8/Component_Function_3/NAND4_in[1] ,
         \SB1_2_8/Component_Function_3/NAND4_in[0] ,
         \SB1_2_8/Component_Function_4/NAND4_in[3] ,
         \SB1_2_8/Component_Function_4/NAND4_in[2] ,
         \SB1_2_8/Component_Function_4/NAND4_in[1] ,
         \SB1_2_8/Component_Function_4/NAND4_in[0] ,
         \SB1_2_9/Component_Function_2/NAND4_in[2] ,
         \SB1_2_9/Component_Function_2/NAND4_in[1] ,
         \SB1_2_9/Component_Function_2/NAND4_in[0] ,
         \SB1_2_9/Component_Function_3/NAND4_in[3] ,
         \SB1_2_9/Component_Function_3/NAND4_in[2] ,
         \SB1_2_9/Component_Function_3/NAND4_in[1] ,
         \SB1_2_9/Component_Function_3/NAND4_in[0] ,
         \SB1_2_9/Component_Function_4/NAND4_in[3] ,
         \SB1_2_9/Component_Function_4/NAND4_in[2] ,
         \SB1_2_9/Component_Function_4/NAND4_in[1] ,
         \SB1_2_9/Component_Function_4/NAND4_in[0] ,
         \SB1_2_10/Component_Function_2/NAND4_in[2] ,
         \SB1_2_10/Component_Function_2/NAND4_in[1] ,
         \SB1_2_10/Component_Function_2/NAND4_in[0] ,
         \SB1_2_10/Component_Function_3/NAND4_in[3] ,
         \SB1_2_10/Component_Function_3/NAND4_in[2] ,
         \SB1_2_10/Component_Function_3/NAND4_in[1] ,
         \SB1_2_10/Component_Function_3/NAND4_in[0] ,
         \SB1_2_10/Component_Function_4/NAND4_in[3] ,
         \SB1_2_10/Component_Function_4/NAND4_in[2] ,
         \SB1_2_10/Component_Function_4/NAND4_in[1] ,
         \SB1_2_10/Component_Function_4/NAND4_in[0] ,
         \SB1_2_11/Component_Function_2/NAND4_in[2] ,
         \SB1_2_11/Component_Function_2/NAND4_in[1] ,
         \SB1_2_11/Component_Function_2/NAND4_in[0] ,
         \SB1_2_11/Component_Function_3/NAND4_in[3] ,
         \SB1_2_11/Component_Function_3/NAND4_in[2] ,
         \SB1_2_11/Component_Function_3/NAND4_in[1] ,
         \SB1_2_11/Component_Function_3/NAND4_in[0] ,
         \SB1_2_11/Component_Function_4/NAND4_in[3] ,
         \SB1_2_11/Component_Function_4/NAND4_in[2] ,
         \SB1_2_11/Component_Function_4/NAND4_in[1] ,
         \SB1_2_11/Component_Function_4/NAND4_in[0] ,
         \SB1_2_12/Component_Function_2/NAND4_in[3] ,
         \SB1_2_12/Component_Function_2/NAND4_in[2] ,
         \SB1_2_12/Component_Function_2/NAND4_in[1] ,
         \SB1_2_12/Component_Function_2/NAND4_in[0] ,
         \SB1_2_12/Component_Function_3/NAND4_in[3] ,
         \SB1_2_12/Component_Function_3/NAND4_in[2] ,
         \SB1_2_12/Component_Function_3/NAND4_in[1] ,
         \SB1_2_12/Component_Function_3/NAND4_in[0] ,
         \SB1_2_12/Component_Function_4/NAND4_in[3] ,
         \SB1_2_12/Component_Function_4/NAND4_in[2] ,
         \SB1_2_12/Component_Function_4/NAND4_in[1] ,
         \SB1_2_12/Component_Function_4/NAND4_in[0] ,
         \SB1_2_13/Component_Function_2/NAND4_in[2] ,
         \SB1_2_13/Component_Function_2/NAND4_in[1] ,
         \SB1_2_13/Component_Function_2/NAND4_in[0] ,
         \SB1_2_13/Component_Function_3/NAND4_in[3] ,
         \SB1_2_13/Component_Function_3/NAND4_in[2] ,
         \SB1_2_13/Component_Function_3/NAND4_in[1] ,
         \SB1_2_13/Component_Function_3/NAND4_in[0] ,
         \SB1_2_13/Component_Function_4/NAND4_in[3] ,
         \SB1_2_13/Component_Function_4/NAND4_in[2] ,
         \SB1_2_13/Component_Function_4/NAND4_in[1] ,
         \SB1_2_13/Component_Function_4/NAND4_in[0] ,
         \SB1_2_14/Component_Function_2/NAND4_in[2] ,
         \SB1_2_14/Component_Function_2/NAND4_in[1] ,
         \SB1_2_14/Component_Function_2/NAND4_in[0] ,
         \SB1_2_14/Component_Function_3/NAND4_in[3] ,
         \SB1_2_14/Component_Function_3/NAND4_in[2] ,
         \SB1_2_14/Component_Function_3/NAND4_in[1] ,
         \SB1_2_14/Component_Function_3/NAND4_in[0] ,
         \SB1_2_14/Component_Function_4/NAND4_in[3] ,
         \SB1_2_14/Component_Function_4/NAND4_in[1] ,
         \SB1_2_14/Component_Function_4/NAND4_in[0] ,
         \SB1_2_15/Component_Function_2/NAND4_in[2] ,
         \SB1_2_15/Component_Function_2/NAND4_in[1] ,
         \SB1_2_15/Component_Function_2/NAND4_in[0] ,
         \SB1_2_15/Component_Function_3/NAND4_in[3] ,
         \SB1_2_15/Component_Function_3/NAND4_in[2] ,
         \SB1_2_15/Component_Function_3/NAND4_in[1] ,
         \SB1_2_15/Component_Function_3/NAND4_in[0] ,
         \SB1_2_15/Component_Function_4/NAND4_in[3] ,
         \SB1_2_15/Component_Function_4/NAND4_in[2] ,
         \SB1_2_15/Component_Function_4/NAND4_in[1] ,
         \SB1_2_15/Component_Function_4/NAND4_in[0] ,
         \SB1_2_16/Component_Function_2/NAND4_in[2] ,
         \SB1_2_16/Component_Function_2/NAND4_in[1] ,
         \SB1_2_16/Component_Function_2/NAND4_in[0] ,
         \SB1_2_16/Component_Function_3/NAND4_in[3] ,
         \SB1_2_16/Component_Function_3/NAND4_in[2] ,
         \SB1_2_16/Component_Function_3/NAND4_in[1] ,
         \SB1_2_16/Component_Function_3/NAND4_in[0] ,
         \SB1_2_16/Component_Function_4/NAND4_in[3] ,
         \SB1_2_16/Component_Function_4/NAND4_in[2] ,
         \SB1_2_16/Component_Function_4/NAND4_in[1] ,
         \SB1_2_16/Component_Function_4/NAND4_in[0] ,
         \SB1_2_17/Component_Function_2/NAND4_in[3] ,
         \SB1_2_17/Component_Function_2/NAND4_in[2] ,
         \SB1_2_17/Component_Function_2/NAND4_in[1] ,
         \SB1_2_17/Component_Function_2/NAND4_in[0] ,
         \SB1_2_17/Component_Function_3/NAND4_in[3] ,
         \SB1_2_17/Component_Function_3/NAND4_in[2] ,
         \SB1_2_17/Component_Function_3/NAND4_in[1] ,
         \SB1_2_17/Component_Function_3/NAND4_in[0] ,
         \SB1_2_17/Component_Function_4/NAND4_in[3] ,
         \SB1_2_17/Component_Function_4/NAND4_in[2] ,
         \SB1_2_17/Component_Function_4/NAND4_in[1] ,
         \SB1_2_17/Component_Function_4/NAND4_in[0] ,
         \SB1_2_18/Component_Function_2/NAND4_in[2] ,
         \SB1_2_18/Component_Function_2/NAND4_in[1] ,
         \SB1_2_18/Component_Function_2/NAND4_in[0] ,
         \SB1_2_18/Component_Function_3/NAND4_in[3] ,
         \SB1_2_18/Component_Function_3/NAND4_in[2] ,
         \SB1_2_18/Component_Function_3/NAND4_in[1] ,
         \SB1_2_18/Component_Function_3/NAND4_in[0] ,
         \SB1_2_18/Component_Function_4/NAND4_in[3] ,
         \SB1_2_18/Component_Function_4/NAND4_in[2] ,
         \SB1_2_18/Component_Function_4/NAND4_in[1] ,
         \SB1_2_18/Component_Function_4/NAND4_in[0] ,
         \SB1_2_19/Component_Function_2/NAND4_in[2] ,
         \SB1_2_19/Component_Function_2/NAND4_in[1] ,
         \SB1_2_19/Component_Function_2/NAND4_in[0] ,
         \SB1_2_19/Component_Function_3/NAND4_in[3] ,
         \SB1_2_19/Component_Function_3/NAND4_in[2] ,
         \SB1_2_19/Component_Function_3/NAND4_in[1] ,
         \SB1_2_19/Component_Function_3/NAND4_in[0] ,
         \SB1_2_19/Component_Function_4/NAND4_in[3] ,
         \SB1_2_19/Component_Function_4/NAND4_in[1] ,
         \SB1_2_19/Component_Function_4/NAND4_in[0] ,
         \SB1_2_20/Component_Function_2/NAND4_in[3] ,
         \SB1_2_20/Component_Function_2/NAND4_in[2] ,
         \SB1_2_20/Component_Function_2/NAND4_in[1] ,
         \SB1_2_20/Component_Function_2/NAND4_in[0] ,
         \SB1_2_20/Component_Function_3/NAND4_in[3] ,
         \SB1_2_20/Component_Function_3/NAND4_in[2] ,
         \SB1_2_20/Component_Function_3/NAND4_in[1] ,
         \SB1_2_20/Component_Function_3/NAND4_in[0] ,
         \SB1_2_20/Component_Function_4/NAND4_in[3] ,
         \SB1_2_20/Component_Function_4/NAND4_in[2] ,
         \SB1_2_20/Component_Function_4/NAND4_in[1] ,
         \SB1_2_20/Component_Function_4/NAND4_in[0] ,
         \SB1_2_21/Component_Function_2/NAND4_in[2] ,
         \SB1_2_21/Component_Function_2/NAND4_in[1] ,
         \SB1_2_21/Component_Function_2/NAND4_in[0] ,
         \SB1_2_21/Component_Function_3/NAND4_in[3] ,
         \SB1_2_21/Component_Function_3/NAND4_in[2] ,
         \SB1_2_21/Component_Function_3/NAND4_in[1] ,
         \SB1_2_21/Component_Function_3/NAND4_in[0] ,
         \SB1_2_21/Component_Function_4/NAND4_in[3] ,
         \SB1_2_21/Component_Function_4/NAND4_in[2] ,
         \SB1_2_21/Component_Function_4/NAND4_in[1] ,
         \SB1_2_21/Component_Function_4/NAND4_in[0] ,
         \SB1_2_22/Component_Function_2/NAND4_in[3] ,
         \SB1_2_22/Component_Function_2/NAND4_in[2] ,
         \SB1_2_22/Component_Function_2/NAND4_in[1] ,
         \SB1_2_22/Component_Function_2/NAND4_in[0] ,
         \SB1_2_22/Component_Function_3/NAND4_in[3] ,
         \SB1_2_22/Component_Function_3/NAND4_in[2] ,
         \SB1_2_22/Component_Function_3/NAND4_in[1] ,
         \SB1_2_22/Component_Function_3/NAND4_in[0] ,
         \SB1_2_22/Component_Function_4/NAND4_in[3] ,
         \SB1_2_22/Component_Function_4/NAND4_in[1] ,
         \SB1_2_22/Component_Function_4/NAND4_in[0] ,
         \SB1_2_23/Component_Function_2/NAND4_in[2] ,
         \SB1_2_23/Component_Function_2/NAND4_in[1] ,
         \SB1_2_23/Component_Function_2/NAND4_in[0] ,
         \SB1_2_23/Component_Function_3/NAND4_in[3] ,
         \SB1_2_23/Component_Function_3/NAND4_in[2] ,
         \SB1_2_23/Component_Function_3/NAND4_in[1] ,
         \SB1_2_23/Component_Function_3/NAND4_in[0] ,
         \SB1_2_23/Component_Function_4/NAND4_in[3] ,
         \SB1_2_23/Component_Function_4/NAND4_in[2] ,
         \SB1_2_23/Component_Function_4/NAND4_in[1] ,
         \SB1_2_23/Component_Function_4/NAND4_in[0] ,
         \SB1_2_24/Component_Function_2/NAND4_in[2] ,
         \SB1_2_24/Component_Function_2/NAND4_in[1] ,
         \SB1_2_24/Component_Function_2/NAND4_in[0] ,
         \SB1_2_24/Component_Function_3/NAND4_in[3] ,
         \SB1_2_24/Component_Function_3/NAND4_in[2] ,
         \SB1_2_24/Component_Function_3/NAND4_in[1] ,
         \SB1_2_24/Component_Function_3/NAND4_in[0] ,
         \SB1_2_24/Component_Function_4/NAND4_in[3] ,
         \SB1_2_24/Component_Function_4/NAND4_in[1] ,
         \SB1_2_24/Component_Function_4/NAND4_in[0] ,
         \SB1_2_25/Component_Function_2/NAND4_in[2] ,
         \SB1_2_25/Component_Function_2/NAND4_in[1] ,
         \SB1_2_25/Component_Function_2/NAND4_in[0] ,
         \SB1_2_25/Component_Function_3/NAND4_in[3] ,
         \SB1_2_25/Component_Function_3/NAND4_in[2] ,
         \SB1_2_25/Component_Function_3/NAND4_in[1] ,
         \SB1_2_25/Component_Function_3/NAND4_in[0] ,
         \SB1_2_25/Component_Function_4/NAND4_in[3] ,
         \SB1_2_25/Component_Function_4/NAND4_in[1] ,
         \SB1_2_25/Component_Function_4/NAND4_in[0] ,
         \SB1_2_26/Component_Function_2/NAND4_in[2] ,
         \SB1_2_26/Component_Function_2/NAND4_in[1] ,
         \SB1_2_26/Component_Function_2/NAND4_in[0] ,
         \SB1_2_26/Component_Function_3/NAND4_in[3] ,
         \SB1_2_26/Component_Function_3/NAND4_in[2] ,
         \SB1_2_26/Component_Function_3/NAND4_in[1] ,
         \SB1_2_26/Component_Function_3/NAND4_in[0] ,
         \SB1_2_26/Component_Function_4/NAND4_in[3] ,
         \SB1_2_26/Component_Function_4/NAND4_in[2] ,
         \SB1_2_26/Component_Function_4/NAND4_in[1] ,
         \SB1_2_26/Component_Function_4/NAND4_in[0] ,
         \SB1_2_27/Component_Function_2/NAND4_in[2] ,
         \SB1_2_27/Component_Function_2/NAND4_in[1] ,
         \SB1_2_27/Component_Function_2/NAND4_in[0] ,
         \SB1_2_27/Component_Function_3/NAND4_in[3] ,
         \SB1_2_27/Component_Function_3/NAND4_in[2] ,
         \SB1_2_27/Component_Function_3/NAND4_in[1] ,
         \SB1_2_27/Component_Function_3/NAND4_in[0] ,
         \SB1_2_27/Component_Function_4/NAND4_in[3] ,
         \SB1_2_27/Component_Function_4/NAND4_in[2] ,
         \SB1_2_27/Component_Function_4/NAND4_in[1] ,
         \SB1_2_27/Component_Function_4/NAND4_in[0] ,
         \SB1_2_28/Component_Function_2/NAND4_in[2] ,
         \SB1_2_28/Component_Function_2/NAND4_in[1] ,
         \SB1_2_28/Component_Function_2/NAND4_in[0] ,
         \SB1_2_28/Component_Function_3/NAND4_in[3] ,
         \SB1_2_28/Component_Function_3/NAND4_in[2] ,
         \SB1_2_28/Component_Function_3/NAND4_in[1] ,
         \SB1_2_28/Component_Function_3/NAND4_in[0] ,
         \SB1_2_28/Component_Function_4/NAND4_in[3] ,
         \SB1_2_28/Component_Function_4/NAND4_in[2] ,
         \SB1_2_28/Component_Function_4/NAND4_in[1] ,
         \SB1_2_28/Component_Function_4/NAND4_in[0] ,
         \SB1_2_29/Component_Function_2/NAND4_in[3] ,
         \SB1_2_29/Component_Function_2/NAND4_in[2] ,
         \SB1_2_29/Component_Function_2/NAND4_in[1] ,
         \SB1_2_29/Component_Function_2/NAND4_in[0] ,
         \SB1_2_29/Component_Function_3/NAND4_in[3] ,
         \SB1_2_29/Component_Function_3/NAND4_in[2] ,
         \SB1_2_29/Component_Function_3/NAND4_in[1] ,
         \SB1_2_29/Component_Function_3/NAND4_in[0] ,
         \SB1_2_29/Component_Function_4/NAND4_in[3] ,
         \SB1_2_29/Component_Function_4/NAND4_in[2] ,
         \SB1_2_29/Component_Function_4/NAND4_in[1] ,
         \SB1_2_29/Component_Function_4/NAND4_in[0] ,
         \SB1_2_30/Component_Function_2/NAND4_in[2] ,
         \SB1_2_30/Component_Function_2/NAND4_in[1] ,
         \SB1_2_30/Component_Function_2/NAND4_in[0] ,
         \SB1_2_30/Component_Function_3/NAND4_in[3] ,
         \SB1_2_30/Component_Function_3/NAND4_in[2] ,
         \SB1_2_30/Component_Function_3/NAND4_in[1] ,
         \SB1_2_30/Component_Function_3/NAND4_in[0] ,
         \SB1_2_30/Component_Function_4/NAND4_in[3] ,
         \SB1_2_30/Component_Function_4/NAND4_in[2] ,
         \SB1_2_30/Component_Function_4/NAND4_in[1] ,
         \SB1_2_30/Component_Function_4/NAND4_in[0] ,
         \SB1_2_31/Component_Function_2/NAND4_in[3] ,
         \SB1_2_31/Component_Function_2/NAND4_in[1] ,
         \SB1_2_31/Component_Function_2/NAND4_in[0] ,
         \SB1_2_31/Component_Function_3/NAND4_in[2] ,
         \SB1_2_31/Component_Function_3/NAND4_in[1] ,
         \SB1_2_31/Component_Function_3/NAND4_in[0] ,
         \SB1_2_31/Component_Function_4/NAND4_in[3] ,
         \SB1_2_31/Component_Function_4/NAND4_in[2] ,
         \SB1_2_31/Component_Function_4/NAND4_in[1] ,
         \SB1_2_31/Component_Function_4/NAND4_in[0] ,
         \SB2_2_0/Component_Function_2/NAND4_in[2] ,
         \SB2_2_0/Component_Function_2/NAND4_in[1] ,
         \SB2_2_0/Component_Function_2/NAND4_in[0] ,
         \SB2_2_0/Component_Function_3/NAND4_in[3] ,
         \SB2_2_0/Component_Function_3/NAND4_in[2] ,
         \SB2_2_0/Component_Function_3/NAND4_in[1] ,
         \SB2_2_0/Component_Function_3/NAND4_in[0] ,
         \SB2_2_0/Component_Function_4/NAND4_in[3] ,
         \SB2_2_0/Component_Function_4/NAND4_in[1] ,
         \SB2_2_0/Component_Function_4/NAND4_in[0] ,
         \SB2_2_1/Component_Function_2/NAND4_in[2] ,
         \SB2_2_1/Component_Function_2/NAND4_in[1] ,
         \SB2_2_1/Component_Function_2/NAND4_in[0] ,
         \SB2_2_1/Component_Function_3/NAND4_in[2] ,
         \SB2_2_1/Component_Function_3/NAND4_in[1] ,
         \SB2_2_1/Component_Function_3/NAND4_in[0] ,
         \SB2_2_1/Component_Function_4/NAND4_in[2] ,
         \SB2_2_1/Component_Function_4/NAND4_in[1] ,
         \SB2_2_1/Component_Function_4/NAND4_in[0] ,
         \SB2_2_2/Component_Function_2/NAND4_in[2] ,
         \SB2_2_2/Component_Function_2/NAND4_in[1] ,
         \SB2_2_2/Component_Function_2/NAND4_in[0] ,
         \SB2_2_2/Component_Function_3/NAND4_in[2] ,
         \SB2_2_2/Component_Function_3/NAND4_in[1] ,
         \SB2_2_2/Component_Function_3/NAND4_in[0] ,
         \SB2_2_2/Component_Function_4/NAND4_in[2] ,
         \SB2_2_2/Component_Function_4/NAND4_in[1] ,
         \SB2_2_2/Component_Function_4/NAND4_in[0] ,
         \SB2_2_3/Component_Function_2/NAND4_in[3] ,
         \SB2_2_3/Component_Function_2/NAND4_in[1] ,
         \SB2_2_3/Component_Function_2/NAND4_in[0] ,
         \SB2_2_3/Component_Function_3/NAND4_in[3] ,
         \SB2_2_3/Component_Function_3/NAND4_in[2] ,
         \SB2_2_3/Component_Function_3/NAND4_in[1] ,
         \SB2_2_3/Component_Function_3/NAND4_in[0] ,
         \SB2_2_3/Component_Function_4/NAND4_in[3] ,
         \SB2_2_3/Component_Function_4/NAND4_in[1] ,
         \SB2_2_3/Component_Function_4/NAND4_in[0] ,
         \SB2_2_4/Component_Function_2/NAND4_in[3] ,
         \SB2_2_4/Component_Function_2/NAND4_in[2] ,
         \SB2_2_4/Component_Function_2/NAND4_in[1] ,
         \SB2_2_4/Component_Function_2/NAND4_in[0] ,
         \SB2_2_4/Component_Function_3/NAND4_in[3] ,
         \SB2_2_4/Component_Function_3/NAND4_in[2] ,
         \SB2_2_4/Component_Function_3/NAND4_in[1] ,
         \SB2_2_4/Component_Function_3/NAND4_in[0] ,
         \SB2_2_4/Component_Function_4/NAND4_in[3] ,
         \SB2_2_4/Component_Function_4/NAND4_in[1] ,
         \SB2_2_4/Component_Function_4/NAND4_in[0] ,
         \SB2_2_5/Component_Function_2/NAND4_in[3] ,
         \SB2_2_5/Component_Function_2/NAND4_in[2] ,
         \SB2_2_5/Component_Function_2/NAND4_in[1] ,
         \SB2_2_5/Component_Function_2/NAND4_in[0] ,
         \SB2_2_5/Component_Function_3/NAND4_in[3] ,
         \SB2_2_5/Component_Function_3/NAND4_in[2] ,
         \SB2_2_5/Component_Function_3/NAND4_in[1] ,
         \SB2_2_5/Component_Function_3/NAND4_in[0] ,
         \SB2_2_5/Component_Function_4/NAND4_in[2] ,
         \SB2_2_5/Component_Function_4/NAND4_in[1] ,
         \SB2_2_5/Component_Function_4/NAND4_in[0] ,
         \SB2_2_6/Component_Function_2/NAND4_in[1] ,
         \SB2_2_6/Component_Function_2/NAND4_in[0] ,
         \SB2_2_6/Component_Function_3/NAND4_in[3] ,
         \SB2_2_6/Component_Function_3/NAND4_in[2] ,
         \SB2_2_6/Component_Function_3/NAND4_in[1] ,
         \SB2_2_6/Component_Function_3/NAND4_in[0] ,
         \SB2_2_6/Component_Function_4/NAND4_in[2] ,
         \SB2_2_6/Component_Function_4/NAND4_in[1] ,
         \SB2_2_6/Component_Function_4/NAND4_in[0] ,
         \SB2_2_7/Component_Function_2/NAND4_in[3] ,
         \SB2_2_7/Component_Function_2/NAND4_in[2] ,
         \SB2_2_7/Component_Function_2/NAND4_in[1] ,
         \SB2_2_7/Component_Function_2/NAND4_in[0] ,
         \SB2_2_7/Component_Function_3/NAND4_in[3] ,
         \SB2_2_7/Component_Function_3/NAND4_in[2] ,
         \SB2_2_7/Component_Function_3/NAND4_in[1] ,
         \SB2_2_7/Component_Function_3/NAND4_in[0] ,
         \SB2_2_7/Component_Function_4/NAND4_in[3] ,
         \SB2_2_7/Component_Function_4/NAND4_in[2] ,
         \SB2_2_7/Component_Function_4/NAND4_in[1] ,
         \SB2_2_7/Component_Function_4/NAND4_in[0] ,
         \SB2_2_8/Component_Function_2/NAND4_in[2] ,
         \SB2_2_8/Component_Function_2/NAND4_in[1] ,
         \SB2_2_8/Component_Function_2/NAND4_in[0] ,
         \SB2_2_8/Component_Function_3/NAND4_in[1] ,
         \SB2_2_8/Component_Function_3/NAND4_in[0] ,
         \SB2_2_8/Component_Function_4/NAND4_in[2] ,
         \SB2_2_8/Component_Function_4/NAND4_in[1] ,
         \SB2_2_8/Component_Function_4/NAND4_in[0] ,
         \SB2_2_9/Component_Function_2/NAND4_in[2] ,
         \SB2_2_9/Component_Function_2/NAND4_in[1] ,
         \SB2_2_9/Component_Function_2/NAND4_in[0] ,
         \SB2_2_9/Component_Function_3/NAND4_in[3] ,
         \SB2_2_9/Component_Function_3/NAND4_in[2] ,
         \SB2_2_9/Component_Function_3/NAND4_in[1] ,
         \SB2_2_9/Component_Function_3/NAND4_in[0] ,
         \SB2_2_9/Component_Function_4/NAND4_in[2] ,
         \SB2_2_9/Component_Function_4/NAND4_in[1] ,
         \SB2_2_9/Component_Function_4/NAND4_in[0] ,
         \SB2_2_10/Component_Function_2/NAND4_in[2] ,
         \SB2_2_10/Component_Function_2/NAND4_in[1] ,
         \SB2_2_10/Component_Function_2/NAND4_in[0] ,
         \SB2_2_10/Component_Function_3/NAND4_in[2] ,
         \SB2_2_10/Component_Function_3/NAND4_in[1] ,
         \SB2_2_10/Component_Function_3/NAND4_in[0] ,
         \SB2_2_10/Component_Function_4/NAND4_in[2] ,
         \SB2_2_10/Component_Function_4/NAND4_in[1] ,
         \SB2_2_10/Component_Function_4/NAND4_in[0] ,
         \SB2_2_11/Component_Function_2/NAND4_in[1] ,
         \SB2_2_11/Component_Function_2/NAND4_in[0] ,
         \SB2_2_11/Component_Function_3/NAND4_in[2] ,
         \SB2_2_11/Component_Function_3/NAND4_in[1] ,
         \SB2_2_11/Component_Function_3/NAND4_in[0] ,
         \SB2_2_11/Component_Function_4/NAND4_in[2] ,
         \SB2_2_11/Component_Function_4/NAND4_in[1] ,
         \SB2_2_11/Component_Function_4/NAND4_in[0] ,
         \SB2_2_12/Component_Function_2/NAND4_in[3] ,
         \SB2_2_12/Component_Function_2/NAND4_in[2] ,
         \SB2_2_12/Component_Function_2/NAND4_in[1] ,
         \SB2_2_12/Component_Function_2/NAND4_in[0] ,
         \SB2_2_12/Component_Function_3/NAND4_in[3] ,
         \SB2_2_12/Component_Function_3/NAND4_in[2] ,
         \SB2_2_12/Component_Function_3/NAND4_in[1] ,
         \SB2_2_12/Component_Function_3/NAND4_in[0] ,
         \SB2_2_12/Component_Function_4/NAND4_in[2] ,
         \SB2_2_12/Component_Function_4/NAND4_in[1] ,
         \SB2_2_12/Component_Function_4/NAND4_in[0] ,
         \SB2_2_13/Component_Function_2/NAND4_in[3] ,
         \SB2_2_13/Component_Function_2/NAND4_in[2] ,
         \SB2_2_13/Component_Function_2/NAND4_in[1] ,
         \SB2_2_13/Component_Function_2/NAND4_in[0] ,
         \SB2_2_13/Component_Function_3/NAND4_in[3] ,
         \SB2_2_13/Component_Function_3/NAND4_in[2] ,
         \SB2_2_13/Component_Function_3/NAND4_in[1] ,
         \SB2_2_13/Component_Function_3/NAND4_in[0] ,
         \SB2_2_13/Component_Function_4/NAND4_in[3] ,
         \SB2_2_13/Component_Function_4/NAND4_in[2] ,
         \SB2_2_13/Component_Function_4/NAND4_in[0] ,
         \SB2_2_14/Component_Function_2/NAND4_in[3] ,
         \SB2_2_14/Component_Function_2/NAND4_in[2] ,
         \SB2_2_14/Component_Function_2/NAND4_in[1] ,
         \SB2_2_14/Component_Function_2/NAND4_in[0] ,
         \SB2_2_14/Component_Function_3/NAND4_in[3] ,
         \SB2_2_14/Component_Function_3/NAND4_in[2] ,
         \SB2_2_14/Component_Function_3/NAND4_in[1] ,
         \SB2_2_14/Component_Function_3/NAND4_in[0] ,
         \SB2_2_14/Component_Function_4/NAND4_in[2] ,
         \SB2_2_14/Component_Function_4/NAND4_in[1] ,
         \SB2_2_14/Component_Function_4/NAND4_in[0] ,
         \SB2_2_15/Component_Function_2/NAND4_in[2] ,
         \SB2_2_15/Component_Function_2/NAND4_in[1] ,
         \SB2_2_15/Component_Function_2/NAND4_in[0] ,
         \SB2_2_15/Component_Function_3/NAND4_in[3] ,
         \SB2_2_15/Component_Function_3/NAND4_in[2] ,
         \SB2_2_15/Component_Function_3/NAND4_in[1] ,
         \SB2_2_15/Component_Function_3/NAND4_in[0] ,
         \SB2_2_15/Component_Function_4/NAND4_in[2] ,
         \SB2_2_15/Component_Function_4/NAND4_in[1] ,
         \SB2_2_15/Component_Function_4/NAND4_in[0] ,
         \SB2_2_16/Component_Function_2/NAND4_in[3] ,
         \SB2_2_16/Component_Function_2/NAND4_in[2] ,
         \SB2_2_16/Component_Function_2/NAND4_in[1] ,
         \SB2_2_16/Component_Function_2/NAND4_in[0] ,
         \SB2_2_16/Component_Function_3/NAND4_in[2] ,
         \SB2_2_16/Component_Function_3/NAND4_in[1] ,
         \SB2_2_16/Component_Function_3/NAND4_in[0] ,
         \SB2_2_16/Component_Function_4/NAND4_in[3] ,
         \SB2_2_16/Component_Function_4/NAND4_in[2] ,
         \SB2_2_16/Component_Function_4/NAND4_in[1] ,
         \SB2_2_16/Component_Function_4/NAND4_in[0] ,
         \SB2_2_17/Component_Function_2/NAND4_in[3] ,
         \SB2_2_17/Component_Function_2/NAND4_in[1] ,
         \SB2_2_17/Component_Function_2/NAND4_in[0] ,
         \SB2_2_17/Component_Function_3/NAND4_in[2] ,
         \SB2_2_17/Component_Function_3/NAND4_in[1] ,
         \SB2_2_17/Component_Function_3/NAND4_in[0] ,
         \SB2_2_17/Component_Function_4/NAND4_in[2] ,
         \SB2_2_17/Component_Function_4/NAND4_in[1] ,
         \SB2_2_17/Component_Function_4/NAND4_in[0] ,
         \SB2_2_18/Component_Function_2/NAND4_in[2] ,
         \SB2_2_18/Component_Function_2/NAND4_in[1] ,
         \SB2_2_18/Component_Function_2/NAND4_in[0] ,
         \SB2_2_18/Component_Function_3/NAND4_in[2] ,
         \SB2_2_18/Component_Function_3/NAND4_in[1] ,
         \SB2_2_18/Component_Function_3/NAND4_in[0] ,
         \SB2_2_18/Component_Function_4/NAND4_in[2] ,
         \SB2_2_18/Component_Function_4/NAND4_in[1] ,
         \SB2_2_18/Component_Function_4/NAND4_in[0] ,
         \SB2_2_19/Component_Function_2/NAND4_in[3] ,
         \SB2_2_19/Component_Function_2/NAND4_in[2] ,
         \SB2_2_19/Component_Function_2/NAND4_in[1] ,
         \SB2_2_19/Component_Function_2/NAND4_in[0] ,
         \SB2_2_19/Component_Function_3/NAND4_in[3] ,
         \SB2_2_19/Component_Function_3/NAND4_in[2] ,
         \SB2_2_19/Component_Function_3/NAND4_in[1] ,
         \SB2_2_19/Component_Function_3/NAND4_in[0] ,
         \SB2_2_19/Component_Function_4/NAND4_in[3] ,
         \SB2_2_19/Component_Function_4/NAND4_in[1] ,
         \SB2_2_19/Component_Function_4/NAND4_in[0] ,
         \SB2_2_20/Component_Function_2/NAND4_in[2] ,
         \SB2_2_20/Component_Function_2/NAND4_in[1] ,
         \SB2_2_20/Component_Function_2/NAND4_in[0] ,
         \SB2_2_20/Component_Function_3/NAND4_in[2] ,
         \SB2_2_20/Component_Function_3/NAND4_in[0] ,
         \SB2_2_20/Component_Function_4/NAND4_in[3] ,
         \SB2_2_20/Component_Function_4/NAND4_in[1] ,
         \SB2_2_20/Component_Function_4/NAND4_in[0] ,
         \SB2_2_21/Component_Function_2/NAND4_in[3] ,
         \SB2_2_21/Component_Function_2/NAND4_in[1] ,
         \SB2_2_21/Component_Function_2/NAND4_in[0] ,
         \SB2_2_21/Component_Function_3/NAND4_in[3] ,
         \SB2_2_21/Component_Function_3/NAND4_in[2] ,
         \SB2_2_21/Component_Function_3/NAND4_in[1] ,
         \SB2_2_21/Component_Function_3/NAND4_in[0] ,
         \SB2_2_21/Component_Function_4/NAND4_in[2] ,
         \SB2_2_21/Component_Function_4/NAND4_in[1] ,
         \SB2_2_21/Component_Function_4/NAND4_in[0] ,
         \SB2_2_22/Component_Function_2/NAND4_in[3] ,
         \SB2_2_22/Component_Function_2/NAND4_in[2] ,
         \SB2_2_22/Component_Function_2/NAND4_in[1] ,
         \SB2_2_22/Component_Function_2/NAND4_in[0] ,
         \SB2_2_22/Component_Function_3/NAND4_in[3] ,
         \SB2_2_22/Component_Function_3/NAND4_in[2] ,
         \SB2_2_22/Component_Function_3/NAND4_in[1] ,
         \SB2_2_22/Component_Function_3/NAND4_in[0] ,
         \SB2_2_22/Component_Function_4/NAND4_in[3] ,
         \SB2_2_22/Component_Function_4/NAND4_in[1] ,
         \SB2_2_22/Component_Function_4/NAND4_in[0] ,
         \SB2_2_23/Component_Function_2/NAND4_in[3] ,
         \SB2_2_23/Component_Function_2/NAND4_in[2] ,
         \SB2_2_23/Component_Function_2/NAND4_in[1] ,
         \SB2_2_23/Component_Function_2/NAND4_in[0] ,
         \SB2_2_23/Component_Function_3/NAND4_in[2] ,
         \SB2_2_23/Component_Function_3/NAND4_in[1] ,
         \SB2_2_23/Component_Function_4/NAND4_in[3] ,
         \SB2_2_23/Component_Function_4/NAND4_in[2] ,
         \SB2_2_23/Component_Function_4/NAND4_in[1] ,
         \SB2_2_23/Component_Function_4/NAND4_in[0] ,
         \SB2_2_24/Component_Function_2/NAND4_in[2] ,
         \SB2_2_24/Component_Function_2/NAND4_in[1] ,
         \SB2_2_24/Component_Function_2/NAND4_in[0] ,
         \SB2_2_24/Component_Function_3/NAND4_in[2] ,
         \SB2_2_24/Component_Function_3/NAND4_in[1] ,
         \SB2_2_24/Component_Function_3/NAND4_in[0] ,
         \SB2_2_24/Component_Function_4/NAND4_in[3] ,
         \SB2_2_24/Component_Function_4/NAND4_in[2] ,
         \SB2_2_24/Component_Function_4/NAND4_in[1] ,
         \SB2_2_24/Component_Function_4/NAND4_in[0] ,
         \SB2_2_25/Component_Function_2/NAND4_in[2] ,
         \SB2_2_25/Component_Function_2/NAND4_in[1] ,
         \SB2_2_25/Component_Function_2/NAND4_in[0] ,
         \SB2_2_25/Component_Function_3/NAND4_in[3] ,
         \SB2_2_25/Component_Function_3/NAND4_in[2] ,
         \SB2_2_25/Component_Function_3/NAND4_in[1] ,
         \SB2_2_25/Component_Function_3/NAND4_in[0] ,
         \SB2_2_25/Component_Function_4/NAND4_in[2] ,
         \SB2_2_25/Component_Function_4/NAND4_in[1] ,
         \SB2_2_25/Component_Function_4/NAND4_in[0] ,
         \SB2_2_26/Component_Function_2/NAND4_in[1] ,
         \SB2_2_26/Component_Function_2/NAND4_in[0] ,
         \SB2_2_26/Component_Function_3/NAND4_in[2] ,
         \SB2_2_26/Component_Function_3/NAND4_in[1] ,
         \SB2_2_26/Component_Function_3/NAND4_in[0] ,
         \SB2_2_26/Component_Function_4/NAND4_in[2] ,
         \SB2_2_26/Component_Function_4/NAND4_in[1] ,
         \SB2_2_26/Component_Function_4/NAND4_in[0] ,
         \SB2_2_27/Component_Function_2/NAND4_in[2] ,
         \SB2_2_27/Component_Function_2/NAND4_in[1] ,
         \SB2_2_27/Component_Function_2/NAND4_in[0] ,
         \SB2_2_27/Component_Function_3/NAND4_in[3] ,
         \SB2_2_27/Component_Function_3/NAND4_in[2] ,
         \SB2_2_27/Component_Function_3/NAND4_in[1] ,
         \SB2_2_27/Component_Function_3/NAND4_in[0] ,
         \SB2_2_27/Component_Function_4/NAND4_in[2] ,
         \SB2_2_27/Component_Function_4/NAND4_in[1] ,
         \SB2_2_27/Component_Function_4/NAND4_in[0] ,
         \SB2_2_28/Component_Function_2/NAND4_in[3] ,
         \SB2_2_28/Component_Function_2/NAND4_in[0] ,
         \SB2_2_28/Component_Function_3/NAND4_in[3] ,
         \SB2_2_28/Component_Function_3/NAND4_in[2] ,
         \SB2_2_28/Component_Function_3/NAND4_in[1] ,
         \SB2_2_28/Component_Function_3/NAND4_in[0] ,
         \SB2_2_28/Component_Function_4/NAND4_in[3] ,
         \SB2_2_28/Component_Function_4/NAND4_in[1] ,
         \SB2_2_28/Component_Function_4/NAND4_in[0] ,
         \SB2_2_29/Component_Function_2/NAND4_in[2] ,
         \SB2_2_29/Component_Function_2/NAND4_in[1] ,
         \SB2_2_29/Component_Function_2/NAND4_in[0] ,
         \SB2_2_29/Component_Function_3/NAND4_in[3] ,
         \SB2_2_29/Component_Function_3/NAND4_in[1] ,
         \SB2_2_29/Component_Function_3/NAND4_in[0] ,
         \SB2_2_29/Component_Function_4/NAND4_in[2] ,
         \SB2_2_29/Component_Function_4/NAND4_in[1] ,
         \SB2_2_29/Component_Function_4/NAND4_in[0] ,
         \SB2_2_30/Component_Function_2/NAND4_in[3] ,
         \SB2_2_30/Component_Function_2/NAND4_in[2] ,
         \SB2_2_30/Component_Function_2/NAND4_in[1] ,
         \SB2_2_30/Component_Function_2/NAND4_in[0] ,
         \SB2_2_30/Component_Function_3/NAND4_in[3] ,
         \SB2_2_30/Component_Function_3/NAND4_in[2] ,
         \SB2_2_30/Component_Function_3/NAND4_in[1] ,
         \SB2_2_30/Component_Function_3/NAND4_in[0] ,
         \SB2_2_30/Component_Function_4/NAND4_in[3] ,
         \SB2_2_30/Component_Function_4/NAND4_in[2] ,
         \SB2_2_30/Component_Function_4/NAND4_in[1] ,
         \SB2_2_30/Component_Function_4/NAND4_in[0] ,
         \SB2_2_31/Component_Function_2/NAND4_in[3] ,
         \SB2_2_31/Component_Function_2/NAND4_in[1] ,
         \SB2_2_31/Component_Function_2/NAND4_in[0] ,
         \SB2_2_31/Component_Function_3/NAND4_in[3] ,
         \SB2_2_31/Component_Function_3/NAND4_in[2] ,
         \SB2_2_31/Component_Function_3/NAND4_in[1] ,
         \SB2_2_31/Component_Function_3/NAND4_in[0] ,
         \SB2_2_31/Component_Function_4/NAND4_in[3] ,
         \SB2_2_31/Component_Function_4/NAND4_in[2] ,
         \SB2_2_31/Component_Function_4/NAND4_in[1] ,
         \SB2_2_31/Component_Function_4/NAND4_in[0] ,
         \SB1_3_0/Component_Function_2/NAND4_in[3] ,
         \SB1_3_0/Component_Function_2/NAND4_in[2] ,
         \SB1_3_0/Component_Function_2/NAND4_in[1] ,
         \SB1_3_0/Component_Function_2/NAND4_in[0] ,
         \SB1_3_0/Component_Function_3/NAND4_in[3] ,
         \SB1_3_0/Component_Function_3/NAND4_in[2] ,
         \SB1_3_0/Component_Function_3/NAND4_in[1] ,
         \SB1_3_0/Component_Function_3/NAND4_in[0] ,
         \SB1_3_0/Component_Function_4/NAND4_in[3] ,
         \SB1_3_0/Component_Function_4/NAND4_in[2] ,
         \SB1_3_0/Component_Function_4/NAND4_in[1] ,
         \SB1_3_0/Component_Function_4/NAND4_in[0] ,
         \SB1_3_1/Component_Function_2/NAND4_in[3] ,
         \SB1_3_1/Component_Function_2/NAND4_in[2] ,
         \SB1_3_1/Component_Function_2/NAND4_in[1] ,
         \SB1_3_1/Component_Function_2/NAND4_in[0] ,
         \SB1_3_1/Component_Function_3/NAND4_in[3] ,
         \SB1_3_1/Component_Function_3/NAND4_in[1] ,
         \SB1_3_1/Component_Function_3/NAND4_in[0] ,
         \SB1_3_1/Component_Function_4/NAND4_in[3] ,
         \SB1_3_1/Component_Function_4/NAND4_in[2] ,
         \SB1_3_1/Component_Function_4/NAND4_in[1] ,
         \SB1_3_1/Component_Function_4/NAND4_in[0] ,
         \SB1_3_2/Component_Function_2/NAND4_in[2] ,
         \SB1_3_2/Component_Function_2/NAND4_in[1] ,
         \SB1_3_2/Component_Function_2/NAND4_in[0] ,
         \SB1_3_2/Component_Function_3/NAND4_in[3] ,
         \SB1_3_2/Component_Function_3/NAND4_in[2] ,
         \SB1_3_2/Component_Function_3/NAND4_in[1] ,
         \SB1_3_2/Component_Function_3/NAND4_in[0] ,
         \SB1_3_2/Component_Function_4/NAND4_in[3] ,
         \SB1_3_2/Component_Function_4/NAND4_in[1] ,
         \SB1_3_2/Component_Function_4/NAND4_in[0] ,
         \SB1_3_3/Component_Function_2/NAND4_in[2] ,
         \SB1_3_3/Component_Function_2/NAND4_in[1] ,
         \SB1_3_3/Component_Function_2/NAND4_in[0] ,
         \SB1_3_3/Component_Function_3/NAND4_in[3] ,
         \SB1_3_3/Component_Function_3/NAND4_in[2] ,
         \SB1_3_3/Component_Function_3/NAND4_in[1] ,
         \SB1_3_3/Component_Function_3/NAND4_in[0] ,
         \SB1_3_3/Component_Function_4/NAND4_in[3] ,
         \SB1_3_3/Component_Function_4/NAND4_in[2] ,
         \SB1_3_3/Component_Function_4/NAND4_in[1] ,
         \SB1_3_3/Component_Function_4/NAND4_in[0] ,
         \SB1_3_4/Component_Function_2/NAND4_in[3] ,
         \SB1_3_4/Component_Function_2/NAND4_in[2] ,
         \SB1_3_4/Component_Function_2/NAND4_in[1] ,
         \SB1_3_4/Component_Function_2/NAND4_in[0] ,
         \SB1_3_4/Component_Function_3/NAND4_in[3] ,
         \SB1_3_4/Component_Function_3/NAND4_in[2] ,
         \SB1_3_4/Component_Function_3/NAND4_in[1] ,
         \SB1_3_4/Component_Function_3/NAND4_in[0] ,
         \SB1_3_4/Component_Function_4/NAND4_in[3] ,
         \SB1_3_4/Component_Function_4/NAND4_in[2] ,
         \SB1_3_4/Component_Function_4/NAND4_in[1] ,
         \SB1_3_4/Component_Function_4/NAND4_in[0] ,
         \SB1_3_5/Component_Function_2/NAND4_in[2] ,
         \SB1_3_5/Component_Function_2/NAND4_in[1] ,
         \SB1_3_5/Component_Function_2/NAND4_in[0] ,
         \SB1_3_5/Component_Function_3/NAND4_in[3] ,
         \SB1_3_5/Component_Function_3/NAND4_in[2] ,
         \SB1_3_5/Component_Function_3/NAND4_in[1] ,
         \SB1_3_5/Component_Function_3/NAND4_in[0] ,
         \SB1_3_5/Component_Function_4/NAND4_in[3] ,
         \SB1_3_5/Component_Function_4/NAND4_in[1] ,
         \SB1_3_5/Component_Function_4/NAND4_in[0] ,
         \SB1_3_6/Component_Function_2/NAND4_in[3] ,
         \SB1_3_6/Component_Function_2/NAND4_in[2] ,
         \SB1_3_6/Component_Function_2/NAND4_in[1] ,
         \SB1_3_6/Component_Function_2/NAND4_in[0] ,
         \SB1_3_6/Component_Function_3/NAND4_in[3] ,
         \SB1_3_6/Component_Function_3/NAND4_in[2] ,
         \SB1_3_6/Component_Function_3/NAND4_in[1] ,
         \SB1_3_6/Component_Function_3/NAND4_in[0] ,
         \SB1_3_6/Component_Function_4/NAND4_in[3] ,
         \SB1_3_6/Component_Function_4/NAND4_in[2] ,
         \SB1_3_6/Component_Function_4/NAND4_in[1] ,
         \SB1_3_6/Component_Function_4/NAND4_in[0] ,
         \SB1_3_7/Component_Function_2/NAND4_in[2] ,
         \SB1_3_7/Component_Function_2/NAND4_in[1] ,
         \SB1_3_7/Component_Function_2/NAND4_in[0] ,
         \SB1_3_7/Component_Function_3/NAND4_in[3] ,
         \SB1_3_7/Component_Function_3/NAND4_in[2] ,
         \SB1_3_7/Component_Function_3/NAND4_in[1] ,
         \SB1_3_7/Component_Function_3/NAND4_in[0] ,
         \SB1_3_7/Component_Function_4/NAND4_in[3] ,
         \SB1_3_7/Component_Function_4/NAND4_in[2] ,
         \SB1_3_7/Component_Function_4/NAND4_in[1] ,
         \SB1_3_7/Component_Function_4/NAND4_in[0] ,
         \SB1_3_8/Component_Function_2/NAND4_in[2] ,
         \SB1_3_8/Component_Function_2/NAND4_in[1] ,
         \SB1_3_8/Component_Function_2/NAND4_in[0] ,
         \SB1_3_8/Component_Function_3/NAND4_in[3] ,
         \SB1_3_8/Component_Function_3/NAND4_in[2] ,
         \SB1_3_8/Component_Function_3/NAND4_in[1] ,
         \SB1_3_8/Component_Function_3/NAND4_in[0] ,
         \SB1_3_8/Component_Function_4/NAND4_in[3] ,
         \SB1_3_8/Component_Function_4/NAND4_in[2] ,
         \SB1_3_8/Component_Function_4/NAND4_in[1] ,
         \SB1_3_8/Component_Function_4/NAND4_in[0] ,
         \SB1_3_9/Component_Function_2/NAND4_in[3] ,
         \SB1_3_9/Component_Function_2/NAND4_in[2] ,
         \SB1_3_9/Component_Function_2/NAND4_in[1] ,
         \SB1_3_9/Component_Function_2/NAND4_in[0] ,
         \SB1_3_9/Component_Function_3/NAND4_in[2] ,
         \SB1_3_9/Component_Function_3/NAND4_in[1] ,
         \SB1_3_9/Component_Function_3/NAND4_in[0] ,
         \SB1_3_9/Component_Function_4/NAND4_in[3] ,
         \SB1_3_9/Component_Function_4/NAND4_in[2] ,
         \SB1_3_9/Component_Function_4/NAND4_in[1] ,
         \SB1_3_9/Component_Function_4/NAND4_in[0] ,
         \SB1_3_10/Component_Function_2/NAND4_in[3] ,
         \SB1_3_10/Component_Function_2/NAND4_in[2] ,
         \SB1_3_10/Component_Function_2/NAND4_in[1] ,
         \SB1_3_10/Component_Function_2/NAND4_in[0] ,
         \SB1_3_10/Component_Function_3/NAND4_in[3] ,
         \SB1_3_10/Component_Function_3/NAND4_in[2] ,
         \SB1_3_10/Component_Function_3/NAND4_in[1] ,
         \SB1_3_10/Component_Function_3/NAND4_in[0] ,
         \SB1_3_10/Component_Function_4/NAND4_in[3] ,
         \SB1_3_10/Component_Function_4/NAND4_in[2] ,
         \SB1_3_10/Component_Function_4/NAND4_in[1] ,
         \SB1_3_10/Component_Function_4/NAND4_in[0] ,
         \SB1_3_11/Component_Function_2/NAND4_in[3] ,
         \SB1_3_11/Component_Function_2/NAND4_in[2] ,
         \SB1_3_11/Component_Function_2/NAND4_in[1] ,
         \SB1_3_11/Component_Function_2/NAND4_in[0] ,
         \SB1_3_11/Component_Function_3/NAND4_in[2] ,
         \SB1_3_11/Component_Function_3/NAND4_in[1] ,
         \SB1_3_11/Component_Function_3/NAND4_in[0] ,
         \SB1_3_11/Component_Function_4/NAND4_in[3] ,
         \SB1_3_11/Component_Function_4/NAND4_in[2] ,
         \SB1_3_11/Component_Function_4/NAND4_in[1] ,
         \SB1_3_11/Component_Function_4/NAND4_in[0] ,
         \SB1_3_12/Component_Function_2/NAND4_in[3] ,
         \SB1_3_12/Component_Function_2/NAND4_in[2] ,
         \SB1_3_12/Component_Function_2/NAND4_in[1] ,
         \SB1_3_12/Component_Function_2/NAND4_in[0] ,
         \SB1_3_12/Component_Function_3/NAND4_in[2] ,
         \SB1_3_12/Component_Function_3/NAND4_in[1] ,
         \SB1_3_12/Component_Function_3/NAND4_in[0] ,
         \SB1_3_12/Component_Function_4/NAND4_in[3] ,
         \SB1_3_12/Component_Function_4/NAND4_in[2] ,
         \SB1_3_12/Component_Function_4/NAND4_in[1] ,
         \SB1_3_12/Component_Function_4/NAND4_in[0] ,
         \SB1_3_13/Component_Function_2/NAND4_in[3] ,
         \SB1_3_13/Component_Function_2/NAND4_in[2] ,
         \SB1_3_13/Component_Function_2/NAND4_in[1] ,
         \SB1_3_13/Component_Function_2/NAND4_in[0] ,
         \SB1_3_13/Component_Function_3/NAND4_in[3] ,
         \SB1_3_13/Component_Function_3/NAND4_in[2] ,
         \SB1_3_13/Component_Function_3/NAND4_in[1] ,
         \SB1_3_13/Component_Function_3/NAND4_in[0] ,
         \SB1_3_13/Component_Function_4/NAND4_in[3] ,
         \SB1_3_13/Component_Function_4/NAND4_in[1] ,
         \SB1_3_13/Component_Function_4/NAND4_in[0] ,
         \SB1_3_14/Component_Function_2/NAND4_in[3] ,
         \SB1_3_14/Component_Function_2/NAND4_in[2] ,
         \SB1_3_14/Component_Function_2/NAND4_in[1] ,
         \SB1_3_14/Component_Function_2/NAND4_in[0] ,
         \SB1_3_14/Component_Function_3/NAND4_in[3] ,
         \SB1_3_14/Component_Function_3/NAND4_in[2] ,
         \SB1_3_14/Component_Function_3/NAND4_in[1] ,
         \SB1_3_14/Component_Function_3/NAND4_in[0] ,
         \SB1_3_14/Component_Function_4/NAND4_in[3] ,
         \SB1_3_14/Component_Function_4/NAND4_in[1] ,
         \SB1_3_14/Component_Function_4/NAND4_in[0] ,
         \SB1_3_15/Component_Function_2/NAND4_in[2] ,
         \SB1_3_15/Component_Function_2/NAND4_in[1] ,
         \SB1_3_15/Component_Function_2/NAND4_in[0] ,
         \SB1_3_15/Component_Function_3/NAND4_in[3] ,
         \SB1_3_15/Component_Function_3/NAND4_in[2] ,
         \SB1_3_15/Component_Function_3/NAND4_in[1] ,
         \SB1_3_15/Component_Function_3/NAND4_in[0] ,
         \SB1_3_15/Component_Function_4/NAND4_in[3] ,
         \SB1_3_15/Component_Function_4/NAND4_in[2] ,
         \SB1_3_15/Component_Function_4/NAND4_in[1] ,
         \SB1_3_15/Component_Function_4/NAND4_in[0] ,
         \SB1_3_16/Component_Function_2/NAND4_in[3] ,
         \SB1_3_16/Component_Function_2/NAND4_in[2] ,
         \SB1_3_16/Component_Function_2/NAND4_in[1] ,
         \SB1_3_16/Component_Function_2/NAND4_in[0] ,
         \SB1_3_16/Component_Function_3/NAND4_in[3] ,
         \SB1_3_16/Component_Function_3/NAND4_in[2] ,
         \SB1_3_16/Component_Function_3/NAND4_in[1] ,
         \SB1_3_16/Component_Function_3/NAND4_in[0] ,
         \SB1_3_16/Component_Function_4/NAND4_in[3] ,
         \SB1_3_16/Component_Function_4/NAND4_in[2] ,
         \SB1_3_16/Component_Function_4/NAND4_in[1] ,
         \SB1_3_16/Component_Function_4/NAND4_in[0] ,
         \SB1_3_17/Component_Function_2/NAND4_in[3] ,
         \SB1_3_17/Component_Function_2/NAND4_in[2] ,
         \SB1_3_17/Component_Function_2/NAND4_in[1] ,
         \SB1_3_17/Component_Function_2/NAND4_in[0] ,
         \SB1_3_17/Component_Function_3/NAND4_in[3] ,
         \SB1_3_17/Component_Function_3/NAND4_in[2] ,
         \SB1_3_17/Component_Function_3/NAND4_in[1] ,
         \SB1_3_17/Component_Function_3/NAND4_in[0] ,
         \SB1_3_17/Component_Function_4/NAND4_in[3] ,
         \SB1_3_17/Component_Function_4/NAND4_in[1] ,
         \SB1_3_17/Component_Function_4/NAND4_in[0] ,
         \SB1_3_18/Component_Function_2/NAND4_in[2] ,
         \SB1_3_18/Component_Function_2/NAND4_in[1] ,
         \SB1_3_18/Component_Function_2/NAND4_in[0] ,
         \SB1_3_18/Component_Function_3/NAND4_in[3] ,
         \SB1_3_18/Component_Function_3/NAND4_in[2] ,
         \SB1_3_18/Component_Function_3/NAND4_in[1] ,
         \SB1_3_18/Component_Function_3/NAND4_in[0] ,
         \SB1_3_18/Component_Function_4/NAND4_in[3] ,
         \SB1_3_18/Component_Function_4/NAND4_in[2] ,
         \SB1_3_18/Component_Function_4/NAND4_in[1] ,
         \SB1_3_18/Component_Function_4/NAND4_in[0] ,
         \SB1_3_19/Component_Function_2/NAND4_in[3] ,
         \SB1_3_19/Component_Function_2/NAND4_in[2] ,
         \SB1_3_19/Component_Function_2/NAND4_in[1] ,
         \SB1_3_19/Component_Function_2/NAND4_in[0] ,
         \SB1_3_19/Component_Function_3/NAND4_in[2] ,
         \SB1_3_19/Component_Function_3/NAND4_in[1] ,
         \SB1_3_19/Component_Function_3/NAND4_in[0] ,
         \SB1_3_19/Component_Function_4/NAND4_in[3] ,
         \SB1_3_19/Component_Function_4/NAND4_in[2] ,
         \SB1_3_19/Component_Function_4/NAND4_in[1] ,
         \SB1_3_19/Component_Function_4/NAND4_in[0] ,
         \SB1_3_20/Component_Function_2/NAND4_in[2] ,
         \SB1_3_20/Component_Function_2/NAND4_in[1] ,
         \SB1_3_20/Component_Function_2/NAND4_in[0] ,
         \SB1_3_20/Component_Function_3/NAND4_in[3] ,
         \SB1_3_20/Component_Function_3/NAND4_in[2] ,
         \SB1_3_20/Component_Function_3/NAND4_in[1] ,
         \SB1_3_20/Component_Function_3/NAND4_in[0] ,
         \SB1_3_20/Component_Function_4/NAND4_in[3] ,
         \SB1_3_20/Component_Function_4/NAND4_in[2] ,
         \SB1_3_20/Component_Function_4/NAND4_in[1] ,
         \SB1_3_20/Component_Function_4/NAND4_in[0] ,
         \SB1_3_21/Component_Function_2/NAND4_in[3] ,
         \SB1_3_21/Component_Function_2/NAND4_in[2] ,
         \SB1_3_21/Component_Function_2/NAND4_in[1] ,
         \SB1_3_21/Component_Function_2/NAND4_in[0] ,
         \SB1_3_21/Component_Function_3/NAND4_in[3] ,
         \SB1_3_21/Component_Function_3/NAND4_in[2] ,
         \SB1_3_21/Component_Function_3/NAND4_in[1] ,
         \SB1_3_21/Component_Function_3/NAND4_in[0] ,
         \SB1_3_21/Component_Function_4/NAND4_in[3] ,
         \SB1_3_21/Component_Function_4/NAND4_in[2] ,
         \SB1_3_21/Component_Function_4/NAND4_in[1] ,
         \SB1_3_21/Component_Function_4/NAND4_in[0] ,
         \SB1_3_22/Component_Function_2/NAND4_in[3] ,
         \SB1_3_22/Component_Function_2/NAND4_in[2] ,
         \SB1_3_22/Component_Function_2/NAND4_in[1] ,
         \SB1_3_22/Component_Function_2/NAND4_in[0] ,
         \SB1_3_22/Component_Function_3/NAND4_in[3] ,
         \SB1_3_22/Component_Function_3/NAND4_in[2] ,
         \SB1_3_22/Component_Function_3/NAND4_in[1] ,
         \SB1_3_22/Component_Function_3/NAND4_in[0] ,
         \SB1_3_22/Component_Function_4/NAND4_in[2] ,
         \SB1_3_22/Component_Function_4/NAND4_in[1] ,
         \SB1_3_22/Component_Function_4/NAND4_in[0] ,
         \SB1_3_23/Component_Function_2/NAND4_in[3] ,
         \SB1_3_23/Component_Function_2/NAND4_in[2] ,
         \SB1_3_23/Component_Function_2/NAND4_in[1] ,
         \SB1_3_23/Component_Function_2/NAND4_in[0] ,
         \SB1_3_23/Component_Function_3/NAND4_in[3] ,
         \SB1_3_23/Component_Function_3/NAND4_in[2] ,
         \SB1_3_23/Component_Function_3/NAND4_in[1] ,
         \SB1_3_23/Component_Function_3/NAND4_in[0] ,
         \SB1_3_23/Component_Function_4/NAND4_in[3] ,
         \SB1_3_23/Component_Function_4/NAND4_in[1] ,
         \SB1_3_23/Component_Function_4/NAND4_in[0] ,
         \SB1_3_24/Component_Function_2/NAND4_in[2] ,
         \SB1_3_24/Component_Function_2/NAND4_in[1] ,
         \SB1_3_24/Component_Function_2/NAND4_in[0] ,
         \SB1_3_24/Component_Function_3/NAND4_in[3] ,
         \SB1_3_24/Component_Function_3/NAND4_in[2] ,
         \SB1_3_24/Component_Function_3/NAND4_in[1] ,
         \SB1_3_24/Component_Function_3/NAND4_in[0] ,
         \SB1_3_24/Component_Function_4/NAND4_in[3] ,
         \SB1_3_24/Component_Function_4/NAND4_in[2] ,
         \SB1_3_24/Component_Function_4/NAND4_in[1] ,
         \SB1_3_24/Component_Function_4/NAND4_in[0] ,
         \SB1_3_25/Component_Function_2/NAND4_in[2] ,
         \SB1_3_25/Component_Function_2/NAND4_in[1] ,
         \SB1_3_25/Component_Function_2/NAND4_in[0] ,
         \SB1_3_25/Component_Function_3/NAND4_in[3] ,
         \SB1_3_25/Component_Function_3/NAND4_in[2] ,
         \SB1_3_25/Component_Function_3/NAND4_in[1] ,
         \SB1_3_25/Component_Function_3/NAND4_in[0] ,
         \SB1_3_25/Component_Function_4/NAND4_in[3] ,
         \SB1_3_25/Component_Function_4/NAND4_in[1] ,
         \SB1_3_25/Component_Function_4/NAND4_in[0] ,
         \SB1_3_26/Component_Function_2/NAND4_in[2] ,
         \SB1_3_26/Component_Function_2/NAND4_in[1] ,
         \SB1_3_26/Component_Function_2/NAND4_in[0] ,
         \SB1_3_26/Component_Function_3/NAND4_in[3] ,
         \SB1_3_26/Component_Function_3/NAND4_in[2] ,
         \SB1_3_26/Component_Function_3/NAND4_in[1] ,
         \SB1_3_26/Component_Function_3/NAND4_in[0] ,
         \SB1_3_26/Component_Function_4/NAND4_in[2] ,
         \SB1_3_26/Component_Function_4/NAND4_in[1] ,
         \SB1_3_26/Component_Function_4/NAND4_in[0] ,
         \SB1_3_27/Component_Function_2/NAND4_in[2] ,
         \SB1_3_27/Component_Function_2/NAND4_in[1] ,
         \SB1_3_27/Component_Function_2/NAND4_in[0] ,
         \SB1_3_27/Component_Function_3/NAND4_in[3] ,
         \SB1_3_27/Component_Function_3/NAND4_in[2] ,
         \SB1_3_27/Component_Function_3/NAND4_in[1] ,
         \SB1_3_27/Component_Function_3/NAND4_in[0] ,
         \SB1_3_27/Component_Function_4/NAND4_in[3] ,
         \SB1_3_27/Component_Function_4/NAND4_in[2] ,
         \SB1_3_27/Component_Function_4/NAND4_in[1] ,
         \SB1_3_27/Component_Function_4/NAND4_in[0] ,
         \SB1_3_28/Component_Function_2/NAND4_in[3] ,
         \SB1_3_28/Component_Function_2/NAND4_in[2] ,
         \SB1_3_28/Component_Function_2/NAND4_in[1] ,
         \SB1_3_28/Component_Function_2/NAND4_in[0] ,
         \SB1_3_28/Component_Function_3/NAND4_in[3] ,
         \SB1_3_28/Component_Function_3/NAND4_in[2] ,
         \SB1_3_28/Component_Function_3/NAND4_in[1] ,
         \SB1_3_28/Component_Function_3/NAND4_in[0] ,
         \SB1_3_28/Component_Function_4/NAND4_in[3] ,
         \SB1_3_28/Component_Function_4/NAND4_in[2] ,
         \SB1_3_28/Component_Function_4/NAND4_in[1] ,
         \SB1_3_28/Component_Function_4/NAND4_in[0] ,
         \SB1_3_29/Component_Function_2/NAND4_in[3] ,
         \SB1_3_29/Component_Function_2/NAND4_in[2] ,
         \SB1_3_29/Component_Function_2/NAND4_in[1] ,
         \SB1_3_29/Component_Function_2/NAND4_in[0] ,
         \SB1_3_29/Component_Function_3/NAND4_in[3] ,
         \SB1_3_29/Component_Function_3/NAND4_in[2] ,
         \SB1_3_29/Component_Function_3/NAND4_in[1] ,
         \SB1_3_29/Component_Function_3/NAND4_in[0] ,
         \SB1_3_29/Component_Function_4/NAND4_in[3] ,
         \SB1_3_29/Component_Function_4/NAND4_in[2] ,
         \SB1_3_29/Component_Function_4/NAND4_in[1] ,
         \SB1_3_29/Component_Function_4/NAND4_in[0] ,
         \SB1_3_30/Component_Function_2/NAND4_in[2] ,
         \SB1_3_30/Component_Function_2/NAND4_in[1] ,
         \SB1_3_30/Component_Function_2/NAND4_in[0] ,
         \SB1_3_30/Component_Function_3/NAND4_in[2] ,
         \SB1_3_30/Component_Function_3/NAND4_in[1] ,
         \SB1_3_30/Component_Function_3/NAND4_in[0] ,
         \SB1_3_30/Component_Function_4/NAND4_in[3] ,
         \SB1_3_30/Component_Function_4/NAND4_in[2] ,
         \SB1_3_30/Component_Function_4/NAND4_in[1] ,
         \SB1_3_30/Component_Function_4/NAND4_in[0] ,
         \SB1_3_31/Component_Function_2/NAND4_in[2] ,
         \SB1_3_31/Component_Function_2/NAND4_in[1] ,
         \SB1_3_31/Component_Function_2/NAND4_in[0] ,
         \SB1_3_31/Component_Function_3/NAND4_in[3] ,
         \SB1_3_31/Component_Function_3/NAND4_in[2] ,
         \SB1_3_31/Component_Function_3/NAND4_in[1] ,
         \SB1_3_31/Component_Function_3/NAND4_in[0] ,
         \SB1_3_31/Component_Function_4/NAND4_in[3] ,
         \SB1_3_31/Component_Function_4/NAND4_in[1] ,
         \SB1_3_31/Component_Function_4/NAND4_in[0] ,
         \SB2_3_0/Component_Function_2/NAND4_in[2] ,
         \SB2_3_0/Component_Function_2/NAND4_in[1] ,
         \SB2_3_0/Component_Function_2/NAND4_in[0] ,
         \SB2_3_0/Component_Function_3/NAND4_in[3] ,
         \SB2_3_0/Component_Function_3/NAND4_in[2] ,
         \SB2_3_0/Component_Function_3/NAND4_in[1] ,
         \SB2_3_0/Component_Function_3/NAND4_in[0] ,
         \SB2_3_0/Component_Function_4/NAND4_in[3] ,
         \SB2_3_0/Component_Function_4/NAND4_in[2] ,
         \SB2_3_0/Component_Function_4/NAND4_in[1] ,
         \SB2_3_0/Component_Function_4/NAND4_in[0] ,
         \SB2_3_1/Component_Function_2/NAND4_in[3] ,
         \SB2_3_1/Component_Function_2/NAND4_in[2] ,
         \SB2_3_1/Component_Function_2/NAND4_in[1] ,
         \SB2_3_1/Component_Function_2/NAND4_in[0] ,
         \SB2_3_1/Component_Function_3/NAND4_in[3] ,
         \SB2_3_1/Component_Function_3/NAND4_in[2] ,
         \SB2_3_1/Component_Function_3/NAND4_in[1] ,
         \SB2_3_1/Component_Function_3/NAND4_in[0] ,
         \SB2_3_1/Component_Function_4/NAND4_in[3] ,
         \SB2_3_1/Component_Function_4/NAND4_in[2] ,
         \SB2_3_1/Component_Function_4/NAND4_in[1] ,
         \SB2_3_1/Component_Function_4/NAND4_in[0] ,
         \SB2_3_2/Component_Function_2/NAND4_in[2] ,
         \SB2_3_2/Component_Function_2/NAND4_in[1] ,
         \SB2_3_2/Component_Function_2/NAND4_in[0] ,
         \SB2_3_2/Component_Function_3/NAND4_in[3] ,
         \SB2_3_2/Component_Function_3/NAND4_in[2] ,
         \SB2_3_2/Component_Function_3/NAND4_in[1] ,
         \SB2_3_2/Component_Function_3/NAND4_in[0] ,
         \SB2_3_2/Component_Function_4/NAND4_in[3] ,
         \SB2_3_2/Component_Function_4/NAND4_in[2] ,
         \SB2_3_2/Component_Function_4/NAND4_in[1] ,
         \SB2_3_2/Component_Function_4/NAND4_in[0] ,
         \SB2_3_3/Component_Function_2/NAND4_in[3] ,
         \SB2_3_3/Component_Function_2/NAND4_in[2] ,
         \SB2_3_3/Component_Function_2/NAND4_in[1] ,
         \SB2_3_3/Component_Function_2/NAND4_in[0] ,
         \SB2_3_3/Component_Function_3/NAND4_in[3] ,
         \SB2_3_3/Component_Function_3/NAND4_in[2] ,
         \SB2_3_3/Component_Function_3/NAND4_in[1] ,
         \SB2_3_3/Component_Function_3/NAND4_in[0] ,
         \SB2_3_3/Component_Function_4/NAND4_in[3] ,
         \SB2_3_3/Component_Function_4/NAND4_in[2] ,
         \SB2_3_3/Component_Function_4/NAND4_in[1] ,
         \SB2_3_3/Component_Function_4/NAND4_in[0] ,
         \SB2_3_4/Component_Function_2/NAND4_in[3] ,
         \SB2_3_4/Component_Function_2/NAND4_in[2] ,
         \SB2_3_4/Component_Function_2/NAND4_in[1] ,
         \SB2_3_4/Component_Function_2/NAND4_in[0] ,
         \SB2_3_4/Component_Function_3/NAND4_in[3] ,
         \SB2_3_4/Component_Function_3/NAND4_in[2] ,
         \SB2_3_4/Component_Function_3/NAND4_in[1] ,
         \SB2_3_4/Component_Function_3/NAND4_in[0] ,
         \SB2_3_4/Component_Function_4/NAND4_in[3] ,
         \SB2_3_4/Component_Function_4/NAND4_in[2] ,
         \SB2_3_4/Component_Function_4/NAND4_in[1] ,
         \SB2_3_4/Component_Function_4/NAND4_in[0] ,
         \SB2_3_5/Component_Function_2/NAND4_in[3] ,
         \SB2_3_5/Component_Function_2/NAND4_in[2] ,
         \SB2_3_5/Component_Function_2/NAND4_in[1] ,
         \SB2_3_5/Component_Function_2/NAND4_in[0] ,
         \SB2_3_5/Component_Function_3/NAND4_in[3] ,
         \SB2_3_5/Component_Function_3/NAND4_in[2] ,
         \SB2_3_5/Component_Function_3/NAND4_in[1] ,
         \SB2_3_5/Component_Function_3/NAND4_in[0] ,
         \SB2_3_5/Component_Function_4/NAND4_in[3] ,
         \SB2_3_5/Component_Function_4/NAND4_in[2] ,
         \SB2_3_5/Component_Function_4/NAND4_in[1] ,
         \SB2_3_5/Component_Function_4/NAND4_in[0] ,
         \SB2_3_6/Component_Function_2/NAND4_in[2] ,
         \SB2_3_6/Component_Function_2/NAND4_in[1] ,
         \SB2_3_6/Component_Function_2/NAND4_in[0] ,
         \SB2_3_6/Component_Function_3/NAND4_in[3] ,
         \SB2_3_6/Component_Function_3/NAND4_in[2] ,
         \SB2_3_6/Component_Function_3/NAND4_in[1] ,
         \SB2_3_6/Component_Function_3/NAND4_in[0] ,
         \SB2_3_6/Component_Function_4/NAND4_in[3] ,
         \SB2_3_6/Component_Function_4/NAND4_in[2] ,
         \SB2_3_6/Component_Function_4/NAND4_in[1] ,
         \SB2_3_6/Component_Function_4/NAND4_in[0] ,
         \SB2_3_7/Component_Function_2/NAND4_in[3] ,
         \SB2_3_7/Component_Function_2/NAND4_in[2] ,
         \SB2_3_7/Component_Function_2/NAND4_in[1] ,
         \SB2_3_7/Component_Function_2/NAND4_in[0] ,
         \SB2_3_7/Component_Function_3/NAND4_in[3] ,
         \SB2_3_7/Component_Function_3/NAND4_in[2] ,
         \SB2_3_7/Component_Function_3/NAND4_in[1] ,
         \SB2_3_7/Component_Function_3/NAND4_in[0] ,
         \SB2_3_7/Component_Function_4/NAND4_in[3] ,
         \SB2_3_7/Component_Function_4/NAND4_in[2] ,
         \SB2_3_7/Component_Function_4/NAND4_in[1] ,
         \SB2_3_7/Component_Function_4/NAND4_in[0] ,
         \SB2_3_8/Component_Function_2/NAND4_in[3] ,
         \SB2_3_8/Component_Function_2/NAND4_in[2] ,
         \SB2_3_8/Component_Function_2/NAND4_in[1] ,
         \SB2_3_8/Component_Function_2/NAND4_in[0] ,
         \SB2_3_8/Component_Function_3/NAND4_in[3] ,
         \SB2_3_8/Component_Function_3/NAND4_in[2] ,
         \SB2_3_8/Component_Function_3/NAND4_in[1] ,
         \SB2_3_8/Component_Function_3/NAND4_in[0] ,
         \SB2_3_8/Component_Function_4/NAND4_in[3] ,
         \SB2_3_8/Component_Function_4/NAND4_in[2] ,
         \SB2_3_8/Component_Function_4/NAND4_in[1] ,
         \SB2_3_8/Component_Function_4/NAND4_in[0] ,
         \SB2_3_9/Component_Function_2/NAND4_in[3] ,
         \SB2_3_9/Component_Function_2/NAND4_in[2] ,
         \SB2_3_9/Component_Function_2/NAND4_in[1] ,
         \SB2_3_9/Component_Function_2/NAND4_in[0] ,
         \SB2_3_9/Component_Function_3/NAND4_in[3] ,
         \SB2_3_9/Component_Function_3/NAND4_in[2] ,
         \SB2_3_9/Component_Function_3/NAND4_in[1] ,
         \SB2_3_9/Component_Function_3/NAND4_in[0] ,
         \SB2_3_9/Component_Function_4/NAND4_in[3] ,
         \SB2_3_9/Component_Function_4/NAND4_in[2] ,
         \SB2_3_9/Component_Function_4/NAND4_in[1] ,
         \SB2_3_9/Component_Function_4/NAND4_in[0] ,
         \SB2_3_10/Component_Function_2/NAND4_in[3] ,
         \SB2_3_10/Component_Function_2/NAND4_in[2] ,
         \SB2_3_10/Component_Function_2/NAND4_in[1] ,
         \SB2_3_10/Component_Function_2/NAND4_in[0] ,
         \SB2_3_10/Component_Function_3/NAND4_in[3] ,
         \SB2_3_10/Component_Function_3/NAND4_in[2] ,
         \SB2_3_10/Component_Function_3/NAND4_in[1] ,
         \SB2_3_10/Component_Function_3/NAND4_in[0] ,
         \SB2_3_10/Component_Function_4/NAND4_in[2] ,
         \SB2_3_10/Component_Function_4/NAND4_in[1] ,
         \SB2_3_10/Component_Function_4/NAND4_in[0] ,
         \SB2_3_11/Component_Function_2/NAND4_in[3] ,
         \SB2_3_11/Component_Function_2/NAND4_in[2] ,
         \SB2_3_11/Component_Function_2/NAND4_in[1] ,
         \SB2_3_11/Component_Function_2/NAND4_in[0] ,
         \SB2_3_11/Component_Function_3/NAND4_in[3] ,
         \SB2_3_11/Component_Function_3/NAND4_in[2] ,
         \SB2_3_11/Component_Function_3/NAND4_in[1] ,
         \SB2_3_11/Component_Function_3/NAND4_in[0] ,
         \SB2_3_11/Component_Function_4/NAND4_in[3] ,
         \SB2_3_11/Component_Function_4/NAND4_in[2] ,
         \SB2_3_11/Component_Function_4/NAND4_in[1] ,
         \SB2_3_11/Component_Function_4/NAND4_in[0] ,
         \SB2_3_12/Component_Function_2/NAND4_in[3] ,
         \SB2_3_12/Component_Function_2/NAND4_in[2] ,
         \SB2_3_12/Component_Function_2/NAND4_in[1] ,
         \SB2_3_12/Component_Function_2/NAND4_in[0] ,
         \SB2_3_12/Component_Function_3/NAND4_in[3] ,
         \SB2_3_12/Component_Function_3/NAND4_in[2] ,
         \SB2_3_12/Component_Function_3/NAND4_in[1] ,
         \SB2_3_12/Component_Function_3/NAND4_in[0] ,
         \SB2_3_12/Component_Function_4/NAND4_in[3] ,
         \SB2_3_12/Component_Function_4/NAND4_in[2] ,
         \SB2_3_12/Component_Function_4/NAND4_in[1] ,
         \SB2_3_12/Component_Function_4/NAND4_in[0] ,
         \SB2_3_13/Component_Function_2/NAND4_in[2] ,
         \SB2_3_13/Component_Function_2/NAND4_in[1] ,
         \SB2_3_13/Component_Function_2/NAND4_in[0] ,
         \SB2_3_13/Component_Function_3/NAND4_in[3] ,
         \SB2_3_13/Component_Function_3/NAND4_in[2] ,
         \SB2_3_13/Component_Function_3/NAND4_in[1] ,
         \SB2_3_13/Component_Function_3/NAND4_in[0] ,
         \SB2_3_13/Component_Function_4/NAND4_in[3] ,
         \SB2_3_13/Component_Function_4/NAND4_in[2] ,
         \SB2_3_13/Component_Function_4/NAND4_in[1] ,
         \SB2_3_13/Component_Function_4/NAND4_in[0] ,
         \SB2_3_14/Component_Function_2/NAND4_in[3] ,
         \SB2_3_14/Component_Function_2/NAND4_in[2] ,
         \SB2_3_14/Component_Function_2/NAND4_in[1] ,
         \SB2_3_14/Component_Function_2/NAND4_in[0] ,
         \SB2_3_14/Component_Function_3/NAND4_in[3] ,
         \SB2_3_14/Component_Function_3/NAND4_in[2] ,
         \SB2_3_14/Component_Function_3/NAND4_in[1] ,
         \SB2_3_14/Component_Function_3/NAND4_in[0] ,
         \SB2_3_14/Component_Function_4/NAND4_in[3] ,
         \SB2_3_14/Component_Function_4/NAND4_in[2] ,
         \SB2_3_14/Component_Function_4/NAND4_in[1] ,
         \SB2_3_14/Component_Function_4/NAND4_in[0] ,
         \SB2_3_15/Component_Function_2/NAND4_in[2] ,
         \SB2_3_15/Component_Function_2/NAND4_in[1] ,
         \SB2_3_15/Component_Function_2/NAND4_in[0] ,
         \SB2_3_15/Component_Function_3/NAND4_in[3] ,
         \SB2_3_15/Component_Function_3/NAND4_in[2] ,
         \SB2_3_15/Component_Function_3/NAND4_in[1] ,
         \SB2_3_15/Component_Function_3/NAND4_in[0] ,
         \SB2_3_15/Component_Function_4/NAND4_in[3] ,
         \SB2_3_15/Component_Function_4/NAND4_in[1] ,
         \SB2_3_15/Component_Function_4/NAND4_in[0] ,
         \SB2_3_16/Component_Function_2/NAND4_in[3] ,
         \SB2_3_16/Component_Function_2/NAND4_in[1] ,
         \SB2_3_16/Component_Function_2/NAND4_in[0] ,
         \SB2_3_16/Component_Function_3/NAND4_in[3] ,
         \SB2_3_16/Component_Function_3/NAND4_in[2] ,
         \SB2_3_16/Component_Function_3/NAND4_in[1] ,
         \SB2_3_16/Component_Function_3/NAND4_in[0] ,
         \SB2_3_16/Component_Function_4/NAND4_in[3] ,
         \SB2_3_16/Component_Function_4/NAND4_in[2] ,
         \SB2_3_16/Component_Function_4/NAND4_in[1] ,
         \SB2_3_16/Component_Function_4/NAND4_in[0] ,
         \SB2_3_17/Component_Function_2/NAND4_in[3] ,
         \SB2_3_17/Component_Function_2/NAND4_in[2] ,
         \SB2_3_17/Component_Function_2/NAND4_in[1] ,
         \SB2_3_17/Component_Function_2/NAND4_in[0] ,
         \SB2_3_17/Component_Function_3/NAND4_in[3] ,
         \SB2_3_17/Component_Function_3/NAND4_in[2] ,
         \SB2_3_17/Component_Function_3/NAND4_in[1] ,
         \SB2_3_17/Component_Function_3/NAND4_in[0] ,
         \SB2_3_17/Component_Function_4/NAND4_in[3] ,
         \SB2_3_17/Component_Function_4/NAND4_in[2] ,
         \SB2_3_17/Component_Function_4/NAND4_in[1] ,
         \SB2_3_17/Component_Function_4/NAND4_in[0] ,
         \SB2_3_18/Component_Function_2/NAND4_in[2] ,
         \SB2_3_18/Component_Function_2/NAND4_in[1] ,
         \SB2_3_18/Component_Function_2/NAND4_in[0] ,
         \SB2_3_18/Component_Function_3/NAND4_in[3] ,
         \SB2_3_18/Component_Function_3/NAND4_in[2] ,
         \SB2_3_18/Component_Function_3/NAND4_in[1] ,
         \SB2_3_18/Component_Function_3/NAND4_in[0] ,
         \SB2_3_18/Component_Function_4/NAND4_in[3] ,
         \SB2_3_18/Component_Function_4/NAND4_in[2] ,
         \SB2_3_18/Component_Function_4/NAND4_in[1] ,
         \SB2_3_18/Component_Function_4/NAND4_in[0] ,
         \SB2_3_19/Component_Function_2/NAND4_in[3] ,
         \SB2_3_19/Component_Function_2/NAND4_in[2] ,
         \SB2_3_19/Component_Function_2/NAND4_in[1] ,
         \SB2_3_19/Component_Function_2/NAND4_in[0] ,
         \SB2_3_19/Component_Function_3/NAND4_in[3] ,
         \SB2_3_19/Component_Function_3/NAND4_in[2] ,
         \SB2_3_19/Component_Function_3/NAND4_in[1] ,
         \SB2_3_19/Component_Function_3/NAND4_in[0] ,
         \SB2_3_19/Component_Function_4/NAND4_in[3] ,
         \SB2_3_19/Component_Function_4/NAND4_in[2] ,
         \SB2_3_19/Component_Function_4/NAND4_in[1] ,
         \SB2_3_19/Component_Function_4/NAND4_in[0] ,
         \SB2_3_20/Component_Function_2/NAND4_in[3] ,
         \SB2_3_20/Component_Function_2/NAND4_in[2] ,
         \SB2_3_20/Component_Function_2/NAND4_in[1] ,
         \SB2_3_20/Component_Function_2/NAND4_in[0] ,
         \SB2_3_20/Component_Function_3/NAND4_in[3] ,
         \SB2_3_20/Component_Function_3/NAND4_in[2] ,
         \SB2_3_20/Component_Function_3/NAND4_in[1] ,
         \SB2_3_20/Component_Function_3/NAND4_in[0] ,
         \SB2_3_20/Component_Function_4/NAND4_in[3] ,
         \SB2_3_20/Component_Function_4/NAND4_in[2] ,
         \SB2_3_20/Component_Function_4/NAND4_in[1] ,
         \SB2_3_20/Component_Function_4/NAND4_in[0] ,
         \SB2_3_21/Component_Function_2/NAND4_in[3] ,
         \SB2_3_21/Component_Function_2/NAND4_in[2] ,
         \SB2_3_21/Component_Function_2/NAND4_in[1] ,
         \SB2_3_21/Component_Function_2/NAND4_in[0] ,
         \SB2_3_21/Component_Function_3/NAND4_in[2] ,
         \SB2_3_21/Component_Function_3/NAND4_in[1] ,
         \SB2_3_21/Component_Function_3/NAND4_in[0] ,
         \SB2_3_21/Component_Function_4/NAND4_in[2] ,
         \SB2_3_21/Component_Function_4/NAND4_in[1] ,
         \SB2_3_21/Component_Function_4/NAND4_in[0] ,
         \SB2_3_22/Component_Function_2/NAND4_in[3] ,
         \SB2_3_22/Component_Function_2/NAND4_in[2] ,
         \SB2_3_22/Component_Function_2/NAND4_in[1] ,
         \SB2_3_22/Component_Function_2/NAND4_in[0] ,
         \SB2_3_22/Component_Function_3/NAND4_in[3] ,
         \SB2_3_22/Component_Function_3/NAND4_in[2] ,
         \SB2_3_22/Component_Function_3/NAND4_in[1] ,
         \SB2_3_22/Component_Function_3/NAND4_in[0] ,
         \SB2_3_22/Component_Function_4/NAND4_in[3] ,
         \SB2_3_22/Component_Function_4/NAND4_in[2] ,
         \SB2_3_22/Component_Function_4/NAND4_in[1] ,
         \SB2_3_22/Component_Function_4/NAND4_in[0] ,
         \SB2_3_23/Component_Function_2/NAND4_in[3] ,
         \SB2_3_23/Component_Function_2/NAND4_in[2] ,
         \SB2_3_23/Component_Function_2/NAND4_in[1] ,
         \SB2_3_23/Component_Function_2/NAND4_in[0] ,
         \SB2_3_23/Component_Function_3/NAND4_in[3] ,
         \SB2_3_23/Component_Function_3/NAND4_in[2] ,
         \SB2_3_23/Component_Function_3/NAND4_in[1] ,
         \SB2_3_23/Component_Function_3/NAND4_in[0] ,
         \SB2_3_23/Component_Function_4/NAND4_in[3] ,
         \SB2_3_23/Component_Function_4/NAND4_in[2] ,
         \SB2_3_23/Component_Function_4/NAND4_in[1] ,
         \SB2_3_23/Component_Function_4/NAND4_in[0] ,
         \SB2_3_24/Component_Function_2/NAND4_in[3] ,
         \SB2_3_24/Component_Function_2/NAND4_in[2] ,
         \SB2_3_24/Component_Function_2/NAND4_in[1] ,
         \SB2_3_24/Component_Function_2/NAND4_in[0] ,
         \SB2_3_24/Component_Function_3/NAND4_in[3] ,
         \SB2_3_24/Component_Function_3/NAND4_in[2] ,
         \SB2_3_24/Component_Function_3/NAND4_in[1] ,
         \SB2_3_24/Component_Function_3/NAND4_in[0] ,
         \SB2_3_24/Component_Function_4/NAND4_in[3] ,
         \SB2_3_24/Component_Function_4/NAND4_in[2] ,
         \SB2_3_24/Component_Function_4/NAND4_in[1] ,
         \SB2_3_24/Component_Function_4/NAND4_in[0] ,
         \SB2_3_25/Component_Function_2/NAND4_in[3] ,
         \SB2_3_25/Component_Function_2/NAND4_in[2] ,
         \SB2_3_25/Component_Function_2/NAND4_in[1] ,
         \SB2_3_25/Component_Function_2/NAND4_in[0] ,
         \SB2_3_25/Component_Function_3/NAND4_in[3] ,
         \SB2_3_25/Component_Function_3/NAND4_in[2] ,
         \SB2_3_25/Component_Function_3/NAND4_in[1] ,
         \SB2_3_25/Component_Function_3/NAND4_in[0] ,
         \SB2_3_25/Component_Function_4/NAND4_in[3] ,
         \SB2_3_25/Component_Function_4/NAND4_in[2] ,
         \SB2_3_25/Component_Function_4/NAND4_in[1] ,
         \SB2_3_25/Component_Function_4/NAND4_in[0] ,
         \SB2_3_26/Component_Function_2/NAND4_in[3] ,
         \SB2_3_26/Component_Function_2/NAND4_in[2] ,
         \SB2_3_26/Component_Function_2/NAND4_in[1] ,
         \SB2_3_26/Component_Function_2/NAND4_in[0] ,
         \SB2_3_26/Component_Function_3/NAND4_in[3] ,
         \SB2_3_26/Component_Function_3/NAND4_in[2] ,
         \SB2_3_26/Component_Function_3/NAND4_in[1] ,
         \SB2_3_26/Component_Function_3/NAND4_in[0] ,
         \SB2_3_26/Component_Function_4/NAND4_in[3] ,
         \SB2_3_26/Component_Function_4/NAND4_in[2] ,
         \SB2_3_26/Component_Function_4/NAND4_in[1] ,
         \SB2_3_26/Component_Function_4/NAND4_in[0] ,
         \SB2_3_27/Component_Function_2/NAND4_in[3] ,
         \SB2_3_27/Component_Function_2/NAND4_in[2] ,
         \SB2_3_27/Component_Function_2/NAND4_in[1] ,
         \SB2_3_27/Component_Function_2/NAND4_in[0] ,
         \SB2_3_27/Component_Function_3/NAND4_in[3] ,
         \SB2_3_27/Component_Function_3/NAND4_in[2] ,
         \SB2_3_27/Component_Function_3/NAND4_in[1] ,
         \SB2_3_27/Component_Function_3/NAND4_in[0] ,
         \SB2_3_27/Component_Function_4/NAND4_in[3] ,
         \SB2_3_27/Component_Function_4/NAND4_in[2] ,
         \SB2_3_27/Component_Function_4/NAND4_in[1] ,
         \SB2_3_27/Component_Function_4/NAND4_in[0] ,
         \SB2_3_28/Component_Function_2/NAND4_in[3] ,
         \SB2_3_28/Component_Function_2/NAND4_in[2] ,
         \SB2_3_28/Component_Function_2/NAND4_in[1] ,
         \SB2_3_28/Component_Function_2/NAND4_in[0] ,
         \SB2_3_28/Component_Function_3/NAND4_in[3] ,
         \SB2_3_28/Component_Function_3/NAND4_in[2] ,
         \SB2_3_28/Component_Function_3/NAND4_in[1] ,
         \SB2_3_28/Component_Function_3/NAND4_in[0] ,
         \SB2_3_28/Component_Function_4/NAND4_in[3] ,
         \SB2_3_28/Component_Function_4/NAND4_in[2] ,
         \SB2_3_28/Component_Function_4/NAND4_in[1] ,
         \SB2_3_28/Component_Function_4/NAND4_in[0] ,
         \SB2_3_29/Component_Function_2/NAND4_in[3] ,
         \SB2_3_29/Component_Function_2/NAND4_in[2] ,
         \SB2_3_29/Component_Function_2/NAND4_in[1] ,
         \SB2_3_29/Component_Function_2/NAND4_in[0] ,
         \SB2_3_29/Component_Function_3/NAND4_in[3] ,
         \SB2_3_29/Component_Function_3/NAND4_in[2] ,
         \SB2_3_29/Component_Function_3/NAND4_in[1] ,
         \SB2_3_29/Component_Function_3/NAND4_in[0] ,
         \SB2_3_29/Component_Function_4/NAND4_in[3] ,
         \SB2_3_29/Component_Function_4/NAND4_in[2] ,
         \SB2_3_29/Component_Function_4/NAND4_in[1] ,
         \SB2_3_29/Component_Function_4/NAND4_in[0] ,
         \SB2_3_30/Component_Function_2/NAND4_in[3] ,
         \SB2_3_30/Component_Function_2/NAND4_in[1] ,
         \SB2_3_30/Component_Function_2/NAND4_in[0] ,
         \SB2_3_30/Component_Function_3/NAND4_in[3] ,
         \SB2_3_30/Component_Function_3/NAND4_in[2] ,
         \SB2_3_30/Component_Function_3/NAND4_in[1] ,
         \SB2_3_30/Component_Function_3/NAND4_in[0] ,
         \SB2_3_30/Component_Function_4/NAND4_in[3] ,
         \SB2_3_30/Component_Function_4/NAND4_in[2] ,
         \SB2_3_30/Component_Function_4/NAND4_in[1] ,
         \SB2_3_30/Component_Function_4/NAND4_in[0] ,
         \SB2_3_31/Component_Function_2/NAND4_in[3] ,
         \SB2_3_31/Component_Function_2/NAND4_in[2] ,
         \SB2_3_31/Component_Function_2/NAND4_in[1] ,
         \SB2_3_31/Component_Function_2/NAND4_in[0] ,
         \SB2_3_31/Component_Function_3/NAND4_in[3] ,
         \SB2_3_31/Component_Function_3/NAND4_in[2] ,
         \SB2_3_31/Component_Function_3/NAND4_in[1] ,
         \SB2_3_31/Component_Function_3/NAND4_in[0] ,
         \SB2_3_31/Component_Function_4/NAND4_in[3] ,
         \SB2_3_31/Component_Function_4/NAND4_in[2] ,
         \SB2_3_31/Component_Function_4/NAND4_in[1] ,
         \SB2_3_31/Component_Function_4/NAND4_in[0] ,
         \SB3_0/Component_Function_2/NAND4_in[2] ,
         \SB3_0/Component_Function_2/NAND4_in[1] ,
         \SB3_0/Component_Function_2/NAND4_in[0] ,
         \SB3_0/Component_Function_3/NAND4_in[2] ,
         \SB3_0/Component_Function_3/NAND4_in[1] ,
         \SB3_0/Component_Function_3/NAND4_in[0] ,
         \SB3_0/Component_Function_4/NAND4_in[2] ,
         \SB3_0/Component_Function_4/NAND4_in[1] ,
         \SB3_0/Component_Function_4/NAND4_in[0] ,
         \SB3_1/Component_Function_2/NAND4_in[3] ,
         \SB3_1/Component_Function_2/NAND4_in[2] ,
         \SB3_1/Component_Function_2/NAND4_in[1] ,
         \SB3_1/Component_Function_2/NAND4_in[0] ,
         \SB3_1/Component_Function_3/NAND4_in[3] ,
         \SB3_1/Component_Function_3/NAND4_in[2] ,
         \SB3_1/Component_Function_3/NAND4_in[1] ,
         \SB3_1/Component_Function_3/NAND4_in[0] ,
         \SB3_1/Component_Function_4/NAND4_in[3] ,
         \SB3_1/Component_Function_4/NAND4_in[2] ,
         \SB3_1/Component_Function_4/NAND4_in[1] ,
         \SB3_1/Component_Function_4/NAND4_in[0] ,
         \SB3_2/Component_Function_2/NAND4_in[2] ,
         \SB3_2/Component_Function_2/NAND4_in[1] ,
         \SB3_2/Component_Function_2/NAND4_in[0] ,
         \SB3_2/Component_Function_3/NAND4_in[3] ,
         \SB3_2/Component_Function_3/NAND4_in[2] ,
         \SB3_2/Component_Function_3/NAND4_in[1] ,
         \SB3_2/Component_Function_3/NAND4_in[0] ,
         \SB3_2/Component_Function_4/NAND4_in[2] ,
         \SB3_2/Component_Function_4/NAND4_in[1] ,
         \SB3_2/Component_Function_4/NAND4_in[0] ,
         \SB3_3/Component_Function_2/NAND4_in[2] ,
         \SB3_3/Component_Function_2/NAND4_in[1] ,
         \SB3_3/Component_Function_2/NAND4_in[0] ,
         \SB3_3/Component_Function_3/NAND4_in[3] ,
         \SB3_3/Component_Function_3/NAND4_in[2] ,
         \SB3_3/Component_Function_3/NAND4_in[1] ,
         \SB3_3/Component_Function_3/NAND4_in[0] ,
         \SB3_3/Component_Function_4/NAND4_in[3] ,
         \SB3_3/Component_Function_4/NAND4_in[2] ,
         \SB3_3/Component_Function_4/NAND4_in[1] ,
         \SB3_3/Component_Function_4/NAND4_in[0] ,
         \SB3_4/Component_Function_2/NAND4_in[3] ,
         \SB3_4/Component_Function_2/NAND4_in[1] ,
         \SB3_4/Component_Function_2/NAND4_in[0] ,
         \SB3_4/Component_Function_3/NAND4_in[3] ,
         \SB3_4/Component_Function_3/NAND4_in[2] ,
         \SB3_4/Component_Function_3/NAND4_in[1] ,
         \SB3_4/Component_Function_3/NAND4_in[0] ,
         \SB3_4/Component_Function_4/NAND4_in[3] ,
         \SB3_4/Component_Function_4/NAND4_in[2] ,
         \SB3_4/Component_Function_4/NAND4_in[1] ,
         \SB3_4/Component_Function_4/NAND4_in[0] ,
         \SB3_5/Component_Function_2/NAND4_in[3] ,
         \SB3_5/Component_Function_2/NAND4_in[2] ,
         \SB3_5/Component_Function_2/NAND4_in[1] ,
         \SB3_5/Component_Function_2/NAND4_in[0] ,
         \SB3_5/Component_Function_3/NAND4_in[2] ,
         \SB3_5/Component_Function_3/NAND4_in[1] ,
         \SB3_5/Component_Function_3/NAND4_in[0] ,
         \SB3_5/Component_Function_4/NAND4_in[3] ,
         \SB3_5/Component_Function_4/NAND4_in[2] ,
         \SB3_5/Component_Function_4/NAND4_in[1] ,
         \SB3_5/Component_Function_4/NAND4_in[0] ,
         \SB3_6/Component_Function_2/NAND4_in[3] ,
         \SB3_6/Component_Function_2/NAND4_in[2] ,
         \SB3_6/Component_Function_2/NAND4_in[1] ,
         \SB3_6/Component_Function_2/NAND4_in[0] ,
         \SB3_6/Component_Function_3/NAND4_in[3] ,
         \SB3_6/Component_Function_3/NAND4_in[2] ,
         \SB3_6/Component_Function_3/NAND4_in[1] ,
         \SB3_6/Component_Function_3/NAND4_in[0] ,
         \SB3_6/Component_Function_4/NAND4_in[3] ,
         \SB3_6/Component_Function_4/NAND4_in[2] ,
         \SB3_6/Component_Function_4/NAND4_in[1] ,
         \SB3_6/Component_Function_4/NAND4_in[0] ,
         \SB3_7/Component_Function_2/NAND4_in[3] ,
         \SB3_7/Component_Function_2/NAND4_in[2] ,
         \SB3_7/Component_Function_2/NAND4_in[1] ,
         \SB3_7/Component_Function_2/NAND4_in[0] ,
         \SB3_7/Component_Function_3/NAND4_in[3] ,
         \SB3_7/Component_Function_3/NAND4_in[1] ,
         \SB3_7/Component_Function_3/NAND4_in[0] ,
         \SB3_7/Component_Function_4/NAND4_in[3] ,
         \SB3_7/Component_Function_4/NAND4_in[2] ,
         \SB3_7/Component_Function_4/NAND4_in[1] ,
         \SB3_7/Component_Function_4/NAND4_in[0] ,
         \SB3_8/Component_Function_2/NAND4_in[3] ,
         \SB3_8/Component_Function_2/NAND4_in[2] ,
         \SB3_8/Component_Function_2/NAND4_in[1] ,
         \SB3_8/Component_Function_2/NAND4_in[0] ,
         \SB3_8/Component_Function_3/NAND4_in[3] ,
         \SB3_8/Component_Function_3/NAND4_in[2] ,
         \SB3_8/Component_Function_3/NAND4_in[1] ,
         \SB3_8/Component_Function_3/NAND4_in[0] ,
         \SB3_8/Component_Function_4/NAND4_in[3] ,
         \SB3_8/Component_Function_4/NAND4_in[1] ,
         \SB3_8/Component_Function_4/NAND4_in[0] ,
         \SB3_9/Component_Function_2/NAND4_in[3] ,
         \SB3_9/Component_Function_2/NAND4_in[2] ,
         \SB3_9/Component_Function_2/NAND4_in[1] ,
         \SB3_9/Component_Function_2/NAND4_in[0] ,
         \SB3_9/Component_Function_3/NAND4_in[3] ,
         \SB3_9/Component_Function_3/NAND4_in[2] ,
         \SB3_9/Component_Function_3/NAND4_in[1] ,
         \SB3_9/Component_Function_3/NAND4_in[0] ,
         \SB3_9/Component_Function_4/NAND4_in[3] ,
         \SB3_9/Component_Function_4/NAND4_in[2] ,
         \SB3_9/Component_Function_4/NAND4_in[1] ,
         \SB3_9/Component_Function_4/NAND4_in[0] ,
         \SB3_10/Component_Function_2/NAND4_in[3] ,
         \SB3_10/Component_Function_2/NAND4_in[2] ,
         \SB3_10/Component_Function_2/NAND4_in[1] ,
         \SB3_10/Component_Function_2/NAND4_in[0] ,
         \SB3_10/Component_Function_3/NAND4_in[3] ,
         \SB3_10/Component_Function_3/NAND4_in[2] ,
         \SB3_10/Component_Function_3/NAND4_in[1] ,
         \SB3_10/Component_Function_3/NAND4_in[0] ,
         \SB3_10/Component_Function_4/NAND4_in[3] ,
         \SB3_10/Component_Function_4/NAND4_in[1] ,
         \SB3_10/Component_Function_4/NAND4_in[0] ,
         \SB3_11/Component_Function_2/NAND4_in[3] ,
         \SB3_11/Component_Function_2/NAND4_in[2] ,
         \SB3_11/Component_Function_2/NAND4_in[1] ,
         \SB3_11/Component_Function_2/NAND4_in[0] ,
         \SB3_11/Component_Function_3/NAND4_in[2] ,
         \SB3_11/Component_Function_3/NAND4_in[1] ,
         \SB3_11/Component_Function_3/NAND4_in[0] ,
         \SB3_11/Component_Function_4/NAND4_in[3] ,
         \SB3_11/Component_Function_4/NAND4_in[2] ,
         \SB3_11/Component_Function_4/NAND4_in[1] ,
         \SB3_11/Component_Function_4/NAND4_in[0] ,
         \SB3_12/Component_Function_2/NAND4_in[3] ,
         \SB3_12/Component_Function_2/NAND4_in[1] ,
         \SB3_12/Component_Function_2/NAND4_in[0] ,
         \SB3_12/Component_Function_3/NAND4_in[3] ,
         \SB3_12/Component_Function_3/NAND4_in[2] ,
         \SB3_12/Component_Function_3/NAND4_in[1] ,
         \SB3_12/Component_Function_3/NAND4_in[0] ,
         \SB3_12/Component_Function_4/NAND4_in[3] ,
         \SB3_12/Component_Function_4/NAND4_in[2] ,
         \SB3_12/Component_Function_4/NAND4_in[1] ,
         \SB3_12/Component_Function_4/NAND4_in[0] ,
         \SB3_13/Component_Function_2/NAND4_in[3] ,
         \SB3_13/Component_Function_2/NAND4_in[2] ,
         \SB3_13/Component_Function_2/NAND4_in[1] ,
         \SB3_13/Component_Function_2/NAND4_in[0] ,
         \SB3_13/Component_Function_3/NAND4_in[3] ,
         \SB3_13/Component_Function_3/NAND4_in[2] ,
         \SB3_13/Component_Function_3/NAND4_in[1] ,
         \SB3_13/Component_Function_3/NAND4_in[0] ,
         \SB3_13/Component_Function_4/NAND4_in[3] ,
         \SB3_13/Component_Function_4/NAND4_in[2] ,
         \SB3_13/Component_Function_4/NAND4_in[1] ,
         \SB3_13/Component_Function_4/NAND4_in[0] ,
         \SB3_14/Component_Function_2/NAND4_in[3] ,
         \SB3_14/Component_Function_2/NAND4_in[2] ,
         \SB3_14/Component_Function_2/NAND4_in[1] ,
         \SB3_14/Component_Function_2/NAND4_in[0] ,
         \SB3_14/Component_Function_3/NAND4_in[2] ,
         \SB3_14/Component_Function_3/NAND4_in[1] ,
         \SB3_14/Component_Function_3/NAND4_in[0] ,
         \SB3_14/Component_Function_4/NAND4_in[3] ,
         \SB3_14/Component_Function_4/NAND4_in[2] ,
         \SB3_14/Component_Function_4/NAND4_in[1] ,
         \SB3_14/Component_Function_4/NAND4_in[0] ,
         \SB3_15/Component_Function_2/NAND4_in[2] ,
         \SB3_15/Component_Function_2/NAND4_in[1] ,
         \SB3_15/Component_Function_2/NAND4_in[0] ,
         \SB3_15/Component_Function_3/NAND4_in[3] ,
         \SB3_15/Component_Function_3/NAND4_in[2] ,
         \SB3_15/Component_Function_3/NAND4_in[1] ,
         \SB3_15/Component_Function_3/NAND4_in[0] ,
         \SB3_15/Component_Function_4/NAND4_in[3] ,
         \SB3_15/Component_Function_4/NAND4_in[2] ,
         \SB3_15/Component_Function_4/NAND4_in[1] ,
         \SB3_15/Component_Function_4/NAND4_in[0] ,
         \SB3_16/Component_Function_2/NAND4_in[3] ,
         \SB3_16/Component_Function_2/NAND4_in[2] ,
         \SB3_16/Component_Function_2/NAND4_in[1] ,
         \SB3_16/Component_Function_2/NAND4_in[0] ,
         \SB3_16/Component_Function_3/NAND4_in[3] ,
         \SB3_16/Component_Function_3/NAND4_in[2] ,
         \SB3_16/Component_Function_3/NAND4_in[1] ,
         \SB3_16/Component_Function_3/NAND4_in[0] ,
         \SB3_16/Component_Function_4/NAND4_in[3] ,
         \SB3_16/Component_Function_4/NAND4_in[1] ,
         \SB3_16/Component_Function_4/NAND4_in[0] ,
         \SB3_17/Component_Function_2/NAND4_in[3] ,
         \SB3_17/Component_Function_2/NAND4_in[2] ,
         \SB3_17/Component_Function_2/NAND4_in[1] ,
         \SB3_17/Component_Function_2/NAND4_in[0] ,
         \SB3_17/Component_Function_3/NAND4_in[3] ,
         \SB3_17/Component_Function_3/NAND4_in[2] ,
         \SB3_17/Component_Function_3/NAND4_in[1] ,
         \SB3_17/Component_Function_3/NAND4_in[0] ,
         \SB3_17/Component_Function_4/NAND4_in[3] ,
         \SB3_17/Component_Function_4/NAND4_in[2] ,
         \SB3_17/Component_Function_4/NAND4_in[1] ,
         \SB3_17/Component_Function_4/NAND4_in[0] ,
         \SB3_18/Component_Function_2/NAND4_in[3] ,
         \SB3_18/Component_Function_2/NAND4_in[2] ,
         \SB3_18/Component_Function_2/NAND4_in[1] ,
         \SB3_18/Component_Function_2/NAND4_in[0] ,
         \SB3_18/Component_Function_3/NAND4_in[3] ,
         \SB3_18/Component_Function_3/NAND4_in[2] ,
         \SB3_18/Component_Function_3/NAND4_in[1] ,
         \SB3_18/Component_Function_3/NAND4_in[0] ,
         \SB3_18/Component_Function_4/NAND4_in[3] ,
         \SB3_18/Component_Function_4/NAND4_in[2] ,
         \SB3_18/Component_Function_4/NAND4_in[1] ,
         \SB3_18/Component_Function_4/NAND4_in[0] ,
         \SB3_19/Component_Function_2/NAND4_in[3] ,
         \SB3_19/Component_Function_2/NAND4_in[2] ,
         \SB3_19/Component_Function_2/NAND4_in[1] ,
         \SB3_19/Component_Function_2/NAND4_in[0] ,
         \SB3_19/Component_Function_3/NAND4_in[3] ,
         \SB3_19/Component_Function_3/NAND4_in[2] ,
         \SB3_19/Component_Function_3/NAND4_in[1] ,
         \SB3_19/Component_Function_3/NAND4_in[0] ,
         \SB3_19/Component_Function_4/NAND4_in[3] ,
         \SB3_19/Component_Function_4/NAND4_in[2] ,
         \SB3_19/Component_Function_4/NAND4_in[1] ,
         \SB3_19/Component_Function_4/NAND4_in[0] ,
         \SB3_20/Component_Function_2/NAND4_in[3] ,
         \SB3_20/Component_Function_2/NAND4_in[2] ,
         \SB3_20/Component_Function_2/NAND4_in[1] ,
         \SB3_20/Component_Function_2/NAND4_in[0] ,
         \SB3_20/Component_Function_3/NAND4_in[2] ,
         \SB3_20/Component_Function_3/NAND4_in[1] ,
         \SB3_20/Component_Function_3/NAND4_in[0] ,
         \SB3_20/Component_Function_4/NAND4_in[3] ,
         \SB3_20/Component_Function_4/NAND4_in[2] ,
         \SB3_20/Component_Function_4/NAND4_in[1] ,
         \SB3_20/Component_Function_4/NAND4_in[0] ,
         \SB3_21/Component_Function_2/NAND4_in[3] ,
         \SB3_21/Component_Function_2/NAND4_in[2] ,
         \SB3_21/Component_Function_2/NAND4_in[1] ,
         \SB3_21/Component_Function_2/NAND4_in[0] ,
         \SB3_21/Component_Function_3/NAND4_in[3] ,
         \SB3_21/Component_Function_3/NAND4_in[2] ,
         \SB3_21/Component_Function_3/NAND4_in[1] ,
         \SB3_21/Component_Function_3/NAND4_in[0] ,
         \SB3_21/Component_Function_4/NAND4_in[3] ,
         \SB3_21/Component_Function_4/NAND4_in[2] ,
         \SB3_21/Component_Function_4/NAND4_in[1] ,
         \SB3_21/Component_Function_4/NAND4_in[0] ,
         \SB3_22/Component_Function_2/NAND4_in[2] ,
         \SB3_22/Component_Function_2/NAND4_in[1] ,
         \SB3_22/Component_Function_2/NAND4_in[0] ,
         \SB3_22/Component_Function_3/NAND4_in[3] ,
         \SB3_22/Component_Function_3/NAND4_in[2] ,
         \SB3_22/Component_Function_3/NAND4_in[1] ,
         \SB3_22/Component_Function_3/NAND4_in[0] ,
         \SB3_22/Component_Function_4/NAND4_in[3] ,
         \SB3_22/Component_Function_4/NAND4_in[2] ,
         \SB3_22/Component_Function_4/NAND4_in[1] ,
         \SB3_22/Component_Function_4/NAND4_in[0] ,
         \SB3_23/Component_Function_2/NAND4_in[3] ,
         \SB3_23/Component_Function_2/NAND4_in[2] ,
         \SB3_23/Component_Function_2/NAND4_in[1] ,
         \SB3_23/Component_Function_2/NAND4_in[0] ,
         \SB3_23/Component_Function_3/NAND4_in[2] ,
         \SB3_23/Component_Function_3/NAND4_in[1] ,
         \SB3_23/Component_Function_3/NAND4_in[0] ,
         \SB3_23/Component_Function_4/NAND4_in[3] ,
         \SB3_23/Component_Function_4/NAND4_in[1] ,
         \SB3_23/Component_Function_4/NAND4_in[0] ,
         \SB3_24/Component_Function_2/NAND4_in[3] ,
         \SB3_24/Component_Function_2/NAND4_in[2] ,
         \SB3_24/Component_Function_2/NAND4_in[1] ,
         \SB3_24/Component_Function_2/NAND4_in[0] ,
         \SB3_24/Component_Function_3/NAND4_in[2] ,
         \SB3_24/Component_Function_3/NAND4_in[1] ,
         \SB3_24/Component_Function_4/NAND4_in[3] ,
         \SB3_24/Component_Function_4/NAND4_in[2] ,
         \SB3_24/Component_Function_4/NAND4_in[1] ,
         \SB3_24/Component_Function_4/NAND4_in[0] ,
         \SB3_25/Component_Function_2/NAND4_in[3] ,
         \SB3_25/Component_Function_2/NAND4_in[2] ,
         \SB3_25/Component_Function_2/NAND4_in[1] ,
         \SB3_25/Component_Function_2/NAND4_in[0] ,
         \SB3_25/Component_Function_3/NAND4_in[3] ,
         \SB3_25/Component_Function_3/NAND4_in[2] ,
         \SB3_25/Component_Function_3/NAND4_in[1] ,
         \SB3_25/Component_Function_3/NAND4_in[0] ,
         \SB3_25/Component_Function_4/NAND4_in[3] ,
         \SB3_25/Component_Function_4/NAND4_in[2] ,
         \SB3_25/Component_Function_4/NAND4_in[1] ,
         \SB3_25/Component_Function_4/NAND4_in[0] ,
         \SB3_26/Component_Function_2/NAND4_in[2] ,
         \SB3_26/Component_Function_2/NAND4_in[1] ,
         \SB3_26/Component_Function_2/NAND4_in[0] ,
         \SB3_26/Component_Function_3/NAND4_in[3] ,
         \SB3_26/Component_Function_3/NAND4_in[2] ,
         \SB3_26/Component_Function_3/NAND4_in[1] ,
         \SB3_26/Component_Function_3/NAND4_in[0] ,
         \SB3_26/Component_Function_4/NAND4_in[3] ,
         \SB3_26/Component_Function_4/NAND4_in[2] ,
         \SB3_26/Component_Function_4/NAND4_in[1] ,
         \SB3_26/Component_Function_4/NAND4_in[0] ,
         \SB3_27/Component_Function_2/NAND4_in[3] ,
         \SB3_27/Component_Function_2/NAND4_in[2] ,
         \SB3_27/Component_Function_2/NAND4_in[1] ,
         \SB3_27/Component_Function_2/NAND4_in[0] ,
         \SB3_27/Component_Function_3/NAND4_in[3] ,
         \SB3_27/Component_Function_3/NAND4_in[2] ,
         \SB3_27/Component_Function_3/NAND4_in[1] ,
         \SB3_27/Component_Function_3/NAND4_in[0] ,
         \SB3_27/Component_Function_4/NAND4_in[3] ,
         \SB3_27/Component_Function_4/NAND4_in[2] ,
         \SB3_27/Component_Function_4/NAND4_in[1] ,
         \SB3_27/Component_Function_4/NAND4_in[0] ,
         \SB3_28/Component_Function_2/NAND4_in[3] ,
         \SB3_28/Component_Function_2/NAND4_in[2] ,
         \SB3_28/Component_Function_2/NAND4_in[1] ,
         \SB3_28/Component_Function_2/NAND4_in[0] ,
         \SB3_28/Component_Function_3/NAND4_in[3] ,
         \SB3_28/Component_Function_3/NAND4_in[1] ,
         \SB3_28/Component_Function_3/NAND4_in[0] ,
         \SB3_28/Component_Function_4/NAND4_in[3] ,
         \SB3_28/Component_Function_4/NAND4_in[2] ,
         \SB3_28/Component_Function_4/NAND4_in[1] ,
         \SB3_28/Component_Function_4/NAND4_in[0] ,
         \SB3_29/Component_Function_2/NAND4_in[3] ,
         \SB3_29/Component_Function_2/NAND4_in[1] ,
         \SB3_29/Component_Function_2/NAND4_in[0] ,
         \SB3_29/Component_Function_3/NAND4_in[2] ,
         \SB3_29/Component_Function_3/NAND4_in[1] ,
         \SB3_29/Component_Function_3/NAND4_in[0] ,
         \SB3_29/Component_Function_4/NAND4_in[3] ,
         \SB3_29/Component_Function_4/NAND4_in[2] ,
         \SB3_29/Component_Function_4/NAND4_in[1] ,
         \SB3_29/Component_Function_4/NAND4_in[0] ,
         \SB3_30/Component_Function_2/NAND4_in[2] ,
         \SB3_30/Component_Function_2/NAND4_in[1] ,
         \SB3_30/Component_Function_2/NAND4_in[0] ,
         \SB3_30/Component_Function_3/NAND4_in[3] ,
         \SB3_30/Component_Function_3/NAND4_in[2] ,
         \SB3_30/Component_Function_3/NAND4_in[1] ,
         \SB3_30/Component_Function_3/NAND4_in[0] ,
         \SB3_30/Component_Function_4/NAND4_in[3] ,
         \SB3_30/Component_Function_4/NAND4_in[2] ,
         \SB3_30/Component_Function_4/NAND4_in[1] ,
         \SB3_30/Component_Function_4/NAND4_in[0] ,
         \SB3_31/Component_Function_2/NAND4_in[2] ,
         \SB3_31/Component_Function_2/NAND4_in[1] ,
         \SB3_31/Component_Function_2/NAND4_in[0] ,
         \SB3_31/Component_Function_3/NAND4_in[3] ,
         \SB3_31/Component_Function_3/NAND4_in[2] ,
         \SB3_31/Component_Function_3/NAND4_in[1] ,
         \SB3_31/Component_Function_3/NAND4_in[0] ,
         \SB3_31/Component_Function_4/NAND4_in[3] ,
         \SB3_31/Component_Function_4/NAND4_in[2] ,
         \SB3_31/Component_Function_4/NAND4_in[1] ,
         \SB3_31/Component_Function_4/NAND4_in[0] ,
         \SB4_0/Component_Function_2/NAND4_in[3] ,
         \SB4_0/Component_Function_2/NAND4_in[2] ,
         \SB4_0/Component_Function_2/NAND4_in[1] ,
         \SB4_0/Component_Function_2/NAND4_in[0] ,
         \SB4_0/Component_Function_3/NAND4_in[1] ,
         \SB4_0/Component_Function_3/NAND4_in[0] ,
         \SB4_0/Component_Function_4/NAND4_in[3] ,
         \SB4_0/Component_Function_4/NAND4_in[2] ,
         \SB4_0/Component_Function_4/NAND4_in[1] ,
         \SB4_0/Component_Function_4/NAND4_in[0] ,
         \SB4_1/Component_Function_2/NAND4_in[3] ,
         \SB4_1/Component_Function_2/NAND4_in[2] ,
         \SB4_1/Component_Function_2/NAND4_in[1] ,
         \SB4_1/Component_Function_3/NAND4_in[3] ,
         \SB4_1/Component_Function_3/NAND4_in[1] ,
         \SB4_1/Component_Function_3/NAND4_in[0] ,
         \SB4_1/Component_Function_4/NAND4_in[3] ,
         \SB4_1/Component_Function_4/NAND4_in[2] ,
         \SB4_2/Component_Function_2/NAND4_in[3] ,
         \SB4_2/Component_Function_2/NAND4_in[2] ,
         \SB4_2/Component_Function_2/NAND4_in[1] ,
         \SB4_2/Component_Function_2/NAND4_in[0] ,
         \SB4_2/Component_Function_3/NAND4_in[3] ,
         \SB4_2/Component_Function_3/NAND4_in[1] ,
         \SB4_2/Component_Function_3/NAND4_in[0] ,
         \SB4_2/Component_Function_4/NAND4_in[2] ,
         \SB4_2/Component_Function_4/NAND4_in[1] ,
         \SB4_2/Component_Function_4/NAND4_in[0] ,
         \SB4_3/Component_Function_2/NAND4_in[2] ,
         \SB4_3/Component_Function_2/NAND4_in[1] ,
         \SB4_3/Component_Function_3/NAND4_in[3] ,
         \SB4_3/Component_Function_3/NAND4_in[2] ,
         \SB4_3/Component_Function_3/NAND4_in[1] ,
         \SB4_3/Component_Function_3/NAND4_in[0] ,
         \SB4_3/Component_Function_4/NAND4_in[3] ,
         \SB4_3/Component_Function_4/NAND4_in[2] ,
         \SB4_3/Component_Function_4/NAND4_in[1] ,
         \SB4_3/Component_Function_4/NAND4_in[0] ,
         \SB4_4/Component_Function_2/NAND4_in[2] ,
         \SB4_4/Component_Function_2/NAND4_in[1] ,
         \SB4_4/Component_Function_2/NAND4_in[0] ,
         \SB4_4/Component_Function_3/NAND4_in[3] ,
         \SB4_4/Component_Function_3/NAND4_in[1] ,
         \SB4_4/Component_Function_3/NAND4_in[0] ,
         \SB4_4/Component_Function_4/NAND4_in[3] ,
         \SB4_4/Component_Function_4/NAND4_in[2] ,
         \SB4_4/Component_Function_4/NAND4_in[0] ,
         \SB4_5/Component_Function_2/NAND4_in[3] ,
         \SB4_5/Component_Function_2/NAND4_in[2] ,
         \SB4_5/Component_Function_2/NAND4_in[1] ,
         \SB4_5/Component_Function_2/NAND4_in[0] ,
         \SB4_5/Component_Function_3/NAND4_in[3] ,
         \SB4_5/Component_Function_3/NAND4_in[2] ,
         \SB4_5/Component_Function_3/NAND4_in[1] ,
         \SB4_5/Component_Function_3/NAND4_in[0] ,
         \SB4_5/Component_Function_4/NAND4_in[2] ,
         \SB4_5/Component_Function_4/NAND4_in[0] ,
         \SB4_6/Component_Function_2/NAND4_in[3] ,
         \SB4_6/Component_Function_2/NAND4_in[2] ,
         \SB4_6/Component_Function_2/NAND4_in[1] ,
         \SB4_6/Component_Function_3/NAND4_in[3] ,
         \SB4_6/Component_Function_3/NAND4_in[2] ,
         \SB4_6/Component_Function_3/NAND4_in[1] ,
         \SB4_6/Component_Function_3/NAND4_in[0] ,
         \SB4_6/Component_Function_4/NAND4_in[3] ,
         \SB4_6/Component_Function_4/NAND4_in[2] ,
         \SB4_6/Component_Function_4/NAND4_in[0] ,
         \SB4_7/Component_Function_2/NAND4_in[2] ,
         \SB4_7/Component_Function_2/NAND4_in[1] ,
         \SB4_7/Component_Function_3/NAND4_in[3] ,
         \SB4_7/Component_Function_3/NAND4_in[2] ,
         \SB4_7/Component_Function_3/NAND4_in[1] ,
         \SB4_7/Component_Function_3/NAND4_in[0] ,
         \SB4_7/Component_Function_4/NAND4_in[2] ,
         \SB4_7/Component_Function_4/NAND4_in[1] ,
         \SB4_7/Component_Function_4/NAND4_in[0] ,
         \SB4_8/Component_Function_2/NAND4_in[2] ,
         \SB4_8/Component_Function_2/NAND4_in[1] ,
         \SB4_8/Component_Function_2/NAND4_in[0] ,
         \SB4_8/Component_Function_3/NAND4_in[3] ,
         \SB4_8/Component_Function_3/NAND4_in[1] ,
         \SB4_8/Component_Function_3/NAND4_in[0] ,
         \SB4_8/Component_Function_4/NAND4_in[3] ,
         \SB4_8/Component_Function_4/NAND4_in[2] ,
         \SB4_8/Component_Function_4/NAND4_in[1] ,
         \SB4_8/Component_Function_4/NAND4_in[0] ,
         \SB4_9/Component_Function_2/NAND4_in[3] ,
         \SB4_9/Component_Function_2/NAND4_in[2] ,
         \SB4_9/Component_Function_2/NAND4_in[1] ,
         \SB4_9/Component_Function_2/NAND4_in[0] ,
         \SB4_9/Component_Function_3/NAND4_in[3] ,
         \SB4_9/Component_Function_3/NAND4_in[2] ,
         \SB4_9/Component_Function_3/NAND4_in[1] ,
         \SB4_9/Component_Function_3/NAND4_in[0] ,
         \SB4_9/Component_Function_4/NAND4_in[3] ,
         \SB4_9/Component_Function_4/NAND4_in[0] ,
         \SB4_10/Component_Function_2/NAND4_in[2] ,
         \SB4_10/Component_Function_2/NAND4_in[1] ,
         \SB4_10/Component_Function_3/NAND4_in[3] ,
         \SB4_10/Component_Function_3/NAND4_in[0] ,
         \SB4_10/Component_Function_4/NAND4_in[3] ,
         \SB4_10/Component_Function_4/NAND4_in[2] ,
         \SB4_10/Component_Function_4/NAND4_in[1] ,
         \SB4_10/Component_Function_4/NAND4_in[0] ,
         \SB4_11/Component_Function_2/NAND4_in[2] ,
         \SB4_11/Component_Function_2/NAND4_in[1] ,
         \SB4_11/Component_Function_2/NAND4_in[0] ,
         \SB4_11/Component_Function_3/NAND4_in[3] ,
         \SB4_11/Component_Function_3/NAND4_in[0] ,
         \SB4_11/Component_Function_4/NAND4_in[2] ,
         \SB4_11/Component_Function_4/NAND4_in[1] ,
         \SB4_11/Component_Function_4/NAND4_in[0] ,
         \SB4_12/Component_Function_2/NAND4_in[2] ,
         \SB4_12/Component_Function_2/NAND4_in[1] ,
         \SB4_12/Component_Function_2/NAND4_in[0] ,
         \SB4_12/Component_Function_3/NAND4_in[3] ,
         \SB4_12/Component_Function_3/NAND4_in[2] ,
         \SB4_12/Component_Function_3/NAND4_in[1] ,
         \SB4_12/Component_Function_3/NAND4_in[0] ,
         \SB4_12/Component_Function_4/NAND4_in[3] ,
         \SB4_12/Component_Function_4/NAND4_in[2] ,
         \SB4_12/Component_Function_4/NAND4_in[1] ,
         \SB4_12/Component_Function_4/NAND4_in[0] ,
         \SB4_13/Component_Function_2/NAND4_in[3] ,
         \SB4_13/Component_Function_2/NAND4_in[2] ,
         \SB4_13/Component_Function_2/NAND4_in[1] ,
         \SB4_13/Component_Function_3/NAND4_in[3] ,
         \SB4_13/Component_Function_3/NAND4_in[1] ,
         \SB4_13/Component_Function_3/NAND4_in[0] ,
         \SB4_13/Component_Function_4/NAND4_in[3] ,
         \SB4_13/Component_Function_4/NAND4_in[2] ,
         \SB4_13/Component_Function_4/NAND4_in[1] ,
         \SB4_13/Component_Function_4/NAND4_in[0] ,
         \SB4_14/Component_Function_2/NAND4_in[2] ,
         \SB4_14/Component_Function_2/NAND4_in[1] ,
         \SB4_14/Component_Function_2/NAND4_in[0] ,
         \SB4_14/Component_Function_3/NAND4_in[3] ,
         \SB4_14/Component_Function_3/NAND4_in[2] ,
         \SB4_14/Component_Function_3/NAND4_in[1] ,
         \SB4_14/Component_Function_3/NAND4_in[0] ,
         \SB4_14/Component_Function_4/NAND4_in[2] ,
         \SB4_14/Component_Function_4/NAND4_in[1] ,
         \SB4_14/Component_Function_4/NAND4_in[0] ,
         \SB4_15/Component_Function_2/NAND4_in[2] ,
         \SB4_15/Component_Function_2/NAND4_in[1] ,
         \SB4_15/Component_Function_2/NAND4_in[0] ,
         \SB4_15/Component_Function_3/NAND4_in[3] ,
         \SB4_15/Component_Function_3/NAND4_in[2] ,
         \SB4_15/Component_Function_3/NAND4_in[1] ,
         \SB4_15/Component_Function_3/NAND4_in[0] ,
         \SB4_15/Component_Function_4/NAND4_in[3] ,
         \SB4_15/Component_Function_4/NAND4_in[2] ,
         \SB4_15/Component_Function_4/NAND4_in[1] ,
         \SB4_15/Component_Function_4/NAND4_in[0] ,
         \SB4_16/Component_Function_2/NAND4_in[3] ,
         \SB4_16/Component_Function_2/NAND4_in[2] ,
         \SB4_16/Component_Function_2/NAND4_in[1] ,
         \SB4_16/Component_Function_3/NAND4_in[3] ,
         \SB4_16/Component_Function_3/NAND4_in[2] ,
         \SB4_16/Component_Function_3/NAND4_in[1] ,
         \SB4_16/Component_Function_3/NAND4_in[0] ,
         \SB4_16/Component_Function_4/NAND4_in[3] ,
         \SB4_16/Component_Function_4/NAND4_in[2] ,
         \SB4_16/Component_Function_4/NAND4_in[1] ,
         \SB4_17/Component_Function_2/NAND4_in[2] ,
         \SB4_17/Component_Function_2/NAND4_in[1] ,
         \SB4_17/Component_Function_3/NAND4_in[3] ,
         \SB4_17/Component_Function_3/NAND4_in[0] ,
         \SB4_17/Component_Function_4/NAND4_in[3] ,
         \SB4_17/Component_Function_4/NAND4_in[2] ,
         \SB4_18/Component_Function_2/NAND4_in[2] ,
         \SB4_18/Component_Function_2/NAND4_in[1] ,
         \SB4_18/Component_Function_2/NAND4_in[0] ,
         \SB4_18/Component_Function_3/NAND4_in[3] ,
         \SB4_18/Component_Function_3/NAND4_in[2] ,
         \SB4_18/Component_Function_3/NAND4_in[1] ,
         \SB4_18/Component_Function_3/NAND4_in[0] ,
         \SB4_18/Component_Function_4/NAND4_in[2] ,
         \SB4_18/Component_Function_4/NAND4_in[1] ,
         \SB4_18/Component_Function_4/NAND4_in[0] ,
         \SB4_19/Component_Function_2/NAND4_in[2] ,
         \SB4_19/Component_Function_2/NAND4_in[1] ,
         \SB4_19/Component_Function_2/NAND4_in[0] ,
         \SB4_19/Component_Function_3/NAND4_in[3] ,
         \SB4_19/Component_Function_3/NAND4_in[2] ,
         \SB4_19/Component_Function_3/NAND4_in[1] ,
         \SB4_19/Component_Function_3/NAND4_in[0] ,
         \SB4_19/Component_Function_4/NAND4_in[3] ,
         \SB4_19/Component_Function_4/NAND4_in[2] ,
         \SB4_19/Component_Function_4/NAND4_in[0] ,
         \SB4_20/Component_Function_2/NAND4_in[3] ,
         \SB4_20/Component_Function_2/NAND4_in[2] ,
         \SB4_20/Component_Function_2/NAND4_in[1] ,
         \SB4_20/Component_Function_2/NAND4_in[0] ,
         \SB4_20/Component_Function_3/NAND4_in[3] ,
         \SB4_20/Component_Function_3/NAND4_in[1] ,
         \SB4_20/Component_Function_3/NAND4_in[0] ,
         \SB4_20/Component_Function_4/NAND4_in[3] ,
         \SB4_20/Component_Function_4/NAND4_in[2] ,
         \SB4_20/Component_Function_4/NAND4_in[1] ,
         \SB4_20/Component_Function_4/NAND4_in[0] ,
         \SB4_21/Component_Function_2/NAND4_in[2] ,
         \SB4_21/Component_Function_2/NAND4_in[1] ,
         \SB4_21/Component_Function_2/NAND4_in[0] ,
         \SB4_21/Component_Function_3/NAND4_in[3] ,
         \SB4_21/Component_Function_3/NAND4_in[1] ,
         \SB4_21/Component_Function_3/NAND4_in[0] ,
         \SB4_21/Component_Function_4/NAND4_in[2] ,
         \SB4_21/Component_Function_4/NAND4_in[1] ,
         \SB4_21/Component_Function_4/NAND4_in[0] ,
         \SB4_22/Component_Function_2/NAND4_in[2] ,
         \SB4_22/Component_Function_2/NAND4_in[1] ,
         \SB4_22/Component_Function_3/NAND4_in[3] ,
         \SB4_22/Component_Function_3/NAND4_in[2] ,
         \SB4_22/Component_Function_3/NAND4_in[1] ,
         \SB4_22/Component_Function_3/NAND4_in[0] ,
         \SB4_22/Component_Function_4/NAND4_in[2] ,
         \SB4_22/Component_Function_4/NAND4_in[1] ,
         \SB4_22/Component_Function_4/NAND4_in[0] ,
         \SB4_23/Component_Function_2/NAND4_in[2] ,
         \SB4_23/Component_Function_2/NAND4_in[1] ,
         \SB4_23/Component_Function_2/NAND4_in[0] ,
         \SB4_23/Component_Function_3/NAND4_in[3] ,
         \SB4_23/Component_Function_3/NAND4_in[2] ,
         \SB4_23/Component_Function_3/NAND4_in[1] ,
         \SB4_23/Component_Function_3/NAND4_in[0] ,
         \SB4_23/Component_Function_4/NAND4_in[3] ,
         \SB4_23/Component_Function_4/NAND4_in[2] ,
         \SB4_23/Component_Function_4/NAND4_in[1] ,
         \SB4_23/Component_Function_4/NAND4_in[0] ,
         \SB4_24/Component_Function_2/NAND4_in[3] ,
         \SB4_24/Component_Function_2/NAND4_in[2] ,
         \SB4_24/Component_Function_2/NAND4_in[1] ,
         \SB4_24/Component_Function_3/NAND4_in[3] ,
         \SB4_24/Component_Function_3/NAND4_in[1] ,
         \SB4_24/Component_Function_3/NAND4_in[0] ,
         \SB4_24/Component_Function_4/NAND4_in[3] ,
         \SB4_24/Component_Function_4/NAND4_in[2] ,
         \SB4_24/Component_Function_4/NAND4_in[1] ,
         \SB4_24/Component_Function_4/NAND4_in[0] ,
         \SB4_25/Component_Function_2/NAND4_in[3] ,
         \SB4_25/Component_Function_2/NAND4_in[2] ,
         \SB4_25/Component_Function_2/NAND4_in[1] ,
         \SB4_25/Component_Function_2/NAND4_in[0] ,
         \SB4_25/Component_Function_3/NAND4_in[3] ,
         \SB4_25/Component_Function_3/NAND4_in[1] ,
         \SB4_25/Component_Function_3/NAND4_in[0] ,
         \SB4_25/Component_Function_4/NAND4_in[2] ,
         \SB4_25/Component_Function_4/NAND4_in[1] ,
         \SB4_25/Component_Function_4/NAND4_in[0] ,
         \SB4_26/Component_Function_2/NAND4_in[2] ,
         \SB4_26/Component_Function_2/NAND4_in[1] ,
         \SB4_26/Component_Function_3/NAND4_in[3] ,
         \SB4_26/Component_Function_3/NAND4_in[1] ,
         \SB4_26/Component_Function_3/NAND4_in[0] ,
         \SB4_26/Component_Function_4/NAND4_in[3] ,
         \SB4_26/Component_Function_4/NAND4_in[2] ,
         \SB4_27/Component_Function_2/NAND4_in[2] ,
         \SB4_27/Component_Function_2/NAND4_in[1] ,
         \SB4_27/Component_Function_3/NAND4_in[3] ,
         \SB4_27/Component_Function_3/NAND4_in[2] ,
         \SB4_27/Component_Function_3/NAND4_in[1] ,
         \SB4_27/Component_Function_3/NAND4_in[0] ,
         \SB4_27/Component_Function_4/NAND4_in[3] ,
         \SB4_27/Component_Function_4/NAND4_in[2] ,
         \SB4_27/Component_Function_4/NAND4_in[1] ,
         \SB4_27/Component_Function_4/NAND4_in[0] ,
         \SB4_28/Component_Function_2/NAND4_in[2] ,
         \SB4_28/Component_Function_2/NAND4_in[1] ,
         \SB4_28/Component_Function_2/NAND4_in[0] ,
         \SB4_28/Component_Function_3/NAND4_in[3] ,
         \SB4_28/Component_Function_3/NAND4_in[1] ,
         \SB4_28/Component_Function_3/NAND4_in[0] ,
         \SB4_28/Component_Function_4/NAND4_in[3] ,
         \SB4_28/Component_Function_4/NAND4_in[2] ,
         \SB4_28/Component_Function_4/NAND4_in[1] ,
         \SB4_28/Component_Function_4/NAND4_in[0] ,
         \SB4_29/Component_Function_2/NAND4_in[2] ,
         \SB4_29/Component_Function_2/NAND4_in[1] ,
         \SB4_29/Component_Function_3/NAND4_in[3] ,
         \SB4_29/Component_Function_3/NAND4_in[1] ,
         \SB4_29/Component_Function_3/NAND4_in[0] ,
         \SB4_29/Component_Function_4/NAND4_in[2] ,
         \SB4_29/Component_Function_4/NAND4_in[1] ,
         \SB4_30/Component_Function_2/NAND4_in[2] ,
         \SB4_30/Component_Function_2/NAND4_in[1] ,
         \SB4_30/Component_Function_3/NAND4_in[3] ,
         \SB4_30/Component_Function_3/NAND4_in[2] ,
         \SB4_30/Component_Function_3/NAND4_in[1] ,
         \SB4_30/Component_Function_3/NAND4_in[0] ,
         \SB4_30/Component_Function_4/NAND4_in[3] ,
         \SB4_30/Component_Function_4/NAND4_in[2] ,
         \SB4_30/Component_Function_4/NAND4_in[1] ,
         \SB4_30/Component_Function_4/NAND4_in[0] ,
         \SB4_31/Component_Function_2/NAND4_in[3] ,
         \SB4_31/Component_Function_2/NAND4_in[2] ,
         \SB4_31/Component_Function_2/NAND4_in[1] ,
         \SB4_31/Component_Function_3/NAND4_in[3] ,
         \SB4_31/Component_Function_3/NAND4_in[2] ,
         \SB4_31/Component_Function_3/NAND4_in[1] ,
         \SB4_31/Component_Function_3/NAND4_in[0] ,
         \SB4_31/Component_Function_4/NAND4_in[2] ,
         \SB4_31/Component_Function_4/NAND4_in[1] ,
         \SB4_31/Component_Function_4/NAND4_in[0] ,
         \SB1_0_0/Component_Function_0/NAND4_in[3] ,
         \SB1_0_0/Component_Function_0/NAND4_in[2] ,
         \SB1_0_0/Component_Function_0/NAND4_in[1] ,
         \SB1_0_0/Component_Function_0/NAND4_in[0] ,
         \SB1_0_0/Component_Function_1/NAND4_in[3] ,
         \SB1_0_0/Component_Function_1/NAND4_in[2] ,
         \SB1_0_0/Component_Function_1/NAND4_in[1] ,
         \SB1_0_0/Component_Function_1/NAND4_in[0] ,
         \SB1_0_0/Component_Function_5/NAND4_in[3] ,
         \SB1_0_0/Component_Function_5/NAND4_in[2] ,
         \SB1_0_0/Component_Function_5/NAND4_in[1] ,
         \SB1_0_0/Component_Function_5/NAND4_in[0] ,
         \SB1_0_1/Component_Function_0/NAND4_in[3] ,
         \SB1_0_1/Component_Function_0/NAND4_in[2] ,
         \SB1_0_1/Component_Function_0/NAND4_in[1] ,
         \SB1_0_1/Component_Function_0/NAND4_in[0] ,
         \SB1_0_1/Component_Function_1/NAND4_in[3] ,
         \SB1_0_1/Component_Function_1/NAND4_in[1] ,
         \SB1_0_1/Component_Function_1/NAND4_in[0] ,
         \SB1_0_1/Component_Function_5/NAND4_in[3] ,
         \SB1_0_1/Component_Function_5/NAND4_in[2] ,
         \SB1_0_1/Component_Function_5/NAND4_in[1] ,
         \SB1_0_1/Component_Function_5/NAND4_in[0] ,
         \SB1_0_2/Component_Function_0/NAND4_in[3] ,
         \SB1_0_2/Component_Function_0/NAND4_in[2] ,
         \SB1_0_2/Component_Function_0/NAND4_in[1] ,
         \SB1_0_2/Component_Function_0/NAND4_in[0] ,
         \SB1_0_2/Component_Function_1/NAND4_in[3] ,
         \SB1_0_2/Component_Function_1/NAND4_in[2] ,
         \SB1_0_2/Component_Function_1/NAND4_in[1] ,
         \SB1_0_2/Component_Function_1/NAND4_in[0] ,
         \SB1_0_2/Component_Function_5/NAND4_in[3] ,
         \SB1_0_2/Component_Function_5/NAND4_in[1] ,
         \SB1_0_2/Component_Function_5/NAND4_in[0] ,
         \SB1_0_3/Component_Function_0/NAND4_in[3] ,
         \SB1_0_3/Component_Function_0/NAND4_in[2] ,
         \SB1_0_3/Component_Function_0/NAND4_in[1] ,
         \SB1_0_3/Component_Function_0/NAND4_in[0] ,
         \SB1_0_3/Component_Function_1/NAND4_in[3] ,
         \SB1_0_3/Component_Function_1/NAND4_in[2] ,
         \SB1_0_3/Component_Function_1/NAND4_in[1] ,
         \SB1_0_3/Component_Function_1/NAND4_in[0] ,
         \SB1_0_3/Component_Function_5/NAND4_in[3] ,
         \SB1_0_3/Component_Function_5/NAND4_in[2] ,
         \SB1_0_3/Component_Function_5/NAND4_in[1] ,
         \SB1_0_3/Component_Function_5/NAND4_in[0] ,
         \SB1_0_4/Component_Function_0/NAND4_in[3] ,
         \SB1_0_4/Component_Function_0/NAND4_in[2] ,
         \SB1_0_4/Component_Function_0/NAND4_in[1] ,
         \SB1_0_4/Component_Function_0/NAND4_in[0] ,
         \SB1_0_4/Component_Function_1/NAND4_in[3] ,
         \SB1_0_4/Component_Function_1/NAND4_in[2] ,
         \SB1_0_4/Component_Function_1/NAND4_in[1] ,
         \SB1_0_4/Component_Function_1/NAND4_in[0] ,
         \SB1_0_4/Component_Function_5/NAND4_in[3] ,
         \SB1_0_4/Component_Function_5/NAND4_in[2] ,
         \SB1_0_4/Component_Function_5/NAND4_in[1] ,
         \SB1_0_4/Component_Function_5/NAND4_in[0] ,
         \SB1_0_5/Component_Function_0/NAND4_in[3] ,
         \SB1_0_5/Component_Function_0/NAND4_in[2] ,
         \SB1_0_5/Component_Function_0/NAND4_in[1] ,
         \SB1_0_5/Component_Function_0/NAND4_in[0] ,
         \SB1_0_5/Component_Function_1/NAND4_in[3] ,
         \SB1_0_5/Component_Function_1/NAND4_in[2] ,
         \SB1_0_5/Component_Function_1/NAND4_in[1] ,
         \SB1_0_5/Component_Function_1/NAND4_in[0] ,
         \SB1_0_5/Component_Function_5/NAND4_in[3] ,
         \SB1_0_5/Component_Function_5/NAND4_in[1] ,
         \SB1_0_5/Component_Function_5/NAND4_in[0] ,
         \SB1_0_6/Component_Function_0/NAND4_in[3] ,
         \SB1_0_6/Component_Function_0/NAND4_in[2] ,
         \SB1_0_6/Component_Function_0/NAND4_in[1] ,
         \SB1_0_6/Component_Function_0/NAND4_in[0] ,
         \SB1_0_6/Component_Function_1/NAND4_in[3] ,
         \SB1_0_6/Component_Function_1/NAND4_in[2] ,
         \SB1_0_6/Component_Function_1/NAND4_in[1] ,
         \SB1_0_6/Component_Function_1/NAND4_in[0] ,
         \SB1_0_6/Component_Function_5/NAND4_in[3] ,
         \SB1_0_6/Component_Function_5/NAND4_in[1] ,
         \SB1_0_6/Component_Function_5/NAND4_in[0] ,
         \SB1_0_7/Component_Function_0/NAND4_in[3] ,
         \SB1_0_7/Component_Function_0/NAND4_in[2] ,
         \SB1_0_7/Component_Function_0/NAND4_in[1] ,
         \SB1_0_7/Component_Function_0/NAND4_in[0] ,
         \SB1_0_7/Component_Function_1/NAND4_in[3] ,
         \SB1_0_7/Component_Function_1/NAND4_in[2] ,
         \SB1_0_7/Component_Function_1/NAND4_in[1] ,
         \SB1_0_7/Component_Function_1/NAND4_in[0] ,
         \SB1_0_7/Component_Function_5/NAND4_in[3] ,
         \SB1_0_7/Component_Function_5/NAND4_in[2] ,
         \SB1_0_7/Component_Function_5/NAND4_in[1] ,
         \SB1_0_7/Component_Function_5/NAND4_in[0] ,
         \SB1_0_8/Component_Function_0/NAND4_in[3] ,
         \SB1_0_8/Component_Function_0/NAND4_in[2] ,
         \SB1_0_8/Component_Function_0/NAND4_in[1] ,
         \SB1_0_8/Component_Function_0/NAND4_in[0] ,
         \SB1_0_8/Component_Function_1/NAND4_in[3] ,
         \SB1_0_8/Component_Function_1/NAND4_in[2] ,
         \SB1_0_8/Component_Function_1/NAND4_in[1] ,
         \SB1_0_8/Component_Function_1/NAND4_in[0] ,
         \SB1_0_8/Component_Function_5/NAND4_in[3] ,
         \SB1_0_8/Component_Function_5/NAND4_in[1] ,
         \SB1_0_8/Component_Function_5/NAND4_in[0] ,
         \SB1_0_9/Component_Function_0/NAND4_in[3] ,
         \SB1_0_9/Component_Function_0/NAND4_in[2] ,
         \SB1_0_9/Component_Function_0/NAND4_in[1] ,
         \SB1_0_9/Component_Function_0/NAND4_in[0] ,
         \SB1_0_9/Component_Function_1/NAND4_in[3] ,
         \SB1_0_9/Component_Function_1/NAND4_in[2] ,
         \SB1_0_9/Component_Function_1/NAND4_in[1] ,
         \SB1_0_9/Component_Function_1/NAND4_in[0] ,
         \SB1_0_9/Component_Function_5/NAND4_in[3] ,
         \SB1_0_9/Component_Function_5/NAND4_in[2] ,
         \SB1_0_9/Component_Function_5/NAND4_in[1] ,
         \SB1_0_9/Component_Function_5/NAND4_in[0] ,
         \SB1_0_10/Component_Function_0/NAND4_in[3] ,
         \SB1_0_10/Component_Function_0/NAND4_in[2] ,
         \SB1_0_10/Component_Function_0/NAND4_in[1] ,
         \SB1_0_10/Component_Function_0/NAND4_in[0] ,
         \SB1_0_10/Component_Function_1/NAND4_in[3] ,
         \SB1_0_10/Component_Function_1/NAND4_in[2] ,
         \SB1_0_10/Component_Function_1/NAND4_in[1] ,
         \SB1_0_10/Component_Function_1/NAND4_in[0] ,
         \SB1_0_10/Component_Function_5/NAND4_in[3] ,
         \SB1_0_10/Component_Function_5/NAND4_in[2] ,
         \SB1_0_10/Component_Function_5/NAND4_in[1] ,
         \SB1_0_10/Component_Function_5/NAND4_in[0] ,
         \SB1_0_11/Component_Function_0/NAND4_in[3] ,
         \SB1_0_11/Component_Function_0/NAND4_in[2] ,
         \SB1_0_11/Component_Function_0/NAND4_in[1] ,
         \SB1_0_11/Component_Function_0/NAND4_in[0] ,
         \SB1_0_11/Component_Function_1/NAND4_in[3] ,
         \SB1_0_11/Component_Function_1/NAND4_in[2] ,
         \SB1_0_11/Component_Function_1/NAND4_in[1] ,
         \SB1_0_11/Component_Function_1/NAND4_in[0] ,
         \SB1_0_11/Component_Function_5/NAND4_in[3] ,
         \SB1_0_11/Component_Function_5/NAND4_in[1] ,
         \SB1_0_11/Component_Function_5/NAND4_in[0] ,
         \SB1_0_12/Component_Function_0/NAND4_in[3] ,
         \SB1_0_12/Component_Function_0/NAND4_in[2] ,
         \SB1_0_12/Component_Function_0/NAND4_in[1] ,
         \SB1_0_12/Component_Function_0/NAND4_in[0] ,
         \SB1_0_12/Component_Function_1/NAND4_in[3] ,
         \SB1_0_12/Component_Function_1/NAND4_in[2] ,
         \SB1_0_12/Component_Function_1/NAND4_in[1] ,
         \SB1_0_12/Component_Function_1/NAND4_in[0] ,
         \SB1_0_12/Component_Function_5/NAND4_in[3] ,
         \SB1_0_12/Component_Function_5/NAND4_in[2] ,
         \SB1_0_12/Component_Function_5/NAND4_in[1] ,
         \SB1_0_12/Component_Function_5/NAND4_in[0] ,
         \SB1_0_13/Component_Function_0/NAND4_in[3] ,
         \SB1_0_13/Component_Function_0/NAND4_in[2] ,
         \SB1_0_13/Component_Function_0/NAND4_in[1] ,
         \SB1_0_13/Component_Function_0/NAND4_in[0] ,
         \SB1_0_13/Component_Function_1/NAND4_in[3] ,
         \SB1_0_13/Component_Function_1/NAND4_in[2] ,
         \SB1_0_13/Component_Function_1/NAND4_in[1] ,
         \SB1_0_13/Component_Function_1/NAND4_in[0] ,
         \SB1_0_13/Component_Function_5/NAND4_in[3] ,
         \SB1_0_13/Component_Function_5/NAND4_in[2] ,
         \SB1_0_13/Component_Function_5/NAND4_in[1] ,
         \SB1_0_13/Component_Function_5/NAND4_in[0] ,
         \SB1_0_14/Component_Function_0/NAND4_in[3] ,
         \SB1_0_14/Component_Function_0/NAND4_in[2] ,
         \SB1_0_14/Component_Function_0/NAND4_in[1] ,
         \SB1_0_14/Component_Function_0/NAND4_in[0] ,
         \SB1_0_14/Component_Function_1/NAND4_in[3] ,
         \SB1_0_14/Component_Function_1/NAND4_in[2] ,
         \SB1_0_14/Component_Function_1/NAND4_in[1] ,
         \SB1_0_14/Component_Function_1/NAND4_in[0] ,
         \SB1_0_14/Component_Function_5/NAND4_in[3] ,
         \SB1_0_14/Component_Function_5/NAND4_in[2] ,
         \SB1_0_14/Component_Function_5/NAND4_in[1] ,
         \SB1_0_14/Component_Function_5/NAND4_in[0] ,
         \SB1_0_15/Component_Function_0/NAND4_in[3] ,
         \SB1_0_15/Component_Function_0/NAND4_in[2] ,
         \SB1_0_15/Component_Function_0/NAND4_in[1] ,
         \SB1_0_15/Component_Function_0/NAND4_in[0] ,
         \SB1_0_15/Component_Function_1/NAND4_in[3] ,
         \SB1_0_15/Component_Function_1/NAND4_in[2] ,
         \SB1_0_15/Component_Function_1/NAND4_in[1] ,
         \SB1_0_15/Component_Function_1/NAND4_in[0] ,
         \SB1_0_15/Component_Function_5/NAND4_in[3] ,
         \SB1_0_15/Component_Function_5/NAND4_in[1] ,
         \SB1_0_15/Component_Function_5/NAND4_in[0] ,
         \SB1_0_16/Component_Function_0/NAND4_in[3] ,
         \SB1_0_16/Component_Function_0/NAND4_in[2] ,
         \SB1_0_16/Component_Function_0/NAND4_in[1] ,
         \SB1_0_16/Component_Function_0/NAND4_in[0] ,
         \SB1_0_16/Component_Function_1/NAND4_in[3] ,
         \SB1_0_16/Component_Function_1/NAND4_in[2] ,
         \SB1_0_16/Component_Function_1/NAND4_in[1] ,
         \SB1_0_16/Component_Function_1/NAND4_in[0] ,
         \SB1_0_16/Component_Function_5/NAND4_in[3] ,
         \SB1_0_16/Component_Function_5/NAND4_in[1] ,
         \SB1_0_16/Component_Function_5/NAND4_in[0] ,
         \SB1_0_17/Component_Function_0/NAND4_in[3] ,
         \SB1_0_17/Component_Function_0/NAND4_in[2] ,
         \SB1_0_17/Component_Function_0/NAND4_in[1] ,
         \SB1_0_17/Component_Function_0/NAND4_in[0] ,
         \SB1_0_17/Component_Function_1/NAND4_in[3] ,
         \SB1_0_17/Component_Function_1/NAND4_in[2] ,
         \SB1_0_17/Component_Function_1/NAND4_in[1] ,
         \SB1_0_17/Component_Function_1/NAND4_in[0] ,
         \SB1_0_17/Component_Function_5/NAND4_in[3] ,
         \SB1_0_17/Component_Function_5/NAND4_in[2] ,
         \SB1_0_17/Component_Function_5/NAND4_in[1] ,
         \SB1_0_17/Component_Function_5/NAND4_in[0] ,
         \SB1_0_18/Component_Function_0/NAND4_in[3] ,
         \SB1_0_18/Component_Function_0/NAND4_in[1] ,
         \SB1_0_18/Component_Function_0/NAND4_in[0] ,
         \SB1_0_18/Component_Function_1/NAND4_in[3] ,
         \SB1_0_18/Component_Function_1/NAND4_in[2] ,
         \SB1_0_18/Component_Function_1/NAND4_in[1] ,
         \SB1_0_18/Component_Function_1/NAND4_in[0] ,
         \SB1_0_18/Component_Function_5/NAND4_in[3] ,
         \SB1_0_18/Component_Function_5/NAND4_in[1] ,
         \SB1_0_18/Component_Function_5/NAND4_in[0] ,
         \SB1_0_19/Component_Function_0/NAND4_in[3] ,
         \SB1_0_19/Component_Function_0/NAND4_in[2] ,
         \SB1_0_19/Component_Function_0/NAND4_in[1] ,
         \SB1_0_19/Component_Function_0/NAND4_in[0] ,
         \SB1_0_19/Component_Function_1/NAND4_in[3] ,
         \SB1_0_19/Component_Function_1/NAND4_in[1] ,
         \SB1_0_19/Component_Function_1/NAND4_in[0] ,
         \SB1_0_19/Component_Function_5/NAND4_in[3] ,
         \SB1_0_19/Component_Function_5/NAND4_in[2] ,
         \SB1_0_19/Component_Function_5/NAND4_in[1] ,
         \SB1_0_19/Component_Function_5/NAND4_in[0] ,
         \SB1_0_20/Component_Function_0/NAND4_in[3] ,
         \SB1_0_20/Component_Function_0/NAND4_in[2] ,
         \SB1_0_20/Component_Function_0/NAND4_in[1] ,
         \SB1_0_20/Component_Function_0/NAND4_in[0] ,
         \SB1_0_20/Component_Function_1/NAND4_in[3] ,
         \SB1_0_20/Component_Function_1/NAND4_in[2] ,
         \SB1_0_20/Component_Function_1/NAND4_in[1] ,
         \SB1_0_20/Component_Function_1/NAND4_in[0] ,
         \SB1_0_20/Component_Function_5/NAND4_in[3] ,
         \SB1_0_20/Component_Function_5/NAND4_in[1] ,
         \SB1_0_20/Component_Function_5/NAND4_in[0] ,
         \SB1_0_21/Component_Function_0/NAND4_in[3] ,
         \SB1_0_21/Component_Function_0/NAND4_in[2] ,
         \SB1_0_21/Component_Function_0/NAND4_in[1] ,
         \SB1_0_21/Component_Function_0/NAND4_in[0] ,
         \SB1_0_21/Component_Function_1/NAND4_in[3] ,
         \SB1_0_21/Component_Function_1/NAND4_in[2] ,
         \SB1_0_21/Component_Function_1/NAND4_in[1] ,
         \SB1_0_21/Component_Function_1/NAND4_in[0] ,
         \SB1_0_21/Component_Function_5/NAND4_in[3] ,
         \SB1_0_21/Component_Function_5/NAND4_in[1] ,
         \SB1_0_21/Component_Function_5/NAND4_in[0] ,
         \SB1_0_22/Component_Function_0/NAND4_in[3] ,
         \SB1_0_22/Component_Function_0/NAND4_in[2] ,
         \SB1_0_22/Component_Function_0/NAND4_in[1] ,
         \SB1_0_22/Component_Function_0/NAND4_in[0] ,
         \SB1_0_22/Component_Function_1/NAND4_in[2] ,
         \SB1_0_22/Component_Function_1/NAND4_in[1] ,
         \SB1_0_22/Component_Function_1/NAND4_in[0] ,
         \SB1_0_22/Component_Function_5/NAND4_in[3] ,
         \SB1_0_22/Component_Function_5/NAND4_in[2] ,
         \SB1_0_22/Component_Function_5/NAND4_in[1] ,
         \SB1_0_22/Component_Function_5/NAND4_in[0] ,
         \SB1_0_23/Component_Function_0/NAND4_in[3] ,
         \SB1_0_23/Component_Function_0/NAND4_in[2] ,
         \SB1_0_23/Component_Function_0/NAND4_in[1] ,
         \SB1_0_23/Component_Function_0/NAND4_in[0] ,
         \SB1_0_23/Component_Function_1/NAND4_in[3] ,
         \SB1_0_23/Component_Function_1/NAND4_in[2] ,
         \SB1_0_23/Component_Function_1/NAND4_in[1] ,
         \SB1_0_23/Component_Function_1/NAND4_in[0] ,
         \SB1_0_23/Component_Function_5/NAND4_in[3] ,
         \SB1_0_23/Component_Function_5/NAND4_in[1] ,
         \SB1_0_24/Component_Function_0/NAND4_in[3] ,
         \SB1_0_24/Component_Function_0/NAND4_in[2] ,
         \SB1_0_24/Component_Function_0/NAND4_in[1] ,
         \SB1_0_24/Component_Function_0/NAND4_in[0] ,
         \SB1_0_24/Component_Function_1/NAND4_in[3] ,
         \SB1_0_24/Component_Function_1/NAND4_in[2] ,
         \SB1_0_24/Component_Function_1/NAND4_in[1] ,
         \SB1_0_24/Component_Function_1/NAND4_in[0] ,
         \SB1_0_24/Component_Function_5/NAND4_in[3] ,
         \SB1_0_24/Component_Function_5/NAND4_in[2] ,
         \SB1_0_24/Component_Function_5/NAND4_in[1] ,
         \SB1_0_24/Component_Function_5/NAND4_in[0] ,
         \SB1_0_25/Component_Function_0/NAND4_in[2] ,
         \SB1_0_25/Component_Function_0/NAND4_in[1] ,
         \SB1_0_25/Component_Function_0/NAND4_in[0] ,
         \SB1_0_25/Component_Function_1/NAND4_in[3] ,
         \SB1_0_25/Component_Function_1/NAND4_in[2] ,
         \SB1_0_25/Component_Function_1/NAND4_in[1] ,
         \SB1_0_25/Component_Function_1/NAND4_in[0] ,
         \SB1_0_25/Component_Function_5/NAND4_in[3] ,
         \SB1_0_25/Component_Function_5/NAND4_in[1] ,
         \SB1_0_25/Component_Function_5/NAND4_in[0] ,
         \SB1_0_26/Component_Function_0/NAND4_in[3] ,
         \SB1_0_26/Component_Function_0/NAND4_in[2] ,
         \SB1_0_26/Component_Function_0/NAND4_in[1] ,
         \SB1_0_26/Component_Function_0/NAND4_in[0] ,
         \SB1_0_26/Component_Function_1/NAND4_in[3] ,
         \SB1_0_26/Component_Function_1/NAND4_in[2] ,
         \SB1_0_26/Component_Function_1/NAND4_in[1] ,
         \SB1_0_26/Component_Function_1/NAND4_in[0] ,
         \SB1_0_26/Component_Function_5/NAND4_in[3] ,
         \SB1_0_26/Component_Function_5/NAND4_in[1] ,
         \SB1_0_26/Component_Function_5/NAND4_in[0] ,
         \SB1_0_27/Component_Function_0/NAND4_in[3] ,
         \SB1_0_27/Component_Function_0/NAND4_in[2] ,
         \SB1_0_27/Component_Function_0/NAND4_in[1] ,
         \SB1_0_27/Component_Function_0/NAND4_in[0] ,
         \SB1_0_27/Component_Function_1/NAND4_in[3] ,
         \SB1_0_27/Component_Function_1/NAND4_in[2] ,
         \SB1_0_27/Component_Function_1/NAND4_in[1] ,
         \SB1_0_27/Component_Function_1/NAND4_in[0] ,
         \SB1_0_27/Component_Function_5/NAND4_in[3] ,
         \SB1_0_27/Component_Function_5/NAND4_in[2] ,
         \SB1_0_27/Component_Function_5/NAND4_in[1] ,
         \SB1_0_27/Component_Function_5/NAND4_in[0] ,
         \SB1_0_28/Component_Function_0/NAND4_in[3] ,
         \SB1_0_28/Component_Function_0/NAND4_in[2] ,
         \SB1_0_28/Component_Function_0/NAND4_in[1] ,
         \SB1_0_28/Component_Function_0/NAND4_in[0] ,
         \SB1_0_28/Component_Function_1/NAND4_in[3] ,
         \SB1_0_28/Component_Function_1/NAND4_in[2] ,
         \SB1_0_28/Component_Function_1/NAND4_in[1] ,
         \SB1_0_28/Component_Function_1/NAND4_in[0] ,
         \SB1_0_28/Component_Function_5/NAND4_in[3] ,
         \SB1_0_28/Component_Function_5/NAND4_in[2] ,
         \SB1_0_28/Component_Function_5/NAND4_in[1] ,
         \SB1_0_28/Component_Function_5/NAND4_in[0] ,
         \SB1_0_29/Component_Function_0/NAND4_in[3] ,
         \SB1_0_29/Component_Function_0/NAND4_in[2] ,
         \SB1_0_29/Component_Function_0/NAND4_in[1] ,
         \SB1_0_29/Component_Function_0/NAND4_in[0] ,
         \SB1_0_29/Component_Function_1/NAND4_in[3] ,
         \SB1_0_29/Component_Function_1/NAND4_in[2] ,
         \SB1_0_29/Component_Function_1/NAND4_in[1] ,
         \SB1_0_29/Component_Function_1/NAND4_in[0] ,
         \SB1_0_29/Component_Function_5/NAND4_in[3] ,
         \SB1_0_29/Component_Function_5/NAND4_in[2] ,
         \SB1_0_29/Component_Function_5/NAND4_in[1] ,
         \SB1_0_29/Component_Function_5/NAND4_in[0] ,
         \SB1_0_30/Component_Function_0/NAND4_in[3] ,
         \SB1_0_30/Component_Function_0/NAND4_in[2] ,
         \SB1_0_30/Component_Function_0/NAND4_in[1] ,
         \SB1_0_30/Component_Function_0/NAND4_in[0] ,
         \SB1_0_30/Component_Function_1/NAND4_in[3] ,
         \SB1_0_30/Component_Function_1/NAND4_in[2] ,
         \SB1_0_30/Component_Function_1/NAND4_in[1] ,
         \SB1_0_30/Component_Function_1/NAND4_in[0] ,
         \SB1_0_30/Component_Function_5/NAND4_in[3] ,
         \SB1_0_30/Component_Function_5/NAND4_in[2] ,
         \SB1_0_30/Component_Function_5/NAND4_in[1] ,
         \SB1_0_30/Component_Function_5/NAND4_in[0] ,
         \SB1_0_31/Component_Function_0/NAND4_in[3] ,
         \SB1_0_31/Component_Function_0/NAND4_in[2] ,
         \SB1_0_31/Component_Function_0/NAND4_in[1] ,
         \SB1_0_31/Component_Function_0/NAND4_in[0] ,
         \SB1_0_31/Component_Function_1/NAND4_in[3] ,
         \SB1_0_31/Component_Function_1/NAND4_in[2] ,
         \SB1_0_31/Component_Function_1/NAND4_in[1] ,
         \SB1_0_31/Component_Function_1/NAND4_in[0] ,
         \SB1_0_31/Component_Function_5/NAND4_in[3] ,
         \SB1_0_31/Component_Function_5/NAND4_in[2] ,
         \SB1_0_31/Component_Function_5/NAND4_in[1] ,
         \SB1_0_31/Component_Function_5/NAND4_in[0] ,
         \SB2_0_0/Component_Function_0/NAND4_in[3] ,
         \SB2_0_0/Component_Function_0/NAND4_in[2] ,
         \SB2_0_0/Component_Function_0/NAND4_in[1] ,
         \SB2_0_0/Component_Function_0/NAND4_in[0] ,
         \SB2_0_0/Component_Function_1/NAND4_in[3] ,
         \SB2_0_0/Component_Function_1/NAND4_in[2] ,
         \SB2_0_0/Component_Function_1/NAND4_in[1] ,
         \SB2_0_0/Component_Function_1/NAND4_in[0] ,
         \SB2_0_0/Component_Function_5/NAND4_in[2] ,
         \SB2_0_0/Component_Function_5/NAND4_in[1] ,
         \SB2_0_0/Component_Function_5/NAND4_in[0] ,
         \SB2_0_1/Component_Function_0/NAND4_in[3] ,
         \SB2_0_1/Component_Function_0/NAND4_in[2] ,
         \SB2_0_1/Component_Function_0/NAND4_in[1] ,
         \SB2_0_1/Component_Function_0/NAND4_in[0] ,
         \SB2_0_1/Component_Function_1/NAND4_in[3] ,
         \SB2_0_1/Component_Function_1/NAND4_in[2] ,
         \SB2_0_1/Component_Function_1/NAND4_in[1] ,
         \SB2_0_1/Component_Function_1/NAND4_in[0] ,
         \SB2_0_1/Component_Function_5/NAND4_in[3] ,
         \SB2_0_1/Component_Function_5/NAND4_in[1] ,
         \SB2_0_1/Component_Function_5/NAND4_in[0] ,
         \SB2_0_2/Component_Function_0/NAND4_in[3] ,
         \SB2_0_2/Component_Function_0/NAND4_in[2] ,
         \SB2_0_2/Component_Function_0/NAND4_in[1] ,
         \SB2_0_2/Component_Function_0/NAND4_in[0] ,
         \SB2_0_2/Component_Function_1/NAND4_in[3] ,
         \SB2_0_2/Component_Function_1/NAND4_in[2] ,
         \SB2_0_2/Component_Function_1/NAND4_in[1] ,
         \SB2_0_2/Component_Function_1/NAND4_in[0] ,
         \SB2_0_2/Component_Function_5/NAND4_in[3] ,
         \SB2_0_2/Component_Function_5/NAND4_in[2] ,
         \SB2_0_2/Component_Function_5/NAND4_in[1] ,
         \SB2_0_3/Component_Function_0/NAND4_in[3] ,
         \SB2_0_3/Component_Function_0/NAND4_in[2] ,
         \SB2_0_3/Component_Function_0/NAND4_in[1] ,
         \SB2_0_3/Component_Function_0/NAND4_in[0] ,
         \SB2_0_3/Component_Function_1/NAND4_in[3] ,
         \SB2_0_3/Component_Function_1/NAND4_in[2] ,
         \SB2_0_3/Component_Function_1/NAND4_in[1] ,
         \SB2_0_3/Component_Function_1/NAND4_in[0] ,
         \SB2_0_3/Component_Function_5/NAND4_in[3] ,
         \SB2_0_3/Component_Function_5/NAND4_in[2] ,
         \SB2_0_3/Component_Function_5/NAND4_in[1] ,
         \SB2_0_3/Component_Function_5/NAND4_in[0] ,
         \SB2_0_4/Component_Function_0/NAND4_in[3] ,
         \SB2_0_4/Component_Function_0/NAND4_in[2] ,
         \SB2_0_4/Component_Function_0/NAND4_in[1] ,
         \SB2_0_4/Component_Function_0/NAND4_in[0] ,
         \SB2_0_4/Component_Function_1/NAND4_in[3] ,
         \SB2_0_4/Component_Function_1/NAND4_in[2] ,
         \SB2_0_4/Component_Function_1/NAND4_in[1] ,
         \SB2_0_4/Component_Function_1/NAND4_in[0] ,
         \SB2_0_4/Component_Function_5/NAND4_in[3] ,
         \SB2_0_4/Component_Function_5/NAND4_in[2] ,
         \SB2_0_4/Component_Function_5/NAND4_in[1] ,
         \SB2_0_4/Component_Function_5/NAND4_in[0] ,
         \SB2_0_5/Component_Function_0/NAND4_in[3] ,
         \SB2_0_5/Component_Function_0/NAND4_in[2] ,
         \SB2_0_5/Component_Function_0/NAND4_in[1] ,
         \SB2_0_5/Component_Function_0/NAND4_in[0] ,
         \SB2_0_5/Component_Function_1/NAND4_in[3] ,
         \SB2_0_5/Component_Function_1/NAND4_in[2] ,
         \SB2_0_5/Component_Function_1/NAND4_in[1] ,
         \SB2_0_5/Component_Function_1/NAND4_in[0] ,
         \SB2_0_5/Component_Function_5/NAND4_in[3] ,
         \SB2_0_5/Component_Function_5/NAND4_in[2] ,
         \SB2_0_5/Component_Function_5/NAND4_in[1] ,
         \SB2_0_5/Component_Function_5/NAND4_in[0] ,
         \SB2_0_6/Component_Function_0/NAND4_in[3] ,
         \SB2_0_6/Component_Function_0/NAND4_in[2] ,
         \SB2_0_6/Component_Function_0/NAND4_in[1] ,
         \SB2_0_6/Component_Function_0/NAND4_in[0] ,
         \SB2_0_6/Component_Function_1/NAND4_in[3] ,
         \SB2_0_6/Component_Function_1/NAND4_in[2] ,
         \SB2_0_6/Component_Function_1/NAND4_in[1] ,
         \SB2_0_6/Component_Function_1/NAND4_in[0] ,
         \SB2_0_6/Component_Function_5/NAND4_in[3] ,
         \SB2_0_6/Component_Function_5/NAND4_in[1] ,
         \SB2_0_6/Component_Function_5/NAND4_in[0] ,
         \SB2_0_7/Component_Function_0/NAND4_in[3] ,
         \SB2_0_7/Component_Function_0/NAND4_in[2] ,
         \SB2_0_7/Component_Function_0/NAND4_in[1] ,
         \SB2_0_7/Component_Function_0/NAND4_in[0] ,
         \SB2_0_7/Component_Function_1/NAND4_in[3] ,
         \SB2_0_7/Component_Function_1/NAND4_in[2] ,
         \SB2_0_7/Component_Function_1/NAND4_in[1] ,
         \SB2_0_7/Component_Function_1/NAND4_in[0] ,
         \SB2_0_7/Component_Function_5/NAND4_in[3] ,
         \SB2_0_7/Component_Function_5/NAND4_in[2] ,
         \SB2_0_7/Component_Function_5/NAND4_in[1] ,
         \SB2_0_8/Component_Function_0/NAND4_in[3] ,
         \SB2_0_8/Component_Function_0/NAND4_in[2] ,
         \SB2_0_8/Component_Function_0/NAND4_in[1] ,
         \SB2_0_8/Component_Function_0/NAND4_in[0] ,
         \SB2_0_8/Component_Function_1/NAND4_in[3] ,
         \SB2_0_8/Component_Function_1/NAND4_in[2] ,
         \SB2_0_8/Component_Function_1/NAND4_in[1] ,
         \SB2_0_8/Component_Function_1/NAND4_in[0] ,
         \SB2_0_8/Component_Function_5/NAND4_in[3] ,
         \SB2_0_8/Component_Function_5/NAND4_in[1] ,
         \SB2_0_8/Component_Function_5/NAND4_in[0] ,
         \SB2_0_9/Component_Function_0/NAND4_in[3] ,
         \SB2_0_9/Component_Function_0/NAND4_in[2] ,
         \SB2_0_9/Component_Function_0/NAND4_in[1] ,
         \SB2_0_9/Component_Function_0/NAND4_in[0] ,
         \SB2_0_9/Component_Function_1/NAND4_in[3] ,
         \SB2_0_9/Component_Function_1/NAND4_in[2] ,
         \SB2_0_9/Component_Function_1/NAND4_in[1] ,
         \SB2_0_9/Component_Function_1/NAND4_in[0] ,
         \SB2_0_9/Component_Function_5/NAND4_in[3] ,
         \SB2_0_9/Component_Function_5/NAND4_in[1] ,
         \SB2_0_9/Component_Function_5/NAND4_in[0] ,
         \SB2_0_10/Component_Function_0/NAND4_in[3] ,
         \SB2_0_10/Component_Function_0/NAND4_in[2] ,
         \SB2_0_10/Component_Function_0/NAND4_in[1] ,
         \SB2_0_10/Component_Function_0/NAND4_in[0] ,
         \SB2_0_10/Component_Function_1/NAND4_in[3] ,
         \SB2_0_10/Component_Function_1/NAND4_in[2] ,
         \SB2_0_10/Component_Function_1/NAND4_in[1] ,
         \SB2_0_10/Component_Function_1/NAND4_in[0] ,
         \SB2_0_10/Component_Function_5/NAND4_in[3] ,
         \SB2_0_10/Component_Function_5/NAND4_in[2] ,
         \SB2_0_10/Component_Function_5/NAND4_in[1] ,
         \SB2_0_11/Component_Function_0/NAND4_in[3] ,
         \SB2_0_11/Component_Function_0/NAND4_in[2] ,
         \SB2_0_11/Component_Function_0/NAND4_in[1] ,
         \SB2_0_11/Component_Function_0/NAND4_in[0] ,
         \SB2_0_11/Component_Function_1/NAND4_in[3] ,
         \SB2_0_11/Component_Function_1/NAND4_in[2] ,
         \SB2_0_11/Component_Function_1/NAND4_in[1] ,
         \SB2_0_11/Component_Function_1/NAND4_in[0] ,
         \SB2_0_11/Component_Function_5/NAND4_in[3] ,
         \SB2_0_11/Component_Function_5/NAND4_in[2] ,
         \SB2_0_11/Component_Function_5/NAND4_in[1] ,
         \SB2_0_11/Component_Function_5/NAND4_in[0] ,
         \SB2_0_12/Component_Function_0/NAND4_in[3] ,
         \SB2_0_12/Component_Function_0/NAND4_in[2] ,
         \SB2_0_12/Component_Function_0/NAND4_in[1] ,
         \SB2_0_12/Component_Function_0/NAND4_in[0] ,
         \SB2_0_12/Component_Function_1/NAND4_in[3] ,
         \SB2_0_12/Component_Function_1/NAND4_in[2] ,
         \SB2_0_12/Component_Function_1/NAND4_in[1] ,
         \SB2_0_12/Component_Function_1/NAND4_in[0] ,
         \SB2_0_12/Component_Function_5/NAND4_in[3] ,
         \SB2_0_12/Component_Function_5/NAND4_in[2] ,
         \SB2_0_12/Component_Function_5/NAND4_in[1] ,
         \SB2_0_12/Component_Function_5/NAND4_in[0] ,
         \SB2_0_13/Component_Function_0/NAND4_in[3] ,
         \SB2_0_13/Component_Function_0/NAND4_in[2] ,
         \SB2_0_13/Component_Function_0/NAND4_in[1] ,
         \SB2_0_13/Component_Function_0/NAND4_in[0] ,
         \SB2_0_13/Component_Function_1/NAND4_in[3] ,
         \SB2_0_13/Component_Function_1/NAND4_in[2] ,
         \SB2_0_13/Component_Function_1/NAND4_in[1] ,
         \SB2_0_13/Component_Function_1/NAND4_in[0] ,
         \SB2_0_13/Component_Function_5/NAND4_in[3] ,
         \SB2_0_13/Component_Function_5/NAND4_in[1] ,
         \SB2_0_13/Component_Function_5/NAND4_in[0] ,
         \SB2_0_14/Component_Function_0/NAND4_in[3] ,
         \SB2_0_14/Component_Function_0/NAND4_in[2] ,
         \SB2_0_14/Component_Function_0/NAND4_in[1] ,
         \SB2_0_14/Component_Function_0/NAND4_in[0] ,
         \SB2_0_14/Component_Function_1/NAND4_in[3] ,
         \SB2_0_14/Component_Function_1/NAND4_in[2] ,
         \SB2_0_14/Component_Function_1/NAND4_in[1] ,
         \SB2_0_14/Component_Function_1/NAND4_in[0] ,
         \SB2_0_14/Component_Function_5/NAND4_in[3] ,
         \SB2_0_14/Component_Function_5/NAND4_in[2] ,
         \SB2_0_14/Component_Function_5/NAND4_in[1] ,
         \SB2_0_14/Component_Function_5/NAND4_in[0] ,
         \SB2_0_15/Component_Function_0/NAND4_in[3] ,
         \SB2_0_15/Component_Function_0/NAND4_in[2] ,
         \SB2_0_15/Component_Function_0/NAND4_in[1] ,
         \SB2_0_15/Component_Function_0/NAND4_in[0] ,
         \SB2_0_15/Component_Function_1/NAND4_in[3] ,
         \SB2_0_15/Component_Function_1/NAND4_in[2] ,
         \SB2_0_15/Component_Function_1/NAND4_in[1] ,
         \SB2_0_15/Component_Function_1/NAND4_in[0] ,
         \SB2_0_15/Component_Function_5/NAND4_in[3] ,
         \SB2_0_15/Component_Function_5/NAND4_in[2] ,
         \SB2_0_15/Component_Function_5/NAND4_in[1] ,
         \SB2_0_15/Component_Function_5/NAND4_in[0] ,
         \SB2_0_16/Component_Function_0/NAND4_in[3] ,
         \SB2_0_16/Component_Function_0/NAND4_in[2] ,
         \SB2_0_16/Component_Function_0/NAND4_in[1] ,
         \SB2_0_16/Component_Function_0/NAND4_in[0] ,
         \SB2_0_16/Component_Function_1/NAND4_in[3] ,
         \SB2_0_16/Component_Function_1/NAND4_in[2] ,
         \SB2_0_16/Component_Function_1/NAND4_in[1] ,
         \SB2_0_16/Component_Function_1/NAND4_in[0] ,
         \SB2_0_16/Component_Function_5/NAND4_in[3] ,
         \SB2_0_16/Component_Function_5/NAND4_in[2] ,
         \SB2_0_16/Component_Function_5/NAND4_in[1] ,
         \SB2_0_16/Component_Function_5/NAND4_in[0] ,
         \SB2_0_17/Component_Function_0/NAND4_in[3] ,
         \SB2_0_17/Component_Function_0/NAND4_in[2] ,
         \SB2_0_17/Component_Function_0/NAND4_in[1] ,
         \SB2_0_17/Component_Function_0/NAND4_in[0] ,
         \SB2_0_17/Component_Function_1/NAND4_in[3] ,
         \SB2_0_17/Component_Function_1/NAND4_in[2] ,
         \SB2_0_17/Component_Function_1/NAND4_in[1] ,
         \SB2_0_17/Component_Function_1/NAND4_in[0] ,
         \SB2_0_17/Component_Function_5/NAND4_in[2] ,
         \SB2_0_17/Component_Function_5/NAND4_in[1] ,
         \SB2_0_17/Component_Function_5/NAND4_in[0] ,
         \SB2_0_18/Component_Function_0/NAND4_in[3] ,
         \SB2_0_18/Component_Function_0/NAND4_in[2] ,
         \SB2_0_18/Component_Function_0/NAND4_in[1] ,
         \SB2_0_18/Component_Function_0/NAND4_in[0] ,
         \SB2_0_18/Component_Function_1/NAND4_in[3] ,
         \SB2_0_18/Component_Function_1/NAND4_in[2] ,
         \SB2_0_18/Component_Function_1/NAND4_in[1] ,
         \SB2_0_18/Component_Function_1/NAND4_in[0] ,
         \SB2_0_18/Component_Function_5/NAND4_in[3] ,
         \SB2_0_18/Component_Function_5/NAND4_in[2] ,
         \SB2_0_18/Component_Function_5/NAND4_in[1] ,
         \SB2_0_18/Component_Function_5/NAND4_in[0] ,
         \SB2_0_19/Component_Function_0/NAND4_in[3] ,
         \SB2_0_19/Component_Function_0/NAND4_in[2] ,
         \SB2_0_19/Component_Function_0/NAND4_in[1] ,
         \SB2_0_19/Component_Function_0/NAND4_in[0] ,
         \SB2_0_19/Component_Function_1/NAND4_in[3] ,
         \SB2_0_19/Component_Function_1/NAND4_in[2] ,
         \SB2_0_19/Component_Function_1/NAND4_in[1] ,
         \SB2_0_19/Component_Function_1/NAND4_in[0] ,
         \SB2_0_19/Component_Function_5/NAND4_in[3] ,
         \SB2_0_19/Component_Function_5/NAND4_in[2] ,
         \SB2_0_19/Component_Function_5/NAND4_in[1] ,
         \SB2_0_19/Component_Function_5/NAND4_in[0] ,
         \SB2_0_20/Component_Function_0/NAND4_in[3] ,
         \SB2_0_20/Component_Function_0/NAND4_in[2] ,
         \SB2_0_20/Component_Function_0/NAND4_in[1] ,
         \SB2_0_20/Component_Function_0/NAND4_in[0] ,
         \SB2_0_20/Component_Function_1/NAND4_in[3] ,
         \SB2_0_20/Component_Function_1/NAND4_in[2] ,
         \SB2_0_20/Component_Function_1/NAND4_in[1] ,
         \SB2_0_20/Component_Function_1/NAND4_in[0] ,
         \SB2_0_20/Component_Function_5/NAND4_in[1] ,
         \SB2_0_21/Component_Function_0/NAND4_in[3] ,
         \SB2_0_21/Component_Function_0/NAND4_in[2] ,
         \SB2_0_21/Component_Function_0/NAND4_in[1] ,
         \SB2_0_21/Component_Function_0/NAND4_in[0] ,
         \SB2_0_21/Component_Function_1/NAND4_in[3] ,
         \SB2_0_21/Component_Function_1/NAND4_in[2] ,
         \SB2_0_21/Component_Function_1/NAND4_in[1] ,
         \SB2_0_21/Component_Function_1/NAND4_in[0] ,
         \SB2_0_21/Component_Function_5/NAND4_in[3] ,
         \SB2_0_21/Component_Function_5/NAND4_in[2] ,
         \SB2_0_21/Component_Function_5/NAND4_in[1] ,
         \SB2_0_21/Component_Function_5/NAND4_in[0] ,
         \SB2_0_22/Component_Function_0/NAND4_in[3] ,
         \SB2_0_22/Component_Function_0/NAND4_in[2] ,
         \SB2_0_22/Component_Function_0/NAND4_in[1] ,
         \SB2_0_22/Component_Function_0/NAND4_in[0] ,
         \SB2_0_22/Component_Function_1/NAND4_in[3] ,
         \SB2_0_22/Component_Function_1/NAND4_in[2] ,
         \SB2_0_22/Component_Function_1/NAND4_in[1] ,
         \SB2_0_22/Component_Function_1/NAND4_in[0] ,
         \SB2_0_22/Component_Function_5/NAND4_in[3] ,
         \SB2_0_22/Component_Function_5/NAND4_in[2] ,
         \SB2_0_22/Component_Function_5/NAND4_in[1] ,
         \SB2_0_22/Component_Function_5/NAND4_in[0] ,
         \SB2_0_23/Component_Function_0/NAND4_in[3] ,
         \SB2_0_23/Component_Function_0/NAND4_in[1] ,
         \SB2_0_23/Component_Function_0/NAND4_in[0] ,
         \SB2_0_23/Component_Function_1/NAND4_in[3] ,
         \SB2_0_23/Component_Function_1/NAND4_in[2] ,
         \SB2_0_23/Component_Function_1/NAND4_in[1] ,
         \SB2_0_23/Component_Function_1/NAND4_in[0] ,
         \SB2_0_23/Component_Function_5/NAND4_in[3] ,
         \SB2_0_23/Component_Function_5/NAND4_in[1] ,
         \SB2_0_23/Component_Function_5/NAND4_in[0] ,
         \SB2_0_24/Component_Function_0/NAND4_in[3] ,
         \SB2_0_24/Component_Function_0/NAND4_in[2] ,
         \SB2_0_24/Component_Function_0/NAND4_in[1] ,
         \SB2_0_24/Component_Function_0/NAND4_in[0] ,
         \SB2_0_24/Component_Function_1/NAND4_in[3] ,
         \SB2_0_24/Component_Function_1/NAND4_in[2] ,
         \SB2_0_24/Component_Function_1/NAND4_in[1] ,
         \SB2_0_24/Component_Function_1/NAND4_in[0] ,
         \SB2_0_24/Component_Function_5/NAND4_in[3] ,
         \SB2_0_24/Component_Function_5/NAND4_in[2] ,
         \SB2_0_24/Component_Function_5/NAND4_in[1] ,
         \SB2_0_24/Component_Function_5/NAND4_in[0] ,
         \SB2_0_25/Component_Function_0/NAND4_in[2] ,
         \SB2_0_25/Component_Function_0/NAND4_in[1] ,
         \SB2_0_25/Component_Function_0/NAND4_in[0] ,
         \SB2_0_25/Component_Function_1/NAND4_in[3] ,
         \SB2_0_25/Component_Function_1/NAND4_in[2] ,
         \SB2_0_25/Component_Function_1/NAND4_in[1] ,
         \SB2_0_25/Component_Function_1/NAND4_in[0] ,
         \SB2_0_25/Component_Function_5/NAND4_in[3] ,
         \SB2_0_25/Component_Function_5/NAND4_in[1] ,
         \SB2_0_25/Component_Function_5/NAND4_in[0] ,
         \SB2_0_26/Component_Function_0/NAND4_in[3] ,
         \SB2_0_26/Component_Function_0/NAND4_in[2] ,
         \SB2_0_26/Component_Function_0/NAND4_in[1] ,
         \SB2_0_26/Component_Function_0/NAND4_in[0] ,
         \SB2_0_26/Component_Function_1/NAND4_in[3] ,
         \SB2_0_26/Component_Function_1/NAND4_in[2] ,
         \SB2_0_26/Component_Function_1/NAND4_in[1] ,
         \SB2_0_26/Component_Function_1/NAND4_in[0] ,
         \SB2_0_26/Component_Function_5/NAND4_in[2] ,
         \SB2_0_26/Component_Function_5/NAND4_in[0] ,
         \SB2_0_27/Component_Function_0/NAND4_in[3] ,
         \SB2_0_27/Component_Function_0/NAND4_in[2] ,
         \SB2_0_27/Component_Function_0/NAND4_in[1] ,
         \SB2_0_27/Component_Function_0/NAND4_in[0] ,
         \SB2_0_27/Component_Function_1/NAND4_in[3] ,
         \SB2_0_27/Component_Function_1/NAND4_in[2] ,
         \SB2_0_27/Component_Function_1/NAND4_in[1] ,
         \SB2_0_27/Component_Function_1/NAND4_in[0] ,
         \SB2_0_27/Component_Function_5/NAND4_in[3] ,
         \SB2_0_27/Component_Function_5/NAND4_in[2] ,
         \SB2_0_27/Component_Function_5/NAND4_in[1] ,
         \SB2_0_27/Component_Function_5/NAND4_in[0] ,
         \SB2_0_28/Component_Function_0/NAND4_in[3] ,
         \SB2_0_28/Component_Function_0/NAND4_in[2] ,
         \SB2_0_28/Component_Function_0/NAND4_in[1] ,
         \SB2_0_28/Component_Function_0/NAND4_in[0] ,
         \SB2_0_28/Component_Function_1/NAND4_in[3] ,
         \SB2_0_28/Component_Function_1/NAND4_in[2] ,
         \SB2_0_28/Component_Function_1/NAND4_in[1] ,
         \SB2_0_28/Component_Function_1/NAND4_in[0] ,
         \SB2_0_28/Component_Function_5/NAND4_in[3] ,
         \SB2_0_28/Component_Function_5/NAND4_in[1] ,
         \SB2_0_28/Component_Function_5/NAND4_in[0] ,
         \SB2_0_29/Component_Function_0/NAND4_in[3] ,
         \SB2_0_29/Component_Function_0/NAND4_in[2] ,
         \SB2_0_29/Component_Function_0/NAND4_in[1] ,
         \SB2_0_29/Component_Function_0/NAND4_in[0] ,
         \SB2_0_29/Component_Function_1/NAND4_in[3] ,
         \SB2_0_29/Component_Function_1/NAND4_in[2] ,
         \SB2_0_29/Component_Function_1/NAND4_in[1] ,
         \SB2_0_29/Component_Function_1/NAND4_in[0] ,
         \SB2_0_29/Component_Function_5/NAND4_in[3] ,
         \SB2_0_29/Component_Function_5/NAND4_in[2] ,
         \SB2_0_29/Component_Function_5/NAND4_in[1] ,
         \SB2_0_30/Component_Function_0/NAND4_in[3] ,
         \SB2_0_30/Component_Function_0/NAND4_in[2] ,
         \SB2_0_30/Component_Function_0/NAND4_in[1] ,
         \SB2_0_30/Component_Function_0/NAND4_in[0] ,
         \SB2_0_30/Component_Function_1/NAND4_in[3] ,
         \SB2_0_30/Component_Function_1/NAND4_in[2] ,
         \SB2_0_30/Component_Function_1/NAND4_in[1] ,
         \SB2_0_30/Component_Function_1/NAND4_in[0] ,
         \SB2_0_30/Component_Function_5/NAND4_in[2] ,
         \SB2_0_30/Component_Function_5/NAND4_in[1] ,
         \SB2_0_31/Component_Function_0/NAND4_in[3] ,
         \SB2_0_31/Component_Function_0/NAND4_in[2] ,
         \SB2_0_31/Component_Function_0/NAND4_in[1] ,
         \SB2_0_31/Component_Function_0/NAND4_in[0] ,
         \SB2_0_31/Component_Function_1/NAND4_in[3] ,
         \SB2_0_31/Component_Function_1/NAND4_in[2] ,
         \SB2_0_31/Component_Function_1/NAND4_in[1] ,
         \SB2_0_31/Component_Function_1/NAND4_in[0] ,
         \SB2_0_31/Component_Function_5/NAND4_in[3] ,
         \SB2_0_31/Component_Function_5/NAND4_in[2] ,
         \SB2_0_31/Component_Function_5/NAND4_in[1] ,
         \SB2_0_31/Component_Function_5/NAND4_in[0] ,
         \SB1_1_0/Component_Function_0/NAND4_in[3] ,
         \SB1_1_0/Component_Function_0/NAND4_in[2] ,
         \SB1_1_0/Component_Function_0/NAND4_in[1] ,
         \SB1_1_0/Component_Function_0/NAND4_in[0] ,
         \SB1_1_0/Component_Function_1/NAND4_in[3] ,
         \SB1_1_0/Component_Function_1/NAND4_in[2] ,
         \SB1_1_0/Component_Function_1/NAND4_in[1] ,
         \SB1_1_0/Component_Function_1/NAND4_in[0] ,
         \SB1_1_0/Component_Function_5/NAND4_in[3] ,
         \SB1_1_0/Component_Function_5/NAND4_in[1] ,
         \SB1_1_0/Component_Function_5/NAND4_in[0] ,
         \SB1_1_1/Component_Function_0/NAND4_in[2] ,
         \SB1_1_1/Component_Function_0/NAND4_in[1] ,
         \SB1_1_1/Component_Function_0/NAND4_in[0] ,
         \SB1_1_1/Component_Function_1/NAND4_in[3] ,
         \SB1_1_1/Component_Function_1/NAND4_in[2] ,
         \SB1_1_1/Component_Function_1/NAND4_in[1] ,
         \SB1_1_1/Component_Function_1/NAND4_in[0] ,
         \SB1_1_1/Component_Function_5/NAND4_in[3] ,
         \SB1_1_1/Component_Function_5/NAND4_in[1] ,
         \SB1_1_1/Component_Function_5/NAND4_in[0] ,
         \SB1_1_2/Component_Function_0/NAND4_in[3] ,
         \SB1_1_2/Component_Function_0/NAND4_in[2] ,
         \SB1_1_2/Component_Function_0/NAND4_in[1] ,
         \SB1_1_2/Component_Function_0/NAND4_in[0] ,
         \SB1_1_2/Component_Function_1/NAND4_in[2] ,
         \SB1_1_2/Component_Function_1/NAND4_in[1] ,
         \SB1_1_2/Component_Function_1/NAND4_in[0] ,
         \SB1_1_2/Component_Function_5/NAND4_in[3] ,
         \SB1_1_2/Component_Function_5/NAND4_in[1] ,
         \SB1_1_2/Component_Function_5/NAND4_in[0] ,
         \SB1_1_3/Component_Function_0/NAND4_in[3] ,
         \SB1_1_3/Component_Function_0/NAND4_in[2] ,
         \SB1_1_3/Component_Function_0/NAND4_in[1] ,
         \SB1_1_3/Component_Function_0/NAND4_in[0] ,
         \SB1_1_3/Component_Function_1/NAND4_in[3] ,
         \SB1_1_3/Component_Function_1/NAND4_in[2] ,
         \SB1_1_3/Component_Function_1/NAND4_in[1] ,
         \SB1_1_3/Component_Function_1/NAND4_in[0] ,
         \SB1_1_3/Component_Function_5/NAND4_in[2] ,
         \SB1_1_3/Component_Function_5/NAND4_in[1] ,
         \SB1_1_3/Component_Function_5/NAND4_in[0] ,
         \SB1_1_4/Component_Function_0/NAND4_in[3] ,
         \SB1_1_4/Component_Function_0/NAND4_in[2] ,
         \SB1_1_4/Component_Function_0/NAND4_in[1] ,
         \SB1_1_4/Component_Function_0/NAND4_in[0] ,
         \SB1_1_4/Component_Function_1/NAND4_in[3] ,
         \SB1_1_4/Component_Function_1/NAND4_in[2] ,
         \SB1_1_4/Component_Function_1/NAND4_in[1] ,
         \SB1_1_4/Component_Function_1/NAND4_in[0] ,
         \SB1_1_4/Component_Function_5/NAND4_in[3] ,
         \SB1_1_4/Component_Function_5/NAND4_in[1] ,
         \SB1_1_4/Component_Function_5/NAND4_in[0] ,
         \SB1_1_5/Component_Function_0/NAND4_in[3] ,
         \SB1_1_5/Component_Function_0/NAND4_in[2] ,
         \SB1_1_5/Component_Function_0/NAND4_in[1] ,
         \SB1_1_5/Component_Function_0/NAND4_in[0] ,
         \SB1_1_5/Component_Function_1/NAND4_in[3] ,
         \SB1_1_5/Component_Function_1/NAND4_in[2] ,
         \SB1_1_5/Component_Function_1/NAND4_in[1] ,
         \SB1_1_5/Component_Function_1/NAND4_in[0] ,
         \SB1_1_5/Component_Function_5/NAND4_in[3] ,
         \SB1_1_5/Component_Function_5/NAND4_in[1] ,
         \SB1_1_5/Component_Function_5/NAND4_in[0] ,
         \SB1_1_6/Component_Function_0/NAND4_in[3] ,
         \SB1_1_6/Component_Function_0/NAND4_in[2] ,
         \SB1_1_6/Component_Function_0/NAND4_in[1] ,
         \SB1_1_6/Component_Function_0/NAND4_in[0] ,
         \SB1_1_6/Component_Function_1/NAND4_in[3] ,
         \SB1_1_6/Component_Function_1/NAND4_in[2] ,
         \SB1_1_6/Component_Function_1/NAND4_in[1] ,
         \SB1_1_6/Component_Function_1/NAND4_in[0] ,
         \SB1_1_6/Component_Function_5/NAND4_in[3] ,
         \SB1_1_6/Component_Function_5/NAND4_in[1] ,
         \SB1_1_6/Component_Function_5/NAND4_in[0] ,
         \SB1_1_7/Component_Function_0/NAND4_in[3] ,
         \SB1_1_7/Component_Function_0/NAND4_in[2] ,
         \SB1_1_7/Component_Function_0/NAND4_in[1] ,
         \SB1_1_7/Component_Function_0/NAND4_in[0] ,
         \SB1_1_7/Component_Function_1/NAND4_in[3] ,
         \SB1_1_7/Component_Function_1/NAND4_in[2] ,
         \SB1_1_7/Component_Function_1/NAND4_in[1] ,
         \SB1_1_7/Component_Function_1/NAND4_in[0] ,
         \SB1_1_7/Component_Function_5/NAND4_in[3] ,
         \SB1_1_7/Component_Function_5/NAND4_in[1] ,
         \SB1_1_7/Component_Function_5/NAND4_in[0] ,
         \SB1_1_8/Component_Function_0/NAND4_in[3] ,
         \SB1_1_8/Component_Function_0/NAND4_in[2] ,
         \SB1_1_8/Component_Function_0/NAND4_in[1] ,
         \SB1_1_8/Component_Function_0/NAND4_in[0] ,
         \SB1_1_8/Component_Function_1/NAND4_in[3] ,
         \SB1_1_8/Component_Function_1/NAND4_in[2] ,
         \SB1_1_8/Component_Function_1/NAND4_in[1] ,
         \SB1_1_8/Component_Function_1/NAND4_in[0] ,
         \SB1_1_8/Component_Function_5/NAND4_in[3] ,
         \SB1_1_8/Component_Function_5/NAND4_in[1] ,
         \SB1_1_8/Component_Function_5/NAND4_in[0] ,
         \SB1_1_9/Component_Function_0/NAND4_in[3] ,
         \SB1_1_9/Component_Function_0/NAND4_in[2] ,
         \SB1_1_9/Component_Function_0/NAND4_in[1] ,
         \SB1_1_9/Component_Function_0/NAND4_in[0] ,
         \SB1_1_9/Component_Function_1/NAND4_in[3] ,
         \SB1_1_9/Component_Function_1/NAND4_in[2] ,
         \SB1_1_9/Component_Function_1/NAND4_in[1] ,
         \SB1_1_9/Component_Function_1/NAND4_in[0] ,
         \SB1_1_9/Component_Function_5/NAND4_in[3] ,
         \SB1_1_9/Component_Function_5/NAND4_in[2] ,
         \SB1_1_9/Component_Function_5/NAND4_in[1] ,
         \SB1_1_9/Component_Function_5/NAND4_in[0] ,
         \SB1_1_10/Component_Function_0/NAND4_in[3] ,
         \SB1_1_10/Component_Function_0/NAND4_in[2] ,
         \SB1_1_10/Component_Function_0/NAND4_in[1] ,
         \SB1_1_10/Component_Function_0/NAND4_in[0] ,
         \SB1_1_10/Component_Function_1/NAND4_in[3] ,
         \SB1_1_10/Component_Function_1/NAND4_in[2] ,
         \SB1_1_10/Component_Function_1/NAND4_in[1] ,
         \SB1_1_10/Component_Function_1/NAND4_in[0] ,
         \SB1_1_10/Component_Function_5/NAND4_in[3] ,
         \SB1_1_10/Component_Function_5/NAND4_in[1] ,
         \SB1_1_10/Component_Function_5/NAND4_in[0] ,
         \SB1_1_11/Component_Function_0/NAND4_in[3] ,
         \SB1_1_11/Component_Function_0/NAND4_in[2] ,
         \SB1_1_11/Component_Function_0/NAND4_in[1] ,
         \SB1_1_11/Component_Function_0/NAND4_in[0] ,
         \SB1_1_11/Component_Function_1/NAND4_in[3] ,
         \SB1_1_11/Component_Function_1/NAND4_in[2] ,
         \SB1_1_11/Component_Function_1/NAND4_in[1] ,
         \SB1_1_11/Component_Function_1/NAND4_in[0] ,
         \SB1_1_11/Component_Function_5/NAND4_in[3] ,
         \SB1_1_11/Component_Function_5/NAND4_in[1] ,
         \SB1_1_11/Component_Function_5/NAND4_in[0] ,
         \SB1_1_12/Component_Function_0/NAND4_in[3] ,
         \SB1_1_12/Component_Function_0/NAND4_in[1] ,
         \SB1_1_12/Component_Function_0/NAND4_in[0] ,
         \SB1_1_12/Component_Function_1/NAND4_in[2] ,
         \SB1_1_12/Component_Function_1/NAND4_in[1] ,
         \SB1_1_12/Component_Function_1/NAND4_in[0] ,
         \SB1_1_12/Component_Function_5/NAND4_in[3] ,
         \SB1_1_12/Component_Function_5/NAND4_in[1] ,
         \SB1_1_12/Component_Function_5/NAND4_in[0] ,
         \SB1_1_13/Component_Function_0/NAND4_in[3] ,
         \SB1_1_13/Component_Function_0/NAND4_in[2] ,
         \SB1_1_13/Component_Function_0/NAND4_in[1] ,
         \SB1_1_13/Component_Function_0/NAND4_in[0] ,
         \SB1_1_13/Component_Function_1/NAND4_in[3] ,
         \SB1_1_13/Component_Function_1/NAND4_in[2] ,
         \SB1_1_13/Component_Function_1/NAND4_in[1] ,
         \SB1_1_13/Component_Function_1/NAND4_in[0] ,
         \SB1_1_13/Component_Function_5/NAND4_in[3] ,
         \SB1_1_13/Component_Function_5/NAND4_in[1] ,
         \SB1_1_13/Component_Function_5/NAND4_in[0] ,
         \SB1_1_14/Component_Function_0/NAND4_in[3] ,
         \SB1_1_14/Component_Function_0/NAND4_in[2] ,
         \SB1_1_14/Component_Function_0/NAND4_in[1] ,
         \SB1_1_14/Component_Function_0/NAND4_in[0] ,
         \SB1_1_14/Component_Function_1/NAND4_in[3] ,
         \SB1_1_14/Component_Function_1/NAND4_in[2] ,
         \SB1_1_14/Component_Function_1/NAND4_in[1] ,
         \SB1_1_14/Component_Function_1/NAND4_in[0] ,
         \SB1_1_14/Component_Function_5/NAND4_in[3] ,
         \SB1_1_14/Component_Function_5/NAND4_in[1] ,
         \SB1_1_14/Component_Function_5/NAND4_in[0] ,
         \SB1_1_15/Component_Function_0/NAND4_in[3] ,
         \SB1_1_15/Component_Function_0/NAND4_in[1] ,
         \SB1_1_15/Component_Function_0/NAND4_in[0] ,
         \SB1_1_15/Component_Function_1/NAND4_in[3] ,
         \SB1_1_15/Component_Function_1/NAND4_in[2] ,
         \SB1_1_15/Component_Function_1/NAND4_in[1] ,
         \SB1_1_15/Component_Function_1/NAND4_in[0] ,
         \SB1_1_15/Component_Function_5/NAND4_in[3] ,
         \SB1_1_15/Component_Function_5/NAND4_in[1] ,
         \SB1_1_15/Component_Function_5/NAND4_in[0] ,
         \SB1_1_16/Component_Function_0/NAND4_in[3] ,
         \SB1_1_16/Component_Function_0/NAND4_in[2] ,
         \SB1_1_16/Component_Function_0/NAND4_in[1] ,
         \SB1_1_16/Component_Function_0/NAND4_in[0] ,
         \SB1_1_16/Component_Function_1/NAND4_in[3] ,
         \SB1_1_16/Component_Function_1/NAND4_in[2] ,
         \SB1_1_16/Component_Function_1/NAND4_in[1] ,
         \SB1_1_16/Component_Function_1/NAND4_in[0] ,
         \SB1_1_16/Component_Function_5/NAND4_in[2] ,
         \SB1_1_16/Component_Function_5/NAND4_in[1] ,
         \SB1_1_16/Component_Function_5/NAND4_in[0] ,
         \SB1_1_17/Component_Function_0/NAND4_in[3] ,
         \SB1_1_17/Component_Function_0/NAND4_in[2] ,
         \SB1_1_17/Component_Function_0/NAND4_in[1] ,
         \SB1_1_17/Component_Function_0/NAND4_in[0] ,
         \SB1_1_17/Component_Function_1/NAND4_in[3] ,
         \SB1_1_17/Component_Function_1/NAND4_in[2] ,
         \SB1_1_17/Component_Function_1/NAND4_in[1] ,
         \SB1_1_17/Component_Function_1/NAND4_in[0] ,
         \SB1_1_17/Component_Function_5/NAND4_in[3] ,
         \SB1_1_17/Component_Function_5/NAND4_in[1] ,
         \SB1_1_17/Component_Function_5/NAND4_in[0] ,
         \SB1_1_18/Component_Function_0/NAND4_in[3] ,
         \SB1_1_18/Component_Function_0/NAND4_in[2] ,
         \SB1_1_18/Component_Function_0/NAND4_in[1] ,
         \SB1_1_18/Component_Function_0/NAND4_in[0] ,
         \SB1_1_18/Component_Function_1/NAND4_in[3] ,
         \SB1_1_18/Component_Function_1/NAND4_in[2] ,
         \SB1_1_18/Component_Function_1/NAND4_in[0] ,
         \SB1_1_18/Component_Function_5/NAND4_in[3] ,
         \SB1_1_18/Component_Function_5/NAND4_in[1] ,
         \SB1_1_18/Component_Function_5/NAND4_in[0] ,
         \SB1_1_19/Component_Function_0/NAND4_in[3] ,
         \SB1_1_19/Component_Function_0/NAND4_in[2] ,
         \SB1_1_19/Component_Function_0/NAND4_in[1] ,
         \SB1_1_19/Component_Function_0/NAND4_in[0] ,
         \SB1_1_19/Component_Function_1/NAND4_in[3] ,
         \SB1_1_19/Component_Function_1/NAND4_in[2] ,
         \SB1_1_19/Component_Function_1/NAND4_in[1] ,
         \SB1_1_19/Component_Function_1/NAND4_in[0] ,
         \SB1_1_19/Component_Function_5/NAND4_in[3] ,
         \SB1_1_19/Component_Function_5/NAND4_in[1] ,
         \SB1_1_19/Component_Function_5/NAND4_in[0] ,
         \SB1_1_20/Component_Function_0/NAND4_in[3] ,
         \SB1_1_20/Component_Function_0/NAND4_in[2] ,
         \SB1_1_20/Component_Function_0/NAND4_in[1] ,
         \SB1_1_20/Component_Function_0/NAND4_in[0] ,
         \SB1_1_20/Component_Function_1/NAND4_in[3] ,
         \SB1_1_20/Component_Function_1/NAND4_in[2] ,
         \SB1_1_20/Component_Function_1/NAND4_in[1] ,
         \SB1_1_20/Component_Function_1/NAND4_in[0] ,
         \SB1_1_20/Component_Function_5/NAND4_in[2] ,
         \SB1_1_20/Component_Function_5/NAND4_in[1] ,
         \SB1_1_20/Component_Function_5/NAND4_in[0] ,
         \SB1_1_21/Component_Function_0/NAND4_in[3] ,
         \SB1_1_21/Component_Function_0/NAND4_in[2] ,
         \SB1_1_21/Component_Function_0/NAND4_in[1] ,
         \SB1_1_21/Component_Function_0/NAND4_in[0] ,
         \SB1_1_21/Component_Function_1/NAND4_in[3] ,
         \SB1_1_21/Component_Function_1/NAND4_in[1] ,
         \SB1_1_21/Component_Function_1/NAND4_in[0] ,
         \SB1_1_21/Component_Function_5/NAND4_in[2] ,
         \SB1_1_21/Component_Function_5/NAND4_in[1] ,
         \SB1_1_21/Component_Function_5/NAND4_in[0] ,
         \SB1_1_22/Component_Function_0/NAND4_in[3] ,
         \SB1_1_22/Component_Function_0/NAND4_in[2] ,
         \SB1_1_22/Component_Function_0/NAND4_in[1] ,
         \SB1_1_22/Component_Function_0/NAND4_in[0] ,
         \SB1_1_22/Component_Function_1/NAND4_in[3] ,
         \SB1_1_22/Component_Function_1/NAND4_in[2] ,
         \SB1_1_22/Component_Function_1/NAND4_in[1] ,
         \SB1_1_22/Component_Function_1/NAND4_in[0] ,
         \SB1_1_22/Component_Function_5/NAND4_in[3] ,
         \SB1_1_22/Component_Function_5/NAND4_in[1] ,
         \SB1_1_22/Component_Function_5/NAND4_in[0] ,
         \SB1_1_23/Component_Function_0/NAND4_in[3] ,
         \SB1_1_23/Component_Function_0/NAND4_in[2] ,
         \SB1_1_23/Component_Function_0/NAND4_in[1] ,
         \SB1_1_23/Component_Function_0/NAND4_in[0] ,
         \SB1_1_23/Component_Function_1/NAND4_in[3] ,
         \SB1_1_23/Component_Function_1/NAND4_in[2] ,
         \SB1_1_23/Component_Function_1/NAND4_in[1] ,
         \SB1_1_23/Component_Function_1/NAND4_in[0] ,
         \SB1_1_23/Component_Function_5/NAND4_in[3] ,
         \SB1_1_23/Component_Function_5/NAND4_in[1] ,
         \SB1_1_23/Component_Function_5/NAND4_in[0] ,
         \SB1_1_24/Component_Function_0/NAND4_in[3] ,
         \SB1_1_24/Component_Function_0/NAND4_in[2] ,
         \SB1_1_24/Component_Function_0/NAND4_in[1] ,
         \SB1_1_24/Component_Function_0/NAND4_in[0] ,
         \SB1_1_24/Component_Function_1/NAND4_in[2] ,
         \SB1_1_24/Component_Function_1/NAND4_in[1] ,
         \SB1_1_24/Component_Function_1/NAND4_in[0] ,
         \SB1_1_24/Component_Function_5/NAND4_in[3] ,
         \SB1_1_24/Component_Function_5/NAND4_in[1] ,
         \SB1_1_24/Component_Function_5/NAND4_in[0] ,
         \SB1_1_25/Component_Function_0/NAND4_in[3] ,
         \SB1_1_25/Component_Function_0/NAND4_in[2] ,
         \SB1_1_25/Component_Function_0/NAND4_in[1] ,
         \SB1_1_25/Component_Function_0/NAND4_in[0] ,
         \SB1_1_25/Component_Function_1/NAND4_in[3] ,
         \SB1_1_25/Component_Function_1/NAND4_in[2] ,
         \SB1_1_25/Component_Function_1/NAND4_in[1] ,
         \SB1_1_25/Component_Function_1/NAND4_in[0] ,
         \SB1_1_25/Component_Function_5/NAND4_in[3] ,
         \SB1_1_25/Component_Function_5/NAND4_in[1] ,
         \SB1_1_25/Component_Function_5/NAND4_in[0] ,
         \SB1_1_26/Component_Function_0/NAND4_in[3] ,
         \SB1_1_26/Component_Function_0/NAND4_in[2] ,
         \SB1_1_26/Component_Function_0/NAND4_in[1] ,
         \SB1_1_26/Component_Function_0/NAND4_in[0] ,
         \SB1_1_26/Component_Function_1/NAND4_in[3] ,
         \SB1_1_26/Component_Function_1/NAND4_in[2] ,
         \SB1_1_26/Component_Function_1/NAND4_in[1] ,
         \SB1_1_26/Component_Function_1/NAND4_in[0] ,
         \SB1_1_26/Component_Function_5/NAND4_in[3] ,
         \SB1_1_26/Component_Function_5/NAND4_in[1] ,
         \SB1_1_26/Component_Function_5/NAND4_in[0] ,
         \SB1_1_27/Component_Function_0/NAND4_in[3] ,
         \SB1_1_27/Component_Function_0/NAND4_in[2] ,
         \SB1_1_27/Component_Function_0/NAND4_in[1] ,
         \SB1_1_27/Component_Function_0/NAND4_in[0] ,
         \SB1_1_27/Component_Function_1/NAND4_in[3] ,
         \SB1_1_27/Component_Function_1/NAND4_in[2] ,
         \SB1_1_27/Component_Function_1/NAND4_in[1] ,
         \SB1_1_27/Component_Function_1/NAND4_in[0] ,
         \SB1_1_27/Component_Function_5/NAND4_in[3] ,
         \SB1_1_27/Component_Function_5/NAND4_in[1] ,
         \SB1_1_27/Component_Function_5/NAND4_in[0] ,
         \SB1_1_28/Component_Function_0/NAND4_in[3] ,
         \SB1_1_28/Component_Function_0/NAND4_in[2] ,
         \SB1_1_28/Component_Function_0/NAND4_in[1] ,
         \SB1_1_28/Component_Function_0/NAND4_in[0] ,
         \SB1_1_28/Component_Function_1/NAND4_in[3] ,
         \SB1_1_28/Component_Function_1/NAND4_in[2] ,
         \SB1_1_28/Component_Function_1/NAND4_in[1] ,
         \SB1_1_28/Component_Function_1/NAND4_in[0] ,
         \SB1_1_28/Component_Function_5/NAND4_in[3] ,
         \SB1_1_28/Component_Function_5/NAND4_in[1] ,
         \SB1_1_28/Component_Function_5/NAND4_in[0] ,
         \SB1_1_29/Component_Function_0/NAND4_in[3] ,
         \SB1_1_29/Component_Function_0/NAND4_in[2] ,
         \SB1_1_29/Component_Function_0/NAND4_in[1] ,
         \SB1_1_29/Component_Function_0/NAND4_in[0] ,
         \SB1_1_29/Component_Function_1/NAND4_in[3] ,
         \SB1_1_29/Component_Function_1/NAND4_in[2] ,
         \SB1_1_29/Component_Function_1/NAND4_in[1] ,
         \SB1_1_29/Component_Function_1/NAND4_in[0] ,
         \SB1_1_29/Component_Function_5/NAND4_in[3] ,
         \SB1_1_29/Component_Function_5/NAND4_in[1] ,
         \SB1_1_29/Component_Function_5/NAND4_in[0] ,
         \SB1_1_30/Component_Function_0/NAND4_in[3] ,
         \SB1_1_30/Component_Function_0/NAND4_in[2] ,
         \SB1_1_30/Component_Function_0/NAND4_in[1] ,
         \SB1_1_30/Component_Function_0/NAND4_in[0] ,
         \SB1_1_30/Component_Function_1/NAND4_in[2] ,
         \SB1_1_30/Component_Function_1/NAND4_in[1] ,
         \SB1_1_30/Component_Function_1/NAND4_in[0] ,
         \SB1_1_30/Component_Function_5/NAND4_in[2] ,
         \SB1_1_30/Component_Function_5/NAND4_in[1] ,
         \SB1_1_30/Component_Function_5/NAND4_in[0] ,
         \SB1_1_31/Component_Function_0/NAND4_in[3] ,
         \SB1_1_31/Component_Function_0/NAND4_in[2] ,
         \SB1_1_31/Component_Function_0/NAND4_in[1] ,
         \SB1_1_31/Component_Function_0/NAND4_in[0] ,
         \SB1_1_31/Component_Function_1/NAND4_in[3] ,
         \SB1_1_31/Component_Function_1/NAND4_in[2] ,
         \SB1_1_31/Component_Function_1/NAND4_in[1] ,
         \SB1_1_31/Component_Function_1/NAND4_in[0] ,
         \SB1_1_31/Component_Function_5/NAND4_in[3] ,
         \SB1_1_31/Component_Function_5/NAND4_in[1] ,
         \SB1_1_31/Component_Function_5/NAND4_in[0] ,
         \SB2_1_0/Component_Function_0/NAND4_in[3] ,
         \SB2_1_0/Component_Function_0/NAND4_in[2] ,
         \SB2_1_0/Component_Function_0/NAND4_in[1] ,
         \SB2_1_0/Component_Function_0/NAND4_in[0] ,
         \SB2_1_0/Component_Function_1/NAND4_in[3] ,
         \SB2_1_0/Component_Function_1/NAND4_in[2] ,
         \SB2_1_0/Component_Function_1/NAND4_in[1] ,
         \SB2_1_0/Component_Function_1/NAND4_in[0] ,
         \SB2_1_0/Component_Function_5/NAND4_in[2] ,
         \SB2_1_0/Component_Function_5/NAND4_in[1] ,
         \SB2_1_0/Component_Function_5/NAND4_in[0] ,
         \SB2_1_1/Component_Function_0/NAND4_in[3] ,
         \SB2_1_1/Component_Function_0/NAND4_in[2] ,
         \SB2_1_1/Component_Function_0/NAND4_in[1] ,
         \SB2_1_1/Component_Function_0/NAND4_in[0] ,
         \SB2_1_1/Component_Function_1/NAND4_in[3] ,
         \SB2_1_1/Component_Function_1/NAND4_in[2] ,
         \SB2_1_1/Component_Function_1/NAND4_in[1] ,
         \SB2_1_1/Component_Function_1/NAND4_in[0] ,
         \SB2_1_1/Component_Function_5/NAND4_in[3] ,
         \SB2_1_1/Component_Function_5/NAND4_in[1] ,
         \SB2_1_1/Component_Function_5/NAND4_in[0] ,
         \SB2_1_2/Component_Function_0/NAND4_in[3] ,
         \SB2_1_2/Component_Function_0/NAND4_in[2] ,
         \SB2_1_2/Component_Function_0/NAND4_in[1] ,
         \SB2_1_2/Component_Function_0/NAND4_in[0] ,
         \SB2_1_2/Component_Function_1/NAND4_in[3] ,
         \SB2_1_2/Component_Function_1/NAND4_in[2] ,
         \SB2_1_2/Component_Function_1/NAND4_in[1] ,
         \SB2_1_2/Component_Function_1/NAND4_in[0] ,
         \SB2_1_2/Component_Function_5/NAND4_in[2] ,
         \SB2_1_2/Component_Function_5/NAND4_in[1] ,
         \SB2_1_2/Component_Function_5/NAND4_in[0] ,
         \SB2_1_3/Component_Function_0/NAND4_in[3] ,
         \SB2_1_3/Component_Function_0/NAND4_in[2] ,
         \SB2_1_3/Component_Function_0/NAND4_in[1] ,
         \SB2_1_3/Component_Function_0/NAND4_in[0] ,
         \SB2_1_3/Component_Function_1/NAND4_in[2] ,
         \SB2_1_3/Component_Function_1/NAND4_in[1] ,
         \SB2_1_3/Component_Function_1/NAND4_in[0] ,
         \SB2_1_3/Component_Function_5/NAND4_in[2] ,
         \SB2_1_3/Component_Function_5/NAND4_in[1] ,
         \SB2_1_4/Component_Function_0/NAND4_in[3] ,
         \SB2_1_4/Component_Function_0/NAND4_in[2] ,
         \SB2_1_4/Component_Function_0/NAND4_in[1] ,
         \SB2_1_4/Component_Function_0/NAND4_in[0] ,
         \SB2_1_4/Component_Function_1/NAND4_in[3] ,
         \SB2_1_4/Component_Function_1/NAND4_in[2] ,
         \SB2_1_4/Component_Function_1/NAND4_in[1] ,
         \SB2_1_4/Component_Function_1/NAND4_in[0] ,
         \SB2_1_4/Component_Function_5/NAND4_in[3] ,
         \SB2_1_4/Component_Function_5/NAND4_in[2] ,
         \SB2_1_4/Component_Function_5/NAND4_in[1] ,
         \SB2_1_4/Component_Function_5/NAND4_in[0] ,
         \SB2_1_5/Component_Function_0/NAND4_in[3] ,
         \SB2_1_5/Component_Function_0/NAND4_in[2] ,
         \SB2_1_5/Component_Function_0/NAND4_in[1] ,
         \SB2_1_5/Component_Function_0/NAND4_in[0] ,
         \SB2_1_5/Component_Function_1/NAND4_in[3] ,
         \SB2_1_5/Component_Function_1/NAND4_in[2] ,
         \SB2_1_5/Component_Function_1/NAND4_in[1] ,
         \SB2_1_5/Component_Function_1/NAND4_in[0] ,
         \SB2_1_5/Component_Function_5/NAND4_in[2] ,
         \SB2_1_5/Component_Function_5/NAND4_in[1] ,
         \SB2_1_6/Component_Function_0/NAND4_in[3] ,
         \SB2_1_6/Component_Function_0/NAND4_in[2] ,
         \SB2_1_6/Component_Function_0/NAND4_in[1] ,
         \SB2_1_6/Component_Function_0/NAND4_in[0] ,
         \SB2_1_6/Component_Function_1/NAND4_in[3] ,
         \SB2_1_6/Component_Function_1/NAND4_in[2] ,
         \SB2_1_6/Component_Function_1/NAND4_in[1] ,
         \SB2_1_6/Component_Function_1/NAND4_in[0] ,
         \SB2_1_6/Component_Function_5/NAND4_in[3] ,
         \SB2_1_6/Component_Function_5/NAND4_in[2] ,
         \SB2_1_6/Component_Function_5/NAND4_in[1] ,
         \SB2_1_6/Component_Function_5/NAND4_in[0] ,
         \SB2_1_7/Component_Function_0/NAND4_in[3] ,
         \SB2_1_7/Component_Function_0/NAND4_in[2] ,
         \SB2_1_7/Component_Function_0/NAND4_in[1] ,
         \SB2_1_7/Component_Function_0/NAND4_in[0] ,
         \SB2_1_7/Component_Function_1/NAND4_in[3] ,
         \SB2_1_7/Component_Function_1/NAND4_in[2] ,
         \SB2_1_7/Component_Function_1/NAND4_in[1] ,
         \SB2_1_7/Component_Function_1/NAND4_in[0] ,
         \SB2_1_7/Component_Function_5/NAND4_in[3] ,
         \SB2_1_7/Component_Function_5/NAND4_in[2] ,
         \SB2_1_7/Component_Function_5/NAND4_in[1] ,
         \SB2_1_7/Component_Function_5/NAND4_in[0] ,
         \SB2_1_8/Component_Function_0/NAND4_in[3] ,
         \SB2_1_8/Component_Function_0/NAND4_in[2] ,
         \SB2_1_8/Component_Function_0/NAND4_in[1] ,
         \SB2_1_8/Component_Function_0/NAND4_in[0] ,
         \SB2_1_8/Component_Function_1/NAND4_in[3] ,
         \SB2_1_8/Component_Function_1/NAND4_in[2] ,
         \SB2_1_8/Component_Function_1/NAND4_in[1] ,
         \SB2_1_8/Component_Function_1/NAND4_in[0] ,
         \SB2_1_8/Component_Function_5/NAND4_in[3] ,
         \SB2_1_8/Component_Function_5/NAND4_in[2] ,
         \SB2_1_8/Component_Function_5/NAND4_in[1] ,
         \SB2_1_8/Component_Function_5/NAND4_in[0] ,
         \SB2_1_9/Component_Function_0/NAND4_in[3] ,
         \SB2_1_9/Component_Function_0/NAND4_in[2] ,
         \SB2_1_9/Component_Function_0/NAND4_in[1] ,
         \SB2_1_9/Component_Function_0/NAND4_in[0] ,
         \SB2_1_9/Component_Function_1/NAND4_in[3] ,
         \SB2_1_9/Component_Function_1/NAND4_in[2] ,
         \SB2_1_9/Component_Function_1/NAND4_in[1] ,
         \SB2_1_9/Component_Function_1/NAND4_in[0] ,
         \SB2_1_9/Component_Function_5/NAND4_in[3] ,
         \SB2_1_9/Component_Function_5/NAND4_in[2] ,
         \SB2_1_9/Component_Function_5/NAND4_in[1] ,
         \SB2_1_9/Component_Function_5/NAND4_in[0] ,
         \SB2_1_10/Component_Function_0/NAND4_in[3] ,
         \SB2_1_10/Component_Function_0/NAND4_in[2] ,
         \SB2_1_10/Component_Function_0/NAND4_in[1] ,
         \SB2_1_10/Component_Function_0/NAND4_in[0] ,
         \SB2_1_10/Component_Function_1/NAND4_in[3] ,
         \SB2_1_10/Component_Function_1/NAND4_in[2] ,
         \SB2_1_10/Component_Function_1/NAND4_in[1] ,
         \SB2_1_10/Component_Function_1/NAND4_in[0] ,
         \SB2_1_10/Component_Function_5/NAND4_in[3] ,
         \SB2_1_10/Component_Function_5/NAND4_in[1] ,
         \SB2_1_10/Component_Function_5/NAND4_in[0] ,
         \SB2_1_11/Component_Function_0/NAND4_in[3] ,
         \SB2_1_11/Component_Function_0/NAND4_in[2] ,
         \SB2_1_11/Component_Function_0/NAND4_in[1] ,
         \SB2_1_11/Component_Function_0/NAND4_in[0] ,
         \SB2_1_11/Component_Function_1/NAND4_in[3] ,
         \SB2_1_11/Component_Function_1/NAND4_in[2] ,
         \SB2_1_11/Component_Function_1/NAND4_in[1] ,
         \SB2_1_11/Component_Function_1/NAND4_in[0] ,
         \SB2_1_11/Component_Function_5/NAND4_in[3] ,
         \SB2_1_11/Component_Function_5/NAND4_in[2] ,
         \SB2_1_11/Component_Function_5/NAND4_in[1] ,
         \SB2_1_12/Component_Function_0/NAND4_in[3] ,
         \SB2_1_12/Component_Function_0/NAND4_in[2] ,
         \SB2_1_12/Component_Function_0/NAND4_in[1] ,
         \SB2_1_12/Component_Function_0/NAND4_in[0] ,
         \SB2_1_12/Component_Function_1/NAND4_in[3] ,
         \SB2_1_12/Component_Function_1/NAND4_in[2] ,
         \SB2_1_12/Component_Function_1/NAND4_in[1] ,
         \SB2_1_12/Component_Function_1/NAND4_in[0] ,
         \SB2_1_12/Component_Function_5/NAND4_in[3] ,
         \SB2_1_12/Component_Function_5/NAND4_in[2] ,
         \SB2_1_12/Component_Function_5/NAND4_in[1] ,
         \SB2_1_13/Component_Function_0/NAND4_in[3] ,
         \SB2_1_13/Component_Function_0/NAND4_in[2] ,
         \SB2_1_13/Component_Function_0/NAND4_in[1] ,
         \SB2_1_13/Component_Function_0/NAND4_in[0] ,
         \SB2_1_13/Component_Function_1/NAND4_in[3] ,
         \SB2_1_13/Component_Function_1/NAND4_in[2] ,
         \SB2_1_13/Component_Function_1/NAND4_in[1] ,
         \SB2_1_13/Component_Function_1/NAND4_in[0] ,
         \SB2_1_13/Component_Function_5/NAND4_in[3] ,
         \SB2_1_13/Component_Function_5/NAND4_in[2] ,
         \SB2_1_13/Component_Function_5/NAND4_in[1] ,
         \SB2_1_13/Component_Function_5/NAND4_in[0] ,
         \SB2_1_14/Component_Function_0/NAND4_in[3] ,
         \SB2_1_14/Component_Function_0/NAND4_in[2] ,
         \SB2_1_14/Component_Function_0/NAND4_in[1] ,
         \SB2_1_14/Component_Function_0/NAND4_in[0] ,
         \SB2_1_14/Component_Function_1/NAND4_in[2] ,
         \SB2_1_14/Component_Function_1/NAND4_in[1] ,
         \SB2_1_14/Component_Function_1/NAND4_in[0] ,
         \SB2_1_14/Component_Function_5/NAND4_in[3] ,
         \SB2_1_14/Component_Function_5/NAND4_in[2] ,
         \SB2_1_14/Component_Function_5/NAND4_in[1] ,
         \SB2_1_14/Component_Function_5/NAND4_in[0] ,
         \SB2_1_15/Component_Function_0/NAND4_in[3] ,
         \SB2_1_15/Component_Function_0/NAND4_in[2] ,
         \SB2_1_15/Component_Function_0/NAND4_in[1] ,
         \SB2_1_15/Component_Function_0/NAND4_in[0] ,
         \SB2_1_15/Component_Function_1/NAND4_in[2] ,
         \SB2_1_15/Component_Function_1/NAND4_in[1] ,
         \SB2_1_15/Component_Function_1/NAND4_in[0] ,
         \SB2_1_15/Component_Function_5/NAND4_in[3] ,
         \SB2_1_15/Component_Function_5/NAND4_in[2] ,
         \SB2_1_15/Component_Function_5/NAND4_in[1] ,
         \SB2_1_15/Component_Function_5/NAND4_in[0] ,
         \SB2_1_16/Component_Function_0/NAND4_in[3] ,
         \SB2_1_16/Component_Function_0/NAND4_in[2] ,
         \SB2_1_16/Component_Function_0/NAND4_in[1] ,
         \SB2_1_16/Component_Function_0/NAND4_in[0] ,
         \SB2_1_16/Component_Function_1/NAND4_in[2] ,
         \SB2_1_16/Component_Function_1/NAND4_in[1] ,
         \SB2_1_16/Component_Function_1/NAND4_in[0] ,
         \SB2_1_16/Component_Function_5/NAND4_in[3] ,
         \SB2_1_16/Component_Function_5/NAND4_in[2] ,
         \SB2_1_16/Component_Function_5/NAND4_in[1] ,
         \SB2_1_16/Component_Function_5/NAND4_in[0] ,
         \SB2_1_17/Component_Function_0/NAND4_in[3] ,
         \SB2_1_17/Component_Function_0/NAND4_in[2] ,
         \SB2_1_17/Component_Function_0/NAND4_in[1] ,
         \SB2_1_17/Component_Function_0/NAND4_in[0] ,
         \SB2_1_17/Component_Function_1/NAND4_in[3] ,
         \SB2_1_17/Component_Function_1/NAND4_in[2] ,
         \SB2_1_17/Component_Function_1/NAND4_in[1] ,
         \SB2_1_17/Component_Function_1/NAND4_in[0] ,
         \SB2_1_17/Component_Function_5/NAND4_in[2] ,
         \SB2_1_17/Component_Function_5/NAND4_in[1] ,
         \SB2_1_17/Component_Function_5/NAND4_in[0] ,
         \SB2_1_18/Component_Function_0/NAND4_in[3] ,
         \SB2_1_18/Component_Function_0/NAND4_in[2] ,
         \SB2_1_18/Component_Function_0/NAND4_in[1] ,
         \SB2_1_18/Component_Function_0/NAND4_in[0] ,
         \SB2_1_18/Component_Function_1/NAND4_in[3] ,
         \SB2_1_18/Component_Function_1/NAND4_in[2] ,
         \SB2_1_18/Component_Function_1/NAND4_in[1] ,
         \SB2_1_18/Component_Function_1/NAND4_in[0] ,
         \SB2_1_18/Component_Function_5/NAND4_in[3] ,
         \SB2_1_18/Component_Function_5/NAND4_in[2] ,
         \SB2_1_18/Component_Function_5/NAND4_in[1] ,
         \SB2_1_18/Component_Function_5/NAND4_in[0] ,
         \SB2_1_19/Component_Function_0/NAND4_in[3] ,
         \SB2_1_19/Component_Function_0/NAND4_in[2] ,
         \SB2_1_19/Component_Function_0/NAND4_in[1] ,
         \SB2_1_19/Component_Function_0/NAND4_in[0] ,
         \SB2_1_19/Component_Function_1/NAND4_in[2] ,
         \SB2_1_19/Component_Function_1/NAND4_in[1] ,
         \SB2_1_19/Component_Function_1/NAND4_in[0] ,
         \SB2_1_19/Component_Function_5/NAND4_in[3] ,
         \SB2_1_19/Component_Function_5/NAND4_in[2] ,
         \SB2_1_19/Component_Function_5/NAND4_in[1] ,
         \SB2_1_19/Component_Function_5/NAND4_in[0] ,
         \SB2_1_20/Component_Function_0/NAND4_in[2] ,
         \SB2_1_20/Component_Function_0/NAND4_in[1] ,
         \SB2_1_20/Component_Function_0/NAND4_in[0] ,
         \SB2_1_20/Component_Function_1/NAND4_in[3] ,
         \SB2_1_20/Component_Function_1/NAND4_in[2] ,
         \SB2_1_20/Component_Function_1/NAND4_in[1] ,
         \SB2_1_20/Component_Function_1/NAND4_in[0] ,
         \SB2_1_20/Component_Function_5/NAND4_in[3] ,
         \SB2_1_20/Component_Function_5/NAND4_in[2] ,
         \SB2_1_20/Component_Function_5/NAND4_in[1] ,
         \SB2_1_21/Component_Function_0/NAND4_in[3] ,
         \SB2_1_21/Component_Function_0/NAND4_in[2] ,
         \SB2_1_21/Component_Function_0/NAND4_in[1] ,
         \SB2_1_21/Component_Function_0/NAND4_in[0] ,
         \SB2_1_21/Component_Function_1/NAND4_in[3] ,
         \SB2_1_21/Component_Function_1/NAND4_in[2] ,
         \SB2_1_21/Component_Function_1/NAND4_in[1] ,
         \SB2_1_21/Component_Function_1/NAND4_in[0] ,
         \SB2_1_21/Component_Function_5/NAND4_in[3] ,
         \SB2_1_21/Component_Function_5/NAND4_in[2] ,
         \SB2_1_21/Component_Function_5/NAND4_in[1] ,
         \SB2_1_21/Component_Function_5/NAND4_in[0] ,
         \SB2_1_22/Component_Function_0/NAND4_in[3] ,
         \SB2_1_22/Component_Function_0/NAND4_in[2] ,
         \SB2_1_22/Component_Function_0/NAND4_in[1] ,
         \SB2_1_22/Component_Function_0/NAND4_in[0] ,
         \SB2_1_22/Component_Function_1/NAND4_in[3] ,
         \SB2_1_22/Component_Function_1/NAND4_in[2] ,
         \SB2_1_22/Component_Function_1/NAND4_in[1] ,
         \SB2_1_22/Component_Function_1/NAND4_in[0] ,
         \SB2_1_22/Component_Function_5/NAND4_in[3] ,
         \SB2_1_22/Component_Function_5/NAND4_in[1] ,
         \SB2_1_22/Component_Function_5/NAND4_in[0] ,
         \SB2_1_23/Component_Function_0/NAND4_in[3] ,
         \SB2_1_23/Component_Function_0/NAND4_in[2] ,
         \SB2_1_23/Component_Function_0/NAND4_in[1] ,
         \SB2_1_23/Component_Function_0/NAND4_in[0] ,
         \SB2_1_23/Component_Function_1/NAND4_in[3] ,
         \SB2_1_23/Component_Function_1/NAND4_in[2] ,
         \SB2_1_23/Component_Function_1/NAND4_in[1] ,
         \SB2_1_23/Component_Function_1/NAND4_in[0] ,
         \SB2_1_23/Component_Function_5/NAND4_in[3] ,
         \SB2_1_23/Component_Function_5/NAND4_in[1] ,
         \SB2_1_23/Component_Function_5/NAND4_in[0] ,
         \SB2_1_24/Component_Function_0/NAND4_in[3] ,
         \SB2_1_24/Component_Function_0/NAND4_in[2] ,
         \SB2_1_24/Component_Function_0/NAND4_in[1] ,
         \SB2_1_24/Component_Function_0/NAND4_in[0] ,
         \SB2_1_24/Component_Function_1/NAND4_in[3] ,
         \SB2_1_24/Component_Function_1/NAND4_in[2] ,
         \SB2_1_24/Component_Function_1/NAND4_in[1] ,
         \SB2_1_24/Component_Function_1/NAND4_in[0] ,
         \SB2_1_24/Component_Function_5/NAND4_in[3] ,
         \SB2_1_24/Component_Function_5/NAND4_in[2] ,
         \SB2_1_24/Component_Function_5/NAND4_in[1] ,
         \SB2_1_25/Component_Function_0/NAND4_in[2] ,
         \SB2_1_25/Component_Function_0/NAND4_in[1] ,
         \SB2_1_25/Component_Function_0/NAND4_in[0] ,
         \SB2_1_25/Component_Function_1/NAND4_in[3] ,
         \SB2_1_25/Component_Function_1/NAND4_in[2] ,
         \SB2_1_25/Component_Function_1/NAND4_in[1] ,
         \SB2_1_25/Component_Function_1/NAND4_in[0] ,
         \SB2_1_25/Component_Function_5/NAND4_in[3] ,
         \SB2_1_25/Component_Function_5/NAND4_in[1] ,
         \SB2_1_25/Component_Function_5/NAND4_in[0] ,
         \SB2_1_26/Component_Function_0/NAND4_in[3] ,
         \SB2_1_26/Component_Function_0/NAND4_in[2] ,
         \SB2_1_26/Component_Function_0/NAND4_in[1] ,
         \SB2_1_26/Component_Function_0/NAND4_in[0] ,
         \SB2_1_26/Component_Function_1/NAND4_in[2] ,
         \SB2_1_26/Component_Function_1/NAND4_in[1] ,
         \SB2_1_26/Component_Function_1/NAND4_in[0] ,
         \SB2_1_26/Component_Function_5/NAND4_in[3] ,
         \SB2_1_26/Component_Function_5/NAND4_in[2] ,
         \SB2_1_26/Component_Function_5/NAND4_in[1] ,
         \SB2_1_26/Component_Function_5/NAND4_in[0] ,
         \SB2_1_27/Component_Function_0/NAND4_in[3] ,
         \SB2_1_27/Component_Function_0/NAND4_in[2] ,
         \SB2_1_27/Component_Function_0/NAND4_in[1] ,
         \SB2_1_27/Component_Function_0/NAND4_in[0] ,
         \SB2_1_27/Component_Function_1/NAND4_in[3] ,
         \SB2_1_27/Component_Function_1/NAND4_in[2] ,
         \SB2_1_27/Component_Function_1/NAND4_in[1] ,
         \SB2_1_27/Component_Function_1/NAND4_in[0] ,
         \SB2_1_27/Component_Function_5/NAND4_in[3] ,
         \SB2_1_27/Component_Function_5/NAND4_in[1] ,
         \SB2_1_27/Component_Function_5/NAND4_in[0] ,
         \SB2_1_28/Component_Function_0/NAND4_in[3] ,
         \SB2_1_28/Component_Function_0/NAND4_in[2] ,
         \SB2_1_28/Component_Function_0/NAND4_in[1] ,
         \SB2_1_28/Component_Function_0/NAND4_in[0] ,
         \SB2_1_28/Component_Function_1/NAND4_in[3] ,
         \SB2_1_28/Component_Function_1/NAND4_in[2] ,
         \SB2_1_28/Component_Function_1/NAND4_in[1] ,
         \SB2_1_28/Component_Function_1/NAND4_in[0] ,
         \SB2_1_28/Component_Function_5/NAND4_in[3] ,
         \SB2_1_28/Component_Function_5/NAND4_in[2] ,
         \SB2_1_28/Component_Function_5/NAND4_in[1] ,
         \SB2_1_29/Component_Function_0/NAND4_in[3] ,
         \SB2_1_29/Component_Function_0/NAND4_in[2] ,
         \SB2_1_29/Component_Function_0/NAND4_in[1] ,
         \SB2_1_29/Component_Function_0/NAND4_in[0] ,
         \SB2_1_29/Component_Function_1/NAND4_in[2] ,
         \SB2_1_29/Component_Function_1/NAND4_in[1] ,
         \SB2_1_29/Component_Function_1/NAND4_in[0] ,
         \SB2_1_29/Component_Function_5/NAND4_in[3] ,
         \SB2_1_29/Component_Function_5/NAND4_in[2] ,
         \SB2_1_29/Component_Function_5/NAND4_in[1] ,
         \SB2_1_30/Component_Function_0/NAND4_in[3] ,
         \SB2_1_30/Component_Function_0/NAND4_in[2] ,
         \SB2_1_30/Component_Function_0/NAND4_in[1] ,
         \SB2_1_30/Component_Function_0/NAND4_in[0] ,
         \SB2_1_30/Component_Function_1/NAND4_in[3] ,
         \SB2_1_30/Component_Function_1/NAND4_in[2] ,
         \SB2_1_30/Component_Function_1/NAND4_in[1] ,
         \SB2_1_30/Component_Function_1/NAND4_in[0] ,
         \SB2_1_30/Component_Function_5/NAND4_in[2] ,
         \SB2_1_30/Component_Function_5/NAND4_in[1] ,
         \SB2_1_30/Component_Function_5/NAND4_in[0] ,
         \SB2_1_31/Component_Function_0/NAND4_in[3] ,
         \SB2_1_31/Component_Function_0/NAND4_in[2] ,
         \SB2_1_31/Component_Function_0/NAND4_in[1] ,
         \SB2_1_31/Component_Function_0/NAND4_in[0] ,
         \SB2_1_31/Component_Function_1/NAND4_in[2] ,
         \SB2_1_31/Component_Function_1/NAND4_in[1] ,
         \SB2_1_31/Component_Function_1/NAND4_in[0] ,
         \SB2_1_31/Component_Function_5/NAND4_in[3] ,
         \SB2_1_31/Component_Function_5/NAND4_in[2] ,
         \SB2_1_31/Component_Function_5/NAND4_in[1] ,
         \SB2_1_31/Component_Function_5/NAND4_in[0] ,
         \SB1_2_0/Component_Function_0/NAND4_in[3] ,
         \SB1_2_0/Component_Function_0/NAND4_in[2] ,
         \SB1_2_0/Component_Function_0/NAND4_in[1] ,
         \SB1_2_0/Component_Function_0/NAND4_in[0] ,
         \SB1_2_0/Component_Function_1/NAND4_in[3] ,
         \SB1_2_0/Component_Function_1/NAND4_in[2] ,
         \SB1_2_0/Component_Function_1/NAND4_in[1] ,
         \SB1_2_0/Component_Function_1/NAND4_in[0] ,
         \SB1_2_0/Component_Function_5/NAND4_in[3] ,
         \SB1_2_0/Component_Function_5/NAND4_in[1] ,
         \SB1_2_0/Component_Function_5/NAND4_in[0] ,
         \SB1_2_1/Component_Function_0/NAND4_in[3] ,
         \SB1_2_1/Component_Function_0/NAND4_in[2] ,
         \SB1_2_1/Component_Function_0/NAND4_in[1] ,
         \SB1_2_1/Component_Function_0/NAND4_in[0] ,
         \SB1_2_1/Component_Function_1/NAND4_in[3] ,
         \SB1_2_1/Component_Function_1/NAND4_in[2] ,
         \SB1_2_1/Component_Function_1/NAND4_in[1] ,
         \SB1_2_1/Component_Function_1/NAND4_in[0] ,
         \SB1_2_1/Component_Function_5/NAND4_in[3] ,
         \SB1_2_1/Component_Function_5/NAND4_in[1] ,
         \SB1_2_1/Component_Function_5/NAND4_in[0] ,
         \SB1_2_2/Component_Function_0/NAND4_in[3] ,
         \SB1_2_2/Component_Function_0/NAND4_in[1] ,
         \SB1_2_2/Component_Function_0/NAND4_in[0] ,
         \SB1_2_2/Component_Function_1/NAND4_in[3] ,
         \SB1_2_2/Component_Function_1/NAND4_in[1] ,
         \SB1_2_2/Component_Function_1/NAND4_in[0] ,
         \SB1_2_2/Component_Function_5/NAND4_in[3] ,
         \SB1_2_2/Component_Function_5/NAND4_in[1] ,
         \SB1_2_2/Component_Function_5/NAND4_in[0] ,
         \SB1_2_3/Component_Function_0/NAND4_in[3] ,
         \SB1_2_3/Component_Function_0/NAND4_in[2] ,
         \SB1_2_3/Component_Function_0/NAND4_in[1] ,
         \SB1_2_3/Component_Function_0/NAND4_in[0] ,
         \SB1_2_3/Component_Function_1/NAND4_in[3] ,
         \SB1_2_3/Component_Function_1/NAND4_in[2] ,
         \SB1_2_3/Component_Function_1/NAND4_in[1] ,
         \SB1_2_3/Component_Function_1/NAND4_in[0] ,
         \SB1_2_3/Component_Function_5/NAND4_in[3] ,
         \SB1_2_3/Component_Function_5/NAND4_in[1] ,
         \SB1_2_3/Component_Function_5/NAND4_in[0] ,
         \SB1_2_4/Component_Function_0/NAND4_in[3] ,
         \SB1_2_4/Component_Function_0/NAND4_in[2] ,
         \SB1_2_4/Component_Function_0/NAND4_in[1] ,
         \SB1_2_4/Component_Function_0/NAND4_in[0] ,
         \SB1_2_4/Component_Function_1/NAND4_in[3] ,
         \SB1_2_4/Component_Function_1/NAND4_in[2] ,
         \SB1_2_4/Component_Function_1/NAND4_in[1] ,
         \SB1_2_4/Component_Function_1/NAND4_in[0] ,
         \SB1_2_4/Component_Function_5/NAND4_in[3] ,
         \SB1_2_4/Component_Function_5/NAND4_in[1] ,
         \SB1_2_4/Component_Function_5/NAND4_in[0] ,
         \SB1_2_5/Component_Function_0/NAND4_in[3] ,
         \SB1_2_5/Component_Function_0/NAND4_in[2] ,
         \SB1_2_5/Component_Function_0/NAND4_in[1] ,
         \SB1_2_5/Component_Function_0/NAND4_in[0] ,
         \SB1_2_5/Component_Function_1/NAND4_in[3] ,
         \SB1_2_5/Component_Function_1/NAND4_in[2] ,
         \SB1_2_5/Component_Function_1/NAND4_in[1] ,
         \SB1_2_5/Component_Function_1/NAND4_in[0] ,
         \SB1_2_5/Component_Function_5/NAND4_in[2] ,
         \SB1_2_5/Component_Function_5/NAND4_in[1] ,
         \SB1_2_5/Component_Function_5/NAND4_in[0] ,
         \SB1_2_6/Component_Function_0/NAND4_in[3] ,
         \SB1_2_6/Component_Function_0/NAND4_in[2] ,
         \SB1_2_6/Component_Function_0/NAND4_in[1] ,
         \SB1_2_6/Component_Function_0/NAND4_in[0] ,
         \SB1_2_6/Component_Function_1/NAND4_in[3] ,
         \SB1_2_6/Component_Function_1/NAND4_in[2] ,
         \SB1_2_6/Component_Function_1/NAND4_in[1] ,
         \SB1_2_6/Component_Function_1/NAND4_in[0] ,
         \SB1_2_6/Component_Function_5/NAND4_in[2] ,
         \SB1_2_6/Component_Function_5/NAND4_in[1] ,
         \SB1_2_6/Component_Function_5/NAND4_in[0] ,
         \SB1_2_7/Component_Function_0/NAND4_in[3] ,
         \SB1_2_7/Component_Function_0/NAND4_in[2] ,
         \SB1_2_7/Component_Function_0/NAND4_in[1] ,
         \SB1_2_7/Component_Function_0/NAND4_in[0] ,
         \SB1_2_7/Component_Function_1/NAND4_in[3] ,
         \SB1_2_7/Component_Function_1/NAND4_in[2] ,
         \SB1_2_7/Component_Function_1/NAND4_in[1] ,
         \SB1_2_7/Component_Function_1/NAND4_in[0] ,
         \SB1_2_7/Component_Function_5/NAND4_in[3] ,
         \SB1_2_7/Component_Function_5/NAND4_in[1] ,
         \SB1_2_7/Component_Function_5/NAND4_in[0] ,
         \SB1_2_8/Component_Function_0/NAND4_in[3] ,
         \SB1_2_8/Component_Function_0/NAND4_in[2] ,
         \SB1_2_8/Component_Function_0/NAND4_in[1] ,
         \SB1_2_8/Component_Function_0/NAND4_in[0] ,
         \SB1_2_8/Component_Function_1/NAND4_in[3] ,
         \SB1_2_8/Component_Function_1/NAND4_in[2] ,
         \SB1_2_8/Component_Function_1/NAND4_in[1] ,
         \SB1_2_8/Component_Function_1/NAND4_in[0] ,
         \SB1_2_8/Component_Function_5/NAND4_in[2] ,
         \SB1_2_8/Component_Function_5/NAND4_in[1] ,
         \SB1_2_8/Component_Function_5/NAND4_in[0] ,
         \SB1_2_9/Component_Function_0/NAND4_in[3] ,
         \SB1_2_9/Component_Function_0/NAND4_in[2] ,
         \SB1_2_9/Component_Function_0/NAND4_in[1] ,
         \SB1_2_9/Component_Function_0/NAND4_in[0] ,
         \SB1_2_9/Component_Function_1/NAND4_in[3] ,
         \SB1_2_9/Component_Function_1/NAND4_in[2] ,
         \SB1_2_9/Component_Function_1/NAND4_in[1] ,
         \SB1_2_9/Component_Function_1/NAND4_in[0] ,
         \SB1_2_9/Component_Function_5/NAND4_in[3] ,
         \SB1_2_9/Component_Function_5/NAND4_in[1] ,
         \SB1_2_9/Component_Function_5/NAND4_in[0] ,
         \SB1_2_10/Component_Function_0/NAND4_in[3] ,
         \SB1_2_10/Component_Function_0/NAND4_in[1] ,
         \SB1_2_10/Component_Function_0/NAND4_in[0] ,
         \SB1_2_10/Component_Function_1/NAND4_in[3] ,
         \SB1_2_10/Component_Function_1/NAND4_in[2] ,
         \SB1_2_10/Component_Function_1/NAND4_in[1] ,
         \SB1_2_10/Component_Function_1/NAND4_in[0] ,
         \SB1_2_10/Component_Function_5/NAND4_in[3] ,
         \SB1_2_10/Component_Function_5/NAND4_in[1] ,
         \SB1_2_10/Component_Function_5/NAND4_in[0] ,
         \SB1_2_11/Component_Function_0/NAND4_in[3] ,
         \SB1_2_11/Component_Function_0/NAND4_in[2] ,
         \SB1_2_11/Component_Function_0/NAND4_in[1] ,
         \SB1_2_11/Component_Function_0/NAND4_in[0] ,
         \SB1_2_11/Component_Function_1/NAND4_in[3] ,
         \SB1_2_11/Component_Function_1/NAND4_in[2] ,
         \SB1_2_11/Component_Function_1/NAND4_in[1] ,
         \SB1_2_11/Component_Function_1/NAND4_in[0] ,
         \SB1_2_11/Component_Function_5/NAND4_in[3] ,
         \SB1_2_11/Component_Function_5/NAND4_in[1] ,
         \SB1_2_11/Component_Function_5/NAND4_in[0] ,
         \SB1_2_12/Component_Function_0/NAND4_in[2] ,
         \SB1_2_12/Component_Function_0/NAND4_in[1] ,
         \SB1_2_12/Component_Function_0/NAND4_in[0] ,
         \SB1_2_12/Component_Function_1/NAND4_in[3] ,
         \SB1_2_12/Component_Function_1/NAND4_in[2] ,
         \SB1_2_12/Component_Function_1/NAND4_in[1] ,
         \SB1_2_12/Component_Function_1/NAND4_in[0] ,
         \SB1_2_12/Component_Function_5/NAND4_in[2] ,
         \SB1_2_12/Component_Function_5/NAND4_in[1] ,
         \SB1_2_12/Component_Function_5/NAND4_in[0] ,
         \SB1_2_13/Component_Function_0/NAND4_in[3] ,
         \SB1_2_13/Component_Function_0/NAND4_in[2] ,
         \SB1_2_13/Component_Function_0/NAND4_in[1] ,
         \SB1_2_13/Component_Function_0/NAND4_in[0] ,
         \SB1_2_13/Component_Function_1/NAND4_in[3] ,
         \SB1_2_13/Component_Function_1/NAND4_in[2] ,
         \SB1_2_13/Component_Function_1/NAND4_in[1] ,
         \SB1_2_13/Component_Function_1/NAND4_in[0] ,
         \SB1_2_13/Component_Function_5/NAND4_in[3] ,
         \SB1_2_13/Component_Function_5/NAND4_in[1] ,
         \SB1_2_13/Component_Function_5/NAND4_in[0] ,
         \SB1_2_14/Component_Function_0/NAND4_in[3] ,
         \SB1_2_14/Component_Function_0/NAND4_in[2] ,
         \SB1_2_14/Component_Function_0/NAND4_in[1] ,
         \SB1_2_14/Component_Function_0/NAND4_in[0] ,
         \SB1_2_14/Component_Function_1/NAND4_in[3] ,
         \SB1_2_14/Component_Function_1/NAND4_in[2] ,
         \SB1_2_14/Component_Function_1/NAND4_in[1] ,
         \SB1_2_14/Component_Function_1/NAND4_in[0] ,
         \SB1_2_14/Component_Function_5/NAND4_in[3] ,
         \SB1_2_14/Component_Function_5/NAND4_in[1] ,
         \SB1_2_14/Component_Function_5/NAND4_in[0] ,
         \SB1_2_15/Component_Function_0/NAND4_in[3] ,
         \SB1_2_15/Component_Function_0/NAND4_in[2] ,
         \SB1_2_15/Component_Function_0/NAND4_in[1] ,
         \SB1_2_15/Component_Function_0/NAND4_in[0] ,
         \SB1_2_15/Component_Function_1/NAND4_in[3] ,
         \SB1_2_15/Component_Function_1/NAND4_in[2] ,
         \SB1_2_15/Component_Function_1/NAND4_in[1] ,
         \SB1_2_15/Component_Function_1/NAND4_in[0] ,
         \SB1_2_15/Component_Function_5/NAND4_in[3] ,
         \SB1_2_15/Component_Function_5/NAND4_in[1] ,
         \SB1_2_15/Component_Function_5/NAND4_in[0] ,
         \SB1_2_16/Component_Function_0/NAND4_in[3] ,
         \SB1_2_16/Component_Function_0/NAND4_in[2] ,
         \SB1_2_16/Component_Function_0/NAND4_in[1] ,
         \SB1_2_16/Component_Function_0/NAND4_in[0] ,
         \SB1_2_16/Component_Function_1/NAND4_in[3] ,
         \SB1_2_16/Component_Function_1/NAND4_in[2] ,
         \SB1_2_16/Component_Function_1/NAND4_in[1] ,
         \SB1_2_16/Component_Function_1/NAND4_in[0] ,
         \SB1_2_16/Component_Function_5/NAND4_in[3] ,
         \SB1_2_16/Component_Function_5/NAND4_in[1] ,
         \SB1_2_16/Component_Function_5/NAND4_in[0] ,
         \SB1_2_17/Component_Function_0/NAND4_in[3] ,
         \SB1_2_17/Component_Function_0/NAND4_in[2] ,
         \SB1_2_17/Component_Function_0/NAND4_in[1] ,
         \SB1_2_17/Component_Function_0/NAND4_in[0] ,
         \SB1_2_17/Component_Function_1/NAND4_in[3] ,
         \SB1_2_17/Component_Function_1/NAND4_in[2] ,
         \SB1_2_17/Component_Function_1/NAND4_in[1] ,
         \SB1_2_17/Component_Function_1/NAND4_in[0] ,
         \SB1_2_17/Component_Function_5/NAND4_in[3] ,
         \SB1_2_17/Component_Function_5/NAND4_in[1] ,
         \SB1_2_17/Component_Function_5/NAND4_in[0] ,
         \SB1_2_18/Component_Function_0/NAND4_in[3] ,
         \SB1_2_18/Component_Function_0/NAND4_in[2] ,
         \SB1_2_18/Component_Function_0/NAND4_in[1] ,
         \SB1_2_18/Component_Function_0/NAND4_in[0] ,
         \SB1_2_18/Component_Function_1/NAND4_in[3] ,
         \SB1_2_18/Component_Function_1/NAND4_in[2] ,
         \SB1_2_18/Component_Function_1/NAND4_in[1] ,
         \SB1_2_18/Component_Function_1/NAND4_in[0] ,
         \SB1_2_18/Component_Function_5/NAND4_in[3] ,
         \SB1_2_18/Component_Function_5/NAND4_in[1] ,
         \SB1_2_18/Component_Function_5/NAND4_in[0] ,
         \SB1_2_19/Component_Function_0/NAND4_in[3] ,
         \SB1_2_19/Component_Function_0/NAND4_in[2] ,
         \SB1_2_19/Component_Function_0/NAND4_in[1] ,
         \SB1_2_19/Component_Function_0/NAND4_in[0] ,
         \SB1_2_19/Component_Function_1/NAND4_in[3] ,
         \SB1_2_19/Component_Function_1/NAND4_in[2] ,
         \SB1_2_19/Component_Function_1/NAND4_in[1] ,
         \SB1_2_19/Component_Function_1/NAND4_in[0] ,
         \SB1_2_19/Component_Function_5/NAND4_in[3] ,
         \SB1_2_19/Component_Function_5/NAND4_in[1] ,
         \SB1_2_19/Component_Function_5/NAND4_in[0] ,
         \SB1_2_20/Component_Function_0/NAND4_in[3] ,
         \SB1_2_20/Component_Function_0/NAND4_in[2] ,
         \SB1_2_20/Component_Function_0/NAND4_in[1] ,
         \SB1_2_20/Component_Function_0/NAND4_in[0] ,
         \SB1_2_20/Component_Function_1/NAND4_in[3] ,
         \SB1_2_20/Component_Function_1/NAND4_in[2] ,
         \SB1_2_20/Component_Function_1/NAND4_in[1] ,
         \SB1_2_20/Component_Function_1/NAND4_in[0] ,
         \SB1_2_20/Component_Function_5/NAND4_in[3] ,
         \SB1_2_20/Component_Function_5/NAND4_in[1] ,
         \SB1_2_20/Component_Function_5/NAND4_in[0] ,
         \SB1_2_21/Component_Function_0/NAND4_in[3] ,
         \SB1_2_21/Component_Function_0/NAND4_in[2] ,
         \SB1_2_21/Component_Function_0/NAND4_in[1] ,
         \SB1_2_21/Component_Function_0/NAND4_in[0] ,
         \SB1_2_21/Component_Function_1/NAND4_in[3] ,
         \SB1_2_21/Component_Function_1/NAND4_in[2] ,
         \SB1_2_21/Component_Function_1/NAND4_in[1] ,
         \SB1_2_21/Component_Function_1/NAND4_in[0] ,
         \SB1_2_21/Component_Function_5/NAND4_in[3] ,
         \SB1_2_21/Component_Function_5/NAND4_in[1] ,
         \SB1_2_21/Component_Function_5/NAND4_in[0] ,
         \SB1_2_22/Component_Function_0/NAND4_in[3] ,
         \SB1_2_22/Component_Function_0/NAND4_in[2] ,
         \SB1_2_22/Component_Function_0/NAND4_in[1] ,
         \SB1_2_22/Component_Function_0/NAND4_in[0] ,
         \SB1_2_22/Component_Function_1/NAND4_in[3] ,
         \SB1_2_22/Component_Function_1/NAND4_in[2] ,
         \SB1_2_22/Component_Function_1/NAND4_in[1] ,
         \SB1_2_22/Component_Function_1/NAND4_in[0] ,
         \SB1_2_22/Component_Function_5/NAND4_in[3] ,
         \SB1_2_22/Component_Function_5/NAND4_in[1] ,
         \SB1_2_22/Component_Function_5/NAND4_in[0] ,
         \SB1_2_23/Component_Function_0/NAND4_in[3] ,
         \SB1_2_23/Component_Function_0/NAND4_in[2] ,
         \SB1_2_23/Component_Function_0/NAND4_in[1] ,
         \SB1_2_23/Component_Function_0/NAND4_in[0] ,
         \SB1_2_23/Component_Function_1/NAND4_in[3] ,
         \SB1_2_23/Component_Function_1/NAND4_in[2] ,
         \SB1_2_23/Component_Function_1/NAND4_in[1] ,
         \SB1_2_23/Component_Function_1/NAND4_in[0] ,
         \SB1_2_23/Component_Function_5/NAND4_in[3] ,
         \SB1_2_23/Component_Function_5/NAND4_in[1] ,
         \SB1_2_23/Component_Function_5/NAND4_in[0] ,
         \SB1_2_24/Component_Function_0/NAND4_in[3] ,
         \SB1_2_24/Component_Function_0/NAND4_in[2] ,
         \SB1_2_24/Component_Function_0/NAND4_in[1] ,
         \SB1_2_24/Component_Function_0/NAND4_in[0] ,
         \SB1_2_24/Component_Function_1/NAND4_in[3] ,
         \SB1_2_24/Component_Function_1/NAND4_in[2] ,
         \SB1_2_24/Component_Function_1/NAND4_in[1] ,
         \SB1_2_24/Component_Function_1/NAND4_in[0] ,
         \SB1_2_24/Component_Function_5/NAND4_in[3] ,
         \SB1_2_24/Component_Function_5/NAND4_in[1] ,
         \SB1_2_24/Component_Function_5/NAND4_in[0] ,
         \SB1_2_25/Component_Function_0/NAND4_in[3] ,
         \SB1_2_25/Component_Function_0/NAND4_in[2] ,
         \SB1_2_25/Component_Function_0/NAND4_in[1] ,
         \SB1_2_25/Component_Function_0/NAND4_in[0] ,
         \SB1_2_25/Component_Function_1/NAND4_in[3] ,
         \SB1_2_25/Component_Function_1/NAND4_in[2] ,
         \SB1_2_25/Component_Function_1/NAND4_in[1] ,
         \SB1_2_25/Component_Function_1/NAND4_in[0] ,
         \SB1_2_25/Component_Function_5/NAND4_in[3] ,
         \SB1_2_25/Component_Function_5/NAND4_in[1] ,
         \SB1_2_25/Component_Function_5/NAND4_in[0] ,
         \SB1_2_26/Component_Function_0/NAND4_in[3] ,
         \SB1_2_26/Component_Function_0/NAND4_in[1] ,
         \SB1_2_26/Component_Function_0/NAND4_in[0] ,
         \SB1_2_26/Component_Function_1/NAND4_in[3] ,
         \SB1_2_26/Component_Function_1/NAND4_in[2] ,
         \SB1_2_26/Component_Function_1/NAND4_in[1] ,
         \SB1_2_26/Component_Function_1/NAND4_in[0] ,
         \SB1_2_26/Component_Function_5/NAND4_in[3] ,
         \SB1_2_26/Component_Function_5/NAND4_in[1] ,
         \SB1_2_26/Component_Function_5/NAND4_in[0] ,
         \SB1_2_27/Component_Function_0/NAND4_in[3] ,
         \SB1_2_27/Component_Function_0/NAND4_in[2] ,
         \SB1_2_27/Component_Function_0/NAND4_in[1] ,
         \SB1_2_27/Component_Function_0/NAND4_in[0] ,
         \SB1_2_27/Component_Function_1/NAND4_in[3] ,
         \SB1_2_27/Component_Function_1/NAND4_in[2] ,
         \SB1_2_27/Component_Function_1/NAND4_in[1] ,
         \SB1_2_27/Component_Function_1/NAND4_in[0] ,
         \SB1_2_27/Component_Function_5/NAND4_in[3] ,
         \SB1_2_27/Component_Function_5/NAND4_in[1] ,
         \SB1_2_27/Component_Function_5/NAND4_in[0] ,
         \SB1_2_28/Component_Function_0/NAND4_in[3] ,
         \SB1_2_28/Component_Function_0/NAND4_in[2] ,
         \SB1_2_28/Component_Function_0/NAND4_in[1] ,
         \SB1_2_28/Component_Function_0/NAND4_in[0] ,
         \SB1_2_28/Component_Function_1/NAND4_in[3] ,
         \SB1_2_28/Component_Function_1/NAND4_in[2] ,
         \SB1_2_28/Component_Function_1/NAND4_in[1] ,
         \SB1_2_28/Component_Function_1/NAND4_in[0] ,
         \SB1_2_28/Component_Function_5/NAND4_in[3] ,
         \SB1_2_28/Component_Function_5/NAND4_in[1] ,
         \SB1_2_28/Component_Function_5/NAND4_in[0] ,
         \SB1_2_29/Component_Function_0/NAND4_in[3] ,
         \SB1_2_29/Component_Function_0/NAND4_in[2] ,
         \SB1_2_29/Component_Function_0/NAND4_in[1] ,
         \SB1_2_29/Component_Function_0/NAND4_in[0] ,
         \SB1_2_29/Component_Function_1/NAND4_in[3] ,
         \SB1_2_29/Component_Function_1/NAND4_in[2] ,
         \SB1_2_29/Component_Function_1/NAND4_in[1] ,
         \SB1_2_29/Component_Function_1/NAND4_in[0] ,
         \SB1_2_29/Component_Function_5/NAND4_in[3] ,
         \SB1_2_29/Component_Function_5/NAND4_in[1] ,
         \SB1_2_29/Component_Function_5/NAND4_in[0] ,
         \SB1_2_30/Component_Function_0/NAND4_in[3] ,
         \SB1_2_30/Component_Function_0/NAND4_in[2] ,
         \SB1_2_30/Component_Function_0/NAND4_in[1] ,
         \SB1_2_30/Component_Function_0/NAND4_in[0] ,
         \SB1_2_30/Component_Function_1/NAND4_in[3] ,
         \SB1_2_30/Component_Function_1/NAND4_in[2] ,
         \SB1_2_30/Component_Function_1/NAND4_in[1] ,
         \SB1_2_30/Component_Function_1/NAND4_in[0] ,
         \SB1_2_30/Component_Function_5/NAND4_in[3] ,
         \SB1_2_30/Component_Function_5/NAND4_in[1] ,
         \SB1_2_30/Component_Function_5/NAND4_in[0] ,
         \SB1_2_31/Component_Function_0/NAND4_in[3] ,
         \SB1_2_31/Component_Function_0/NAND4_in[2] ,
         \SB1_2_31/Component_Function_0/NAND4_in[1] ,
         \SB1_2_31/Component_Function_0/NAND4_in[0] ,
         \SB1_2_31/Component_Function_1/NAND4_in[2] ,
         \SB1_2_31/Component_Function_1/NAND4_in[1] ,
         \SB1_2_31/Component_Function_1/NAND4_in[0] ,
         \SB1_2_31/Component_Function_5/NAND4_in[3] ,
         \SB1_2_31/Component_Function_5/NAND4_in[1] ,
         \SB1_2_31/Component_Function_5/NAND4_in[0] ,
         \SB2_2_0/Component_Function_0/NAND4_in[3] ,
         \SB2_2_0/Component_Function_0/NAND4_in[2] ,
         \SB2_2_0/Component_Function_0/NAND4_in[1] ,
         \SB2_2_0/Component_Function_0/NAND4_in[0] ,
         \SB2_2_0/Component_Function_1/NAND4_in[3] ,
         \SB2_2_0/Component_Function_1/NAND4_in[2] ,
         \SB2_2_0/Component_Function_1/NAND4_in[1] ,
         \SB2_2_0/Component_Function_1/NAND4_in[0] ,
         \SB2_2_0/Component_Function_5/NAND4_in[3] ,
         \SB2_2_0/Component_Function_5/NAND4_in[2] ,
         \SB2_2_0/Component_Function_5/NAND4_in[1] ,
         \SB2_2_0/Component_Function_5/NAND4_in[0] ,
         \SB2_2_1/Component_Function_0/NAND4_in[3] ,
         \SB2_2_1/Component_Function_0/NAND4_in[2] ,
         \SB2_2_1/Component_Function_0/NAND4_in[1] ,
         \SB2_2_1/Component_Function_0/NAND4_in[0] ,
         \SB2_2_1/Component_Function_1/NAND4_in[2] ,
         \SB2_2_1/Component_Function_1/NAND4_in[1] ,
         \SB2_2_1/Component_Function_1/NAND4_in[0] ,
         \SB2_2_1/Component_Function_5/NAND4_in[3] ,
         \SB2_2_1/Component_Function_5/NAND4_in[2] ,
         \SB2_2_1/Component_Function_5/NAND4_in[1] ,
         \SB2_2_1/Component_Function_5/NAND4_in[0] ,
         \SB2_2_2/Component_Function_0/NAND4_in[3] ,
         \SB2_2_2/Component_Function_0/NAND4_in[2] ,
         \SB2_2_2/Component_Function_0/NAND4_in[1] ,
         \SB2_2_2/Component_Function_0/NAND4_in[0] ,
         \SB2_2_2/Component_Function_1/NAND4_in[3] ,
         \SB2_2_2/Component_Function_1/NAND4_in[2] ,
         \SB2_2_2/Component_Function_1/NAND4_in[1] ,
         \SB2_2_2/Component_Function_1/NAND4_in[0] ,
         \SB2_2_2/Component_Function_5/NAND4_in[3] ,
         \SB2_2_2/Component_Function_5/NAND4_in[2] ,
         \SB2_2_2/Component_Function_5/NAND4_in[1] ,
         \SB2_2_3/Component_Function_0/NAND4_in[3] ,
         \SB2_2_3/Component_Function_0/NAND4_in[2] ,
         \SB2_2_3/Component_Function_0/NAND4_in[1] ,
         \SB2_2_3/Component_Function_0/NAND4_in[0] ,
         \SB2_2_3/Component_Function_1/NAND4_in[3] ,
         \SB2_2_3/Component_Function_1/NAND4_in[2] ,
         \SB2_2_3/Component_Function_1/NAND4_in[1] ,
         \SB2_2_3/Component_Function_1/NAND4_in[0] ,
         \SB2_2_3/Component_Function_5/NAND4_in[3] ,
         \SB2_2_3/Component_Function_5/NAND4_in[2] ,
         \SB2_2_3/Component_Function_5/NAND4_in[1] ,
         \SB2_2_3/Component_Function_5/NAND4_in[0] ,
         \SB2_2_4/Component_Function_0/NAND4_in[3] ,
         \SB2_2_4/Component_Function_0/NAND4_in[2] ,
         \SB2_2_4/Component_Function_0/NAND4_in[1] ,
         \SB2_2_4/Component_Function_0/NAND4_in[0] ,
         \SB2_2_4/Component_Function_1/NAND4_in[3] ,
         \SB2_2_4/Component_Function_1/NAND4_in[2] ,
         \SB2_2_4/Component_Function_1/NAND4_in[1] ,
         \SB2_2_4/Component_Function_1/NAND4_in[0] ,
         \SB2_2_4/Component_Function_5/NAND4_in[3] ,
         \SB2_2_4/Component_Function_5/NAND4_in[1] ,
         \SB2_2_4/Component_Function_5/NAND4_in[0] ,
         \SB2_2_5/Component_Function_0/NAND4_in[3] ,
         \SB2_2_5/Component_Function_0/NAND4_in[2] ,
         \SB2_2_5/Component_Function_0/NAND4_in[1] ,
         \SB2_2_5/Component_Function_0/NAND4_in[0] ,
         \SB2_2_5/Component_Function_1/NAND4_in[3] ,
         \SB2_2_5/Component_Function_1/NAND4_in[2] ,
         \SB2_2_5/Component_Function_1/NAND4_in[1] ,
         \SB2_2_5/Component_Function_1/NAND4_in[0] ,
         \SB2_2_5/Component_Function_5/NAND4_in[3] ,
         \SB2_2_5/Component_Function_5/NAND4_in[2] ,
         \SB2_2_5/Component_Function_5/NAND4_in[1] ,
         \SB2_2_5/Component_Function_5/NAND4_in[0] ,
         \SB2_2_6/Component_Function_0/NAND4_in[3] ,
         \SB2_2_6/Component_Function_0/NAND4_in[2] ,
         \SB2_2_6/Component_Function_0/NAND4_in[1] ,
         \SB2_2_6/Component_Function_0/NAND4_in[0] ,
         \SB2_2_6/Component_Function_1/NAND4_in[3] ,
         \SB2_2_6/Component_Function_1/NAND4_in[2] ,
         \SB2_2_6/Component_Function_1/NAND4_in[1] ,
         \SB2_2_6/Component_Function_1/NAND4_in[0] ,
         \SB2_2_6/Component_Function_5/NAND4_in[3] ,
         \SB2_2_6/Component_Function_5/NAND4_in[2] ,
         \SB2_2_6/Component_Function_5/NAND4_in[1] ,
         \SB2_2_6/Component_Function_5/NAND4_in[0] ,
         \SB2_2_7/Component_Function_0/NAND4_in[3] ,
         \SB2_2_7/Component_Function_0/NAND4_in[2] ,
         \SB2_2_7/Component_Function_0/NAND4_in[1] ,
         \SB2_2_7/Component_Function_0/NAND4_in[0] ,
         \SB2_2_7/Component_Function_1/NAND4_in[3] ,
         \SB2_2_7/Component_Function_1/NAND4_in[2] ,
         \SB2_2_7/Component_Function_1/NAND4_in[1] ,
         \SB2_2_7/Component_Function_1/NAND4_in[0] ,
         \SB2_2_7/Component_Function_5/NAND4_in[3] ,
         \SB2_2_7/Component_Function_5/NAND4_in[2] ,
         \SB2_2_7/Component_Function_5/NAND4_in[1] ,
         \SB2_2_7/Component_Function_5/NAND4_in[0] ,
         \SB2_2_8/Component_Function_0/NAND4_in[3] ,
         \SB2_2_8/Component_Function_0/NAND4_in[2] ,
         \SB2_2_8/Component_Function_0/NAND4_in[1] ,
         \SB2_2_8/Component_Function_0/NAND4_in[0] ,
         \SB2_2_8/Component_Function_1/NAND4_in[3] ,
         \SB2_2_8/Component_Function_1/NAND4_in[2] ,
         \SB2_2_8/Component_Function_1/NAND4_in[1] ,
         \SB2_2_8/Component_Function_1/NAND4_in[0] ,
         \SB2_2_8/Component_Function_5/NAND4_in[3] ,
         \SB2_2_8/Component_Function_5/NAND4_in[2] ,
         \SB2_2_8/Component_Function_5/NAND4_in[1] ,
         \SB2_2_8/Component_Function_5/NAND4_in[0] ,
         \SB2_2_9/Component_Function_0/NAND4_in[3] ,
         \SB2_2_9/Component_Function_0/NAND4_in[2] ,
         \SB2_2_9/Component_Function_0/NAND4_in[1] ,
         \SB2_2_9/Component_Function_0/NAND4_in[0] ,
         \SB2_2_9/Component_Function_1/NAND4_in[3] ,
         \SB2_2_9/Component_Function_1/NAND4_in[2] ,
         \SB2_2_9/Component_Function_1/NAND4_in[1] ,
         \SB2_2_9/Component_Function_1/NAND4_in[0] ,
         \SB2_2_9/Component_Function_5/NAND4_in[3] ,
         \SB2_2_9/Component_Function_5/NAND4_in[2] ,
         \SB2_2_9/Component_Function_5/NAND4_in[1] ,
         \SB2_2_10/Component_Function_0/NAND4_in[3] ,
         \SB2_2_10/Component_Function_0/NAND4_in[2] ,
         \SB2_2_10/Component_Function_0/NAND4_in[1] ,
         \SB2_2_10/Component_Function_0/NAND4_in[0] ,
         \SB2_2_10/Component_Function_1/NAND4_in[2] ,
         \SB2_2_10/Component_Function_1/NAND4_in[1] ,
         \SB2_2_10/Component_Function_1/NAND4_in[0] ,
         \SB2_2_10/Component_Function_5/NAND4_in[3] ,
         \SB2_2_10/Component_Function_5/NAND4_in[2] ,
         \SB2_2_10/Component_Function_5/NAND4_in[1] ,
         \SB2_2_10/Component_Function_5/NAND4_in[0] ,
         \SB2_2_11/Component_Function_0/NAND4_in[3] ,
         \SB2_2_11/Component_Function_0/NAND4_in[2] ,
         \SB2_2_11/Component_Function_0/NAND4_in[1] ,
         \SB2_2_11/Component_Function_0/NAND4_in[0] ,
         \SB2_2_11/Component_Function_1/NAND4_in[3] ,
         \SB2_2_11/Component_Function_1/NAND4_in[2] ,
         \SB2_2_11/Component_Function_1/NAND4_in[1] ,
         \SB2_2_11/Component_Function_1/NAND4_in[0] ,
         \SB2_2_11/Component_Function_5/NAND4_in[3] ,
         \SB2_2_11/Component_Function_5/NAND4_in[2] ,
         \SB2_2_11/Component_Function_5/NAND4_in[1] ,
         \SB2_2_12/Component_Function_0/NAND4_in[2] ,
         \SB2_2_12/Component_Function_0/NAND4_in[1] ,
         \SB2_2_12/Component_Function_0/NAND4_in[0] ,
         \SB2_2_12/Component_Function_1/NAND4_in[3] ,
         \SB2_2_12/Component_Function_1/NAND4_in[2] ,
         \SB2_2_12/Component_Function_1/NAND4_in[1] ,
         \SB2_2_12/Component_Function_1/NAND4_in[0] ,
         \SB2_2_12/Component_Function_5/NAND4_in[3] ,
         \SB2_2_12/Component_Function_5/NAND4_in[2] ,
         \SB2_2_12/Component_Function_5/NAND4_in[1] ,
         \SB2_2_12/Component_Function_5/NAND4_in[0] ,
         \SB2_2_13/Component_Function_0/NAND4_in[3] ,
         \SB2_2_13/Component_Function_0/NAND4_in[2] ,
         \SB2_2_13/Component_Function_0/NAND4_in[1] ,
         \SB2_2_13/Component_Function_0/NAND4_in[0] ,
         \SB2_2_13/Component_Function_1/NAND4_in[3] ,
         \SB2_2_13/Component_Function_1/NAND4_in[2] ,
         \SB2_2_13/Component_Function_1/NAND4_in[1] ,
         \SB2_2_13/Component_Function_1/NAND4_in[0] ,
         \SB2_2_13/Component_Function_5/NAND4_in[3] ,
         \SB2_2_13/Component_Function_5/NAND4_in[2] ,
         \SB2_2_13/Component_Function_5/NAND4_in[1] ,
         \SB2_2_14/Component_Function_0/NAND4_in[3] ,
         \SB2_2_14/Component_Function_0/NAND4_in[2] ,
         \SB2_2_14/Component_Function_0/NAND4_in[1] ,
         \SB2_2_14/Component_Function_0/NAND4_in[0] ,
         \SB2_2_14/Component_Function_1/NAND4_in[2] ,
         \SB2_2_14/Component_Function_1/NAND4_in[1] ,
         \SB2_2_14/Component_Function_1/NAND4_in[0] ,
         \SB2_2_14/Component_Function_5/NAND4_in[2] ,
         \SB2_2_14/Component_Function_5/NAND4_in[1] ,
         \SB2_2_14/Component_Function_5/NAND4_in[0] ,
         \SB2_2_15/Component_Function_0/NAND4_in[3] ,
         \SB2_2_15/Component_Function_0/NAND4_in[2] ,
         \SB2_2_15/Component_Function_0/NAND4_in[1] ,
         \SB2_2_15/Component_Function_0/NAND4_in[0] ,
         \SB2_2_15/Component_Function_1/NAND4_in[3] ,
         \SB2_2_15/Component_Function_1/NAND4_in[2] ,
         \SB2_2_15/Component_Function_1/NAND4_in[1] ,
         \SB2_2_15/Component_Function_1/NAND4_in[0] ,
         \SB2_2_15/Component_Function_5/NAND4_in[3] ,
         \SB2_2_15/Component_Function_5/NAND4_in[2] ,
         \SB2_2_15/Component_Function_5/NAND4_in[1] ,
         \SB2_2_15/Component_Function_5/NAND4_in[0] ,
         \SB2_2_16/Component_Function_0/NAND4_in[3] ,
         \SB2_2_16/Component_Function_0/NAND4_in[2] ,
         \SB2_2_16/Component_Function_0/NAND4_in[1] ,
         \SB2_2_16/Component_Function_0/NAND4_in[0] ,
         \SB2_2_16/Component_Function_1/NAND4_in[3] ,
         \SB2_2_16/Component_Function_1/NAND4_in[2] ,
         \SB2_2_16/Component_Function_1/NAND4_in[1] ,
         \SB2_2_16/Component_Function_1/NAND4_in[0] ,
         \SB2_2_16/Component_Function_5/NAND4_in[3] ,
         \SB2_2_16/Component_Function_5/NAND4_in[1] ,
         \SB2_2_16/Component_Function_5/NAND4_in[0] ,
         \SB2_2_17/Component_Function_0/NAND4_in[3] ,
         \SB2_2_17/Component_Function_0/NAND4_in[2] ,
         \SB2_2_17/Component_Function_0/NAND4_in[1] ,
         \SB2_2_17/Component_Function_0/NAND4_in[0] ,
         \SB2_2_17/Component_Function_1/NAND4_in[3] ,
         \SB2_2_17/Component_Function_1/NAND4_in[2] ,
         \SB2_2_17/Component_Function_1/NAND4_in[1] ,
         \SB2_2_17/Component_Function_1/NAND4_in[0] ,
         \SB2_2_17/Component_Function_5/NAND4_in[3] ,
         \SB2_2_17/Component_Function_5/NAND4_in[2] ,
         \SB2_2_17/Component_Function_5/NAND4_in[1] ,
         \SB2_2_17/Component_Function_5/NAND4_in[0] ,
         \SB2_2_18/Component_Function_0/NAND4_in[3] ,
         \SB2_2_18/Component_Function_0/NAND4_in[2] ,
         \SB2_2_18/Component_Function_0/NAND4_in[1] ,
         \SB2_2_18/Component_Function_0/NAND4_in[0] ,
         \SB2_2_18/Component_Function_1/NAND4_in[3] ,
         \SB2_2_18/Component_Function_1/NAND4_in[1] ,
         \SB2_2_18/Component_Function_1/NAND4_in[0] ,
         \SB2_2_18/Component_Function_5/NAND4_in[2] ,
         \SB2_2_18/Component_Function_5/NAND4_in[1] ,
         \SB2_2_18/Component_Function_5/NAND4_in[0] ,
         \SB2_2_19/Component_Function_0/NAND4_in[3] ,
         \SB2_2_19/Component_Function_0/NAND4_in[2] ,
         \SB2_2_19/Component_Function_0/NAND4_in[1] ,
         \SB2_2_19/Component_Function_0/NAND4_in[0] ,
         \SB2_2_19/Component_Function_1/NAND4_in[3] ,
         \SB2_2_19/Component_Function_1/NAND4_in[2] ,
         \SB2_2_19/Component_Function_1/NAND4_in[1] ,
         \SB2_2_19/Component_Function_1/NAND4_in[0] ,
         \SB2_2_19/Component_Function_5/NAND4_in[3] ,
         \SB2_2_19/Component_Function_5/NAND4_in[2] ,
         \SB2_2_19/Component_Function_5/NAND4_in[1] ,
         \SB2_2_19/Component_Function_5/NAND4_in[0] ,
         \SB2_2_20/Component_Function_0/NAND4_in[3] ,
         \SB2_2_20/Component_Function_0/NAND4_in[2] ,
         \SB2_2_20/Component_Function_0/NAND4_in[1] ,
         \SB2_2_20/Component_Function_0/NAND4_in[0] ,
         \SB2_2_20/Component_Function_1/NAND4_in[3] ,
         \SB2_2_20/Component_Function_1/NAND4_in[2] ,
         \SB2_2_20/Component_Function_1/NAND4_in[1] ,
         \SB2_2_20/Component_Function_1/NAND4_in[0] ,
         \SB2_2_20/Component_Function_5/NAND4_in[3] ,
         \SB2_2_20/Component_Function_5/NAND4_in[2] ,
         \SB2_2_20/Component_Function_5/NAND4_in[1] ,
         \SB2_2_20/Component_Function_5/NAND4_in[0] ,
         \SB2_2_21/Component_Function_0/NAND4_in[3] ,
         \SB2_2_21/Component_Function_0/NAND4_in[2] ,
         \SB2_2_21/Component_Function_0/NAND4_in[1] ,
         \SB2_2_21/Component_Function_0/NAND4_in[0] ,
         \SB2_2_21/Component_Function_1/NAND4_in[3] ,
         \SB2_2_21/Component_Function_1/NAND4_in[2] ,
         \SB2_2_21/Component_Function_1/NAND4_in[1] ,
         \SB2_2_21/Component_Function_1/NAND4_in[0] ,
         \SB2_2_21/Component_Function_5/NAND4_in[3] ,
         \SB2_2_21/Component_Function_5/NAND4_in[2] ,
         \SB2_2_21/Component_Function_5/NAND4_in[1] ,
         \SB2_2_21/Component_Function_5/NAND4_in[0] ,
         \SB2_2_22/Component_Function_0/NAND4_in[3] ,
         \SB2_2_22/Component_Function_0/NAND4_in[2] ,
         \SB2_2_22/Component_Function_0/NAND4_in[1] ,
         \SB2_2_22/Component_Function_0/NAND4_in[0] ,
         \SB2_2_22/Component_Function_1/NAND4_in[3] ,
         \SB2_2_22/Component_Function_1/NAND4_in[2] ,
         \SB2_2_22/Component_Function_1/NAND4_in[1] ,
         \SB2_2_22/Component_Function_1/NAND4_in[0] ,
         \SB2_2_22/Component_Function_5/NAND4_in[3] ,
         \SB2_2_22/Component_Function_5/NAND4_in[2] ,
         \SB2_2_22/Component_Function_5/NAND4_in[1] ,
         \SB2_2_22/Component_Function_5/NAND4_in[0] ,
         \SB2_2_23/Component_Function_0/NAND4_in[3] ,
         \SB2_2_23/Component_Function_0/NAND4_in[2] ,
         \SB2_2_23/Component_Function_0/NAND4_in[1] ,
         \SB2_2_23/Component_Function_0/NAND4_in[0] ,
         \SB2_2_23/Component_Function_1/NAND4_in[3] ,
         \SB2_2_23/Component_Function_1/NAND4_in[2] ,
         \SB2_2_23/Component_Function_1/NAND4_in[1] ,
         \SB2_2_23/Component_Function_1/NAND4_in[0] ,
         \SB2_2_23/Component_Function_5/NAND4_in[3] ,
         \SB2_2_23/Component_Function_5/NAND4_in[1] ,
         \SB2_2_23/Component_Function_5/NAND4_in[0] ,
         \SB2_2_24/Component_Function_0/NAND4_in[2] ,
         \SB2_2_24/Component_Function_0/NAND4_in[1] ,
         \SB2_2_24/Component_Function_0/NAND4_in[0] ,
         \SB2_2_24/Component_Function_1/NAND4_in[3] ,
         \SB2_2_24/Component_Function_1/NAND4_in[2] ,
         \SB2_2_24/Component_Function_1/NAND4_in[1] ,
         \SB2_2_24/Component_Function_1/NAND4_in[0] ,
         \SB2_2_24/Component_Function_5/NAND4_in[3] ,
         \SB2_2_24/Component_Function_5/NAND4_in[2] ,
         \SB2_2_24/Component_Function_5/NAND4_in[1] ,
         \SB2_2_24/Component_Function_5/NAND4_in[0] ,
         \SB2_2_25/Component_Function_0/NAND4_in[3] ,
         \SB2_2_25/Component_Function_0/NAND4_in[2] ,
         \SB2_2_25/Component_Function_0/NAND4_in[1] ,
         \SB2_2_25/Component_Function_0/NAND4_in[0] ,
         \SB2_2_25/Component_Function_1/NAND4_in[3] ,
         \SB2_2_25/Component_Function_1/NAND4_in[2] ,
         \SB2_2_25/Component_Function_1/NAND4_in[1] ,
         \SB2_2_25/Component_Function_1/NAND4_in[0] ,
         \SB2_2_25/Component_Function_5/NAND4_in[3] ,
         \SB2_2_25/Component_Function_5/NAND4_in[2] ,
         \SB2_2_25/Component_Function_5/NAND4_in[1] ,
         \SB2_2_25/Component_Function_5/NAND4_in[0] ,
         \SB2_2_26/Component_Function_0/NAND4_in[3] ,
         \SB2_2_26/Component_Function_0/NAND4_in[2] ,
         \SB2_2_26/Component_Function_0/NAND4_in[1] ,
         \SB2_2_26/Component_Function_0/NAND4_in[0] ,
         \SB2_2_26/Component_Function_1/NAND4_in[3] ,
         \SB2_2_26/Component_Function_1/NAND4_in[2] ,
         \SB2_2_26/Component_Function_1/NAND4_in[1] ,
         \SB2_2_26/Component_Function_1/NAND4_in[0] ,
         \SB2_2_26/Component_Function_5/NAND4_in[3] ,
         \SB2_2_26/Component_Function_5/NAND4_in[2] ,
         \SB2_2_26/Component_Function_5/NAND4_in[1] ,
         \SB2_2_27/Component_Function_0/NAND4_in[3] ,
         \SB2_2_27/Component_Function_0/NAND4_in[2] ,
         \SB2_2_27/Component_Function_0/NAND4_in[1] ,
         \SB2_2_27/Component_Function_0/NAND4_in[0] ,
         \SB2_2_27/Component_Function_1/NAND4_in[3] ,
         \SB2_2_27/Component_Function_1/NAND4_in[2] ,
         \SB2_2_27/Component_Function_1/NAND4_in[1] ,
         \SB2_2_27/Component_Function_1/NAND4_in[0] ,
         \SB2_2_27/Component_Function_5/NAND4_in[3] ,
         \SB2_2_27/Component_Function_5/NAND4_in[2] ,
         \SB2_2_27/Component_Function_5/NAND4_in[1] ,
         \SB2_2_27/Component_Function_5/NAND4_in[0] ,
         \SB2_2_28/Component_Function_0/NAND4_in[3] ,
         \SB2_2_28/Component_Function_0/NAND4_in[2] ,
         \SB2_2_28/Component_Function_0/NAND4_in[1] ,
         \SB2_2_28/Component_Function_0/NAND4_in[0] ,
         \SB2_2_28/Component_Function_1/NAND4_in[3] ,
         \SB2_2_28/Component_Function_1/NAND4_in[2] ,
         \SB2_2_28/Component_Function_1/NAND4_in[1] ,
         \SB2_2_28/Component_Function_1/NAND4_in[0] ,
         \SB2_2_28/Component_Function_5/NAND4_in[3] ,
         \SB2_2_28/Component_Function_5/NAND4_in[2] ,
         \SB2_2_28/Component_Function_5/NAND4_in[1] ,
         \SB2_2_28/Component_Function_5/NAND4_in[0] ,
         \SB2_2_29/Component_Function_0/NAND4_in[3] ,
         \SB2_2_29/Component_Function_0/NAND4_in[2] ,
         \SB2_2_29/Component_Function_0/NAND4_in[1] ,
         \SB2_2_29/Component_Function_0/NAND4_in[0] ,
         \SB2_2_29/Component_Function_1/NAND4_in[3] ,
         \SB2_2_29/Component_Function_1/NAND4_in[2] ,
         \SB2_2_29/Component_Function_1/NAND4_in[1] ,
         \SB2_2_29/Component_Function_1/NAND4_in[0] ,
         \SB2_2_29/Component_Function_5/NAND4_in[3] ,
         \SB2_2_29/Component_Function_5/NAND4_in[1] ,
         \SB2_2_29/Component_Function_5/NAND4_in[0] ,
         \SB2_2_30/Component_Function_0/NAND4_in[3] ,
         \SB2_2_30/Component_Function_0/NAND4_in[2] ,
         \SB2_2_30/Component_Function_0/NAND4_in[1] ,
         \SB2_2_30/Component_Function_0/NAND4_in[0] ,
         \SB2_2_30/Component_Function_1/NAND4_in[3] ,
         \SB2_2_30/Component_Function_1/NAND4_in[2] ,
         \SB2_2_30/Component_Function_1/NAND4_in[1] ,
         \SB2_2_30/Component_Function_1/NAND4_in[0] ,
         \SB2_2_30/Component_Function_5/NAND4_in[3] ,
         \SB2_2_30/Component_Function_5/NAND4_in[2] ,
         \SB2_2_30/Component_Function_5/NAND4_in[1] ,
         \SB2_2_31/Component_Function_0/NAND4_in[3] ,
         \SB2_2_31/Component_Function_0/NAND4_in[2] ,
         \SB2_2_31/Component_Function_0/NAND4_in[1] ,
         \SB2_2_31/Component_Function_0/NAND4_in[0] ,
         \SB2_2_31/Component_Function_1/NAND4_in[3] ,
         \SB2_2_31/Component_Function_1/NAND4_in[2] ,
         \SB2_2_31/Component_Function_1/NAND4_in[1] ,
         \SB2_2_31/Component_Function_1/NAND4_in[0] ,
         \SB2_2_31/Component_Function_5/NAND4_in[3] ,
         \SB2_2_31/Component_Function_5/NAND4_in[2] ,
         \SB2_2_31/Component_Function_5/NAND4_in[1] ,
         \SB2_2_31/Component_Function_5/NAND4_in[0] ,
         \SB1_3_0/Component_Function_0/NAND4_in[3] ,
         \SB1_3_0/Component_Function_0/NAND4_in[2] ,
         \SB1_3_0/Component_Function_0/NAND4_in[1] ,
         \SB1_3_0/Component_Function_0/NAND4_in[0] ,
         \SB1_3_0/Component_Function_1/NAND4_in[3] ,
         \SB1_3_0/Component_Function_1/NAND4_in[2] ,
         \SB1_3_0/Component_Function_1/NAND4_in[1] ,
         \SB1_3_0/Component_Function_1/NAND4_in[0] ,
         \SB1_3_0/Component_Function_5/NAND4_in[3] ,
         \SB1_3_0/Component_Function_5/NAND4_in[1] ,
         \SB1_3_0/Component_Function_5/NAND4_in[0] ,
         \SB1_3_1/Component_Function_0/NAND4_in[3] ,
         \SB1_3_1/Component_Function_0/NAND4_in[2] ,
         \SB1_3_1/Component_Function_0/NAND4_in[1] ,
         \SB1_3_1/Component_Function_0/NAND4_in[0] ,
         \SB1_3_1/Component_Function_1/NAND4_in[3] ,
         \SB1_3_1/Component_Function_1/NAND4_in[2] ,
         \SB1_3_1/Component_Function_1/NAND4_in[1] ,
         \SB1_3_1/Component_Function_1/NAND4_in[0] ,
         \SB1_3_1/Component_Function_5/NAND4_in[3] ,
         \SB1_3_1/Component_Function_5/NAND4_in[1] ,
         \SB1_3_1/Component_Function_5/NAND4_in[0] ,
         \SB1_3_2/Component_Function_0/NAND4_in[3] ,
         \SB1_3_2/Component_Function_0/NAND4_in[2] ,
         \SB1_3_2/Component_Function_0/NAND4_in[1] ,
         \SB1_3_2/Component_Function_0/NAND4_in[0] ,
         \SB1_3_2/Component_Function_1/NAND4_in[3] ,
         \SB1_3_2/Component_Function_1/NAND4_in[2] ,
         \SB1_3_2/Component_Function_1/NAND4_in[1] ,
         \SB1_3_2/Component_Function_1/NAND4_in[0] ,
         \SB1_3_2/Component_Function_5/NAND4_in[2] ,
         \SB1_3_2/Component_Function_5/NAND4_in[1] ,
         \SB1_3_2/Component_Function_5/NAND4_in[0] ,
         \SB1_3_3/Component_Function_0/NAND4_in[3] ,
         \SB1_3_3/Component_Function_0/NAND4_in[2] ,
         \SB1_3_3/Component_Function_0/NAND4_in[1] ,
         \SB1_3_3/Component_Function_0/NAND4_in[0] ,
         \SB1_3_3/Component_Function_1/NAND4_in[3] ,
         \SB1_3_3/Component_Function_1/NAND4_in[2] ,
         \SB1_3_3/Component_Function_1/NAND4_in[1] ,
         \SB1_3_3/Component_Function_1/NAND4_in[0] ,
         \SB1_3_3/Component_Function_5/NAND4_in[3] ,
         \SB1_3_3/Component_Function_5/NAND4_in[1] ,
         \SB1_3_3/Component_Function_5/NAND4_in[0] ,
         \SB1_3_4/Component_Function_0/NAND4_in[3] ,
         \SB1_3_4/Component_Function_0/NAND4_in[2] ,
         \SB1_3_4/Component_Function_0/NAND4_in[1] ,
         \SB1_3_4/Component_Function_0/NAND4_in[0] ,
         \SB1_3_4/Component_Function_1/NAND4_in[3] ,
         \SB1_3_4/Component_Function_1/NAND4_in[2] ,
         \SB1_3_4/Component_Function_1/NAND4_in[1] ,
         \SB1_3_4/Component_Function_1/NAND4_in[0] ,
         \SB1_3_4/Component_Function_5/NAND4_in[3] ,
         \SB1_3_4/Component_Function_5/NAND4_in[1] ,
         \SB1_3_4/Component_Function_5/NAND4_in[0] ,
         \SB1_3_5/Component_Function_0/NAND4_in[3] ,
         \SB1_3_5/Component_Function_0/NAND4_in[2] ,
         \SB1_3_5/Component_Function_0/NAND4_in[1] ,
         \SB1_3_5/Component_Function_0/NAND4_in[0] ,
         \SB1_3_5/Component_Function_1/NAND4_in[3] ,
         \SB1_3_5/Component_Function_1/NAND4_in[2] ,
         \SB1_3_5/Component_Function_1/NAND4_in[1] ,
         \SB1_3_5/Component_Function_1/NAND4_in[0] ,
         \SB1_3_5/Component_Function_5/NAND4_in[3] ,
         \SB1_3_5/Component_Function_5/NAND4_in[2] ,
         \SB1_3_5/Component_Function_5/NAND4_in[1] ,
         \SB1_3_5/Component_Function_5/NAND4_in[0] ,
         \SB1_3_6/Component_Function_0/NAND4_in[3] ,
         \SB1_3_6/Component_Function_0/NAND4_in[2] ,
         \SB1_3_6/Component_Function_0/NAND4_in[1] ,
         \SB1_3_6/Component_Function_0/NAND4_in[0] ,
         \SB1_3_6/Component_Function_1/NAND4_in[3] ,
         \SB1_3_6/Component_Function_1/NAND4_in[2] ,
         \SB1_3_6/Component_Function_1/NAND4_in[1] ,
         \SB1_3_6/Component_Function_1/NAND4_in[0] ,
         \SB1_3_6/Component_Function_5/NAND4_in[2] ,
         \SB1_3_6/Component_Function_5/NAND4_in[1] ,
         \SB1_3_6/Component_Function_5/NAND4_in[0] ,
         \SB1_3_7/Component_Function_0/NAND4_in[3] ,
         \SB1_3_7/Component_Function_0/NAND4_in[2] ,
         \SB1_3_7/Component_Function_0/NAND4_in[1] ,
         \SB1_3_7/Component_Function_0/NAND4_in[0] ,
         \SB1_3_7/Component_Function_1/NAND4_in[3] ,
         \SB1_3_7/Component_Function_1/NAND4_in[2] ,
         \SB1_3_7/Component_Function_1/NAND4_in[1] ,
         \SB1_3_7/Component_Function_1/NAND4_in[0] ,
         \SB1_3_7/Component_Function_5/NAND4_in[3] ,
         \SB1_3_7/Component_Function_5/NAND4_in[1] ,
         \SB1_3_7/Component_Function_5/NAND4_in[0] ,
         \SB1_3_8/Component_Function_0/NAND4_in[3] ,
         \SB1_3_8/Component_Function_0/NAND4_in[2] ,
         \SB1_3_8/Component_Function_0/NAND4_in[1] ,
         \SB1_3_8/Component_Function_0/NAND4_in[0] ,
         \SB1_3_8/Component_Function_1/NAND4_in[2] ,
         \SB1_3_8/Component_Function_1/NAND4_in[1] ,
         \SB1_3_8/Component_Function_1/NAND4_in[0] ,
         \SB1_3_8/Component_Function_5/NAND4_in[3] ,
         \SB1_3_8/Component_Function_5/NAND4_in[1] ,
         \SB1_3_8/Component_Function_5/NAND4_in[0] ,
         \SB1_3_9/Component_Function_0/NAND4_in[3] ,
         \SB1_3_9/Component_Function_0/NAND4_in[2] ,
         \SB1_3_9/Component_Function_0/NAND4_in[1] ,
         \SB1_3_9/Component_Function_0/NAND4_in[0] ,
         \SB1_3_9/Component_Function_1/NAND4_in[3] ,
         \SB1_3_9/Component_Function_1/NAND4_in[2] ,
         \SB1_3_9/Component_Function_1/NAND4_in[1] ,
         \SB1_3_9/Component_Function_1/NAND4_in[0] ,
         \SB1_3_9/Component_Function_5/NAND4_in[3] ,
         \SB1_3_9/Component_Function_5/NAND4_in[1] ,
         \SB1_3_9/Component_Function_5/NAND4_in[0] ,
         \SB1_3_10/Component_Function_0/NAND4_in[3] ,
         \SB1_3_10/Component_Function_0/NAND4_in[2] ,
         \SB1_3_10/Component_Function_0/NAND4_in[1] ,
         \SB1_3_10/Component_Function_0/NAND4_in[0] ,
         \SB1_3_10/Component_Function_1/NAND4_in[3] ,
         \SB1_3_10/Component_Function_1/NAND4_in[2] ,
         \SB1_3_10/Component_Function_1/NAND4_in[1] ,
         \SB1_3_10/Component_Function_1/NAND4_in[0] ,
         \SB1_3_10/Component_Function_5/NAND4_in[3] ,
         \SB1_3_10/Component_Function_5/NAND4_in[2] ,
         \SB1_3_10/Component_Function_5/NAND4_in[1] ,
         \SB1_3_10/Component_Function_5/NAND4_in[0] ,
         \SB1_3_11/Component_Function_0/NAND4_in[3] ,
         \SB1_3_11/Component_Function_0/NAND4_in[2] ,
         \SB1_3_11/Component_Function_0/NAND4_in[1] ,
         \SB1_3_11/Component_Function_0/NAND4_in[0] ,
         \SB1_3_11/Component_Function_1/NAND4_in[3] ,
         \SB1_3_11/Component_Function_1/NAND4_in[2] ,
         \SB1_3_11/Component_Function_1/NAND4_in[1] ,
         \SB1_3_11/Component_Function_1/NAND4_in[0] ,
         \SB1_3_11/Component_Function_5/NAND4_in[3] ,
         \SB1_3_11/Component_Function_5/NAND4_in[2] ,
         \SB1_3_11/Component_Function_5/NAND4_in[1] ,
         \SB1_3_11/Component_Function_5/NAND4_in[0] ,
         \SB1_3_12/Component_Function_0/NAND4_in[3] ,
         \SB1_3_12/Component_Function_0/NAND4_in[2] ,
         \SB1_3_12/Component_Function_0/NAND4_in[1] ,
         \SB1_3_12/Component_Function_0/NAND4_in[0] ,
         \SB1_3_12/Component_Function_1/NAND4_in[2] ,
         \SB1_3_12/Component_Function_1/NAND4_in[1] ,
         \SB1_3_12/Component_Function_1/NAND4_in[0] ,
         \SB1_3_12/Component_Function_5/NAND4_in[3] ,
         \SB1_3_12/Component_Function_5/NAND4_in[1] ,
         \SB1_3_12/Component_Function_5/NAND4_in[0] ,
         \SB1_3_13/Component_Function_0/NAND4_in[3] ,
         \SB1_3_13/Component_Function_0/NAND4_in[2] ,
         \SB1_3_13/Component_Function_0/NAND4_in[1] ,
         \SB1_3_13/Component_Function_0/NAND4_in[0] ,
         \SB1_3_13/Component_Function_1/NAND4_in[3] ,
         \SB1_3_13/Component_Function_1/NAND4_in[2] ,
         \SB1_3_13/Component_Function_1/NAND4_in[1] ,
         \SB1_3_13/Component_Function_1/NAND4_in[0] ,
         \SB1_3_13/Component_Function_5/NAND4_in[3] ,
         \SB1_3_13/Component_Function_5/NAND4_in[1] ,
         \SB1_3_13/Component_Function_5/NAND4_in[0] ,
         \SB1_3_14/Component_Function_0/NAND4_in[3] ,
         \SB1_3_14/Component_Function_0/NAND4_in[2] ,
         \SB1_3_14/Component_Function_0/NAND4_in[1] ,
         \SB1_3_14/Component_Function_0/NAND4_in[0] ,
         \SB1_3_14/Component_Function_1/NAND4_in[3] ,
         \SB1_3_14/Component_Function_1/NAND4_in[2] ,
         \SB1_3_14/Component_Function_1/NAND4_in[1] ,
         \SB1_3_14/Component_Function_1/NAND4_in[0] ,
         \SB1_3_14/Component_Function_5/NAND4_in[3] ,
         \SB1_3_14/Component_Function_5/NAND4_in[1] ,
         \SB1_3_14/Component_Function_5/NAND4_in[0] ,
         \SB1_3_15/Component_Function_0/NAND4_in[3] ,
         \SB1_3_15/Component_Function_0/NAND4_in[2] ,
         \SB1_3_15/Component_Function_0/NAND4_in[1] ,
         \SB1_3_15/Component_Function_0/NAND4_in[0] ,
         \SB1_3_15/Component_Function_1/NAND4_in[3] ,
         \SB1_3_15/Component_Function_1/NAND4_in[2] ,
         \SB1_3_15/Component_Function_1/NAND4_in[1] ,
         \SB1_3_15/Component_Function_1/NAND4_in[0] ,
         \SB1_3_15/Component_Function_5/NAND4_in[3] ,
         \SB1_3_15/Component_Function_5/NAND4_in[1] ,
         \SB1_3_15/Component_Function_5/NAND4_in[0] ,
         \SB1_3_16/Component_Function_0/NAND4_in[3] ,
         \SB1_3_16/Component_Function_0/NAND4_in[2] ,
         \SB1_3_16/Component_Function_0/NAND4_in[1] ,
         \SB1_3_16/Component_Function_0/NAND4_in[0] ,
         \SB1_3_16/Component_Function_1/NAND4_in[3] ,
         \SB1_3_16/Component_Function_1/NAND4_in[2] ,
         \SB1_3_16/Component_Function_1/NAND4_in[1] ,
         \SB1_3_16/Component_Function_1/NAND4_in[0] ,
         \SB1_3_16/Component_Function_5/NAND4_in[3] ,
         \SB1_3_16/Component_Function_5/NAND4_in[2] ,
         \SB1_3_16/Component_Function_5/NAND4_in[1] ,
         \SB1_3_16/Component_Function_5/NAND4_in[0] ,
         \SB1_3_17/Component_Function_0/NAND4_in[3] ,
         \SB1_3_17/Component_Function_0/NAND4_in[2] ,
         \SB1_3_17/Component_Function_0/NAND4_in[1] ,
         \SB1_3_17/Component_Function_0/NAND4_in[0] ,
         \SB1_3_17/Component_Function_1/NAND4_in[3] ,
         \SB1_3_17/Component_Function_1/NAND4_in[2] ,
         \SB1_3_17/Component_Function_1/NAND4_in[1] ,
         \SB1_3_17/Component_Function_1/NAND4_in[0] ,
         \SB1_3_17/Component_Function_5/NAND4_in[2] ,
         \SB1_3_17/Component_Function_5/NAND4_in[1] ,
         \SB1_3_17/Component_Function_5/NAND4_in[0] ,
         \SB1_3_18/Component_Function_0/NAND4_in[3] ,
         \SB1_3_18/Component_Function_0/NAND4_in[2] ,
         \SB1_3_18/Component_Function_0/NAND4_in[1] ,
         \SB1_3_18/Component_Function_0/NAND4_in[0] ,
         \SB1_3_18/Component_Function_1/NAND4_in[3] ,
         \SB1_3_18/Component_Function_1/NAND4_in[2] ,
         \SB1_3_18/Component_Function_1/NAND4_in[1] ,
         \SB1_3_18/Component_Function_1/NAND4_in[0] ,
         \SB1_3_18/Component_Function_5/NAND4_in[3] ,
         \SB1_3_18/Component_Function_5/NAND4_in[2] ,
         \SB1_3_18/Component_Function_5/NAND4_in[1] ,
         \SB1_3_18/Component_Function_5/NAND4_in[0] ,
         \SB1_3_19/Component_Function_0/NAND4_in[3] ,
         \SB1_3_19/Component_Function_0/NAND4_in[2] ,
         \SB1_3_19/Component_Function_0/NAND4_in[1] ,
         \SB1_3_19/Component_Function_0/NAND4_in[0] ,
         \SB1_3_19/Component_Function_1/NAND4_in[3] ,
         \SB1_3_19/Component_Function_1/NAND4_in[2] ,
         \SB1_3_19/Component_Function_1/NAND4_in[1] ,
         \SB1_3_19/Component_Function_1/NAND4_in[0] ,
         \SB1_3_19/Component_Function_5/NAND4_in[3] ,
         \SB1_3_19/Component_Function_5/NAND4_in[1] ,
         \SB1_3_19/Component_Function_5/NAND4_in[0] ,
         \SB1_3_20/Component_Function_0/NAND4_in[3] ,
         \SB1_3_20/Component_Function_0/NAND4_in[2] ,
         \SB1_3_20/Component_Function_0/NAND4_in[1] ,
         \SB1_3_20/Component_Function_0/NAND4_in[0] ,
         \SB1_3_20/Component_Function_1/NAND4_in[2] ,
         \SB1_3_20/Component_Function_1/NAND4_in[1] ,
         \SB1_3_20/Component_Function_1/NAND4_in[0] ,
         \SB1_3_20/Component_Function_5/NAND4_in[3] ,
         \SB1_3_20/Component_Function_5/NAND4_in[1] ,
         \SB1_3_20/Component_Function_5/NAND4_in[0] ,
         \SB1_3_21/Component_Function_0/NAND4_in[3] ,
         \SB1_3_21/Component_Function_0/NAND4_in[1] ,
         \SB1_3_21/Component_Function_0/NAND4_in[0] ,
         \SB1_3_21/Component_Function_1/NAND4_in[3] ,
         \SB1_3_21/Component_Function_1/NAND4_in[2] ,
         \SB1_3_21/Component_Function_1/NAND4_in[1] ,
         \SB1_3_21/Component_Function_1/NAND4_in[0] ,
         \SB1_3_21/Component_Function_5/NAND4_in[3] ,
         \SB1_3_21/Component_Function_5/NAND4_in[2] ,
         \SB1_3_21/Component_Function_5/NAND4_in[1] ,
         \SB1_3_21/Component_Function_5/NAND4_in[0] ,
         \SB1_3_22/Component_Function_0/NAND4_in[3] ,
         \SB1_3_22/Component_Function_0/NAND4_in[2] ,
         \SB1_3_22/Component_Function_0/NAND4_in[1] ,
         \SB1_3_22/Component_Function_0/NAND4_in[0] ,
         \SB1_3_22/Component_Function_1/NAND4_in[3] ,
         \SB1_3_22/Component_Function_1/NAND4_in[2] ,
         \SB1_3_22/Component_Function_1/NAND4_in[1] ,
         \SB1_3_22/Component_Function_1/NAND4_in[0] ,
         \SB1_3_22/Component_Function_5/NAND4_in[3] ,
         \SB1_3_22/Component_Function_5/NAND4_in[1] ,
         \SB1_3_22/Component_Function_5/NAND4_in[0] ,
         \SB1_3_23/Component_Function_0/NAND4_in[3] ,
         \SB1_3_23/Component_Function_0/NAND4_in[2] ,
         \SB1_3_23/Component_Function_0/NAND4_in[1] ,
         \SB1_3_23/Component_Function_0/NAND4_in[0] ,
         \SB1_3_23/Component_Function_1/NAND4_in[2] ,
         \SB1_3_23/Component_Function_1/NAND4_in[1] ,
         \SB1_3_23/Component_Function_1/NAND4_in[0] ,
         \SB1_3_23/Component_Function_5/NAND4_in[3] ,
         \SB1_3_23/Component_Function_5/NAND4_in[1] ,
         \SB1_3_23/Component_Function_5/NAND4_in[0] ,
         \SB1_3_24/Component_Function_0/NAND4_in[3] ,
         \SB1_3_24/Component_Function_0/NAND4_in[2] ,
         \SB1_3_24/Component_Function_0/NAND4_in[1] ,
         \SB1_3_24/Component_Function_0/NAND4_in[0] ,
         \SB1_3_24/Component_Function_1/NAND4_in[3] ,
         \SB1_3_24/Component_Function_1/NAND4_in[2] ,
         \SB1_3_24/Component_Function_1/NAND4_in[1] ,
         \SB1_3_24/Component_Function_1/NAND4_in[0] ,
         \SB1_3_24/Component_Function_5/NAND4_in[3] ,
         \SB1_3_24/Component_Function_5/NAND4_in[1] ,
         \SB1_3_24/Component_Function_5/NAND4_in[0] ,
         \SB1_3_25/Component_Function_0/NAND4_in[3] ,
         \SB1_3_25/Component_Function_0/NAND4_in[2] ,
         \SB1_3_25/Component_Function_0/NAND4_in[1] ,
         \SB1_3_25/Component_Function_0/NAND4_in[0] ,
         \SB1_3_25/Component_Function_1/NAND4_in[2] ,
         \SB1_3_25/Component_Function_1/NAND4_in[1] ,
         \SB1_3_25/Component_Function_1/NAND4_in[0] ,
         \SB1_3_25/Component_Function_5/NAND4_in[3] ,
         \SB1_3_25/Component_Function_5/NAND4_in[1] ,
         \SB1_3_25/Component_Function_5/NAND4_in[0] ,
         \SB1_3_26/Component_Function_0/NAND4_in[3] ,
         \SB1_3_26/Component_Function_0/NAND4_in[2] ,
         \SB1_3_26/Component_Function_0/NAND4_in[1] ,
         \SB1_3_26/Component_Function_0/NAND4_in[0] ,
         \SB1_3_26/Component_Function_1/NAND4_in[3] ,
         \SB1_3_26/Component_Function_1/NAND4_in[2] ,
         \SB1_3_26/Component_Function_1/NAND4_in[1] ,
         \SB1_3_26/Component_Function_1/NAND4_in[0] ,
         \SB1_3_26/Component_Function_5/NAND4_in[3] ,
         \SB1_3_26/Component_Function_5/NAND4_in[1] ,
         \SB1_3_26/Component_Function_5/NAND4_in[0] ,
         \SB1_3_27/Component_Function_0/NAND4_in[2] ,
         \SB1_3_27/Component_Function_0/NAND4_in[1] ,
         \SB1_3_27/Component_Function_0/NAND4_in[0] ,
         \SB1_3_27/Component_Function_1/NAND4_in[3] ,
         \SB1_3_27/Component_Function_1/NAND4_in[2] ,
         \SB1_3_27/Component_Function_1/NAND4_in[1] ,
         \SB1_3_27/Component_Function_1/NAND4_in[0] ,
         \SB1_3_27/Component_Function_5/NAND4_in[3] ,
         \SB1_3_27/Component_Function_5/NAND4_in[1] ,
         \SB1_3_27/Component_Function_5/NAND4_in[0] ,
         \SB1_3_28/Component_Function_0/NAND4_in[3] ,
         \SB1_3_28/Component_Function_0/NAND4_in[2] ,
         \SB1_3_28/Component_Function_0/NAND4_in[1] ,
         \SB1_3_28/Component_Function_0/NAND4_in[0] ,
         \SB1_3_28/Component_Function_1/NAND4_in[3] ,
         \SB1_3_28/Component_Function_1/NAND4_in[2] ,
         \SB1_3_28/Component_Function_1/NAND4_in[1] ,
         \SB1_3_28/Component_Function_1/NAND4_in[0] ,
         \SB1_3_28/Component_Function_5/NAND4_in[3] ,
         \SB1_3_28/Component_Function_5/NAND4_in[1] ,
         \SB1_3_28/Component_Function_5/NAND4_in[0] ,
         \SB1_3_29/Component_Function_0/NAND4_in[3] ,
         \SB1_3_29/Component_Function_0/NAND4_in[2] ,
         \SB1_3_29/Component_Function_0/NAND4_in[1] ,
         \SB1_3_29/Component_Function_0/NAND4_in[0] ,
         \SB1_3_29/Component_Function_1/NAND4_in[3] ,
         \SB1_3_29/Component_Function_1/NAND4_in[2] ,
         \SB1_3_29/Component_Function_1/NAND4_in[1] ,
         \SB1_3_29/Component_Function_1/NAND4_in[0] ,
         \SB1_3_29/Component_Function_5/NAND4_in[3] ,
         \SB1_3_29/Component_Function_5/NAND4_in[1] ,
         \SB1_3_29/Component_Function_5/NAND4_in[0] ,
         \SB1_3_30/Component_Function_0/NAND4_in[3] ,
         \SB1_3_30/Component_Function_0/NAND4_in[2] ,
         \SB1_3_30/Component_Function_0/NAND4_in[1] ,
         \SB1_3_30/Component_Function_0/NAND4_in[0] ,
         \SB1_3_30/Component_Function_1/NAND4_in[3] ,
         \SB1_3_30/Component_Function_1/NAND4_in[2] ,
         \SB1_3_30/Component_Function_1/NAND4_in[1] ,
         \SB1_3_30/Component_Function_1/NAND4_in[0] ,
         \SB1_3_30/Component_Function_5/NAND4_in[3] ,
         \SB1_3_30/Component_Function_5/NAND4_in[1] ,
         \SB1_3_30/Component_Function_5/NAND4_in[0] ,
         \SB1_3_31/Component_Function_0/NAND4_in[3] ,
         \SB1_3_31/Component_Function_0/NAND4_in[2] ,
         \SB1_3_31/Component_Function_0/NAND4_in[1] ,
         \SB1_3_31/Component_Function_0/NAND4_in[0] ,
         \SB1_3_31/Component_Function_1/NAND4_in[3] ,
         \SB1_3_31/Component_Function_1/NAND4_in[2] ,
         \SB1_3_31/Component_Function_1/NAND4_in[1] ,
         \SB1_3_31/Component_Function_1/NAND4_in[0] ,
         \SB1_3_31/Component_Function_5/NAND4_in[3] ,
         \SB1_3_31/Component_Function_5/NAND4_in[1] ,
         \SB1_3_31/Component_Function_5/NAND4_in[0] ,
         \SB2_3_0/Component_Function_0/NAND4_in[3] ,
         \SB2_3_0/Component_Function_0/NAND4_in[2] ,
         \SB2_3_0/Component_Function_0/NAND4_in[1] ,
         \SB2_3_0/Component_Function_0/NAND4_in[0] ,
         \SB2_3_0/Component_Function_1/NAND4_in[3] ,
         \SB2_3_0/Component_Function_1/NAND4_in[2] ,
         \SB2_3_0/Component_Function_1/NAND4_in[1] ,
         \SB2_3_0/Component_Function_1/NAND4_in[0] ,
         \SB2_3_0/Component_Function_5/NAND4_in[3] ,
         \SB2_3_0/Component_Function_5/NAND4_in[1] ,
         \SB2_3_0/Component_Function_5/NAND4_in[0] ,
         \SB2_3_1/Component_Function_0/NAND4_in[3] ,
         \SB2_3_1/Component_Function_0/NAND4_in[2] ,
         \SB2_3_1/Component_Function_0/NAND4_in[1] ,
         \SB2_3_1/Component_Function_0/NAND4_in[0] ,
         \SB2_3_1/Component_Function_1/NAND4_in[3] ,
         \SB2_3_1/Component_Function_1/NAND4_in[2] ,
         \SB2_3_1/Component_Function_1/NAND4_in[1] ,
         \SB2_3_1/Component_Function_1/NAND4_in[0] ,
         \SB2_3_1/Component_Function_5/NAND4_in[3] ,
         \SB2_3_1/Component_Function_5/NAND4_in[1] ,
         \SB2_3_1/Component_Function_5/NAND4_in[0] ,
         \SB2_3_2/Component_Function_0/NAND4_in[3] ,
         \SB2_3_2/Component_Function_0/NAND4_in[2] ,
         \SB2_3_2/Component_Function_0/NAND4_in[1] ,
         \SB2_3_2/Component_Function_0/NAND4_in[0] ,
         \SB2_3_2/Component_Function_1/NAND4_in[3] ,
         \SB2_3_2/Component_Function_1/NAND4_in[2] ,
         \SB2_3_2/Component_Function_1/NAND4_in[1] ,
         \SB2_3_2/Component_Function_1/NAND4_in[0] ,
         \SB2_3_2/Component_Function_5/NAND4_in[3] ,
         \SB2_3_2/Component_Function_5/NAND4_in[1] ,
         \SB2_3_2/Component_Function_5/NAND4_in[0] ,
         \SB2_3_3/Component_Function_0/NAND4_in[3] ,
         \SB2_3_3/Component_Function_0/NAND4_in[2] ,
         \SB2_3_3/Component_Function_0/NAND4_in[1] ,
         \SB2_3_3/Component_Function_0/NAND4_in[0] ,
         \SB2_3_3/Component_Function_1/NAND4_in[3] ,
         \SB2_3_3/Component_Function_1/NAND4_in[2] ,
         \SB2_3_3/Component_Function_1/NAND4_in[1] ,
         \SB2_3_3/Component_Function_1/NAND4_in[0] ,
         \SB2_3_3/Component_Function_5/NAND4_in[3] ,
         \SB2_3_3/Component_Function_5/NAND4_in[1] ,
         \SB2_3_3/Component_Function_5/NAND4_in[0] ,
         \SB2_3_4/Component_Function_0/NAND4_in[3] ,
         \SB2_3_4/Component_Function_0/NAND4_in[2] ,
         \SB2_3_4/Component_Function_0/NAND4_in[1] ,
         \SB2_3_4/Component_Function_0/NAND4_in[0] ,
         \SB2_3_4/Component_Function_1/NAND4_in[3] ,
         \SB2_3_4/Component_Function_1/NAND4_in[2] ,
         \SB2_3_4/Component_Function_1/NAND4_in[1] ,
         \SB2_3_4/Component_Function_1/NAND4_in[0] ,
         \SB2_3_4/Component_Function_5/NAND4_in[3] ,
         \SB2_3_4/Component_Function_5/NAND4_in[1] ,
         \SB2_3_4/Component_Function_5/NAND4_in[0] ,
         \SB2_3_5/Component_Function_0/NAND4_in[3] ,
         \SB2_3_5/Component_Function_0/NAND4_in[2] ,
         \SB2_3_5/Component_Function_0/NAND4_in[1] ,
         \SB2_3_5/Component_Function_0/NAND4_in[0] ,
         \SB2_3_5/Component_Function_1/NAND4_in[3] ,
         \SB2_3_5/Component_Function_1/NAND4_in[2] ,
         \SB2_3_5/Component_Function_1/NAND4_in[1] ,
         \SB2_3_5/Component_Function_1/NAND4_in[0] ,
         \SB2_3_5/Component_Function_5/NAND4_in[3] ,
         \SB2_3_5/Component_Function_5/NAND4_in[1] ,
         \SB2_3_5/Component_Function_5/NAND4_in[0] ,
         \SB2_3_6/Component_Function_0/NAND4_in[3] ,
         \SB2_3_6/Component_Function_0/NAND4_in[2] ,
         \SB2_3_6/Component_Function_0/NAND4_in[1] ,
         \SB2_3_6/Component_Function_0/NAND4_in[0] ,
         \SB2_3_6/Component_Function_1/NAND4_in[3] ,
         \SB2_3_6/Component_Function_1/NAND4_in[2] ,
         \SB2_3_6/Component_Function_1/NAND4_in[1] ,
         \SB2_3_6/Component_Function_1/NAND4_in[0] ,
         \SB2_3_6/Component_Function_5/NAND4_in[3] ,
         \SB2_3_6/Component_Function_5/NAND4_in[2] ,
         \SB2_3_6/Component_Function_5/NAND4_in[1] ,
         \SB2_3_6/Component_Function_5/NAND4_in[0] ,
         \SB2_3_7/Component_Function_0/NAND4_in[3] ,
         \SB2_3_7/Component_Function_0/NAND4_in[2] ,
         \SB2_3_7/Component_Function_0/NAND4_in[1] ,
         \SB2_3_7/Component_Function_0/NAND4_in[0] ,
         \SB2_3_7/Component_Function_1/NAND4_in[3] ,
         \SB2_3_7/Component_Function_1/NAND4_in[2] ,
         \SB2_3_7/Component_Function_1/NAND4_in[1] ,
         \SB2_3_7/Component_Function_1/NAND4_in[0] ,
         \SB2_3_7/Component_Function_5/NAND4_in[3] ,
         \SB2_3_7/Component_Function_5/NAND4_in[1] ,
         \SB2_3_7/Component_Function_5/NAND4_in[0] ,
         \SB2_3_8/Component_Function_0/NAND4_in[3] ,
         \SB2_3_8/Component_Function_0/NAND4_in[2] ,
         \SB2_3_8/Component_Function_0/NAND4_in[1] ,
         \SB2_3_8/Component_Function_0/NAND4_in[0] ,
         \SB2_3_8/Component_Function_1/NAND4_in[3] ,
         \SB2_3_8/Component_Function_1/NAND4_in[2] ,
         \SB2_3_8/Component_Function_1/NAND4_in[1] ,
         \SB2_3_8/Component_Function_1/NAND4_in[0] ,
         \SB2_3_8/Component_Function_5/NAND4_in[3] ,
         \SB2_3_8/Component_Function_5/NAND4_in[2] ,
         \SB2_3_8/Component_Function_5/NAND4_in[1] ,
         \SB2_3_8/Component_Function_5/NAND4_in[0] ,
         \SB2_3_9/Component_Function_0/NAND4_in[3] ,
         \SB2_3_9/Component_Function_0/NAND4_in[2] ,
         \SB2_3_9/Component_Function_0/NAND4_in[1] ,
         \SB2_3_9/Component_Function_0/NAND4_in[0] ,
         \SB2_3_9/Component_Function_1/NAND4_in[3] ,
         \SB2_3_9/Component_Function_1/NAND4_in[2] ,
         \SB2_3_9/Component_Function_1/NAND4_in[1] ,
         \SB2_3_9/Component_Function_1/NAND4_in[0] ,
         \SB2_3_9/Component_Function_5/NAND4_in[3] ,
         \SB2_3_9/Component_Function_5/NAND4_in[1] ,
         \SB2_3_9/Component_Function_5/NAND4_in[0] ,
         \SB2_3_10/Component_Function_0/NAND4_in[3] ,
         \SB2_3_10/Component_Function_0/NAND4_in[2] ,
         \SB2_3_10/Component_Function_0/NAND4_in[1] ,
         \SB2_3_10/Component_Function_0/NAND4_in[0] ,
         \SB2_3_10/Component_Function_1/NAND4_in[3] ,
         \SB2_3_10/Component_Function_1/NAND4_in[2] ,
         \SB2_3_10/Component_Function_1/NAND4_in[1] ,
         \SB2_3_10/Component_Function_1/NAND4_in[0] ,
         \SB2_3_10/Component_Function_5/NAND4_in[3] ,
         \SB2_3_10/Component_Function_5/NAND4_in[1] ,
         \SB2_3_10/Component_Function_5/NAND4_in[0] ,
         \SB2_3_11/Component_Function_0/NAND4_in[3] ,
         \SB2_3_11/Component_Function_0/NAND4_in[2] ,
         \SB2_3_11/Component_Function_0/NAND4_in[1] ,
         \SB2_3_11/Component_Function_0/NAND4_in[0] ,
         \SB2_3_11/Component_Function_1/NAND4_in[3] ,
         \SB2_3_11/Component_Function_1/NAND4_in[2] ,
         \SB2_3_11/Component_Function_1/NAND4_in[1] ,
         \SB2_3_11/Component_Function_1/NAND4_in[0] ,
         \SB2_3_11/Component_Function_5/NAND4_in[3] ,
         \SB2_3_11/Component_Function_5/NAND4_in[2] ,
         \SB2_3_11/Component_Function_5/NAND4_in[1] ,
         \SB2_3_11/Component_Function_5/NAND4_in[0] ,
         \SB2_3_12/Component_Function_0/NAND4_in[3] ,
         \SB2_3_12/Component_Function_0/NAND4_in[2] ,
         \SB2_3_12/Component_Function_0/NAND4_in[1] ,
         \SB2_3_12/Component_Function_0/NAND4_in[0] ,
         \SB2_3_12/Component_Function_1/NAND4_in[3] ,
         \SB2_3_12/Component_Function_1/NAND4_in[2] ,
         \SB2_3_12/Component_Function_1/NAND4_in[1] ,
         \SB2_3_12/Component_Function_1/NAND4_in[0] ,
         \SB2_3_12/Component_Function_5/NAND4_in[3] ,
         \SB2_3_12/Component_Function_5/NAND4_in[1] ,
         \SB2_3_12/Component_Function_5/NAND4_in[0] ,
         \SB2_3_13/Component_Function_0/NAND4_in[3] ,
         \SB2_3_13/Component_Function_0/NAND4_in[2] ,
         \SB2_3_13/Component_Function_0/NAND4_in[1] ,
         \SB2_3_13/Component_Function_0/NAND4_in[0] ,
         \SB2_3_13/Component_Function_1/NAND4_in[3] ,
         \SB2_3_13/Component_Function_1/NAND4_in[2] ,
         \SB2_3_13/Component_Function_1/NAND4_in[1] ,
         \SB2_3_13/Component_Function_1/NAND4_in[0] ,
         \SB2_3_13/Component_Function_5/NAND4_in[2] ,
         \SB2_3_13/Component_Function_5/NAND4_in[1] ,
         \SB2_3_13/Component_Function_5/NAND4_in[0] ,
         \SB2_3_14/Component_Function_0/NAND4_in[3] ,
         \SB2_3_14/Component_Function_0/NAND4_in[2] ,
         \SB2_3_14/Component_Function_0/NAND4_in[1] ,
         \SB2_3_14/Component_Function_0/NAND4_in[0] ,
         \SB2_3_14/Component_Function_1/NAND4_in[3] ,
         \SB2_3_14/Component_Function_1/NAND4_in[2] ,
         \SB2_3_14/Component_Function_1/NAND4_in[1] ,
         \SB2_3_14/Component_Function_1/NAND4_in[0] ,
         \SB2_3_14/Component_Function_5/NAND4_in[3] ,
         \SB2_3_14/Component_Function_5/NAND4_in[1] ,
         \SB2_3_14/Component_Function_5/NAND4_in[0] ,
         \SB2_3_15/Component_Function_0/NAND4_in[3] ,
         \SB2_3_15/Component_Function_0/NAND4_in[2] ,
         \SB2_3_15/Component_Function_0/NAND4_in[1] ,
         \SB2_3_15/Component_Function_0/NAND4_in[0] ,
         \SB2_3_15/Component_Function_1/NAND4_in[3] ,
         \SB2_3_15/Component_Function_1/NAND4_in[2] ,
         \SB2_3_15/Component_Function_1/NAND4_in[1] ,
         \SB2_3_15/Component_Function_1/NAND4_in[0] ,
         \SB2_3_15/Component_Function_5/NAND4_in[3] ,
         \SB2_3_15/Component_Function_5/NAND4_in[1] ,
         \SB2_3_15/Component_Function_5/NAND4_in[0] ,
         \SB2_3_16/Component_Function_0/NAND4_in[3] ,
         \SB2_3_16/Component_Function_0/NAND4_in[2] ,
         \SB2_3_16/Component_Function_0/NAND4_in[1] ,
         \SB2_3_16/Component_Function_0/NAND4_in[0] ,
         \SB2_3_16/Component_Function_1/NAND4_in[3] ,
         \SB2_3_16/Component_Function_1/NAND4_in[2] ,
         \SB2_3_16/Component_Function_1/NAND4_in[1] ,
         \SB2_3_16/Component_Function_1/NAND4_in[0] ,
         \SB2_3_16/Component_Function_5/NAND4_in[3] ,
         \SB2_3_16/Component_Function_5/NAND4_in[1] ,
         \SB2_3_16/Component_Function_5/NAND4_in[0] ,
         \SB2_3_17/Component_Function_0/NAND4_in[3] ,
         \SB2_3_17/Component_Function_0/NAND4_in[2] ,
         \SB2_3_17/Component_Function_0/NAND4_in[1] ,
         \SB2_3_17/Component_Function_0/NAND4_in[0] ,
         \SB2_3_17/Component_Function_1/NAND4_in[3] ,
         \SB2_3_17/Component_Function_1/NAND4_in[2] ,
         \SB2_3_17/Component_Function_1/NAND4_in[1] ,
         \SB2_3_17/Component_Function_1/NAND4_in[0] ,
         \SB2_3_17/Component_Function_5/NAND4_in[2] ,
         \SB2_3_17/Component_Function_5/NAND4_in[0] ,
         \SB2_3_18/Component_Function_0/NAND4_in[3] ,
         \SB2_3_18/Component_Function_0/NAND4_in[2] ,
         \SB2_3_18/Component_Function_0/NAND4_in[1] ,
         \SB2_3_18/Component_Function_0/NAND4_in[0] ,
         \SB2_3_18/Component_Function_1/NAND4_in[3] ,
         \SB2_3_18/Component_Function_1/NAND4_in[2] ,
         \SB2_3_18/Component_Function_1/NAND4_in[1] ,
         \SB2_3_18/Component_Function_1/NAND4_in[0] ,
         \SB2_3_18/Component_Function_5/NAND4_in[3] ,
         \SB2_3_18/Component_Function_5/NAND4_in[2] ,
         \SB2_3_18/Component_Function_5/NAND4_in[1] ,
         \SB2_3_18/Component_Function_5/NAND4_in[0] ,
         \SB2_3_19/Component_Function_0/NAND4_in[3] ,
         \SB2_3_19/Component_Function_0/NAND4_in[2] ,
         \SB2_3_19/Component_Function_0/NAND4_in[1] ,
         \SB2_3_19/Component_Function_0/NAND4_in[0] ,
         \SB2_3_19/Component_Function_1/NAND4_in[3] ,
         \SB2_3_19/Component_Function_1/NAND4_in[2] ,
         \SB2_3_19/Component_Function_1/NAND4_in[1] ,
         \SB2_3_19/Component_Function_1/NAND4_in[0] ,
         \SB2_3_19/Component_Function_5/NAND4_in[3] ,
         \SB2_3_19/Component_Function_5/NAND4_in[2] ,
         \SB2_3_19/Component_Function_5/NAND4_in[1] ,
         \SB2_3_19/Component_Function_5/NAND4_in[0] ,
         \SB2_3_20/Component_Function_0/NAND4_in[3] ,
         \SB2_3_20/Component_Function_0/NAND4_in[2] ,
         \SB2_3_20/Component_Function_0/NAND4_in[1] ,
         \SB2_3_20/Component_Function_0/NAND4_in[0] ,
         \SB2_3_20/Component_Function_1/NAND4_in[3] ,
         \SB2_3_20/Component_Function_1/NAND4_in[2] ,
         \SB2_3_20/Component_Function_1/NAND4_in[1] ,
         \SB2_3_20/Component_Function_1/NAND4_in[0] ,
         \SB2_3_20/Component_Function_5/NAND4_in[3] ,
         \SB2_3_20/Component_Function_5/NAND4_in[1] ,
         \SB2_3_20/Component_Function_5/NAND4_in[0] ,
         \SB2_3_21/Component_Function_0/NAND4_in[3] ,
         \SB2_3_21/Component_Function_0/NAND4_in[2] ,
         \SB2_3_21/Component_Function_0/NAND4_in[1] ,
         \SB2_3_21/Component_Function_0/NAND4_in[0] ,
         \SB2_3_21/Component_Function_1/NAND4_in[3] ,
         \SB2_3_21/Component_Function_1/NAND4_in[2] ,
         \SB2_3_21/Component_Function_1/NAND4_in[1] ,
         \SB2_3_21/Component_Function_1/NAND4_in[0] ,
         \SB2_3_21/Component_Function_5/NAND4_in[3] ,
         \SB2_3_21/Component_Function_5/NAND4_in[2] ,
         \SB2_3_21/Component_Function_5/NAND4_in[1] ,
         \SB2_3_21/Component_Function_5/NAND4_in[0] ,
         \SB2_3_22/Component_Function_0/NAND4_in[3] ,
         \SB2_3_22/Component_Function_0/NAND4_in[2] ,
         \SB2_3_22/Component_Function_0/NAND4_in[1] ,
         \SB2_3_22/Component_Function_0/NAND4_in[0] ,
         \SB2_3_22/Component_Function_1/NAND4_in[3] ,
         \SB2_3_22/Component_Function_1/NAND4_in[2] ,
         \SB2_3_22/Component_Function_1/NAND4_in[1] ,
         \SB2_3_22/Component_Function_1/NAND4_in[0] ,
         \SB2_3_22/Component_Function_5/NAND4_in[3] ,
         \SB2_3_22/Component_Function_5/NAND4_in[1] ,
         \SB2_3_22/Component_Function_5/NAND4_in[0] ,
         \SB2_3_23/Component_Function_0/NAND4_in[3] ,
         \SB2_3_23/Component_Function_0/NAND4_in[2] ,
         \SB2_3_23/Component_Function_0/NAND4_in[1] ,
         \SB2_3_23/Component_Function_0/NAND4_in[0] ,
         \SB2_3_23/Component_Function_1/NAND4_in[3] ,
         \SB2_3_23/Component_Function_1/NAND4_in[2] ,
         \SB2_3_23/Component_Function_1/NAND4_in[1] ,
         \SB2_3_23/Component_Function_1/NAND4_in[0] ,
         \SB2_3_23/Component_Function_5/NAND4_in[3] ,
         \SB2_3_23/Component_Function_5/NAND4_in[2] ,
         \SB2_3_23/Component_Function_5/NAND4_in[1] ,
         \SB2_3_24/Component_Function_0/NAND4_in[3] ,
         \SB2_3_24/Component_Function_0/NAND4_in[2] ,
         \SB2_3_24/Component_Function_0/NAND4_in[1] ,
         \SB2_3_24/Component_Function_0/NAND4_in[0] ,
         \SB2_3_24/Component_Function_1/NAND4_in[3] ,
         \SB2_3_24/Component_Function_1/NAND4_in[2] ,
         \SB2_3_24/Component_Function_1/NAND4_in[1] ,
         \SB2_3_24/Component_Function_1/NAND4_in[0] ,
         \SB2_3_24/Component_Function_5/NAND4_in[2] ,
         \SB2_3_24/Component_Function_5/NAND4_in[1] ,
         \SB2_3_24/Component_Function_5/NAND4_in[0] ,
         \SB2_3_25/Component_Function_0/NAND4_in[3] ,
         \SB2_3_25/Component_Function_0/NAND4_in[2] ,
         \SB2_3_25/Component_Function_0/NAND4_in[1] ,
         \SB2_3_25/Component_Function_0/NAND4_in[0] ,
         \SB2_3_25/Component_Function_1/NAND4_in[3] ,
         \SB2_3_25/Component_Function_1/NAND4_in[2] ,
         \SB2_3_25/Component_Function_1/NAND4_in[1] ,
         \SB2_3_25/Component_Function_1/NAND4_in[0] ,
         \SB2_3_25/Component_Function_5/NAND4_in[3] ,
         \SB2_3_25/Component_Function_5/NAND4_in[2] ,
         \SB2_3_25/Component_Function_5/NAND4_in[1] ,
         \SB2_3_25/Component_Function_5/NAND4_in[0] ,
         \SB2_3_26/Component_Function_0/NAND4_in[3] ,
         \SB2_3_26/Component_Function_0/NAND4_in[2] ,
         \SB2_3_26/Component_Function_0/NAND4_in[1] ,
         \SB2_3_26/Component_Function_0/NAND4_in[0] ,
         \SB2_3_26/Component_Function_1/NAND4_in[3] ,
         \SB2_3_26/Component_Function_1/NAND4_in[2] ,
         \SB2_3_26/Component_Function_1/NAND4_in[1] ,
         \SB2_3_26/Component_Function_1/NAND4_in[0] ,
         \SB2_3_26/Component_Function_5/NAND4_in[3] ,
         \SB2_3_26/Component_Function_5/NAND4_in[1] ,
         \SB2_3_27/Component_Function_0/NAND4_in[3] ,
         \SB2_3_27/Component_Function_0/NAND4_in[2] ,
         \SB2_3_27/Component_Function_0/NAND4_in[1] ,
         \SB2_3_27/Component_Function_0/NAND4_in[0] ,
         \SB2_3_27/Component_Function_1/NAND4_in[3] ,
         \SB2_3_27/Component_Function_1/NAND4_in[2] ,
         \SB2_3_27/Component_Function_1/NAND4_in[1] ,
         \SB2_3_27/Component_Function_1/NAND4_in[0] ,
         \SB2_3_27/Component_Function_5/NAND4_in[3] ,
         \SB2_3_27/Component_Function_5/NAND4_in[1] ,
         \SB2_3_27/Component_Function_5/NAND4_in[0] ,
         \SB2_3_28/Component_Function_0/NAND4_in[3] ,
         \SB2_3_28/Component_Function_0/NAND4_in[2] ,
         \SB2_3_28/Component_Function_0/NAND4_in[1] ,
         \SB2_3_28/Component_Function_0/NAND4_in[0] ,
         \SB2_3_28/Component_Function_1/NAND4_in[3] ,
         \SB2_3_28/Component_Function_1/NAND4_in[2] ,
         \SB2_3_28/Component_Function_1/NAND4_in[1] ,
         \SB2_3_28/Component_Function_1/NAND4_in[0] ,
         \SB2_3_28/Component_Function_5/NAND4_in[2] ,
         \SB2_3_28/Component_Function_5/NAND4_in[1] ,
         \SB2_3_28/Component_Function_5/NAND4_in[0] ,
         \SB2_3_29/Component_Function_0/NAND4_in[3] ,
         \SB2_3_29/Component_Function_0/NAND4_in[2] ,
         \SB2_3_29/Component_Function_0/NAND4_in[1] ,
         \SB2_3_29/Component_Function_0/NAND4_in[0] ,
         \SB2_3_29/Component_Function_1/NAND4_in[3] ,
         \SB2_3_29/Component_Function_1/NAND4_in[2] ,
         \SB2_3_29/Component_Function_1/NAND4_in[1] ,
         \SB2_3_29/Component_Function_1/NAND4_in[0] ,
         \SB2_3_29/Component_Function_5/NAND4_in[2] ,
         \SB2_3_29/Component_Function_5/NAND4_in[1] ,
         \SB2_3_29/Component_Function_5/NAND4_in[0] ,
         \SB2_3_30/Component_Function_0/NAND4_in[3] ,
         \SB2_3_30/Component_Function_0/NAND4_in[2] ,
         \SB2_3_30/Component_Function_0/NAND4_in[1] ,
         \SB2_3_30/Component_Function_0/NAND4_in[0] ,
         \SB2_3_30/Component_Function_1/NAND4_in[3] ,
         \SB2_3_30/Component_Function_1/NAND4_in[2] ,
         \SB2_3_30/Component_Function_1/NAND4_in[1] ,
         \SB2_3_30/Component_Function_1/NAND4_in[0] ,
         \SB2_3_30/Component_Function_5/NAND4_in[2] ,
         \SB2_3_30/Component_Function_5/NAND4_in[1] ,
         \SB2_3_30/Component_Function_5/NAND4_in[0] ,
         \SB2_3_31/Component_Function_0/NAND4_in[3] ,
         \SB2_3_31/Component_Function_0/NAND4_in[2] ,
         \SB2_3_31/Component_Function_0/NAND4_in[1] ,
         \SB2_3_31/Component_Function_0/NAND4_in[0] ,
         \SB2_3_31/Component_Function_1/NAND4_in[3] ,
         \SB2_3_31/Component_Function_1/NAND4_in[2] ,
         \SB2_3_31/Component_Function_1/NAND4_in[1] ,
         \SB2_3_31/Component_Function_1/NAND4_in[0] ,
         \SB2_3_31/Component_Function_5/NAND4_in[2] ,
         \SB2_3_31/Component_Function_5/NAND4_in[1] ,
         \SB2_3_31/Component_Function_5/NAND4_in[0] ,
         \SB3_0/Component_Function_0/NAND4_in[3] ,
         \SB3_0/Component_Function_0/NAND4_in[2] ,
         \SB3_0/Component_Function_0/NAND4_in[1] ,
         \SB3_0/Component_Function_0/NAND4_in[0] ,
         \SB3_0/Component_Function_1/NAND4_in[3] ,
         \SB3_0/Component_Function_1/NAND4_in[2] ,
         \SB3_0/Component_Function_1/NAND4_in[1] ,
         \SB3_0/Component_Function_1/NAND4_in[0] ,
         \SB3_0/Component_Function_5/NAND4_in[3] ,
         \SB3_0/Component_Function_5/NAND4_in[2] ,
         \SB3_0/Component_Function_5/NAND4_in[1] ,
         \SB3_0/Component_Function_5/NAND4_in[0] ,
         \SB3_1/Component_Function_0/NAND4_in[2] ,
         \SB3_1/Component_Function_0/NAND4_in[1] ,
         \SB3_1/Component_Function_0/NAND4_in[0] ,
         \SB3_1/Component_Function_1/NAND4_in[3] ,
         \SB3_1/Component_Function_1/NAND4_in[2] ,
         \SB3_1/Component_Function_1/NAND4_in[1] ,
         \SB3_1/Component_Function_1/NAND4_in[0] ,
         \SB3_1/Component_Function_5/NAND4_in[3] ,
         \SB3_1/Component_Function_5/NAND4_in[1] ,
         \SB3_1/Component_Function_5/NAND4_in[0] ,
         \SB3_2/Component_Function_0/NAND4_in[2] ,
         \SB3_2/Component_Function_0/NAND4_in[1] ,
         \SB3_2/Component_Function_0/NAND4_in[0] ,
         \SB3_2/Component_Function_1/NAND4_in[3] ,
         \SB3_2/Component_Function_1/NAND4_in[2] ,
         \SB3_2/Component_Function_1/NAND4_in[1] ,
         \SB3_2/Component_Function_1/NAND4_in[0] ,
         \SB3_2/Component_Function_5/NAND4_in[2] ,
         \SB3_2/Component_Function_5/NAND4_in[1] ,
         \SB3_2/Component_Function_5/NAND4_in[0] ,
         \SB3_3/Component_Function_0/NAND4_in[3] ,
         \SB3_3/Component_Function_0/NAND4_in[1] ,
         \SB3_3/Component_Function_0/NAND4_in[0] ,
         \SB3_3/Component_Function_1/NAND4_in[3] ,
         \SB3_3/Component_Function_1/NAND4_in[2] ,
         \SB3_3/Component_Function_1/NAND4_in[1] ,
         \SB3_3/Component_Function_1/NAND4_in[0] ,
         \SB3_3/Component_Function_5/NAND4_in[3] ,
         \SB3_3/Component_Function_5/NAND4_in[1] ,
         \SB3_3/Component_Function_5/NAND4_in[0] ,
         \SB3_4/Component_Function_0/NAND4_in[3] ,
         \SB3_4/Component_Function_0/NAND4_in[2] ,
         \SB3_4/Component_Function_0/NAND4_in[1] ,
         \SB3_4/Component_Function_0/NAND4_in[0] ,
         \SB3_4/Component_Function_1/NAND4_in[3] ,
         \SB3_4/Component_Function_1/NAND4_in[2] ,
         \SB3_4/Component_Function_1/NAND4_in[1] ,
         \SB3_4/Component_Function_1/NAND4_in[0] ,
         \SB3_4/Component_Function_5/NAND4_in[3] ,
         \SB3_4/Component_Function_5/NAND4_in[2] ,
         \SB3_4/Component_Function_5/NAND4_in[1] ,
         \SB3_4/Component_Function_5/NAND4_in[0] ,
         \SB3_5/Component_Function_0/NAND4_in[2] ,
         \SB3_5/Component_Function_0/NAND4_in[1] ,
         \SB3_5/Component_Function_0/NAND4_in[0] ,
         \SB3_5/Component_Function_1/NAND4_in[3] ,
         \SB3_5/Component_Function_1/NAND4_in[2] ,
         \SB3_5/Component_Function_1/NAND4_in[1] ,
         \SB3_5/Component_Function_1/NAND4_in[0] ,
         \SB3_5/Component_Function_5/NAND4_in[3] ,
         \SB3_5/Component_Function_5/NAND4_in[2] ,
         \SB3_5/Component_Function_5/NAND4_in[1] ,
         \SB3_5/Component_Function_5/NAND4_in[0] ,
         \SB3_6/Component_Function_0/NAND4_in[2] ,
         \SB3_6/Component_Function_0/NAND4_in[1] ,
         \SB3_6/Component_Function_0/NAND4_in[0] ,
         \SB3_6/Component_Function_1/NAND4_in[3] ,
         \SB3_6/Component_Function_1/NAND4_in[2] ,
         \SB3_6/Component_Function_1/NAND4_in[1] ,
         \SB3_6/Component_Function_1/NAND4_in[0] ,
         \SB3_6/Component_Function_5/NAND4_in[3] ,
         \SB3_6/Component_Function_5/NAND4_in[2] ,
         \SB3_6/Component_Function_5/NAND4_in[1] ,
         \SB3_6/Component_Function_5/NAND4_in[0] ,
         \SB3_7/Component_Function_0/NAND4_in[2] ,
         \SB3_7/Component_Function_0/NAND4_in[1] ,
         \SB3_7/Component_Function_0/NAND4_in[0] ,
         \SB3_7/Component_Function_1/NAND4_in[3] ,
         \SB3_7/Component_Function_1/NAND4_in[2] ,
         \SB3_7/Component_Function_1/NAND4_in[1] ,
         \SB3_7/Component_Function_1/NAND4_in[0] ,
         \SB3_7/Component_Function_5/NAND4_in[3] ,
         \SB3_7/Component_Function_5/NAND4_in[1] ,
         \SB3_7/Component_Function_5/NAND4_in[0] ,
         \SB3_8/Component_Function_0/NAND4_in[3] ,
         \SB3_8/Component_Function_0/NAND4_in[2] ,
         \SB3_8/Component_Function_0/NAND4_in[1] ,
         \SB3_8/Component_Function_0/NAND4_in[0] ,
         \SB3_8/Component_Function_1/NAND4_in[3] ,
         \SB3_8/Component_Function_1/NAND4_in[2] ,
         \SB3_8/Component_Function_1/NAND4_in[1] ,
         \SB3_8/Component_Function_1/NAND4_in[0] ,
         \SB3_8/Component_Function_5/NAND4_in[3] ,
         \SB3_8/Component_Function_5/NAND4_in[1] ,
         \SB3_8/Component_Function_5/NAND4_in[0] ,
         \SB3_9/Component_Function_0/NAND4_in[3] ,
         \SB3_9/Component_Function_0/NAND4_in[2] ,
         \SB3_9/Component_Function_0/NAND4_in[1] ,
         \SB3_9/Component_Function_0/NAND4_in[0] ,
         \SB3_9/Component_Function_1/NAND4_in[3] ,
         \SB3_9/Component_Function_1/NAND4_in[2] ,
         \SB3_9/Component_Function_1/NAND4_in[1] ,
         \SB3_9/Component_Function_1/NAND4_in[0] ,
         \SB3_9/Component_Function_5/NAND4_in[3] ,
         \SB3_9/Component_Function_5/NAND4_in[1] ,
         \SB3_9/Component_Function_5/NAND4_in[0] ,
         \SB3_10/Component_Function_0/NAND4_in[2] ,
         \SB3_10/Component_Function_0/NAND4_in[1] ,
         \SB3_10/Component_Function_0/NAND4_in[0] ,
         \SB3_10/Component_Function_1/NAND4_in[3] ,
         \SB3_10/Component_Function_1/NAND4_in[2] ,
         \SB3_10/Component_Function_1/NAND4_in[1] ,
         \SB3_10/Component_Function_1/NAND4_in[0] ,
         \SB3_10/Component_Function_5/NAND4_in[3] ,
         \SB3_10/Component_Function_5/NAND4_in[1] ,
         \SB3_10/Component_Function_5/NAND4_in[0] ,
         \SB3_11/Component_Function_0/NAND4_in[3] ,
         \SB3_11/Component_Function_0/NAND4_in[2] ,
         \SB3_11/Component_Function_0/NAND4_in[1] ,
         \SB3_11/Component_Function_0/NAND4_in[0] ,
         \SB3_11/Component_Function_1/NAND4_in[3] ,
         \SB3_11/Component_Function_1/NAND4_in[2] ,
         \SB3_11/Component_Function_1/NAND4_in[1] ,
         \SB3_11/Component_Function_1/NAND4_in[0] ,
         \SB3_11/Component_Function_5/NAND4_in[2] ,
         \SB3_11/Component_Function_5/NAND4_in[1] ,
         \SB3_11/Component_Function_5/NAND4_in[0] ,
         \SB3_12/Component_Function_0/NAND4_in[3] ,
         \SB3_12/Component_Function_0/NAND4_in[2] ,
         \SB3_12/Component_Function_0/NAND4_in[1] ,
         \SB3_12/Component_Function_0/NAND4_in[0] ,
         \SB3_12/Component_Function_1/NAND4_in[3] ,
         \SB3_12/Component_Function_1/NAND4_in[2] ,
         \SB3_12/Component_Function_1/NAND4_in[1] ,
         \SB3_12/Component_Function_1/NAND4_in[0] ,
         \SB3_12/Component_Function_5/NAND4_in[3] ,
         \SB3_12/Component_Function_5/NAND4_in[1] ,
         \SB3_12/Component_Function_5/NAND4_in[0] ,
         \SB3_13/Component_Function_0/NAND4_in[3] ,
         \SB3_13/Component_Function_0/NAND4_in[2] ,
         \SB3_13/Component_Function_0/NAND4_in[1] ,
         \SB3_13/Component_Function_0/NAND4_in[0] ,
         \SB3_13/Component_Function_1/NAND4_in[3] ,
         \SB3_13/Component_Function_1/NAND4_in[2] ,
         \SB3_13/Component_Function_1/NAND4_in[1] ,
         \SB3_13/Component_Function_1/NAND4_in[0] ,
         \SB3_13/Component_Function_5/NAND4_in[3] ,
         \SB3_13/Component_Function_5/NAND4_in[2] ,
         \SB3_13/Component_Function_5/NAND4_in[1] ,
         \SB3_13/Component_Function_5/NAND4_in[0] ,
         \SB3_14/Component_Function_0/NAND4_in[2] ,
         \SB3_14/Component_Function_0/NAND4_in[1] ,
         \SB3_14/Component_Function_0/NAND4_in[0] ,
         \SB3_14/Component_Function_1/NAND4_in[3] ,
         \SB3_14/Component_Function_1/NAND4_in[2] ,
         \SB3_14/Component_Function_1/NAND4_in[1] ,
         \SB3_14/Component_Function_1/NAND4_in[0] ,
         \SB3_14/Component_Function_5/NAND4_in[3] ,
         \SB3_14/Component_Function_5/NAND4_in[1] ,
         \SB3_14/Component_Function_5/NAND4_in[0] ,
         \SB3_15/Component_Function_0/NAND4_in[2] ,
         \SB3_15/Component_Function_0/NAND4_in[1] ,
         \SB3_15/Component_Function_0/NAND4_in[0] ,
         \SB3_15/Component_Function_1/NAND4_in[3] ,
         \SB3_15/Component_Function_1/NAND4_in[2] ,
         \SB3_15/Component_Function_1/NAND4_in[1] ,
         \SB3_15/Component_Function_1/NAND4_in[0] ,
         \SB3_15/Component_Function_5/NAND4_in[3] ,
         \SB3_15/Component_Function_5/NAND4_in[1] ,
         \SB3_15/Component_Function_5/NAND4_in[0] ,
         \SB3_16/Component_Function_0/NAND4_in[3] ,
         \SB3_16/Component_Function_0/NAND4_in[2] ,
         \SB3_16/Component_Function_0/NAND4_in[1] ,
         \SB3_16/Component_Function_0/NAND4_in[0] ,
         \SB3_16/Component_Function_1/NAND4_in[3] ,
         \SB3_16/Component_Function_1/NAND4_in[2] ,
         \SB3_16/Component_Function_1/NAND4_in[1] ,
         \SB3_16/Component_Function_1/NAND4_in[0] ,
         \SB3_16/Component_Function_5/NAND4_in[3] ,
         \SB3_16/Component_Function_5/NAND4_in[1] ,
         \SB3_16/Component_Function_5/NAND4_in[0] ,
         \SB3_17/Component_Function_0/NAND4_in[2] ,
         \SB3_17/Component_Function_0/NAND4_in[1] ,
         \SB3_17/Component_Function_0/NAND4_in[0] ,
         \SB3_17/Component_Function_1/NAND4_in[3] ,
         \SB3_17/Component_Function_1/NAND4_in[2] ,
         \SB3_17/Component_Function_1/NAND4_in[1] ,
         \SB3_17/Component_Function_1/NAND4_in[0] ,
         \SB3_17/Component_Function_5/NAND4_in[3] ,
         \SB3_17/Component_Function_5/NAND4_in[1] ,
         \SB3_17/Component_Function_5/NAND4_in[0] ,
         \SB3_18/Component_Function_0/NAND4_in[2] ,
         \SB3_18/Component_Function_0/NAND4_in[1] ,
         \SB3_18/Component_Function_0/NAND4_in[0] ,
         \SB3_18/Component_Function_1/NAND4_in[3] ,
         \SB3_18/Component_Function_1/NAND4_in[2] ,
         \SB3_18/Component_Function_1/NAND4_in[1] ,
         \SB3_18/Component_Function_1/NAND4_in[0] ,
         \SB3_18/Component_Function_5/NAND4_in[2] ,
         \SB3_18/Component_Function_5/NAND4_in[1] ,
         \SB3_18/Component_Function_5/NAND4_in[0] ,
         \SB3_19/Component_Function_0/NAND4_in[3] ,
         \SB3_19/Component_Function_0/NAND4_in[2] ,
         \SB3_19/Component_Function_0/NAND4_in[1] ,
         \SB3_19/Component_Function_0/NAND4_in[0] ,
         \SB3_19/Component_Function_1/NAND4_in[3] ,
         \SB3_19/Component_Function_1/NAND4_in[2] ,
         \SB3_19/Component_Function_1/NAND4_in[1] ,
         \SB3_19/Component_Function_1/NAND4_in[0] ,
         \SB3_19/Component_Function_5/NAND4_in[2] ,
         \SB3_19/Component_Function_5/NAND4_in[1] ,
         \SB3_19/Component_Function_5/NAND4_in[0] ,
         \SB3_20/Component_Function_0/NAND4_in[3] ,
         \SB3_20/Component_Function_0/NAND4_in[2] ,
         \SB3_20/Component_Function_0/NAND4_in[1] ,
         \SB3_20/Component_Function_0/NAND4_in[0] ,
         \SB3_20/Component_Function_1/NAND4_in[3] ,
         \SB3_20/Component_Function_1/NAND4_in[2] ,
         \SB3_20/Component_Function_1/NAND4_in[1] ,
         \SB3_20/Component_Function_1/NAND4_in[0] ,
         \SB3_20/Component_Function_5/NAND4_in[3] ,
         \SB3_20/Component_Function_5/NAND4_in[1] ,
         \SB3_20/Component_Function_5/NAND4_in[0] ,
         \SB3_21/Component_Function_0/NAND4_in[3] ,
         \SB3_21/Component_Function_0/NAND4_in[2] ,
         \SB3_21/Component_Function_0/NAND4_in[1] ,
         \SB3_21/Component_Function_0/NAND4_in[0] ,
         \SB3_21/Component_Function_1/NAND4_in[2] ,
         \SB3_21/Component_Function_1/NAND4_in[1] ,
         \SB3_21/Component_Function_1/NAND4_in[0] ,
         \SB3_21/Component_Function_5/NAND4_in[3] ,
         \SB3_21/Component_Function_5/NAND4_in[1] ,
         \SB3_21/Component_Function_5/NAND4_in[0] ,
         \SB3_22/Component_Function_0/NAND4_in[2] ,
         \SB3_22/Component_Function_0/NAND4_in[1] ,
         \SB3_22/Component_Function_0/NAND4_in[0] ,
         \SB3_22/Component_Function_1/NAND4_in[3] ,
         \SB3_22/Component_Function_1/NAND4_in[2] ,
         \SB3_22/Component_Function_1/NAND4_in[1] ,
         \SB3_22/Component_Function_1/NAND4_in[0] ,
         \SB3_22/Component_Function_5/NAND4_in[3] ,
         \SB3_22/Component_Function_5/NAND4_in[2] ,
         \SB3_22/Component_Function_5/NAND4_in[1] ,
         \SB3_22/Component_Function_5/NAND4_in[0] ,
         \SB3_23/Component_Function_0/NAND4_in[3] ,
         \SB3_23/Component_Function_0/NAND4_in[2] ,
         \SB3_23/Component_Function_0/NAND4_in[1] ,
         \SB3_23/Component_Function_0/NAND4_in[0] ,
         \SB3_23/Component_Function_1/NAND4_in[3] ,
         \SB3_23/Component_Function_1/NAND4_in[2] ,
         \SB3_23/Component_Function_1/NAND4_in[1] ,
         \SB3_23/Component_Function_1/NAND4_in[0] ,
         \SB3_23/Component_Function_5/NAND4_in[3] ,
         \SB3_23/Component_Function_5/NAND4_in[1] ,
         \SB3_23/Component_Function_5/NAND4_in[0] ,
         \SB3_24/Component_Function_0/NAND4_in[2] ,
         \SB3_24/Component_Function_0/NAND4_in[1] ,
         \SB3_24/Component_Function_0/NAND4_in[0] ,
         \SB3_24/Component_Function_1/NAND4_in[3] ,
         \SB3_24/Component_Function_1/NAND4_in[2] ,
         \SB3_24/Component_Function_1/NAND4_in[1] ,
         \SB3_24/Component_Function_1/NAND4_in[0] ,
         \SB3_24/Component_Function_5/NAND4_in[3] ,
         \SB3_24/Component_Function_5/NAND4_in[1] ,
         \SB3_24/Component_Function_5/NAND4_in[0] ,
         \SB3_25/Component_Function_0/NAND4_in[3] ,
         \SB3_25/Component_Function_0/NAND4_in[2] ,
         \SB3_25/Component_Function_0/NAND4_in[1] ,
         \SB3_25/Component_Function_0/NAND4_in[0] ,
         \SB3_25/Component_Function_1/NAND4_in[3] ,
         \SB3_25/Component_Function_1/NAND4_in[2] ,
         \SB3_25/Component_Function_1/NAND4_in[1] ,
         \SB3_25/Component_Function_1/NAND4_in[0] ,
         \SB3_25/Component_Function_5/NAND4_in[2] ,
         \SB3_25/Component_Function_5/NAND4_in[1] ,
         \SB3_25/Component_Function_5/NAND4_in[0] ,
         \SB3_26/Component_Function_0/NAND4_in[2] ,
         \SB3_26/Component_Function_0/NAND4_in[1] ,
         \SB3_26/Component_Function_0/NAND4_in[0] ,
         \SB3_26/Component_Function_1/NAND4_in[3] ,
         \SB3_26/Component_Function_1/NAND4_in[2] ,
         \SB3_26/Component_Function_1/NAND4_in[1] ,
         \SB3_26/Component_Function_1/NAND4_in[0] ,
         \SB3_26/Component_Function_5/NAND4_in[3] ,
         \SB3_26/Component_Function_5/NAND4_in[1] ,
         \SB3_26/Component_Function_5/NAND4_in[0] ,
         \SB3_27/Component_Function_0/NAND4_in[2] ,
         \SB3_27/Component_Function_0/NAND4_in[1] ,
         \SB3_27/Component_Function_0/NAND4_in[0] ,
         \SB3_27/Component_Function_1/NAND4_in[3] ,
         \SB3_27/Component_Function_1/NAND4_in[2] ,
         \SB3_27/Component_Function_1/NAND4_in[1] ,
         \SB3_27/Component_Function_1/NAND4_in[0] ,
         \SB3_27/Component_Function_5/NAND4_in[3] ,
         \SB3_27/Component_Function_5/NAND4_in[1] ,
         \SB3_27/Component_Function_5/NAND4_in[0] ,
         \SB3_28/Component_Function_0/NAND4_in[3] ,
         \SB3_28/Component_Function_0/NAND4_in[2] ,
         \SB3_28/Component_Function_0/NAND4_in[1] ,
         \SB3_28/Component_Function_0/NAND4_in[0] ,
         \SB3_28/Component_Function_1/NAND4_in[3] ,
         \SB3_28/Component_Function_1/NAND4_in[2] ,
         \SB3_28/Component_Function_1/NAND4_in[1] ,
         \SB3_28/Component_Function_1/NAND4_in[0] ,
         \SB3_28/Component_Function_5/NAND4_in[3] ,
         \SB3_28/Component_Function_5/NAND4_in[1] ,
         \SB3_28/Component_Function_5/NAND4_in[0] ,
         \SB3_29/Component_Function_0/NAND4_in[2] ,
         \SB3_29/Component_Function_0/NAND4_in[1] ,
         \SB3_29/Component_Function_0/NAND4_in[0] ,
         \SB3_29/Component_Function_1/NAND4_in[3] ,
         \SB3_29/Component_Function_1/NAND4_in[2] ,
         \SB3_29/Component_Function_1/NAND4_in[1] ,
         \SB3_29/Component_Function_1/NAND4_in[0] ,
         \SB3_29/Component_Function_5/NAND4_in[3] ,
         \SB3_29/Component_Function_5/NAND4_in[1] ,
         \SB3_29/Component_Function_5/NAND4_in[0] ,
         \SB3_30/Component_Function_0/NAND4_in[3] ,
         \SB3_30/Component_Function_0/NAND4_in[2] ,
         \SB3_30/Component_Function_0/NAND4_in[1] ,
         \SB3_30/Component_Function_0/NAND4_in[0] ,
         \SB3_30/Component_Function_1/NAND4_in[3] ,
         \SB3_30/Component_Function_1/NAND4_in[2] ,
         \SB3_30/Component_Function_1/NAND4_in[1] ,
         \SB3_30/Component_Function_1/NAND4_in[0] ,
         \SB3_30/Component_Function_5/NAND4_in[3] ,
         \SB3_30/Component_Function_5/NAND4_in[1] ,
         \SB3_30/Component_Function_5/NAND4_in[0] ,
         \SB3_31/Component_Function_0/NAND4_in[3] ,
         \SB3_31/Component_Function_0/NAND4_in[2] ,
         \SB3_31/Component_Function_0/NAND4_in[1] ,
         \SB3_31/Component_Function_0/NAND4_in[0] ,
         \SB3_31/Component_Function_1/NAND4_in[3] ,
         \SB3_31/Component_Function_1/NAND4_in[2] ,
         \SB3_31/Component_Function_1/NAND4_in[1] ,
         \SB3_31/Component_Function_1/NAND4_in[0] ,
         \SB3_31/Component_Function_5/NAND4_in[3] ,
         \SB3_31/Component_Function_5/NAND4_in[2] ,
         \SB3_31/Component_Function_5/NAND4_in[1] ,
         \SB3_31/Component_Function_5/NAND4_in[0] ,
         \SB4_0/Component_Function_0/NAND4_in[3] ,
         \SB4_0/Component_Function_0/NAND4_in[2] ,
         \SB4_0/Component_Function_0/NAND4_in[1] ,
         \SB4_0/Component_Function_0/NAND4_in[0] ,
         \SB4_0/Component_Function_1/NAND4_in[3] ,
         \SB4_0/Component_Function_1/NAND4_in[1] ,
         \SB4_0/Component_Function_1/NAND4_in[0] ,
         \SB4_0/Component_Function_5/NAND4_in[3] ,
         \SB4_0/Component_Function_5/NAND4_in[2] ,
         \SB4_0/Component_Function_5/NAND4_in[1] ,
         \SB4_0/Component_Function_5/NAND4_in[0] ,
         \SB4_1/Component_Function_0/NAND4_in[3] ,
         \SB4_1/Component_Function_0/NAND4_in[2] ,
         \SB4_1/Component_Function_0/NAND4_in[1] ,
         \SB4_1/Component_Function_0/NAND4_in[0] ,
         \SB4_1/Component_Function_1/NAND4_in[2] ,
         \SB4_1/Component_Function_1/NAND4_in[1] ,
         \SB4_1/Component_Function_1/NAND4_in[0] ,
         \SB4_1/Component_Function_5/NAND4_in[3] ,
         \SB4_1/Component_Function_5/NAND4_in[2] ,
         \SB4_1/Component_Function_5/NAND4_in[0] ,
         \SB4_2/Component_Function_0/NAND4_in[3] ,
         \SB4_2/Component_Function_0/NAND4_in[2] ,
         \SB4_2/Component_Function_0/NAND4_in[1] ,
         \SB4_2/Component_Function_0/NAND4_in[0] ,
         \SB4_2/Component_Function_1/NAND4_in[2] ,
         \SB4_2/Component_Function_1/NAND4_in[1] ,
         \SB4_2/Component_Function_1/NAND4_in[0] ,
         \SB4_2/Component_Function_5/NAND4_in[3] ,
         \SB4_2/Component_Function_5/NAND4_in[2] ,
         \SB4_2/Component_Function_5/NAND4_in[0] ,
         \SB4_3/Component_Function_0/NAND4_in[3] ,
         \SB4_3/Component_Function_0/NAND4_in[2] ,
         \SB4_3/Component_Function_0/NAND4_in[0] ,
         \SB4_3/Component_Function_1/NAND4_in[1] ,
         \SB4_3/Component_Function_1/NAND4_in[0] ,
         \SB4_3/Component_Function_5/NAND4_in[3] ,
         \SB4_3/Component_Function_5/NAND4_in[2] ,
         \SB4_3/Component_Function_5/NAND4_in[0] ,
         \SB4_4/Component_Function_0/NAND4_in[3] ,
         \SB4_4/Component_Function_0/NAND4_in[2] ,
         \SB4_4/Component_Function_0/NAND4_in[0] ,
         \SB4_4/Component_Function_1/NAND4_in[3] ,
         \SB4_4/Component_Function_1/NAND4_in[1] ,
         \SB4_4/Component_Function_1/NAND4_in[0] ,
         \SB4_4/Component_Function_5/NAND4_in[2] ,
         \SB4_4/Component_Function_5/NAND4_in[1] ,
         \SB4_4/Component_Function_5/NAND4_in[0] ,
         \SB4_5/Component_Function_0/NAND4_in[3] ,
         \SB4_5/Component_Function_0/NAND4_in[2] ,
         \SB4_5/Component_Function_0/NAND4_in[1] ,
         \SB4_5/Component_Function_0/NAND4_in[0] ,
         \SB4_5/Component_Function_1/NAND4_in[2] ,
         \SB4_5/Component_Function_1/NAND4_in[1] ,
         \SB4_5/Component_Function_1/NAND4_in[0] ,
         \SB4_5/Component_Function_5/NAND4_in[3] ,
         \SB4_5/Component_Function_5/NAND4_in[2] ,
         \SB4_5/Component_Function_5/NAND4_in[1] ,
         \SB4_5/Component_Function_5/NAND4_in[0] ,
         \SB4_6/Component_Function_0/NAND4_in[3] ,
         \SB4_6/Component_Function_0/NAND4_in[2] ,
         \SB4_6/Component_Function_0/NAND4_in[1] ,
         \SB4_6/Component_Function_0/NAND4_in[0] ,
         \SB4_6/Component_Function_1/NAND4_in[3] ,
         \SB4_6/Component_Function_1/NAND4_in[2] ,
         \SB4_6/Component_Function_1/NAND4_in[1] ,
         \SB4_6/Component_Function_1/NAND4_in[0] ,
         \SB4_6/Component_Function_5/NAND4_in[3] ,
         \SB4_6/Component_Function_5/NAND4_in[2] ,
         \SB4_6/Component_Function_5/NAND4_in[1] ,
         \SB4_6/Component_Function_5/NAND4_in[0] ,
         \SB4_7/Component_Function_0/NAND4_in[3] ,
         \SB4_7/Component_Function_0/NAND4_in[2] ,
         \SB4_7/Component_Function_0/NAND4_in[1] ,
         \SB4_7/Component_Function_0/NAND4_in[0] ,
         \SB4_7/Component_Function_1/NAND4_in[1] ,
         \SB4_7/Component_Function_1/NAND4_in[0] ,
         \SB4_7/Component_Function_5/NAND4_in[3] ,
         \SB4_7/Component_Function_5/NAND4_in[0] ,
         \SB4_8/Component_Function_0/NAND4_in[3] ,
         \SB4_8/Component_Function_0/NAND4_in[2] ,
         \SB4_8/Component_Function_0/NAND4_in[1] ,
         \SB4_8/Component_Function_0/NAND4_in[0] ,
         \SB4_8/Component_Function_1/NAND4_in[1] ,
         \SB4_8/Component_Function_1/NAND4_in[0] ,
         \SB4_8/Component_Function_5/NAND4_in[3] ,
         \SB4_8/Component_Function_5/NAND4_in[2] ,
         \SB4_8/Component_Function_5/NAND4_in[1] ,
         \SB4_8/Component_Function_5/NAND4_in[0] ,
         \SB4_9/Component_Function_0/NAND4_in[3] ,
         \SB4_9/Component_Function_0/NAND4_in[2] ,
         \SB4_9/Component_Function_0/NAND4_in[1] ,
         \SB4_9/Component_Function_0/NAND4_in[0] ,
         \SB4_9/Component_Function_1/NAND4_in[3] ,
         \SB4_9/Component_Function_1/NAND4_in[2] ,
         \SB4_9/Component_Function_1/NAND4_in[1] ,
         \SB4_9/Component_Function_1/NAND4_in[0] ,
         \SB4_9/Component_Function_5/NAND4_in[3] ,
         \SB4_9/Component_Function_5/NAND4_in[2] ,
         \SB4_9/Component_Function_5/NAND4_in[1] ,
         \SB4_9/Component_Function_5/NAND4_in[0] ,
         \SB4_10/Component_Function_0/NAND4_in[3] ,
         \SB4_10/Component_Function_0/NAND4_in[2] ,
         \SB4_10/Component_Function_0/NAND4_in[1] ,
         \SB4_10/Component_Function_0/NAND4_in[0] ,
         \SB4_10/Component_Function_1/NAND4_in[2] ,
         \SB4_10/Component_Function_1/NAND4_in[1] ,
         \SB4_10/Component_Function_1/NAND4_in[0] ,
         \SB4_10/Component_Function_5/NAND4_in[3] ,
         \SB4_10/Component_Function_5/NAND4_in[2] ,
         \SB4_10/Component_Function_5/NAND4_in[1] ,
         \SB4_10/Component_Function_5/NAND4_in[0] ,
         \SB4_11/Component_Function_0/NAND4_in[3] ,
         \SB4_11/Component_Function_0/NAND4_in[2] ,
         \SB4_11/Component_Function_0/NAND4_in[0] ,
         \SB4_11/Component_Function_1/NAND4_in[2] ,
         \SB4_11/Component_Function_1/NAND4_in[1] ,
         \SB4_11/Component_Function_1/NAND4_in[0] ,
         \SB4_11/Component_Function_5/NAND4_in[3] ,
         \SB4_11/Component_Function_5/NAND4_in[2] ,
         \SB4_11/Component_Function_5/NAND4_in[1] ,
         \SB4_11/Component_Function_5/NAND4_in[0] ,
         \SB4_12/Component_Function_0/NAND4_in[3] ,
         \SB4_12/Component_Function_0/NAND4_in[2] ,
         \SB4_12/Component_Function_0/NAND4_in[1] ,
         \SB4_12/Component_Function_0/NAND4_in[0] ,
         \SB4_12/Component_Function_1/NAND4_in[2] ,
         \SB4_12/Component_Function_1/NAND4_in[1] ,
         \SB4_12/Component_Function_1/NAND4_in[0] ,
         \SB4_12/Component_Function_5/NAND4_in[3] ,
         \SB4_12/Component_Function_5/NAND4_in[2] ,
         \SB4_12/Component_Function_5/NAND4_in[1] ,
         \SB4_12/Component_Function_5/NAND4_in[0] ,
         \SB4_13/Component_Function_0/NAND4_in[3] ,
         \SB4_13/Component_Function_0/NAND4_in[2] ,
         \SB4_13/Component_Function_0/NAND4_in[0] ,
         \SB4_13/Component_Function_1/NAND4_in[3] ,
         \SB4_13/Component_Function_1/NAND4_in[2] ,
         \SB4_13/Component_Function_1/NAND4_in[1] ,
         \SB4_13/Component_Function_1/NAND4_in[0] ,
         \SB4_13/Component_Function_5/NAND4_in[3] ,
         \SB4_13/Component_Function_5/NAND4_in[2] ,
         \SB4_13/Component_Function_5/NAND4_in[1] ,
         \SB4_13/Component_Function_5/NAND4_in[0] ,
         \SB4_14/Component_Function_0/NAND4_in[3] ,
         \SB4_14/Component_Function_0/NAND4_in[2] ,
         \SB4_14/Component_Function_0/NAND4_in[1] ,
         \SB4_14/Component_Function_0/NAND4_in[0] ,
         \SB4_14/Component_Function_1/NAND4_in[2] ,
         \SB4_14/Component_Function_1/NAND4_in[1] ,
         \SB4_14/Component_Function_1/NAND4_in[0] ,
         \SB4_14/Component_Function_5/NAND4_in[3] ,
         \SB4_14/Component_Function_5/NAND4_in[2] ,
         \SB4_14/Component_Function_5/NAND4_in[0] ,
         \SB4_15/Component_Function_0/NAND4_in[3] ,
         \SB4_15/Component_Function_0/NAND4_in[2] ,
         \SB4_15/Component_Function_0/NAND4_in[1] ,
         \SB4_15/Component_Function_0/NAND4_in[0] ,
         \SB4_15/Component_Function_1/NAND4_in[3] ,
         \SB4_15/Component_Function_1/NAND4_in[1] ,
         \SB4_15/Component_Function_1/NAND4_in[0] ,
         \SB4_15/Component_Function_5/NAND4_in[2] ,
         \SB4_15/Component_Function_5/NAND4_in[0] ,
         \SB4_16/Component_Function_0/NAND4_in[3] ,
         \SB4_16/Component_Function_0/NAND4_in[2] ,
         \SB4_16/Component_Function_0/NAND4_in[0] ,
         \SB4_16/Component_Function_1/NAND4_in[2] ,
         \SB4_16/Component_Function_1/NAND4_in[1] ,
         \SB4_16/Component_Function_1/NAND4_in[0] ,
         \SB4_16/Component_Function_5/NAND4_in[3] ,
         \SB4_16/Component_Function_5/NAND4_in[2] ,
         \SB4_16/Component_Function_5/NAND4_in[1] ,
         \SB4_16/Component_Function_5/NAND4_in[0] ,
         \SB4_17/Component_Function_0/NAND4_in[3] ,
         \SB4_17/Component_Function_0/NAND4_in[2] ,
         \SB4_17/Component_Function_0/NAND4_in[1] ,
         \SB4_17/Component_Function_0/NAND4_in[0] ,
         \SB4_17/Component_Function_1/NAND4_in[3] ,
         \SB4_17/Component_Function_1/NAND4_in[2] ,
         \SB4_17/Component_Function_1/NAND4_in[1] ,
         \SB4_17/Component_Function_1/NAND4_in[0] ,
         \SB4_17/Component_Function_5/NAND4_in[3] ,
         \SB4_17/Component_Function_5/NAND4_in[1] ,
         \SB4_17/Component_Function_5/NAND4_in[0] ,
         \SB4_18/Component_Function_0/NAND4_in[3] ,
         \SB4_18/Component_Function_0/NAND4_in[2] ,
         \SB4_18/Component_Function_0/NAND4_in[1] ,
         \SB4_18/Component_Function_0/NAND4_in[0] ,
         \SB4_18/Component_Function_1/NAND4_in[3] ,
         \SB4_18/Component_Function_1/NAND4_in[2] ,
         \SB4_18/Component_Function_1/NAND4_in[1] ,
         \SB4_18/Component_Function_1/NAND4_in[0] ,
         \SB4_18/Component_Function_5/NAND4_in[3] ,
         \SB4_18/Component_Function_5/NAND4_in[2] ,
         \SB4_18/Component_Function_5/NAND4_in[0] ,
         \SB4_19/Component_Function_0/NAND4_in[3] ,
         \SB4_19/Component_Function_0/NAND4_in[2] ,
         \SB4_19/Component_Function_0/NAND4_in[1] ,
         \SB4_19/Component_Function_0/NAND4_in[0] ,
         \SB4_19/Component_Function_1/NAND4_in[3] ,
         \SB4_19/Component_Function_1/NAND4_in[2] ,
         \SB4_19/Component_Function_1/NAND4_in[1] ,
         \SB4_19/Component_Function_1/NAND4_in[0] ,
         \SB4_19/Component_Function_5/NAND4_in[3] ,
         \SB4_19/Component_Function_5/NAND4_in[2] ,
         \SB4_19/Component_Function_5/NAND4_in[1] ,
         \SB4_19/Component_Function_5/NAND4_in[0] ,
         \SB4_20/Component_Function_0/NAND4_in[3] ,
         \SB4_20/Component_Function_0/NAND4_in[2] ,
         \SB4_20/Component_Function_0/NAND4_in[0] ,
         \SB4_20/Component_Function_1/NAND4_in[3] ,
         \SB4_20/Component_Function_1/NAND4_in[1] ,
         \SB4_20/Component_Function_1/NAND4_in[0] ,
         \SB4_20/Component_Function_5/NAND4_in[3] ,
         \SB4_20/Component_Function_5/NAND4_in[2] ,
         \SB4_20/Component_Function_5/NAND4_in[1] ,
         \SB4_20/Component_Function_5/NAND4_in[0] ,
         \SB4_21/Component_Function_0/NAND4_in[3] ,
         \SB4_21/Component_Function_0/NAND4_in[2] ,
         \SB4_21/Component_Function_0/NAND4_in[0] ,
         \SB4_21/Component_Function_1/NAND4_in[1] ,
         \SB4_21/Component_Function_1/NAND4_in[0] ,
         \SB4_21/Component_Function_5/NAND4_in[2] ,
         \SB4_21/Component_Function_5/NAND4_in[1] ,
         \SB4_21/Component_Function_5/NAND4_in[0] ,
         \SB4_22/Component_Function_0/NAND4_in[3] ,
         \SB4_22/Component_Function_0/NAND4_in[2] ,
         \SB4_22/Component_Function_0/NAND4_in[1] ,
         \SB4_22/Component_Function_0/NAND4_in[0] ,
         \SB4_22/Component_Function_1/NAND4_in[3] ,
         \SB4_22/Component_Function_1/NAND4_in[1] ,
         \SB4_22/Component_Function_1/NAND4_in[0] ,
         \SB4_22/Component_Function_5/NAND4_in[3] ,
         \SB4_22/Component_Function_5/NAND4_in[2] ,
         \SB4_22/Component_Function_5/NAND4_in[1] ,
         \SB4_22/Component_Function_5/NAND4_in[0] ,
         \SB4_23/Component_Function_0/NAND4_in[3] ,
         \SB4_23/Component_Function_0/NAND4_in[2] ,
         \SB4_23/Component_Function_0/NAND4_in[1] ,
         \SB4_23/Component_Function_0/NAND4_in[0] ,
         \SB4_23/Component_Function_1/NAND4_in[3] ,
         \SB4_23/Component_Function_1/NAND4_in[2] ,
         \SB4_23/Component_Function_1/NAND4_in[1] ,
         \SB4_23/Component_Function_1/NAND4_in[0] ,
         \SB4_23/Component_Function_5/NAND4_in[3] ,
         \SB4_23/Component_Function_5/NAND4_in[2] ,
         \SB4_23/Component_Function_5/NAND4_in[1] ,
         \SB4_23/Component_Function_5/NAND4_in[0] ,
         \SB4_24/Component_Function_0/NAND4_in[3] ,
         \SB4_24/Component_Function_0/NAND4_in[2] ,
         \SB4_24/Component_Function_0/NAND4_in[0] ,
         \SB4_24/Component_Function_1/NAND4_in[3] ,
         \SB4_24/Component_Function_1/NAND4_in[1] ,
         \SB4_24/Component_Function_1/NAND4_in[0] ,
         \SB4_24/Component_Function_5/NAND4_in[3] ,
         \SB4_24/Component_Function_5/NAND4_in[2] ,
         \SB4_24/Component_Function_5/NAND4_in[1] ,
         \SB4_24/Component_Function_5/NAND4_in[0] ,
         \SB4_25/Component_Function_0/NAND4_in[3] ,
         \SB4_25/Component_Function_0/NAND4_in[2] ,
         \SB4_25/Component_Function_0/NAND4_in[1] ,
         \SB4_25/Component_Function_0/NAND4_in[0] ,
         \SB4_25/Component_Function_1/NAND4_in[3] ,
         \SB4_25/Component_Function_1/NAND4_in[1] ,
         \SB4_25/Component_Function_1/NAND4_in[0] ,
         \SB4_25/Component_Function_5/NAND4_in[3] ,
         \SB4_25/Component_Function_5/NAND4_in[2] ,
         \SB4_25/Component_Function_5/NAND4_in[1] ,
         \SB4_25/Component_Function_5/NAND4_in[0] ,
         \SB4_26/Component_Function_0/NAND4_in[3] ,
         \SB4_26/Component_Function_0/NAND4_in[2] ,
         \SB4_26/Component_Function_0/NAND4_in[0] ,
         \SB4_26/Component_Function_1/NAND4_in[3] ,
         \SB4_26/Component_Function_1/NAND4_in[2] ,
         \SB4_26/Component_Function_1/NAND4_in[1] ,
         \SB4_26/Component_Function_1/NAND4_in[0] ,
         \SB4_26/Component_Function_5/NAND4_in[3] ,
         \SB4_26/Component_Function_5/NAND4_in[2] ,
         \SB4_26/Component_Function_5/NAND4_in[0] ,
         \SB4_27/Component_Function_0/NAND4_in[3] ,
         \SB4_27/Component_Function_0/NAND4_in[2] ,
         \SB4_27/Component_Function_0/NAND4_in[1] ,
         \SB4_27/Component_Function_0/NAND4_in[0] ,
         \SB4_27/Component_Function_1/NAND4_in[2] ,
         \SB4_27/Component_Function_1/NAND4_in[1] ,
         \SB4_27/Component_Function_1/NAND4_in[0] ,
         \SB4_27/Component_Function_5/NAND4_in[3] ,
         \SB4_27/Component_Function_5/NAND4_in[2] ,
         \SB4_27/Component_Function_5/NAND4_in[1] ,
         \SB4_27/Component_Function_5/NAND4_in[0] ,
         \SB4_28/Component_Function_0/NAND4_in[3] ,
         \SB4_28/Component_Function_0/NAND4_in[2] ,
         \SB4_28/Component_Function_0/NAND4_in[1] ,
         \SB4_28/Component_Function_0/NAND4_in[0] ,
         \SB4_28/Component_Function_1/NAND4_in[2] ,
         \SB4_28/Component_Function_1/NAND4_in[1] ,
         \SB4_28/Component_Function_1/NAND4_in[0] ,
         \SB4_28/Component_Function_5/NAND4_in[3] ,
         \SB4_28/Component_Function_5/NAND4_in[2] ,
         \SB4_28/Component_Function_5/NAND4_in[1] ,
         \SB4_28/Component_Function_5/NAND4_in[0] ,
         \SB4_29/Component_Function_0/NAND4_in[3] ,
         \SB4_29/Component_Function_0/NAND4_in[2] ,
         \SB4_29/Component_Function_0/NAND4_in[1] ,
         \SB4_29/Component_Function_0/NAND4_in[0] ,
         \SB4_29/Component_Function_1/NAND4_in[3] ,
         \SB4_29/Component_Function_1/NAND4_in[1] ,
         \SB4_29/Component_Function_1/NAND4_in[0] ,
         \SB4_29/Component_Function_5/NAND4_in[2] ,
         \SB4_29/Component_Function_5/NAND4_in[1] ,
         \SB4_29/Component_Function_5/NAND4_in[0] ,
         \SB4_30/Component_Function_0/NAND4_in[3] ,
         \SB4_30/Component_Function_0/NAND4_in[2] ,
         \SB4_30/Component_Function_0/NAND4_in[0] ,
         \SB4_30/Component_Function_1/NAND4_in[3] ,
         \SB4_30/Component_Function_1/NAND4_in[2] ,
         \SB4_30/Component_Function_1/NAND4_in[1] ,
         \SB4_30/Component_Function_1/NAND4_in[0] ,
         \SB4_30/Component_Function_5/NAND4_in[2] ,
         \SB4_30/Component_Function_5/NAND4_in[1] ,
         \SB4_30/Component_Function_5/NAND4_in[0] ,
         \SB4_31/Component_Function_0/NAND4_in[3] ,
         \SB4_31/Component_Function_0/NAND4_in[0] ,
         \SB4_31/Component_Function_1/NAND4_in[2] ,
         \SB4_31/Component_Function_1/NAND4_in[1] ,
         \SB4_31/Component_Function_1/NAND4_in[0] ,
         \SB4_31/Component_Function_5/NAND4_in[3] ,
         \SB4_31/Component_Function_5/NAND4_in[2] ,
         \SB4_31/Component_Function_5/NAND4_in[1] ,
         \SB4_31/Component_Function_5/NAND4_in[0] , n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n421, n422, n423, n424, n427,
         n428, n430, n431, n432, n433, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n517, n519,
         n520, n521, n546, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n561, n563, n565, n566, n567, n568, n569, n573, n574,
         n578, n579, n580, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n595, n596, n598, n599, n600, n601, n603,
         n604, n605, n609, n611, n613, n615, n616, n617, n618, n619, n620,
         n621, n623, n625, n627, n631, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n644, n645, n646, n647, n650, n652, n653,
         n654, n655, n656, n657, n658, n660, n661, n662, n663, n664, n666,
         n667, n668, n669, n670, n671, n672, n676, n679, n680, n681, n682,
         n683, n684, n685, n686, n688, n689, n690, n691, n693, n695, n696,
         n697, n699, n700, n701, n703, n704, n705, n706, n707, n708, n709,
         n711, n713, n718, n720, n721, n722, n723, n724, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n740, n741, n743,
         n744, n745, n747, n750, n751, n754, n755, n756, n757, n758, n761,
         n762, n763, n764, n765, n767, n769, n771, n772, n773, n774, n776,
         n777, n778, n779, n780, n781, n782, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n821, n822,
         n823, n824, n826, n827, n828, n829, n830, n831, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n880, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n899, n900, n902, n903, n904, n906, n907, n908, n909,
         n912, n914, n915, n917, n919, n920, n922, n923, n924, n925, n926,
         n927, n928, n929, n932, n934, n936, n937, n938, n939, n940, n941,
         n942, n944, n945, n946, n947, n948, n949, n950, n951, n952, n954,
         n955, n956, n957, n958, n959, n960, n961, n963, n964, n965, n966,
         n967, n970, n972, n973, n974, n975, n976, n977, n978, n980, n981,
         n984, n986, n987, n988, n991, n992, n993, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1014, n1015, n1016, n1017, n1020, n1024, n1025, n1026,
         n1028, n1030, n1031, n1032, n1033, n1035, n1036, n1038, n1039, n1040,
         n1041, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1079, n1080, n1081, n1083, n1085, n1086, n1087, n1088,
         n1089, n1090, n1092, n1094, n1095, n1096, n1099, n1100, n1101, n1102,
         n1104, n1105, n1107, n1108, n1109, n1110, n1113, n1114, n1116, n1117,
         n1118, n1119, n1121, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1134, n1135, n1136, n1137, n1138, n1140, n1141,
         n1144, n1145, n1146, n1148, n1151, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1164, n1165, n1166, n1167, n1169,
         n1170, n1171, n1172, n1174, n1175, n1178, n1180, n1182, n1184, n1185,
         n1187, n1188, n1189, n1190, n1191, n1193, n1194, n1196, n1197, n1198,
         n1199, n1200, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1217, n1219, n1220, n1221,
         n1222, n1223, n1225, n1227, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1250, n1252, n1253, n1254, n1255, n1257, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1295, n1296, n1297, n1298, n1299, n1300, n1303, n1304, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1318,
         n1319, n1320, n1322, n1323, n1325, n1326, n1327, n1328, n1329, n1332,
         n1333, n1335, n1336, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1361, n1363, n1364, n1365, n1366, n1367, n1370, n1371,
         n1375, n1376, n1377, n1378, n1380, n1382, n1383, n1385, n1386, n1389,
         n1390, n1391, n1392, n1393, n1394, n1397, n1398, n1399, n1401, n1404,
         n1406, n1407, n1408, n1411, n1414, n1416, n1417, n1418, n1419, n1422,
         n1423, n1424, n1426, n1428, n1429, n1431, n1432, n1434, n1435, n1436,
         n1437, n1438, n1440, n1441, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1453, n1454, n1455, n1457, n1458, n1459, n1460, n1462, n1463,
         n1465, n1466, n1467, n1470, n1473, n1474, n1475, n1480, n1483, n1486,
         n1495, n1497, n1498, n1501, n1502, n1503, n1505, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1522, n1523, n1524, n1525, n1526, n1527, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1569, n1570, n1571, n1572, n1573, n1575,
         n1576, n1577, n1578, n1579, n1581, n1582, n1583, n1584, n1585, n1586,
         n1588, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1604, n1605, n1607, n1608, n1609, n1610, n1611, n1612,
         n1614, n1615, n1616, n1617, n1619, n1620, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1691, n1692, n1693, n1694, n1696, n1697, n1698,
         n1700, n1702, n1703, n1704, n1705, n1706, n1709, n1711, n1712, n1714,
         n1715, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1747, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1761, n1763, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1786, n1787, n1788, n1789, n1790, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1836, n1837, n1838, n1839,
         n1840, n1841, n1843, n1844, n1845, n1846, n1847, n1849, n1850, n1851,
         n1852, n1853, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1884,
         n1885, n1886, n1887, n1888, n1889, n1891, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244;

  NAND3_X1 \SB1_0_0/Component_Function_2/N4  ( .A1(n380), .A2(\SB1_0_0/i0_0 ), 
        .A3(\SB1_0_0/i0_4 ), .ZN(\SB1_0_0/Component_Function_2/NAND4_in[3] )
         );
  NAND3_X1 \SB1_0_0/Component_Function_2/N2  ( .A1(\SB1_0_0/i0_3 ), .A2(
        \SB1_0_0/i0[10] ), .A3(\SB1_0_0/i0[6] ), .ZN(
        \SB1_0_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_0/Component_Function_2/N1  ( .A1(n380), .A2(\SB1_0_0/i0[10] ), .A3(\SB1_0_0/i1[9] ), .ZN(\SB1_0_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_0/Component_Function_3/N4  ( .A1(n380), .A2(\SB1_0_0/i0[8] ), 
        .A3(\SB1_0_0/i3[0] ), .ZN(\SB1_0_0/Component_Function_3/NAND4_in[3] )
         );
  NAND3_X1 \SB1_0_0/Component_Function_3/N1  ( .A1(\SB1_0_0/i1[9] ), .A2(
        \SB1_0_0/i0_3 ), .A3(\SB1_0_0/i0[6] ), .ZN(
        \SB1_0_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_0/Component_Function_4/N4  ( .A1(\SB1_0_0/i1[9] ), .A2(n380), 
        .A3(\SB1_0_0/i0_4 ), .ZN(\SB1_0_0/Component_Function_4/NAND4_in[3] )
         );
  NAND3_X1 \SB1_0_0/Component_Function_4/N2  ( .A1(\SB1_0_0/i3[0] ), .A2(
        \SB1_0_0/i0_0 ), .A3(\SB1_0_0/i1_7 ), .ZN(
        \SB1_0_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_0/Component_Function_4/N1  ( .A1(\SB1_0_0/i0[9] ), .A2(
        \SB1_0_0/i0_0 ), .A3(\SB1_0_0/i0[8] ), .ZN(
        \SB1_0_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N3  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i0[8] ), .A3(\SB1_0_1/i0[9] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N2  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i0[10] ), .A3(\SB1_0_1/i0[6] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N1  ( .A1(\SB1_0_1/i1_5 ), .A2(
        \SB1_0_1/i0[10] ), .A3(\SB1_0_1/i1[9] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N4  ( .A1(\SB1_0_1/i1_5 ), .A2(
        \SB1_0_1/i0[8] ), .A3(\SB1_0_1/i3[0] ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N3  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i1_7 ), .A3(\SB1_0_1/i0[10] ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N1  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i0_3 ), .A3(\SB1_0_1/i0[6] ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N4  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i1_5 ), .A3(\SB1_0_1/i0_4 ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N2  ( .A1(\SB1_0_1/i3[0] ), .A2(
        \SB1_0_1/i0_0 ), .A3(\SB1_0_1/i1_7 ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N1  ( .A1(\SB1_0_1/i0[9] ), .A2(
        \SB1_0_1/i0_0 ), .A3(\SB1_0_1/i0[8] ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_2/N4  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0_0 ), .A3(\SB1_0_2/i0_4 ), .ZN(
        \SB1_0_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_2/N2  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i0[10] ), .A3(\SB1_0_2/i0[6] ), .ZN(
        \SB1_0_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_2/Component_Function_2/N1  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[10] ), .A3(\SB1_0_2/i1[9] ), .ZN(
        \SB1_0_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_3/N4  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[8] ), .A3(\SB1_0_2/i3[0] ), .ZN(
        \SB1_0_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_3/N3  ( .A1(\SB1_0_2/i1[9] ), .A2(
        \SB1_0_2/i1_7 ), .A3(\SB1_0_2/i0[10] ), .ZN(
        \SB1_0_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_2/Component_Function_3/N1  ( .A1(\SB1_0_2/i1[9] ), .A2(
        \SB1_0_2/i0_3 ), .A3(\SB1_0_2/i0[6] ), .ZN(
        \SB1_0_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_4/N4  ( .A1(\SB1_0_2/i1[9] ), .A2(
        \SB1_0_2/i1_5 ), .A3(\SB1_0_2/i0_4 ), .ZN(
        \SB1_0_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_4/N2  ( .A1(\SB1_0_2/i3[0] ), .A2(
        \SB1_0_2/i0_0 ), .A3(\SB1_0_2/i1_7 ), .ZN(
        \SB1_0_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_2/Component_Function_4/N1  ( .A1(\SB1_0_2/i0[9] ), .A2(
        \SB1_0_2/i0_0 ), .A3(\SB1_0_2/i0[8] ), .ZN(
        \SB1_0_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_2/N4  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0_0 ), .A3(\SB1_0_3/i0_4 ), .ZN(
        \SB1_0_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_2/N2  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i0[10] ), .A3(\SB1_0_3/i0[6] ), .ZN(
        \SB1_0_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_3/Component_Function_2/N1  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[10] ), .A3(\SB1_0_3/i1[9] ), .ZN(
        \SB1_0_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_3/N4  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[8] ), .A3(\SB1_0_3/i3[0] ), .ZN(
        \SB1_0_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_3/N1  ( .A1(\SB1_0_3/i1[9] ), .A2(
        \SB1_0_3/i0_3 ), .A3(\SB1_0_3/i0[6] ), .ZN(
        \SB1_0_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N4  ( .A1(\SB1_0_3/i1[9] ), .A2(
        \SB1_0_3/i1_5 ), .A3(\SB1_0_3/i0_4 ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N2  ( .A1(\SB1_0_3/i3[0] ), .A2(
        \SB1_0_3/i0_0 ), .A3(\SB1_0_3/i1_7 ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N1  ( .A1(\SB1_0_3/i0[9] ), .A2(
        \SB1_0_3/i0_0 ), .A3(\SB1_0_3/i0[8] ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N4  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N3  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i0[8] ), .A3(\SB1_0_4/i0[9] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N2  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i0[10] ), .A3(\SB1_0_4/i0[6] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N1  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0[10] ), .A3(\SB1_0_4/i1[9] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_3/N4  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0[8] ), .A3(\SB1_0_4/i3[0] ), .ZN(
        \SB1_0_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_3/N3  ( .A1(\SB1_0_4/i1[9] ), .A2(
        \SB1_0_4/i1_7 ), .A3(\SB1_0_4/i0[10] ), .ZN(
        \SB1_0_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_3/N1  ( .A1(\SB1_0_4/i1[9] ), .A2(
        \SB1_0_4/i0_3 ), .A3(\SB1_0_4/i0[6] ), .ZN(
        \SB1_0_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N4  ( .A1(\SB1_0_4/i1[9] ), .A2(
        \SB1_0_4/i1_5 ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N2  ( .A1(\SB1_0_4/i3[0] ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i1_7 ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N1  ( .A1(\SB1_0_4/i0[9] ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i0[8] ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_2/N3  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i0[8] ), .A3(\SB1_0_5/i0[9] ), .ZN(
        \SB1_0_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_5/Component_Function_2/N2  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i0[10] ), .A3(\SB1_0_5/i0[6] ), .ZN(
        \SB1_0_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_5/Component_Function_2/N1  ( .A1(\SB1_0_5/i1_5 ), .A2(
        \SB1_0_5/i0[10] ), .A3(\SB1_0_5/i1[9] ), .ZN(
        \SB1_0_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_3/N4  ( .A1(\SB1_0_5/i1_5 ), .A2(
        \SB1_0_5/i0[8] ), .A3(\SB1_0_5/i3[0] ), .ZN(
        \SB1_0_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_5/Component_Function_3/N3  ( .A1(\SB1_0_5/i1[9] ), .A2(
        \SB1_0_5/i1_7 ), .A3(\SB1_0_5/i0[10] ), .ZN(
        \SB1_0_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_5/Component_Function_3/N1  ( .A1(\SB1_0_5/i1[9] ), .A2(
        \SB1_0_5/i0_3 ), .A3(\SB1_0_5/i0[6] ), .ZN(
        \SB1_0_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_4/N2  ( .A1(\SB1_0_5/i3[0] ), .A2(
        \SB1_0_5/i0_0 ), .A3(\SB1_0_5/i1_7 ), .ZN(
        \SB1_0_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_5/Component_Function_4/N1  ( .A1(\SB1_0_5/i0[9] ), .A2(
        \SB1_0_5/i0_0 ), .A3(\SB1_0_5/i0[8] ), .ZN(
        \SB1_0_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_2/N4  ( .A1(\SB1_0_6/i1_5 ), .A2(
        \SB1_0_6/i0_0 ), .A3(\SB1_0_6/i0_4 ), .ZN(
        \SB1_0_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_2/N2  ( .A1(n2136), .A2(
        \SB1_0_6/i0[10] ), .A3(\SB1_0_6/i0[6] ), .ZN(
        \SB1_0_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_6/Component_Function_2/N1  ( .A1(\SB1_0_6/i1_5 ), .A2(
        \SB1_0_6/i0[10] ), .A3(\SB1_0_6/i1[9] ), .ZN(
        \SB1_0_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_3/N4  ( .A1(\SB1_0_6/i1_5 ), .A2(
        \SB1_0_6/i0[8] ), .A3(\SB1_0_6/i3[0] ), .ZN(
        \SB1_0_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_3/N3  ( .A1(\SB1_0_6/i1[9] ), .A2(
        \SB1_0_6/i1_7 ), .A3(\SB1_0_6/i0[10] ), .ZN(
        \SB1_0_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_6/Component_Function_3/N1  ( .A1(\SB1_0_6/i1[9] ), .A2(n2136), .A3(\SB1_0_6/i0[6] ), .ZN(\SB1_0_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_4/N4  ( .A1(\SB1_0_6/i1[9] ), .A2(
        \SB1_0_6/i1_5 ), .A3(\SB1_0_6/i0_4 ), .ZN(
        \SB1_0_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_4/N2  ( .A1(\SB1_0_6/i3[0] ), .A2(
        \SB1_0_6/i0_0 ), .A3(\SB1_0_6/i1_7 ), .ZN(
        \SB1_0_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_6/Component_Function_4/N1  ( .A1(\SB1_0_6/i0[9] ), .A2(
        \SB1_0_6/i0_0 ), .A3(\SB1_0_6/i0[8] ), .ZN(
        \SB1_0_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_2/N4  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0_0 ), .A3(\SB1_0_7/i0_4 ), .ZN(
        \SB1_0_7/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_2/N2  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i0[10] ), .A3(\SB1_0_7/i0[6] ), .ZN(
        \SB1_0_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_7/Component_Function_2/N1  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0[10] ), .A3(\SB1_0_7/i1[9] ), .ZN(
        \SB1_0_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_3/N4  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0[8] ), .A3(\SB1_0_7/i3[0] ), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_3/N3  ( .A1(\SB1_0_7/i1[9] ), .A2(
        \SB1_0_7/i1_7 ), .A3(\SB1_0_7/i0[10] ), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_3/N1  ( .A1(\SB1_0_7/i1[9] ), .A2(
        \SB1_0_7/i0_3 ), .A3(\SB1_0_7/i0[6] ), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_4/N4  ( .A1(\SB1_0_7/i1[9] ), .A2(
        \SB1_0_7/i1_5 ), .A3(\SB1_0_7/i0_4 ), .ZN(
        \SB1_0_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_4/N2  ( .A1(\SB1_0_7/i3[0] ), .A2(
        \SB1_0_7/i0_0 ), .A3(\SB1_0_7/i1_7 ), .ZN(
        \SB1_0_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_7/Component_Function_4/N1  ( .A1(\SB1_0_7/i0[9] ), .A2(
        \SB1_0_7/i0_0 ), .A3(\SB1_0_7/i0[8] ), .ZN(
        \SB1_0_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_2/N2  ( .A1(\SB1_0_8/i0_3 ), .A2(
        \SB1_0_8/i0[10] ), .A3(\SB1_0_8/i0[6] ), .ZN(
        \SB1_0_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_8/Component_Function_2/N1  ( .A1(\SB1_0_8/i1_5 ), .A2(
        \SB1_0_8/i0[10] ), .A3(\SB1_0_8/i1[9] ), .ZN(
        \SB1_0_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_3/N4  ( .A1(\SB1_0_8/i1_5 ), .A2(
        \SB1_0_8/i0[8] ), .A3(\SB1_0_8/i3[0] ), .ZN(
        \SB1_0_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_3/N1  ( .A1(\SB1_0_8/i1[9] ), .A2(
        \SB1_0_8/i0_3 ), .A3(\SB1_0_8/i0[6] ), .ZN(
        \SB1_0_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_4/N4  ( .A1(\SB1_0_8/i1[9] ), .A2(
        \SB1_0_8/i1_5 ), .A3(\SB1_0_8/i0_4 ), .ZN(
        \SB1_0_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_4/N1  ( .A1(\SB1_0_8/i0[9] ), .A2(
        \SB1_0_8/i0_0 ), .A3(\SB1_0_8/i0[8] ), .ZN(
        \SB1_0_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N4  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N2  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i0[10] ), .A3(\SB1_0_9/i0[6] ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N1  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0[10] ), .A3(\SB1_0_9/i1[9] ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_3/N4  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i3[0] ), .ZN(
        \SB1_0_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_3/N1  ( .A1(\SB1_0_9/i1[9] ), .A2(
        \SB1_0_9/i0_3 ), .A3(\SB1_0_9/i0[6] ), .ZN(
        \SB1_0_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N4  ( .A1(\SB1_0_9/i1[9] ), .A2(
        \SB1_0_9/i1_5 ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N2  ( .A1(\SB1_0_9/i3[0] ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i1_7 ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N1  ( .A1(\SB1_0_9/i0[9] ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i0[8] ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_2/N4  ( .A1(\SB1_0_10/i1_5 ), .A2(
        \SB1_0_10/i0_0 ), .A3(\SB1_0_10/i0_4 ), .ZN(
        \SB1_0_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_2/N2  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i0[10] ), .A3(\SB1_0_10/i0[6] ), .ZN(
        \SB1_0_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_10/Component_Function_2/N1  ( .A1(\SB1_0_10/i1_5 ), .A2(
        \SB1_0_10/i0[10] ), .A3(\SB1_0_10/i1[9] ), .ZN(
        \SB1_0_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_3/N4  ( .A1(\SB1_0_10/i1_5 ), .A2(
        \SB1_0_10/i0[8] ), .A3(\SB1_0_10/i3[0] ), .ZN(
        \SB1_0_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_3/N3  ( .A1(\SB1_0_10/i1[9] ), .A2(
        \SB1_0_10/i1_7 ), .A3(\SB1_0_10/i0[10] ), .ZN(
        \SB1_0_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_10/Component_Function_3/N1  ( .A1(\SB1_0_10/i1[9] ), .A2(
        \SB1_0_10/i0_3 ), .A3(\SB1_0_10/i0[6] ), .ZN(
        \SB1_0_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_4/N4  ( .A1(\SB1_0_10/i1[9] ), .A2(
        \SB1_0_10/i1_5 ), .A3(\SB1_0_10/i0_4 ), .ZN(
        \SB1_0_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_4/N2  ( .A1(\SB1_0_10/i3[0] ), .A2(
        \SB1_0_10/i0_0 ), .A3(\SB1_0_10/i1_7 ), .ZN(
        \SB1_0_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_10/Component_Function_4/N1  ( .A1(\SB1_0_10/i0[9] ), .A2(
        \SB1_0_10/i0_0 ), .A3(\SB1_0_10/i0[8] ), .ZN(
        \SB1_0_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_2/N4  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0_0 ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_2/N3  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i0[9] ), .ZN(
        \SB1_0_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_2/N2  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i0[10] ), .A3(\SB1_0_11/i0[6] ), .ZN(
        \SB1_0_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_11/Component_Function_2/N1  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0[10] ), .A3(\SB1_0_11/i1[9] ), .ZN(
        \SB1_0_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_3/N4  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i3[0] ), .ZN(
        \SB1_0_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_3/N3  ( .A1(\SB1_0_11/i1[9] ), .A2(
        \SB1_0_11/i1_7 ), .A3(\SB1_0_11/i0[10] ), .ZN(
        \SB1_0_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_3/N1  ( .A1(\SB1_0_11/i1[9] ), .A2(
        \SB1_0_11/i0_3 ), .A3(\SB1_0_11/i0[6] ), .ZN(
        \SB1_0_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_4/N4  ( .A1(\SB1_0_11/i1[9] ), .A2(
        \SB1_0_11/i1_5 ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_4/N3  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i0[10] ), .A3(\SB1_0_11/i0[9] ), .ZN(
        \SB1_0_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_4/N2  ( .A1(\SB1_0_11/i3[0] ), .A2(
        \SB1_0_11/i0_0 ), .A3(\SB1_0_11/i1_7 ), .ZN(
        \SB1_0_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_11/Component_Function_4/N1  ( .A1(\SB1_0_11/i0[9] ), .A2(
        \SB1_0_11/i0_0 ), .A3(\SB1_0_11/i0[8] ), .ZN(
        \SB1_0_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_2/N2  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i0[10] ), .A3(\SB1_0_12/i0[6] ), .ZN(
        \SB1_0_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_12/Component_Function_3/N4  ( .A1(n381), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i3[0] ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_3/N3  ( .A1(\SB1_0_12/i1[9] ), .A2(
        \SB1_0_12/i1_7 ), .A3(\SB1_0_12/i0[10] ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_12/Component_Function_3/N1  ( .A1(\SB1_0_12/i1[9] ), .A2(
        \SB1_0_12/i0_3 ), .A3(\SB1_0_12/i0[6] ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N4  ( .A1(\SB1_0_12/i1[9] ), .A2(
        n381), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N2  ( .A1(\SB1_0_12/i3[0] ), .A2(
        \SB1_0_12/i0_0 ), .A3(\SB1_0_12/i1_7 ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N1  ( .A1(\SB1_0_12/i0[9] ), .A2(
        \SB1_0_12/i0_0 ), .A3(\SB1_0_12/i0[8] ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_2/N3  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i0[8] ), .A3(\SB1_0_13/i0[9] ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_13/Component_Function_2/N2  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i0[10] ), .A3(\SB1_0_13/i0[6] ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_2/N1  ( .A1(\SB1_0_13/i1_5 ), .A2(
        \SB1_0_13/i0[10] ), .A3(\SB1_0_13/i1[9] ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_3/N4  ( .A1(\SB1_0_13/i1_5 ), .A2(
        \SB1_0_13/i0[8] ), .A3(\SB1_0_13/i3[0] ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_3/N3  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i1_7 ), .A3(\SB1_0_13/i0[10] ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_13/Component_Function_3/N1  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i0_3 ), .A3(\SB1_0_13/i0[6] ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N4  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i1_5 ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N2  ( .A1(\SB1_0_13/i3[0] ), .A2(
        \SB1_0_13/i0_0 ), .A3(\SB1_0_13/i1_7 ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N1  ( .A1(\SB1_0_13/i0[9] ), .A2(
        \SB1_0_13/i0_0 ), .A3(\SB1_0_13/i0[8] ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_2/N4  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0_0 ), .A3(\SB1_0_14/i0_4 ), .ZN(
        \SB1_0_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_2/N2  ( .A1(n862), .A2(
        \SB1_0_14/i0[10] ), .A3(\SB1_0_14/i0[6] ), .ZN(
        \SB1_0_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_2/N1  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[10] ), .A3(\SB1_0_14/i1[9] ), .ZN(
        \SB1_0_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N4  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[8] ), .A3(\SB1_0_14/i3[0] ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N3  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i1_7 ), .A3(\SB1_0_14/i0[10] ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N1  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i0_3 ), .A3(\SB1_0_14/i0[6] ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N4  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i1_5 ), .A3(\SB1_0_14/i0_4 ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N3  ( .A1(\SB1_0_14/i0[9] ), .A2(
        \SB1_0_14/i0[10] ), .A3(\SB1_0_14/i0_3 ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N2  ( .A1(\SB1_0_14/i3[0] ), .A2(
        \SB1_0_14/i0_0 ), .A3(\SB1_0_14/i1_7 ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N1  ( .A1(\SB1_0_14/i0[9] ), .A2(
        \SB1_0_14/i0_0 ), .A3(\SB1_0_14/i0[8] ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_2/N4  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0_0 ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_2/N2  ( .A1(\SB1_0_15/i0_3 ), .A2(
        \SB1_0_15/i0[10] ), .A3(\SB1_0_15/i0[6] ), .ZN(
        \SB1_0_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_15/Component_Function_2/N1  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0[10] ), .A3(\SB1_0_15/i1[9] ), .ZN(
        \SB1_0_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_3/N4  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0[8] ), .A3(\SB1_0_15/i3[0] ), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_3/N1  ( .A1(\SB1_0_15/i1[9] ), .A2(
        \SB1_0_15/i0_3 ), .A3(\SB1_0_15/i0[6] ), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N4  ( .A1(\SB1_0_15/i1[9] ), .A2(
        \SB1_0_15/i1_5 ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N2  ( .A1(\SB1_0_15/i3[0] ), .A2(
        \SB1_0_15/i0_0 ), .A3(\SB1_0_15/i1_7 ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N1  ( .A1(\SB1_0_15/i0[9] ), .A2(
        \SB1_0_15/i0_0 ), .A3(\SB1_0_15/i0[8] ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_2/N2  ( .A1(\SB1_0_16/i0_3 ), .A2(
        \SB1_0_16/i0[10] ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_16/Component_Function_2/N1  ( .A1(\SB1_0_16/i1_5 ), .A2(
        \SB1_0_16/i0[10] ), .A3(\SB1_0_16/i1[9] ), .ZN(
        \SB1_0_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_3/N4  ( .A1(\SB1_0_16/i1_5 ), .A2(
        \SB1_0_16/i0[8] ), .A3(\SB1_0_16/i3[0] ), .ZN(
        \SB1_0_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_3/N1  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i0_3 ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_4/N4  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i1_5 ), .A3(\SB1_0_16/i0_4 ), .ZN(
        \SB1_0_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_4/N2  ( .A1(\SB1_0_16/i3[0] ), .A2(
        \SB1_0_16/i0_0 ), .A3(\SB1_0_16/i1_7 ), .ZN(
        \SB1_0_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_16/Component_Function_4/N1  ( .A1(\SB1_0_16/i0[9] ), .A2(
        \SB1_0_16/i0_0 ), .A3(\SB1_0_16/i0[8] ), .ZN(
        \SB1_0_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_2/N4  ( .A1(\SB1_0_17/i1_5 ), .A2(
        \SB1_0_17/i0_0 ), .A3(\SB1_0_17/i0_4 ), .ZN(
        \SB1_0_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_2/N2  ( .A1(\SB1_0_17/i0_3 ), .A2(
        \SB1_0_17/i0[10] ), .A3(\SB1_0_17/i0[6] ), .ZN(
        \SB1_0_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_17/Component_Function_2/N1  ( .A1(\SB1_0_17/i1_5 ), .A2(
        \SB1_0_17/i0[10] ), .A3(\SB1_0_17/i1[9] ), .ZN(
        \SB1_0_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_3/N4  ( .A1(\SB1_0_17/i1_5 ), .A2(
        \SB1_0_17/i0[8] ), .A3(\SB1_0_17/i3[0] ), .ZN(
        \SB1_0_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_3/N3  ( .A1(\SB1_0_17/i1[9] ), .A2(
        \SB1_0_17/i1_7 ), .A3(\SB1_0_17/i0[10] ), .ZN(
        \SB1_0_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_17/Component_Function_3/N1  ( .A1(\SB1_0_17/i1[9] ), .A2(
        \SB1_0_17/i0_3 ), .A3(\SB1_0_17/i0[6] ), .ZN(
        \SB1_0_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_4/N4  ( .A1(\SB1_0_17/i1[9] ), .A2(
        \SB1_0_17/i1_5 ), .A3(\SB1_0_17/i0_4 ), .ZN(
        \SB1_0_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_4/N2  ( .A1(\SB1_0_17/i3[0] ), .A2(
        \SB1_0_17/i0_0 ), .A3(\SB1_0_17/i1_7 ), .ZN(
        \SB1_0_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_17/Component_Function_4/N1  ( .A1(\SB1_0_17/i0[9] ), .A2(
        \SB1_0_17/i0_0 ), .A3(\SB1_0_17/i0[8] ), .ZN(
        \SB1_0_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N4  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0_0 ), .A3(\SB1_0_18/i0_4 ), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N2  ( .A1(\SB1_0_18/i0_3 ), .A2(
        \SB1_0_18/i0[10] ), .A3(\SB1_0_18/i0[6] ), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N1  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0[10] ), .A3(\SB1_0_18/i1[9] ), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_3/N4  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0[8] ), .A3(\SB1_0_18/i3[0] ), .ZN(
        \SB1_0_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_3/N3  ( .A1(\SB1_0_18/i0[10] ), .A2(
        \SB1_0_18/i1_7 ), .A3(\SB1_0_18/i1[9] ), .ZN(
        \SB1_0_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_18/Component_Function_3/N1  ( .A1(\SB1_0_18/i1[9] ), .A2(
        \SB1_0_18/i0_3 ), .A3(\SB1_0_18/i0[6] ), .ZN(
        \SB1_0_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_4/N2  ( .A1(\SB1_0_18/i3[0] ), .A2(
        \SB1_0_18/i0_0 ), .A3(\SB1_0_18/i1_7 ), .ZN(
        \SB1_0_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_19/Component_Function_2/N4  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0_0 ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_2/N2  ( .A1(\SB1_0_19/i0_3 ), .A2(
        \SB1_0_19/i0[10] ), .A3(\SB1_0_19/i0[6] ), .ZN(
        \SB1_0_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_19/Component_Function_2/N1  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0[10] ), .A3(\SB1_0_19/i1[9] ), .ZN(
        \SB1_0_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_3/N4  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0[8] ), .A3(\SB1_0_19/i3[0] ), .ZN(
        \SB1_0_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_3/N1  ( .A1(\SB1_0_19/i1[9] ), .A2(
        \SB1_0_19/i0_3 ), .A3(\SB1_0_19/i0[6] ), .ZN(
        \SB1_0_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N4  ( .A1(\SB1_0_19/i1[9] ), .A2(
        \SB1_0_19/i1_5 ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N2  ( .A1(\SB1_0_19/i3[0] ), .A2(
        \SB1_0_19/i0_0 ), .A3(\SB1_0_19/i1_7 ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N1  ( .A1(\SB1_0_19/i0[9] ), .A2(
        \SB1_0_19/i0_0 ), .A3(\SB1_0_19/i0[8] ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_2/N4  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i0_4 ), .ZN(
        \SB1_0_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_2/N2  ( .A1(\SB1_0_20/i0_3 ), .A2(
        \SB1_0_20/i0[10] ), .A3(\SB1_0_20/i0[6] ), .ZN(
        \SB1_0_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_20/Component_Function_2/N1  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0[10] ), .A3(\SB1_0_20/i1[9] ), .ZN(
        \SB1_0_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_3/N4  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0[8] ), .A3(\SB1_0_20/i3[0] ), .ZN(
        \SB1_0_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_3/N3  ( .A1(\SB1_0_20/i1[9] ), .A2(
        \SB1_0_20/i1_7 ), .A3(\SB1_0_20/i0[10] ), .ZN(
        \SB1_0_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_20/Component_Function_3/N1  ( .A1(\SB1_0_20/i1[9] ), .A2(
        \SB1_0_20/i0_3 ), .A3(\SB1_0_20/i0[6] ), .ZN(
        \SB1_0_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_4/N4  ( .A1(\SB1_0_20/i1[9] ), .A2(
        \SB1_0_20/i1_5 ), .A3(\SB1_0_20/i0_4 ), .ZN(
        \SB1_0_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_4/N2  ( .A1(\SB1_0_20/i3[0] ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i1_7 ), .ZN(
        \SB1_0_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_20/Component_Function_4/N1  ( .A1(\SB1_0_20/i0[9] ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i0[8] ), .ZN(
        \SB1_0_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_2/N4  ( .A1(\SB1_0_21/i1_5 ), .A2(
        \SB1_0_21/i0_0 ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_21/Component_Function_2/N2  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i0[10] ), .A3(\SB1_0_21/i0[6] ), .ZN(
        \SB1_0_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_21/Component_Function_2/N1  ( .A1(\SB1_0_21/i1_5 ), .A2(
        \SB1_0_21/i0[10] ), .A3(\SB1_0_21/i1[9] ), .ZN(
        \SB1_0_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_3/N4  ( .A1(\SB1_0_21/i1_5 ), .A2(
        \SB1_0_21/i0[8] ), .A3(\SB1_0_21/i3[0] ), .ZN(
        \SB1_0_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_21/Component_Function_3/N3  ( .A1(\SB1_0_21/i1[9] ), .A2(
        \SB1_0_21/i1_7 ), .A3(\SB1_0_21/i0[10] ), .ZN(
        \SB1_0_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_21/Component_Function_3/N1  ( .A1(\SB1_0_21/i1[9] ), .A2(
        \SB1_0_21/i0_3 ), .A3(\SB1_0_21/i0[6] ), .ZN(
        \SB1_0_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_4/N4  ( .A1(\SB1_0_21/i1[9] ), .A2(
        \SB1_0_21/i1_5 ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_21/Component_Function_4/N2  ( .A1(\SB1_0_21/i3[0] ), .A2(
        \SB1_0_21/i0_0 ), .A3(\SB1_0_21/i1_7 ), .ZN(
        \SB1_0_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_21/Component_Function_4/N1  ( .A1(\SB1_0_21/i0[9] ), .A2(
        \SB1_0_21/i0_0 ), .A3(\SB1_0_21/i0[8] ), .ZN(
        \SB1_0_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_2/N4  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i0_4 ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_2/N2  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i0[10] ), .A3(\SB1_0_22/i0[6] ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_22/Component_Function_2/N1  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[10] ), .A3(\SB1_0_22/i1[9] ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_3/N4  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[8] ), .A3(\SB1_0_22/i3[0] ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_3/N3  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i1_7 ), .A3(\SB1_0_22/i0[10] ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_22/Component_Function_3/N1  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i0_3 ), .A3(\SB1_0_22/i0[6] ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N4  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i1_5 ), .A3(\SB1_0_22/i0_4 ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N2  ( .A1(\SB1_0_22/i3[0] ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i1_7 ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N1  ( .A1(\SB1_0_22/i0[9] ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i0[8] ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_2/N2  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i0[10] ), .A3(\SB1_0_23/i0[6] ), .ZN(
        \SB1_0_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_2/N1  ( .A1(\SB1_0_23/i1_5 ), .A2(
        \SB1_0_23/i0[10] ), .A3(\SB1_0_23/i1[9] ), .ZN(
        \SB1_0_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_3/N4  ( .A1(\SB1_0_23/i1_5 ), .A2(
        \SB1_0_23/i0[8] ), .A3(\SB1_0_23/i3[0] ), .ZN(
        \SB1_0_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_3/N3  ( .A1(\SB1_0_23/i1[9] ), .A2(
        \SB1_0_23/i1_7 ), .A3(\SB1_0_23/i0[10] ), .ZN(
        \SB1_0_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_23/Component_Function_3/N1  ( .A1(\SB1_0_23/i1[9] ), .A2(
        \SB1_0_23/i0_3 ), .A3(\SB1_0_23/i0[6] ), .ZN(
        \SB1_0_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N2  ( .A1(\SB1_0_23/i3[0] ), .A2(
        \SB1_0_23/i0_0 ), .A3(\SB1_0_23/i1_7 ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N1  ( .A1(\SB1_0_23/i0[9] ), .A2(
        \SB1_0_23/i0_0 ), .A3(\SB1_0_23/i0[8] ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_2/N4  ( .A1(\SB1_0_24/i1_5 ), .A2(
        \SB1_0_24/i0_0 ), .A3(\SB1_0_24/i0_4 ), .ZN(
        \SB1_0_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_2/N2  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i0[10] ), .A3(\SB1_0_24/i0[6] ), .ZN(
        \SB1_0_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_24/Component_Function_2/N1  ( .A1(\SB1_0_24/i1_5 ), .A2(
        \SB1_0_24/i0[10] ), .A3(\SB1_0_24/i1[9] ), .ZN(
        \SB1_0_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_3/N4  ( .A1(\SB1_0_24/i1_5 ), .A2(
        \SB1_0_24/i0[8] ), .A3(\SB1_0_24/i3[0] ), .ZN(
        \SB1_0_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_3/N3  ( .A1(\SB1_0_24/i1[9] ), .A2(
        \SB1_0_24/i1_7 ), .A3(\SB1_0_24/i0[10] ), .ZN(
        \SB1_0_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_24/Component_Function_3/N1  ( .A1(\SB1_0_24/i1[9] ), .A2(
        \SB1_0_24/i0_3 ), .A3(\SB1_0_24/i0[6] ), .ZN(
        \SB1_0_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N4  ( .A1(\SB1_0_24/i1[9] ), .A2(
        \SB1_0_24/i1_5 ), .A3(\SB1_0_24/i0_4 ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N2  ( .A1(\SB1_0_24/i3[0] ), .A2(
        \SB1_0_24/i0_0 ), .A3(\SB1_0_24/i1_7 ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N1  ( .A1(\SB1_0_24/i0[9] ), .A2(
        \SB1_0_24/i0_0 ), .A3(\SB1_0_24/i0[8] ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_2/N4  ( .A1(\SB1_0_25/i1_5 ), .A2(
        \SB1_0_25/i0_0 ), .A3(\SB1_0_25/i0_4 ), .ZN(
        \SB1_0_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_25/Component_Function_2/N2  ( .A1(\SB1_0_25/i0_3 ), .A2(
        \SB1_0_25/i0[10] ), .A3(\SB1_0_25/i0[6] ), .ZN(
        \SB1_0_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_2/N1  ( .A1(\SB1_0_25/i1_5 ), .A2(
        \SB1_0_25/i0[10] ), .A3(\SB1_0_25/i1[9] ), .ZN(
        \SB1_0_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_3/N4  ( .A1(\SB1_0_25/i1_5 ), .A2(
        \SB1_0_25/i0[8] ), .A3(\SB1_0_25/i3[0] ), .ZN(
        \SB1_0_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_25/Component_Function_3/N3  ( .A1(\SB1_0_25/i1[9] ), .A2(
        \SB1_0_25/i1_7 ), .A3(\SB1_0_25/i0[10] ), .ZN(
        \SB1_0_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_25/Component_Function_3/N1  ( .A1(\SB1_0_25/i1[9] ), .A2(
        \SB1_0_25/i0_3 ), .A3(\SB1_0_25/i0[6] ), .ZN(
        \SB1_0_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_4/N4  ( .A1(\SB1_0_25/i1[9] ), .A2(
        \SB1_0_25/i1_5 ), .A3(\SB1_0_25/i0_4 ), .ZN(
        \SB1_0_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_25/Component_Function_4/N2  ( .A1(\SB1_0_25/i3[0] ), .A2(
        \SB1_0_25/i0_0 ), .A3(\SB1_0_25/i1_7 ), .ZN(
        \SB1_0_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_4/N1  ( .A1(\SB1_0_25/i0[9] ), .A2(
        \SB1_0_25/i0_0 ), .A3(\SB1_0_25/i0[8] ), .ZN(
        \SB1_0_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_2/N4  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0_0 ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_2/N2  ( .A1(\SB1_0_26/i0_3 ), .A2(
        \SB1_0_26/i0[10] ), .A3(\SB1_0_26/i0[6] ), .ZN(
        \SB1_0_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_26/Component_Function_2/N1  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0[10] ), .A3(\SB1_0_26/i1[9] ), .ZN(
        \SB1_0_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_3/N4  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0[8] ), .A3(\SB1_0_26/i3[0] ), .ZN(
        \SB1_0_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_3/N3  ( .A1(\SB1_0_26/i1[9] ), .A2(
        \SB1_0_26/i1_7 ), .A3(\SB1_0_26/i0[10] ), .ZN(
        \SB1_0_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_26/Component_Function_3/N1  ( .A1(\SB1_0_26/i1[9] ), .A2(
        \SB1_0_26/i0_3 ), .A3(\SB1_0_26/i0[6] ), .ZN(
        \SB1_0_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_4/N2  ( .A1(\SB1_0_26/i3[0] ), .A2(
        \SB1_0_26/i0_0 ), .A3(\SB1_0_26/i1_7 ), .ZN(
        \SB1_0_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_26/Component_Function_4/N1  ( .A1(\SB1_0_26/i0[9] ), .A2(
        \SB1_0_26/i0_0 ), .A3(\SB1_0_26/i0[8] ), .ZN(
        \SB1_0_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N4  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0_0 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N1  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i1[9] ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_3/N4  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0[8] ), .A3(\SB1_0_27/i3[0] ), .ZN(
        \SB1_0_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_3/N2  ( .A1(\SB1_0_27/i0_0 ), .A2(
        \SB1_0_27/i0_3 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_3/N1  ( .A1(\SB1_0_27/i1[9] ), .A2(
        \SB1_0_27/i0_3 ), .A3(\SB1_0_27/i0[6] ), .ZN(
        \SB1_0_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N4  ( .A1(\SB1_0_27/i1[9] ), .A2(
        \SB1_0_27/i1_5 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N3  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i0_3 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N2  ( .A1(\SB1_0_27/i3[0] ), .A2(
        \SB1_0_27/i0_0 ), .A3(\SB1_0_27/i1_7 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N1  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0_0 ), .A3(\SB1_0_27/i0[8] ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N4  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0_0 ), .A3(\SB1_0_28/i0_4 ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N2  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i0[10] ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N1  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0[10] ), .A3(\SB1_0_28/i1[9] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_3/N4  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0[8] ), .A3(\SB1_0_28/i3[0] ), .ZN(
        \SB1_0_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_3/N1  ( .A1(\SB1_0_28/i1[9] ), .A2(
        \SB1_0_28/i0_3 ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N4  ( .A1(\SB1_0_28/i1[9] ), .A2(
        \SB1_0_28/i1_5 ), .A3(\SB1_0_28/i0_4 ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N2  ( .A1(\SB1_0_28/i3[0] ), .A2(
        \SB1_0_28/i0_0 ), .A3(\SB1_0_28/i1_7 ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N1  ( .A1(\SB1_0_28/i0[9] ), .A2(
        \SB1_0_28/i0_0 ), .A3(\SB1_0_28/i0[8] ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_2/N4  ( .A1(\SB1_0_29/i1_5 ), .A2(
        \SB1_0_29/i0_0 ), .A3(\SB1_0_29/i0_4 ), .ZN(
        \SB1_0_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_2/N2  ( .A1(\SB1_0_29/i0_3 ), .A2(
        \SB1_0_29/i0[10] ), .A3(\SB1_0_29/i0[6] ), .ZN(
        \SB1_0_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_29/Component_Function_2/N1  ( .A1(\SB1_0_29/i1_5 ), .A2(
        \SB1_0_29/i0[10] ), .A3(\SB1_0_29/i1[9] ), .ZN(
        \SB1_0_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_3/N4  ( .A1(\SB1_0_29/i1_5 ), .A2(
        \SB1_0_29/i0[8] ), .A3(\SB1_0_29/i3[0] ), .ZN(
        \SB1_0_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_3/N3  ( .A1(\SB1_0_29/i1[9] ), .A2(
        \SB1_0_29/i1_7 ), .A3(\SB1_0_29/i0[10] ), .ZN(
        \SB1_0_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_29/Component_Function_3/N1  ( .A1(\SB1_0_29/i1[9] ), .A2(
        \SB1_0_29/i0_3 ), .A3(\SB1_0_29/i0[6] ), .ZN(
        \SB1_0_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_4/N4  ( .A1(\SB1_0_29/i1[9] ), .A2(
        \SB1_0_29/i1_5 ), .A3(\SB1_0_29/i0_4 ), .ZN(
        \SB1_0_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_4/N2  ( .A1(\SB1_0_29/i3[0] ), .A2(
        \SB1_0_29/i0_0 ), .A3(\SB1_0_29/i1_7 ), .ZN(
        \SB1_0_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_29/Component_Function_4/N1  ( .A1(\SB1_0_29/i0[9] ), .A2(
        \SB1_0_29/i0_0 ), .A3(\SB1_0_29/i0[8] ), .ZN(
        \SB1_0_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_2/N2  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i0[10] ), .A3(\SB1_0_30/i0[6] ), .ZN(
        \SB1_0_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_30/Component_Function_2/N1  ( .A1(\SB1_0_30/i1_5 ), .A2(
        \SB1_0_30/i0[10] ), .A3(\SB1_0_30/i1[9] ), .ZN(
        \SB1_0_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_3/N1  ( .A1(\SB1_0_30/i1[9] ), .A2(
        \SB1_0_30/i0_3 ), .A3(\SB1_0_30/i0[6] ), .ZN(
        \SB1_0_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N4  ( .A1(\SB1_0_30/i1[9] ), .A2(
        \SB1_0_30/i1_5 ), .A3(\SB1_0_30/i0_4 ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N2  ( .A1(\SB1_0_30/i3[0] ), .A2(
        \SB1_0_30/i0_0 ), .A3(\SB1_0_30/i1_7 ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N1  ( .A1(\SB1_0_30/i0[9] ), .A2(
        \SB1_0_30/i0_0 ), .A3(\SB1_0_30/i0[8] ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_2/N2  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i0[10] ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_31/Component_Function_2/N1  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[10] ), .A3(\SB1_0_31/i1[9] ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_3/N4  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[8] ), .A3(\SB1_0_31/i3[0] ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_3/N3  ( .A1(\SB1_0_31/i1[9] ), .A2(
        \SB1_0_31/i1_7 ), .A3(\SB1_0_31/i0[10] ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_31/Component_Function_3/N2  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_31/Component_Function_3/N1  ( .A1(\SB1_0_31/i1[9] ), .A2(
        \SB1_0_31/i0_3 ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N4  ( .A1(\SB1_0_31/i1[9] ), .A2(
        \SB1_0_31/i1_5 ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N2  ( .A1(\SB1_0_31/i3[0] ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i1_7 ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N1  ( .A1(\SB1_0_31/i0[9] ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i0[8] ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_2/N2  ( .A1(\SB2_0_0/i0_3 ), .A2(
        \SB2_0_0/i0[10] ), .A3(\SB2_0_0/i0[6] ), .ZN(
        \SB2_0_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_0/Component_Function_3/N3  ( .A1(\SB2_0_0/i1[9] ), .A2(
        \SB2_0_0/i1_7 ), .A3(\SB2_0_0/i0[10] ), .ZN(
        \SB2_0_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_0/Component_Function_3/N1  ( .A1(\SB2_0_0/i1[9] ), .A2(
        \SB2_0_0/i0_3 ), .A3(\SB2_0_0/i0[6] ), .ZN(
        \SB2_0_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N3  ( .A1(\SB2_0_0/i0[9] ), .A2(
        \SB2_0_0/i0[10] ), .A3(\SB2_0_0/i0_3 ), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N2  ( .A1(\SB2_0_0/i3[0] ), .A2(
        \SB2_0_0/i0_0 ), .A3(\SB2_0_0/i1_7 ), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N1  ( .A1(\SB2_0_0/i0[9] ), .A2(
        \SB2_0_0/i0_0 ), .A3(\SB2_0_0/i0[8] ), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_2/N2  ( .A1(\SB2_0_1/i0_3 ), .A2(
        \SB2_0_1/i0[10] ), .A3(\SB2_0_1/i0[6] ), .ZN(
        \SB2_0_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_1/Component_Function_2/N1  ( .A1(\SB2_0_1/i1_5 ), .A2(
        \SB2_0_1/i0[10] ), .A3(\SB2_0_1/i1[9] ), .ZN(
        \SB2_0_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_3/N3  ( .A1(\SB2_0_1/i1[9] ), .A2(
        \SB2_0_1/i1_7 ), .A3(\SB2_0_1/i0[10] ), .ZN(
        \SB2_0_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_1/Component_Function_3/N2  ( .A1(\SB2_0_1/i0_0 ), .A2(
        \SB2_0_1/i0_3 ), .A3(\SB2_0_1/i0_4 ), .ZN(
        \SB2_0_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_1/Component_Function_3/N1  ( .A1(\SB2_0_1/i1[9] ), .A2(
        \SB2_0_1/i0_3 ), .A3(\SB2_0_1/i0[6] ), .ZN(
        \SB2_0_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_4/N3  ( .A1(\SB2_0_1/i0[9] ), .A2(
        \SB2_0_1/i0[10] ), .A3(\SB2_0_1/i0_3 ), .ZN(
        \SB2_0_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_1/Component_Function_4/N2  ( .A1(\SB2_0_1/i3[0] ), .A2(
        \SB2_0_1/i0_0 ), .A3(\SB2_0_1/i1_7 ), .ZN(
        \SB2_0_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_1/Component_Function_4/N1  ( .A1(\SB2_0_1/i0[9] ), .A2(
        \SB2_0_1/i0_0 ), .A3(\SB2_0_1/i0[8] ), .ZN(
        \SB2_0_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_2/N3  ( .A1(\SB2_0_2/i0_3 ), .A2(
        \SB2_0_2/i0[8] ), .A3(\SB2_0_2/i0[9] ), .ZN(
        \SB2_0_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_2/N2  ( .A1(\SB2_0_2/i0_3 ), .A2(
        \SB2_0_2/i0[10] ), .A3(\SB2_0_2/i0[6] ), .ZN(
        \SB2_0_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_2/Component_Function_2/N1  ( .A1(\SB2_0_2/i1_5 ), .A2(
        \SB2_0_2/i0[10] ), .A3(\SB2_0_2/i1[9] ), .ZN(
        \SB2_0_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_3/N4  ( .A1(\SB2_0_2/i1_5 ), .A2(
        \SB2_0_2/i0[8] ), .A3(\SB2_0_2/i3[0] ), .ZN(
        \SB2_0_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_2/Component_Function_3/N3  ( .A1(\SB2_0_2/i1[9] ), .A2(
        \SB2_0_2/i1_7 ), .A3(\SB2_0_2/i0[10] ), .ZN(
        \SB2_0_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_3/N2  ( .A1(\SB2_0_2/i0_0 ), .A2(
        \SB2_0_2/i0_3 ), .A3(\SB2_0_2/i0_4 ), .ZN(
        \SB2_0_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_2/Component_Function_3/N1  ( .A1(\SB2_0_2/i1[9] ), .A2(
        \SB2_0_2/i0_3 ), .A3(\SB2_0_2/i0[6] ), .ZN(
        \SB2_0_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N4  ( .A1(\SB2_0_2/i1[9] ), .A2(
        \SB2_0_2/i1_5 ), .A3(\SB2_0_2/i0_4 ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N2  ( .A1(\SB2_0_2/i3[0] ), .A2(
        \SB2_0_2/i0_0 ), .A3(\SB2_0_2/i1_7 ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N1  ( .A1(\SB2_0_2/i0[9] ), .A2(
        \SB2_0_2/i0_0 ), .A3(\SB2_0_2/i0[8] ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_2/N3  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i0[8] ), .A3(\SB2_0_3/i0[9] ), .ZN(
        \SB2_0_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_3/Component_Function_2/N2  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i0[10] ), .A3(\SB2_0_3/i0[6] ), .ZN(
        \SB2_0_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_3/Component_Function_3/N2  ( .A1(\SB2_0_3/i0_0 ), .A2(
        \SB2_0_3/i0_3 ), .A3(\SB2_0_3/i0_4 ), .ZN(
        \SB2_0_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_3/Component_Function_3/N1  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \SB2_0_3/i0_3 ), .A3(\SB2_0_3/i0[6] ), .ZN(
        \SB2_0_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_4/N3  ( .A1(\SB2_0_3/i0[9] ), .A2(
        \SB2_0_3/i0[10] ), .A3(\SB2_0_3/i0_3 ), .ZN(
        \SB2_0_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_3/Component_Function_4/N1  ( .A1(\SB2_0_3/i0[9] ), .A2(
        \SB2_0_3/i0_0 ), .A3(\SB2_0_3/i0[8] ), .ZN(
        \SB2_0_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_2/N4  ( .A1(\SB2_0_4/i1_5 ), .A2(
        \SB2_0_4/i0_0 ), .A3(\SB2_0_4/i0_4 ), .ZN(
        \SB2_0_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_4/Component_Function_2/N2  ( .A1(\SB2_0_4/i0_3 ), .A2(
        \SB2_0_4/i0[10] ), .A3(\SB2_0_4/i0[6] ), .ZN(
        \SB2_0_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_4/Component_Function_2/N1  ( .A1(\SB2_0_4/i1_5 ), .A2(
        \SB2_0_4/i0[10] ), .A3(\SB2_0_4/i1[9] ), .ZN(
        \SB2_0_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_4/N2  ( .A1(\SB2_0_4/i3[0] ), .A2(
        \SB2_0_4/i0_0 ), .A3(\SB2_0_4/i1_7 ), .ZN(
        \SB2_0_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_4/Component_Function_4/N1  ( .A1(\SB2_0_4/i0[9] ), .A2(
        \SB2_0_4/i0_0 ), .A3(\SB2_0_4/i0[8] ), .ZN(
        \SB2_0_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_2/N4  ( .A1(\SB2_0_5/i1_5 ), .A2(
        \SB2_0_5/i0_0 ), .A3(\SB2_0_5/i0_4 ), .ZN(
        \SB2_0_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_5/Component_Function_2/N2  ( .A1(\SB2_0_5/i0_3 ), .A2(
        \SB2_0_5/i0[10] ), .A3(\SB2_0_5/i0[6] ), .ZN(
        \SB2_0_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_5/Component_Function_2/N1  ( .A1(\SB2_0_5/i1_5 ), .A2(
        \SB2_0_5/i0[10] ), .A3(\SB2_0_5/i1[9] ), .ZN(
        \SB2_0_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_3/N3  ( .A1(\SB2_0_5/i1[9] ), .A2(
        \SB2_0_5/i1_7 ), .A3(\SB2_0_5/i0[10] ), .ZN(
        \SB2_0_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_5/Component_Function_3/N1  ( .A1(\SB2_0_5/i1[9] ), .A2(
        \SB2_0_5/i0_3 ), .A3(\SB2_0_5/i0[6] ), .ZN(
        \SB2_0_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_4/N4  ( .A1(\SB2_0_5/i1[9] ), .A2(
        \SB2_0_5/i1_5 ), .A3(\SB2_0_5/i0_4 ), .ZN(
        \SB2_0_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_5/Component_Function_4/N2  ( .A1(\SB2_0_5/i3[0] ), .A2(
        \SB2_0_5/i0_0 ), .A3(\SB2_0_5/i1_7 ), .ZN(
        \SB2_0_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_5/Component_Function_4/N1  ( .A1(\SB2_0_5/i0[9] ), .A2(
        \SB2_0_5/i0_0 ), .A3(\SB2_0_5/i0[8] ), .ZN(
        \SB2_0_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_2/N3  ( .A1(\SB2_0_6/i0_3 ), .A2(
        \SB2_0_6/i0[8] ), .A3(\SB2_0_6/i0[9] ), .ZN(
        \SB2_0_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_6/Component_Function_2/N2  ( .A1(\SB2_0_6/i0_3 ), .A2(
        \SB2_0_6/i0[10] ), .A3(\SB2_0_6/i0[6] ), .ZN(
        \SB2_0_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_6/Component_Function_2/N1  ( .A1(\SB2_0_6/i1_5 ), .A2(
        \SB2_0_6/i0[10] ), .A3(\SB2_0_6/i1[9] ), .ZN(
        \SB2_0_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_3/N3  ( .A1(\SB2_0_6/i1[9] ), .A2(
        \SB2_0_6/i1_7 ), .A3(\SB2_0_6/i0[10] ), .ZN(
        \SB2_0_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_6/Component_Function_3/N1  ( .A1(\SB2_0_6/i1[9] ), .A2(
        \SB2_0_6/i0_3 ), .A3(\SB2_0_6/i0[6] ), .ZN(
        \SB2_0_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_4/N2  ( .A1(\SB2_0_6/i3[0] ), .A2(
        \SB2_0_6/i0_0 ), .A3(\SB2_0_6/i1_7 ), .ZN(
        \SB2_0_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_6/Component_Function_4/N1  ( .A1(\SB2_0_6/i0[9] ), .A2(
        \SB2_0_6/i0_0 ), .A3(\SB2_0_6/i0[8] ), .ZN(
        \SB2_0_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_2/N3  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i0[8] ), .A3(\SB2_0_7/i0[9] ), .ZN(
        \SB2_0_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_2/N2  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i0[10] ), .A3(\SB2_0_7/i0[6] ), .ZN(
        \SB2_0_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_7/Component_Function_3/N3  ( .A1(\SB2_0_7/i1[9] ), .A2(
        \SB2_0_7/i1_7 ), .A3(\SB2_0_7/i0[10] ), .ZN(
        \SB2_0_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_3/N1  ( .A1(\SB2_0_7/i1[9] ), .A2(
        \SB2_0_7/i0_3 ), .A3(\SB2_0_7/i0[6] ), .ZN(
        \SB2_0_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_4/N2  ( .A1(\SB2_0_7/i3[0] ), .A2(
        \SB2_0_7/i0_0 ), .A3(\SB2_0_7/i1_7 ), .ZN(
        \SB2_0_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_7/Component_Function_4/N1  ( .A1(\SB2_0_7/i0[9] ), .A2(
        \SB2_0_7/i0_0 ), .A3(\SB2_0_7/i0[8] ), .ZN(
        \SB2_0_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_2/N4  ( .A1(\SB2_0_8/i1_5 ), .A2(
        \SB2_0_8/i0_0 ), .A3(\SB2_0_8/i0_4 ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_8/Component_Function_2/N2  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i0[10] ), .A3(\SB2_0_8/i0[6] ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_8/Component_Function_2/N1  ( .A1(\SB2_0_8/i1_5 ), .A2(
        \SB2_0_8/i0[10] ), .A3(\SB2_0_8/i1[9] ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_3/N3  ( .A1(\SB2_0_8/i1[9] ), .A2(
        \SB2_0_8/i1_7 ), .A3(\SB2_0_8/i0[10] ), .ZN(
        \SB2_0_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_8/Component_Function_3/N2  ( .A1(\SB2_0_8/i0_0 ), .A2(
        \SB2_0_8/i0_3 ), .A3(\SB2_0_8/i0_4 ), .ZN(
        \SB2_0_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_8/Component_Function_3/N1  ( .A1(\SB2_0_8/i1[9] ), .A2(
        \SB2_0_8/i0_3 ), .A3(\SB2_0_8/i0[6] ), .ZN(
        \SB2_0_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_4/N4  ( .A1(\SB2_0_8/i1[9] ), .A2(
        \SB2_0_8/i1_5 ), .A3(\SB2_0_8/i0_4 ), .ZN(
        \SB2_0_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_8/Component_Function_4/N2  ( .A1(\SB2_0_8/i3[0] ), .A2(
        \SB2_0_8/i0_0 ), .A3(\SB2_0_8/i1_7 ), .ZN(
        \SB2_0_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_8/Component_Function_4/N1  ( .A1(\SB2_0_8/i0[9] ), .A2(
        \SB2_0_8/i0_0 ), .A3(\SB2_0_8/i0[8] ), .ZN(
        \SB2_0_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_2/N3  ( .A1(\SB2_0_9/i0_3 ), .A2(
        \SB2_0_9/i0[8] ), .A3(\SB2_0_9/i0[9] ), .ZN(
        \SB2_0_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_2/N2  ( .A1(\SB2_0_9/i0_3 ), .A2(
        \SB2_0_9/i0[10] ), .A3(\SB2_0_9/i0[6] ), .ZN(
        \SB2_0_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_9/Component_Function_3/N3  ( .A1(\SB2_0_9/i1[9] ), .A2(
        \SB2_0_9/i1_7 ), .A3(\SB2_0_9/i0[10] ), .ZN(
        \SB2_0_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_3/N2  ( .A1(\SB2_0_9/i0_0 ), .A2(
        \SB2_0_9/i0_3 ), .A3(\SB2_0_9/i0_4 ), .ZN(
        \SB2_0_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_9/Component_Function_3/N1  ( .A1(\SB2_0_9/i1[9] ), .A2(
        \SB2_0_9/i0_3 ), .A3(\SB2_0_9/i0[6] ), .ZN(
        \SB2_0_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_4/N2  ( .A1(\SB2_0_9/i3[0] ), .A2(
        \SB2_0_9/i0_0 ), .A3(\SB2_0_9/i1_7 ), .ZN(
        \SB2_0_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_9/Component_Function_4/N1  ( .A1(\SB2_0_9/i0[9] ), .A2(
        \SB2_0_9/i0_0 ), .A3(\SB2_0_9/i0[8] ), .ZN(
        \SB2_0_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_2/N4  ( .A1(\SB2_0_10/i1_5 ), .A2(
        \SB2_0_10/i0_0 ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_2/N2  ( .A1(\SB2_0_10/i0_3 ), .A2(
        \SB2_0_10/i0[10] ), .A3(\SB2_0_10/i0[6] ), .ZN(
        \SB2_0_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_10/Component_Function_3/N3  ( .A1(\SB2_0_10/i1[9] ), .A2(
        \SB2_0_10/i1_7 ), .A3(\SB2_0_10/i0[10] ), .ZN(
        \SB2_0_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_10/Component_Function_3/N1  ( .A1(\SB2_0_10/i1[9] ), .A2(
        \SB2_0_10/i0_3 ), .A3(\SB2_0_10/i0[6] ), .ZN(
        \SB2_0_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_4/N4  ( .A1(\SB2_0_10/i1[9] ), .A2(
        \SB2_0_10/i1_5 ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_4/N2  ( .A1(\SB2_0_10/i3[0] ), .A2(
        \SB2_0_10/i0_0 ), .A3(\SB2_0_10/i1_7 ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_10/Component_Function_4/N1  ( .A1(\SB2_0_10/i0[9] ), .A2(
        \SB2_0_10/i0_0 ), .A3(\SB2_0_10/i0[8] ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_2/N4  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \SB2_0_11/i0_0 ), .A3(\SB2_0_11/i0_4 ), .ZN(
        \SB2_0_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_2/N3  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i0[8] ), .A3(\SB2_0_11/i0[9] ), .ZN(
        \SB2_0_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_2/N2  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i0[10] ), .A3(\SB2_0_11/i0[6] ), .ZN(
        \SB2_0_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_11/Component_Function_2/N1  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \SB2_0_11/i0[10] ), .A3(\SB2_0_11/i1[9] ), .ZN(
        \SB2_0_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_3/N4  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \SB2_0_11/i0[8] ), .A3(\SB2_0_11/i3[0] ), .ZN(
        \SB2_0_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_3/N3  ( .A1(\SB2_0_11/i1[9] ), .A2(
        \SB2_0_11/i1_7 ), .A3(\SB2_0_11/i0[10] ), .ZN(
        \SB2_0_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_3/N1  ( .A1(\SB2_0_11/i1[9] ), .A2(
        \SB2_0_11/i0_3 ), .A3(\SB2_0_11/i0[6] ), .ZN(
        \SB2_0_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_4/N2  ( .A1(\SB2_0_11/i3[0] ), .A2(
        \SB2_0_11/i0_0 ), .A3(\SB2_0_11/i1_7 ), .ZN(
        \SB2_0_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_12/Component_Function_2/N2  ( .A1(\SB2_0_12/i0_3 ), .A2(
        \SB2_0_12/i0[10] ), .A3(\SB2_0_12/i0[6] ), .ZN(
        \SB2_0_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_12/Component_Function_2/N1  ( .A1(\SB2_0_12/i1_5 ), .A2(
        \SB2_0_12/i0[10] ), .A3(\SB2_0_12/i1[9] ), .ZN(
        \SB2_0_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_3/N3  ( .A1(\SB2_0_12/i1[9] ), .A2(
        \SB2_0_12/i1_7 ), .A3(\SB2_0_12/i0[10] ), .ZN(
        \SB2_0_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_3/N2  ( .A1(\SB2_0_12/i0_0 ), .A2(
        \SB2_0_12/i0_3 ), .A3(\SB2_0_12/i0_4 ), .ZN(
        \SB2_0_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N4  ( .A1(\SB2_0_12/i1[9] ), .A2(
        \SB2_0_12/i1_5 ), .A3(\SB2_0_12/i0_4 ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N3  ( .A1(\SB2_0_12/i0[9] ), .A2(
        \SB2_0_12/i0[10] ), .A3(\SB2_0_12/i0_3 ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N2  ( .A1(\SB2_0_12/i3[0] ), .A2(
        \SB2_0_12/i0_0 ), .A3(\SB2_0_12/i1_7 ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N1  ( .A1(\SB2_0_12/i0[9] ), .A2(
        \SB2_0_12/i0_0 ), .A3(\SB2_0_12/i0[8] ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_2/N2  ( .A1(\SB2_0_13/i0_3 ), .A2(
        \SB2_0_13/i0[10] ), .A3(\SB2_0_13/i0[6] ), .ZN(
        \SB2_0_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_13/Component_Function_2/N1  ( .A1(\SB2_0_13/i1_5 ), .A2(
        \SB2_0_13/i0[10] ), .A3(\SB2_0_13/i1[9] ), .ZN(
        \SB2_0_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_3/N4  ( .A1(\SB2_0_13/i1_5 ), .A2(
        \SB2_0_13/i0[8] ), .A3(\SB2_0_13/i3[0] ), .ZN(
        \SB2_0_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_13/Component_Function_3/N3  ( .A1(\SB2_0_13/i1[9] ), .A2(
        \SB2_0_13/i1_7 ), .A3(\SB2_0_13/i0[10] ), .ZN(
        \SB2_0_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_13/Component_Function_3/N1  ( .A1(\SB2_0_13/i1[9] ), .A2(
        \SB2_0_13/i0_3 ), .A3(\SB2_0_13/i0[6] ), .ZN(
        \SB2_0_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N4  ( .A1(\SB2_0_13/i1[9] ), .A2(
        \SB2_0_13/i1_5 ), .A3(\SB2_0_13/i0_4 ), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N2  ( .A1(\SB2_0_13/i3[0] ), .A2(
        \SB2_0_13/i0_0 ), .A3(\SB2_0_13/i1_7 ), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N1  ( .A1(\SB2_0_13/i0[9] ), .A2(
        \SB2_0_13/i0_0 ), .A3(\SB2_0_13/i0[8] ), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_3/N4  ( .A1(\SB2_0_14/i1_5 ), .A2(
        \SB2_0_14/i0[8] ), .A3(\SB2_0_14/i3[0] ), .ZN(
        \SB2_0_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_3/N3  ( .A1(\SB2_0_14/i1[9] ), .A2(
        \SB2_0_14/i1_7 ), .A3(\SB2_0_14/i0[10] ), .ZN(
        \SB2_0_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_14/Component_Function_4/N4  ( .A1(\SB2_0_14/i1[9] ), .A2(
        \SB2_0_14/i1_5 ), .A3(\SB2_0_14/i0_4 ), .ZN(
        \SB2_0_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_4/N2  ( .A1(\SB2_0_14/i3[0] ), .A2(
        \SB2_0_14/i0_0 ), .A3(\SB2_0_14/i1_7 ), .ZN(
        \SB2_0_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_14/Component_Function_4/N1  ( .A1(\SB2_0_14/i0[9] ), .A2(
        \SB2_0_14/i0_0 ), .A3(\SB2_0_14/i0[8] ), .ZN(
        \SB2_0_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_2/N4  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB2_0_15/i0_0 ), .A3(\SB2_0_15/i0_4 ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_15/Component_Function_2/N3  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i0[8] ), .A3(\SB2_0_15/i0[9] ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_15/Component_Function_2/N2  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i0[10] ), .A3(\SB2_0_15/i0[6] ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_15/Component_Function_2/N1  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB2_0_15/i0[10] ), .A3(\SB2_0_15/i1[9] ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_3/N4  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB2_0_15/i0[8] ), .A3(\SB2_0_15/i3[0] ), .ZN(
        \SB2_0_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_15/Component_Function_3/N3  ( .A1(\SB2_0_15/i1[9] ), .A2(
        \SB2_0_15/i1_7 ), .A3(\SB2_0_15/i0[10] ), .ZN(
        \SB2_0_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N4  ( .A1(\SB2_0_15/i1[9] ), .A2(
        \SB2_0_15/i1_5 ), .A3(\SB2_0_15/i0_4 ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N2  ( .A1(\SB2_0_15/i3[0] ), .A2(
        \SB2_0_15/i0_0 ), .A3(\SB2_0_15/i1_7 ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N1  ( .A1(\SB2_0_15/i0[9] ), .A2(
        \SB2_0_15/i0_0 ), .A3(\SB2_0_15/i0[8] ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_2/N1  ( .A1(\SB2_0_16/i1_5 ), .A2(
        \SB2_0_16/i0[10] ), .A3(\SB2_0_16/i1[9] ), .ZN(
        \SB2_0_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_3/N2  ( .A1(\SB2_0_16/i0_0 ), .A2(
        \SB2_0_16/i0_3 ), .A3(\SB2_0_16/i0_4 ), .ZN(
        \SB2_0_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_16/Component_Function_4/N4  ( .A1(\SB2_0_16/i1[9] ), .A2(
        \SB2_0_16/i1_5 ), .A3(\RI3[0][94] ), .ZN(
        \SB2_0_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_4/N1  ( .A1(\SB2_0_16/i0[9] ), .A2(
        \SB2_0_16/i0_0 ), .A3(\SB2_0_16/i0[8] ), .ZN(
        \SB2_0_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_2/N4  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0_0 ), .A3(\SB2_0_17/i0_4 ), .ZN(
        \SB2_0_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_2/N2  ( .A1(\SB2_0_17/i0_3 ), .A2(
        \SB2_0_17/i0[10] ), .A3(\SB2_0_17/i0[6] ), .ZN(
        \SB2_0_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_17/Component_Function_2/N1  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0[10] ), .A3(\SB2_0_17/i1[9] ), .ZN(
        \SB2_0_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_3/N3  ( .A1(\SB2_0_17/i1[9] ), .A2(
        \SB2_0_17/i1_7 ), .A3(\SB2_0_17/i0[10] ), .ZN(
        \SB2_0_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_17/Component_Function_3/N2  ( .A1(\SB2_0_17/i0_0 ), .A2(
        \SB2_0_17/i0_3 ), .A3(\SB2_0_17/i0_4 ), .ZN(
        \SB2_0_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_17/Component_Function_3/N1  ( .A1(\SB2_0_17/i1[9] ), .A2(
        \SB2_0_17/i0_3 ), .A3(\SB2_0_17/i0[6] ), .ZN(
        \SB2_0_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N4  ( .A1(\SB2_0_17/i1[9] ), .A2(
        \SB2_0_17/i1_5 ), .A3(\SB2_0_17/i0_4 ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N3  ( .A1(\SB2_0_17/i0[9] ), .A2(
        \SB2_0_17/i0[10] ), .A3(\SB2_0_17/i0_3 ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N2  ( .A1(\SB2_0_17/i3[0] ), .A2(
        \SB2_0_17/i0_0 ), .A3(\SB2_0_17/i1_7 ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N1  ( .A1(\SB2_0_17/i0[9] ), .A2(
        \SB2_0_17/i0_0 ), .A3(\SB2_0_17/i0[8] ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_18/Component_Function_2/N3  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i0[8] ), .A3(\SB2_0_18/i0[9] ), .ZN(
        \SB2_0_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_18/Component_Function_2/N2  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i0[10] ), .A3(\SB2_0_18/i0[6] ), .ZN(
        \SB2_0_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_18/Component_Function_2/N1  ( .A1(\SB2_0_18/i1_5 ), .A2(
        \SB2_0_18/i0[10] ), .A3(\SB2_0_18/i1[9] ), .ZN(
        \SB2_0_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_18/Component_Function_3/N3  ( .A1(\SB2_0_18/i1[9] ), .A2(
        \SB2_0_18/i1_7 ), .A3(\SB2_0_18/i0[10] ), .ZN(
        \SB2_0_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_18/Component_Function_3/N2  ( .A1(\SB2_0_18/i0_0 ), .A2(
        \SB2_0_18/i0_3 ), .A3(\SB2_0_18/i0_4 ), .ZN(
        \SB2_0_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_18/Component_Function_3/N1  ( .A1(\SB2_0_18/i1[9] ), .A2(
        \SB2_0_18/i0_3 ), .A3(\SB2_0_18/i0[6] ), .ZN(
        \SB2_0_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_18/Component_Function_4/N4  ( .A1(\SB2_0_18/i1[9] ), .A2(
        \SB2_0_18/i1_5 ), .A3(\SB2_0_18/i0_4 ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_18/Component_Function_4/N1  ( .A1(\SB2_0_18/i0[9] ), .A2(
        \SB2_0_18/i0_0 ), .A3(\SB2_0_18/i0[8] ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_2/N3  ( .A1(\SB2_0_19/i0_3 ), .A2(
        \SB2_0_19/i0[8] ), .A3(\SB2_0_19/i0[9] ), .ZN(
        \SB2_0_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_19/Component_Function_2/N2  ( .A1(\SB2_0_19/i0_3 ), .A2(
        \SB2_0_19/i0[10] ), .A3(\SB2_0_19/i0[6] ), .ZN(
        \SB2_0_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_19/Component_Function_2/N1  ( .A1(\SB2_0_19/i1_5 ), .A2(
        \SB2_0_19/i0[10] ), .A3(\SB2_0_19/i1[9] ), .ZN(
        \SB2_0_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_3/N4  ( .A1(\SB2_0_19/i1_5 ), .A2(
        \SB2_0_19/i0[8] ), .A3(\SB2_0_19/i3[0] ), .ZN(
        \SB2_0_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_19/Component_Function_3/N3  ( .A1(\SB2_0_19/i1[9] ), .A2(
        \SB2_0_19/i1_7 ), .A3(\SB2_0_19/i0[10] ), .ZN(
        \SB2_0_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_19/Component_Function_3/N2  ( .A1(\SB2_0_19/i0_0 ), .A2(
        \SB2_0_19/i0_3 ), .A3(\SB2_0_19/i0_4 ), .ZN(
        \SB2_0_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_19/Component_Function_3/N1  ( .A1(\SB2_0_19/i1[9] ), .A2(
        \SB2_0_19/i0_3 ), .A3(\SB2_0_19/i0[6] ), .ZN(
        \SB2_0_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_4/N4  ( .A1(\SB2_0_19/i1[9] ), .A2(
        \SB2_0_19/i1_5 ), .A3(\SB2_0_19/i0_4 ), .ZN(
        \SB2_0_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_19/Component_Function_4/N3  ( .A1(\SB2_0_19/i0[9] ), .A2(
        \SB2_0_19/i0[10] ), .A3(\SB2_0_19/i0_3 ), .ZN(
        \SB2_0_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_19/Component_Function_4/N2  ( .A1(\SB2_0_19/i3[0] ), .A2(
        \SB2_0_19/i0_0 ), .A3(\SB2_0_19/i1_7 ), .ZN(
        \SB2_0_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_19/Component_Function_4/N1  ( .A1(\SB2_0_19/i0[9] ), .A2(
        \SB2_0_19/i0_0 ), .A3(\SB2_0_19/i0[8] ), .ZN(
        \SB2_0_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_20/Component_Function_2/N3  ( .A1(\SB2_0_20/i0_3 ), .A2(
        \SB2_0_20/i0[8] ), .A3(\SB2_0_20/i0[9] ), .ZN(
        \SB2_0_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_20/Component_Function_2/N2  ( .A1(\SB2_0_20/i0_3 ), .A2(
        \SB2_0_20/i0[10] ), .A3(\SB2_0_20/i0[6] ), .ZN(
        \SB2_0_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_20/Component_Function_3/N4  ( .A1(\SB2_0_20/i1_5 ), .A2(
        \SB2_0_20/i0[8] ), .A3(\SB2_0_20/i3[0] ), .ZN(
        \SB2_0_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_20/Component_Function_3/N3  ( .A1(\SB2_0_20/i1[9] ), .A2(
        \SB2_0_20/i1_7 ), .A3(\SB2_0_20/i0[10] ), .ZN(
        \SB2_0_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_20/Component_Function_4/N4  ( .A1(\SB2_0_20/i1[9] ), .A2(
        \SB2_0_20/i1_5 ), .A3(\SB2_0_20/i0_4 ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_20/Component_Function_4/N2  ( .A1(\SB2_0_20/i3[0] ), .A2(
        \SB2_0_20/i0_0 ), .A3(\SB2_0_20/i1_7 ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_20/Component_Function_4/N1  ( .A1(\SB2_0_20/i0[9] ), .A2(
        \SB2_0_20/i0_0 ), .A3(\SB2_0_20/i0[8] ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_21/Component_Function_2/N3  ( .A1(\SB2_0_21/i0_3 ), .A2(
        \SB2_0_21/i0[8] ), .A3(\SB2_0_21/i0[9] ), .ZN(
        \SB2_0_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_21/Component_Function_2/N2  ( .A1(\SB2_0_21/i0_3 ), .A2(
        \SB2_0_21/i0[10] ), .A3(\SB2_0_21/i0[6] ), .ZN(
        \SB2_0_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_21/Component_Function_2/N1  ( .A1(\SB2_0_21/i1_5 ), .A2(
        \SB2_0_21/i0[10] ), .A3(\SB2_0_21/i1[9] ), .ZN(
        \SB2_0_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_21/Component_Function_4/N2  ( .A1(\SB2_0_21/i3[0] ), .A2(
        \SB2_0_21/i0_0 ), .A3(\SB2_0_21/i1_7 ), .ZN(
        \SB2_0_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_21/Component_Function_4/N1  ( .A1(\SB2_0_21/i0[9] ), .A2(
        \SB2_0_21/i0_0 ), .A3(\SB2_0_21/i0[8] ), .ZN(
        \SB2_0_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_22/Component_Function_2/N3  ( .A1(\SB2_0_22/i0_3 ), .A2(
        \SB2_0_22/i0[8] ), .A3(\SB2_0_22/i0[9] ), .ZN(
        \SB2_0_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_22/Component_Function_2/N2  ( .A1(\SB2_0_22/i0_3 ), .A2(
        \SB2_0_22/i0[10] ), .A3(\SB2_0_22/i0[6] ), .ZN(
        \SB2_0_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_22/Component_Function_2/N1  ( .A1(\SB2_0_22/i1_5 ), .A2(
        \SB2_0_22/i0[10] ), .A3(\SB2_0_22/i1[9] ), .ZN(
        \SB2_0_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_22/Component_Function_3/N2  ( .A1(\SB2_0_22/i0_0 ), .A2(
        \SB2_0_22/i0_3 ), .A3(\SB2_0_22/i0_4 ), .ZN(
        \SB2_0_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_22/Component_Function_4/N2  ( .A1(\SB2_0_22/i3[0] ), .A2(
        \SB2_0_22/i0_0 ), .A3(\SB2_0_22/i1_7 ), .ZN(
        \SB2_0_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_22/Component_Function_4/N1  ( .A1(\SB2_0_22/i0[9] ), .A2(
        \SB2_0_22/i0_0 ), .A3(\SB2_0_22/i0[8] ), .ZN(
        \SB2_0_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_2/N2  ( .A1(\SB2_0_23/i0_3 ), .A2(
        \SB2_0_23/i0[10] ), .A3(\SB2_0_23/i0[6] ), .ZN(
        \SB2_0_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_23/Component_Function_2/N1  ( .A1(\SB2_0_23/i1_5 ), .A2(
        \SB2_0_23/i0[10] ), .A3(\SB2_0_23/i1[9] ), .ZN(
        \SB2_0_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_3/N3  ( .A1(\SB2_0_23/i1[9] ), .A2(
        \SB2_0_23/i1_7 ), .A3(\SB2_0_23/i0[10] ), .ZN(
        \SB2_0_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_23/Component_Function_4/N4  ( .A1(\SB2_0_23/i1[9] ), .A2(
        \SB2_0_23/i1_5 ), .A3(\SB2_0_23/i0_4 ), .ZN(
        \SB2_0_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_23/Component_Function_4/N2  ( .A1(\SB2_0_23/i3[0] ), .A2(
        \SB2_0_23/i0_0 ), .A3(\SB2_0_23/i1_7 ), .ZN(
        \SB2_0_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_23/Component_Function_4/N1  ( .A1(\SB2_0_23/i0[9] ), .A2(
        \SB2_0_23/i0_0 ), .A3(\SB2_0_23/i0[8] ), .ZN(
        \SB2_0_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_2/N3  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i0[8] ), .A3(\SB2_0_24/i0[9] ), .ZN(
        \SB2_0_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_2/N2  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i0[10] ), .A3(\SB2_0_24/i0[6] ), .ZN(
        \SB2_0_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_24/Component_Function_3/N3  ( .A1(\SB2_0_24/i1[9] ), .A2(
        \SB2_0_24/i1_7 ), .A3(\SB2_0_24/i0[10] ), .ZN(
        \SB2_0_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_3/N2  ( .A1(\SB2_0_24/i0_0 ), .A2(
        \SB2_0_24/i0_3 ), .A3(\SB2_0_24/i0_4 ), .ZN(
        \SB2_0_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_24/Component_Function_3/N1  ( .A1(\SB2_0_24/i1[9] ), .A2(
        \SB2_0_24/i0_3 ), .A3(\SB2_0_24/i0[6] ), .ZN(
        \SB2_0_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N3  ( .A1(\SB2_0_24/i0[9] ), .A2(
        \SB2_0_24/i0[10] ), .A3(\SB2_0_24/i0_3 ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N2  ( .A1(\SB2_0_24/i3[0] ), .A2(
        \SB2_0_24/i0_0 ), .A3(\SB2_0_24/i1_7 ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N1  ( .A1(\SB2_0_24/i0[9] ), .A2(
        \SB2_0_24/i0_0 ), .A3(\SB2_0_24/i0[8] ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_2/N4  ( .A1(\SB2_0_25/i1_5 ), .A2(
        \SB2_0_25/i0_0 ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_25/Component_Function_2/N3  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i0[8] ), .A3(\SB2_0_25/i0[9] ), .ZN(
        \SB2_0_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_25/Component_Function_2/N2  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i0[10] ), .A3(\SB2_0_25/i0[6] ), .ZN(
        \SB2_0_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_25/Component_Function_2/N1  ( .A1(\SB2_0_25/i1_5 ), .A2(
        \SB2_0_25/i0[10] ), .A3(\SB2_0_25/i1[9] ), .ZN(
        \SB2_0_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_3/N3  ( .A1(\SB2_0_25/i1[9] ), .A2(
        \SB2_0_25/i1_7 ), .A3(\SB2_0_25/i0[10] ), .ZN(
        \SB2_0_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_25/Component_Function_3/N2  ( .A1(\SB2_0_25/i0_0 ), .A2(
        \SB2_0_25/i0_3 ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_25/Component_Function_4/N4  ( .A1(\SB2_0_25/i1[9] ), .A2(
        \SB2_0_25/i1_5 ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_25/Component_Function_4/N2  ( .A1(\SB2_0_25/i3[0] ), .A2(
        \SB2_0_25/i0_0 ), .A3(\SB2_0_25/i1_7 ), .ZN(
        \SB2_0_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_25/Component_Function_4/N1  ( .A1(\SB2_0_25/i0[9] ), .A2(
        \SB2_0_25/i0_0 ), .A3(\SB2_0_25/i0[8] ), .ZN(
        \SB2_0_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_2/N4  ( .A1(\SB2_0_26/i1_5 ), .A2(
        \SB2_0_26/i0_0 ), .A3(\SB2_0_26/i0_4 ), .ZN(
        \SB2_0_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_26/Component_Function_2/N2  ( .A1(\SB2_0_26/i0_3 ), .A2(
        \SB2_0_26/i0[10] ), .A3(\SB2_0_26/i0[6] ), .ZN(
        \SB2_0_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_26/Component_Function_3/N2  ( .A1(\SB2_0_26/i0_0 ), .A2(
        \SB2_0_26/i0_3 ), .A3(\SB2_0_26/i0_4 ), .ZN(
        \SB2_0_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_26/Component_Function_3/N1  ( .A1(\SB2_0_26/i1[9] ), .A2(
        \SB2_0_26/i0_3 ), .A3(\SB2_0_26/i0[6] ), .ZN(
        \SB2_0_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_4/N4  ( .A1(\SB2_0_26/i1[9] ), .A2(
        \SB2_0_26/i1_5 ), .A3(\SB2_0_26/i0_4 ), .ZN(
        \SB2_0_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_26/Component_Function_4/N2  ( .A1(\SB2_0_26/i3[0] ), .A2(
        \SB2_0_26/i0_0 ), .A3(\SB2_0_26/i1_7 ), .ZN(
        \SB2_0_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_26/Component_Function_4/N1  ( .A1(n2132), .A2(
        \SB2_0_26/i0_0 ), .A3(\SB2_0_26/i0[8] ), .ZN(
        \SB2_0_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_2/N4  ( .A1(\SB2_0_27/i1_5 ), .A2(
        \SB2_0_27/i0_0 ), .A3(\SB2_0_27/i0_4 ), .ZN(
        \SB2_0_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_27/Component_Function_2/N2  ( .A1(\SB2_0_27/i0_3 ), .A2(
        \SB2_0_27/i0[10] ), .A3(\SB2_0_27/i0[6] ), .ZN(
        \SB2_0_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_27/Component_Function_4/N4  ( .A1(\SB2_0_27/i1[9] ), .A2(
        \SB2_0_27/i1_5 ), .A3(\SB2_0_27/i0_4 ), .ZN(
        \SB2_0_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_27/Component_Function_4/N1  ( .A1(\SB2_0_27/i0[9] ), .A2(
        \SB2_0_27/i0_0 ), .A3(\SB2_0_27/i0[8] ), .ZN(
        \SB2_0_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_2/N2  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i0[10] ), .A3(\SB2_0_28/i0[6] ), .ZN(
        \SB2_0_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_28/Component_Function_2/N1  ( .A1(\SB2_0_28/i1_5 ), .A2(
        \SB2_0_28/i0[10] ), .A3(\SB2_0_28/i1[9] ), .ZN(
        \SB2_0_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_3/N3  ( .A1(\SB2_0_28/i1[9] ), .A2(
        \SB2_0_28/i1_7 ), .A3(\SB2_0_28/i0[10] ), .ZN(
        \SB2_0_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_28/Component_Function_3/N2  ( .A1(\SB2_0_28/i0_0 ), .A2(
        \SB2_0_28/i0_3 ), .A3(\SB2_0_28/i0_4 ), .ZN(
        \SB2_0_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_28/Component_Function_3/N1  ( .A1(\SB2_0_28/i1[9] ), .A2(
        \SB2_0_28/i0_3 ), .A3(\SB2_0_28/i0[6] ), .ZN(
        \SB2_0_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_4/N4  ( .A1(\SB2_0_28/i1[9] ), .A2(
        \SB2_0_28/i1_5 ), .A3(\SB2_0_28/i0_4 ), .ZN(
        \SB2_0_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_28/Component_Function_4/N2  ( .A1(\SB2_0_28/i3[0] ), .A2(
        \SB2_0_28/i0_0 ), .A3(\SB2_0_28/i1_7 ), .ZN(
        \SB2_0_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_28/Component_Function_4/N1  ( .A1(\SB2_0_28/i0[9] ), .A2(
        \SB2_0_28/i0_0 ), .A3(\SB2_0_28/i0[8] ), .ZN(
        \SB2_0_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_2/N3  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i0[8] ), .A3(\SB2_0_29/i0[9] ), .ZN(
        \SB2_0_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_2/N2  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i0[10] ), .A3(\SB2_0_29/i0[6] ), .ZN(
        \SB2_0_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_29/Component_Function_3/N4  ( .A1(\SB2_0_29/i1_5 ), .A2(
        \SB2_0_29/i0[8] ), .A3(\SB2_0_29/i3[0] ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_3/N3  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i1_7 ), .A3(\SB2_0_29/i0[10] ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_3/N2  ( .A1(\SB2_0_29/i0_0 ), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_29/Component_Function_3/N1  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0[6] ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N4  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i1_5 ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N3  ( .A1(\SB2_0_29/i0[9] ), .A2(
        \SB2_0_29/i0[10] ), .A3(\SB2_0_29/i0_3 ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N2  ( .A1(\SB2_0_29/i3[0] ), .A2(
        \SB2_0_29/i0_0 ), .A3(\SB2_0_29/i1_7 ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N1  ( .A1(\SB2_0_29/i0[9] ), .A2(
        \SB2_0_29/i0_0 ), .A3(\SB2_0_29/i0[8] ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_2/N2  ( .A1(\SB2_0_30/i0_3 ), .A2(
        \SB2_0_30/i0[10] ), .A3(\SB2_0_30/i0[6] ), .ZN(
        \SB2_0_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_30/Component_Function_3/N2  ( .A1(\SB2_0_30/i0_0 ), .A2(
        \SB2_0_30/i0_3 ), .A3(\SB2_0_30/i0_4 ), .ZN(
        \SB2_0_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_30/Component_Function_3/N1  ( .A1(\SB2_0_30/i1[9] ), .A2(
        \SB2_0_30/i0_3 ), .A3(\RI3[0][7] ), .ZN(
        \SB2_0_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N3  ( .A1(\SB2_0_30/i0[9] ), .A2(
        \SB2_0_30/i0[10] ), .A3(\SB2_0_30/i0_3 ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N2  ( .A1(\SB2_0_30/i3[0] ), .A2(
        \SB2_0_30/i0_0 ), .A3(\SB2_0_30/i1_7 ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N1  ( .A1(\SB2_0_30/i0[9] ), .A2(
        \SB2_0_30/i0_0 ), .A3(\SB2_0_30/i0[8] ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_2/N4  ( .A1(\SB2_0_31/i1_5 ), .A2(
        \SB2_0_31/i0_0 ), .A3(\SB2_0_31/i0_4 ), .ZN(
        \SB2_0_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_2/N2  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i0[10] ), .A3(\SB2_0_31/i0[6] ), .ZN(
        \SB2_0_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_31/Component_Function_3/N3  ( .A1(\SB2_0_31/i1[9] ), .A2(
        \SB2_0_31/i1_7 ), .A3(\SB2_0_31/i0[10] ), .ZN(
        \SB2_0_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_3/N1  ( .A1(\SB2_0_31/i1[9] ), .A2(
        \SB2_0_31/i0_3 ), .A3(\SB2_0_31/i0[6] ), .ZN(
        \SB2_0_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_4/N4  ( .A1(\SB2_0_31/i1[9] ), .A2(
        \SB2_0_31/i1_5 ), .A3(\SB2_0_31/i0_4 ), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_4/N2  ( .A1(\SB2_0_31/i3[0] ), .A2(
        \SB2_0_31/i0_0 ), .A3(\SB2_0_31/i1_7 ), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_31/Component_Function_4/N1  ( .A1(\SB2_0_31/i0[9] ), .A2(
        \SB2_0_31/i0_0 ), .A3(\SB2_0_31/i0[8] ), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_2/N2  ( .A1(\SB1_1_0/i0_3 ), .A2(
        \SB1_1_0/i0[10] ), .A3(\SB1_1_0/i0[6] ), .ZN(
        \SB1_1_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_0/Component_Function_2/N1  ( .A1(\SB1_1_0/i1_5 ), .A2(
        \SB1_1_0/i0[10] ), .A3(\SB1_1_0/i1[9] ), .ZN(
        \SB1_1_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_3/N1  ( .A1(\SB1_1_0/i1[9] ), .A2(
        \SB1_1_0/i0_3 ), .A3(\SB1_1_0/i0[6] ), .ZN(
        \SB1_1_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_4/N4  ( .A1(\SB1_1_0/i1[9] ), .A2(
        \SB1_1_0/i1_5 ), .A3(\SB1_1_0/i0_4 ), .ZN(
        \SB1_1_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_0/Component_Function_4/N2  ( .A1(\SB1_1_0/i3[0] ), .A2(
        \SB1_1_0/i0_0 ), .A3(\SB1_1_0/i1_7 ), .ZN(
        \SB1_1_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_0/Component_Function_4/N1  ( .A1(\SB1_1_0/i0[9] ), .A2(
        \SB1_1_0/i0_0 ), .A3(\SB1_1_0/i0[8] ), .ZN(
        \SB1_1_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_2/N2  ( .A1(\SB1_1_1/i0_3 ), .A2(
        \SB1_1_1/i0[10] ), .A3(\SB1_1_1/i0[6] ), .ZN(
        \SB1_1_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_1/Component_Function_2/N1  ( .A1(\SB1_1_1/i1_5 ), .A2(
        \SB1_1_1/i0[10] ), .A3(\SB1_1_1/i1[9] ), .ZN(
        \SB1_1_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_3/N4  ( .A1(\SB1_1_1/i1_5 ), .A2(
        \SB1_1_1/i0[8] ), .A3(\SB1_1_1/i3[0] ), .ZN(
        \SB1_1_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_1/Component_Function_3/N3  ( .A1(\SB1_1_1/i1[9] ), .A2(
        \SB1_1_1/i1_7 ), .A3(\SB1_1_1/i0[10] ), .ZN(
        \SB1_1_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_1/Component_Function_3/N1  ( .A1(\SB1_1_1/i1[9] ), .A2(
        \SB1_1_1/i0_3 ), .A3(\SB1_1_1/i0[6] ), .ZN(
        \SB1_1_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_4/N4  ( .A1(\SB1_1_1/i1[9] ), .A2(
        \SB1_1_1/i1_5 ), .A3(\SB1_1_1/i0_4 ), .ZN(
        \SB1_1_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_1/Component_Function_4/N2  ( .A1(\SB1_1_1/i3[0] ), .A2(
        \SB1_1_1/i0_0 ), .A3(\SB1_1_1/i1_7 ), .ZN(
        \SB1_1_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_1/Component_Function_4/N1  ( .A1(\SB1_1_1/i0[9] ), .A2(
        \SB1_1_1/i0_0 ), .A3(\SB1_1_1/i0[8] ), .ZN(
        \SB1_1_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_2/N2  ( .A1(\SB1_1_2/i0_3 ), .A2(
        \SB1_1_2/i0[10] ), .A3(\SB1_1_2/i0[6] ), .ZN(
        \SB1_1_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_2/Component_Function_2/N1  ( .A1(\SB1_1_2/i1_5 ), .A2(
        \SB1_1_2/i0[10] ), .A3(\SB1_1_2/i1[9] ), .ZN(
        \SB1_1_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_3/N4  ( .A1(\SB1_1_2/i1_5 ), .A2(
        \SB1_1_2/i0[8] ), .A3(\SB1_1_2/i3[0] ), .ZN(
        \SB1_1_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_2/Component_Function_3/N1  ( .A1(\SB1_1_2/i1[9] ), .A2(
        \SB1_1_2/i0_3 ), .A3(\SB1_1_2/i0[6] ), .ZN(
        \SB1_1_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_4/N4  ( .A1(\SB1_1_2/i1[9] ), .A2(
        \SB1_1_2/i1_5 ), .A3(\SB1_1_2/i0_4 ), .ZN(
        \SB1_1_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_2/Component_Function_4/N2  ( .A1(\SB1_1_2/i3[0] ), .A2(
        \SB1_1_2/i0_0 ), .A3(\SB1_1_2/i1_7 ), .ZN(
        \SB1_1_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_3/Component_Function_2/N2  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i0[10] ), .A3(\SB1_1_3/i0[6] ), .ZN(
        \SB1_1_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_3/Component_Function_2/N1  ( .A1(\SB1_1_3/i1_5 ), .A2(
        \SB1_1_3/i0[10] ), .A3(\SB1_1_3/i1[9] ), .ZN(
        \SB1_1_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_3/N4  ( .A1(\SB1_1_3/i1_5 ), .A2(
        \SB1_1_3/i0[8] ), .A3(\SB1_1_3/i3[0] ), .ZN(
        \SB1_1_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_3/Component_Function_3/N1  ( .A1(\SB1_1_3/i1[9] ), .A2(
        \SB1_1_3/i0_3 ), .A3(\SB1_1_3/i0[6] ), .ZN(
        \SB1_1_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_4/N2  ( .A1(\SB1_1_3/i3[0] ), .A2(
        \SB1_1_3/i0_0 ), .A3(\SB1_1_3/i1_7 ), .ZN(
        \SB1_1_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_3/Component_Function_4/N1  ( .A1(\SB1_1_3/i0[9] ), .A2(
        \SB1_1_3/i0_0 ), .A3(\SB1_1_3/i0[8] ), .ZN(
        \SB1_1_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_2/N3  ( .A1(\SB1_1_4/i0_3 ), .A2(
        \SB1_1_4/i0[8] ), .A3(\SB1_1_4/i0[9] ), .ZN(
        \SB1_1_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_4/Component_Function_2/N2  ( .A1(n2149), .A2(
        \SB1_1_4/i0[10] ), .A3(\SB1_1_4/i0[6] ), .ZN(
        \SB1_1_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_4/Component_Function_3/N4  ( .A1(\SB1_1_4/i1_5 ), .A2(
        \SB1_1_4/i0[8] ), .A3(\SB1_1_4/i3[0] ), .ZN(
        \SB1_1_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_4/Component_Function_3/N1  ( .A1(\SB1_1_4/i1[9] ), .A2(n2149), .A3(\SB1_1_4/i0[6] ), .ZN(\SB1_1_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_4/N4  ( .A1(\SB1_1_4/i1[9] ), .A2(
        \SB1_1_4/i1_5 ), .A3(\SB1_1_4/i0_4 ), .ZN(
        \SB1_1_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_4/Component_Function_4/N2  ( .A1(\SB1_1_4/i3[0] ), .A2(
        \SB1_1_4/i0_0 ), .A3(\SB1_1_4/i1_7 ), .ZN(
        \SB1_1_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_4/Component_Function_4/N1  ( .A1(\SB1_1_4/i0[9] ), .A2(
        \SB1_1_4/i0_0 ), .A3(\SB1_1_4/i0[8] ), .ZN(
        \SB1_1_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_2/N2  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i0[10] ), .A3(\SB1_1_5/i0[6] ), .ZN(
        \SB1_1_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_5/Component_Function_2/N1  ( .A1(\SB1_1_5/i1_5 ), .A2(
        \SB1_1_5/i0[10] ), .A3(\SB1_1_5/i1[9] ), .ZN(
        \SB1_1_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_3/N4  ( .A1(\SB1_1_5/i1_5 ), .A2(
        \SB1_1_5/i0[8] ), .A3(\SB1_1_5/i3[0] ), .ZN(
        \SB1_1_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_3/N3  ( .A1(\SB1_1_5/i1[9] ), .A2(
        \SB1_1_5/i1_7 ), .A3(\SB1_1_5/i0[10] ), .ZN(
        \SB1_1_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_5/Component_Function_3/N1  ( .A1(\SB1_1_5/i1[9] ), .A2(
        \SB1_1_5/i0_3 ), .A3(\SB1_1_5/i0[6] ), .ZN(
        \SB1_1_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_4/N4  ( .A1(\SB1_1_5/i1[9] ), .A2(
        \SB1_1_5/i1_5 ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_4/N2  ( .A1(\SB1_1_5/i3[0] ), .A2(
        \SB1_1_5/i0_0 ), .A3(\SB1_1_5/i1_7 ), .ZN(
        \SB1_1_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_5/Component_Function_4/N1  ( .A1(\SB1_1_5/i0[9] ), .A2(
        \SB1_1_5/i0_0 ), .A3(\SB1_1_5/i0[8] ), .ZN(
        \SB1_1_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_2/N2  ( .A1(\SB1_1_6/i0_3 ), .A2(
        \SB1_1_6/i0[10] ), .A3(\SB1_1_6/i0[6] ), .ZN(
        \SB1_1_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_6/Component_Function_2/N1  ( .A1(\SB1_1_6/i1_5 ), .A2(
        \SB1_1_6/i0[10] ), .A3(\SB1_1_6/i1[9] ), .ZN(
        \SB1_1_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_3/N4  ( .A1(\SB1_1_6/i1_5 ), .A2(
        \SB1_1_6/i0[8] ), .A3(\SB1_1_6/i3[0] ), .ZN(
        \SB1_1_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_6/Component_Function_3/N3  ( .A1(\SB1_1_6/i1[9] ), .A2(
        \SB1_1_6/i1_7 ), .A3(\SB1_1_6/i0[10] ), .ZN(
        \SB1_1_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_6/Component_Function_3/N1  ( .A1(\SB1_1_6/i1[9] ), .A2(
        \SB1_1_6/i0_3 ), .A3(\SB1_1_6/i0[6] ), .ZN(
        \SB1_1_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_4/N4  ( .A1(\SB1_1_6/i1[9] ), .A2(
        \SB1_1_6/i1_5 ), .A3(\SB1_1_6/i0_4 ), .ZN(
        \SB1_1_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_6/Component_Function_4/N2  ( .A1(\SB1_1_6/i3[0] ), .A2(
        \SB1_1_6/i0_0 ), .A3(\SB1_1_6/i1_7 ), .ZN(
        \SB1_1_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_6/Component_Function_4/N1  ( .A1(\SB1_1_6/i0[9] ), .A2(
        \SB1_1_6/i0_0 ), .A3(\SB1_1_6/i0[8] ), .ZN(
        \SB1_1_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_2/N2  ( .A1(\SB1_1_7/i0_3 ), .A2(
        \SB1_1_7/i0[10] ), .A3(\SB1_1_7/i0[6] ), .ZN(
        \SB1_1_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_7/Component_Function_2/N1  ( .A1(\SB1_1_7/i1_5 ), .A2(
        \SB1_1_7/i0[10] ), .A3(\SB1_1_7/i1[9] ), .ZN(
        \SB1_1_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_3/N4  ( .A1(\SB1_1_7/i1_5 ), .A2(
        \SB1_1_7/i0[8] ), .A3(\SB1_1_7/i3[0] ), .ZN(
        \SB1_1_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_7/Component_Function_3/N1  ( .A1(\SB1_1_7/i1[9] ), .A2(
        \SB1_1_7/i0_3 ), .A3(\SB1_1_7/i0[6] ), .ZN(
        \SB1_1_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_4/N4  ( .A1(\SB1_1_7/i1[9] ), .A2(
        \SB1_1_7/i1_5 ), .A3(\SB1_1_7/i0_4 ), .ZN(
        \SB1_1_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_7/Component_Function_4/N2  ( .A1(\SB1_1_7/i3[0] ), .A2(
        \SB1_1_7/i0_0 ), .A3(\SB1_1_7/i1_7 ), .ZN(
        \SB1_1_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_7/Component_Function_4/N1  ( .A1(\SB1_1_7/i0[9] ), .A2(
        \SB1_1_7/i0_0 ), .A3(\SB1_1_7/i0[8] ), .ZN(
        \SB1_1_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_8/Component_Function_2/N2  ( .A1(\SB1_1_8/i0_3 ), .A2(
        \SB1_1_8/i0[10] ), .A3(\SB1_1_8/i0[6] ), .ZN(
        \SB1_1_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_2/N1  ( .A1(\SB1_1_8/i1_5 ), .A2(
        \SB1_1_8/i0[10] ), .A3(\SB1_1_8/i1[9] ), .ZN(
        \SB1_1_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_8/Component_Function_3/N3  ( .A1(\SB1_1_8/i1[9] ), .A2(
        \SB1_1_8/i1_7 ), .A3(\SB1_1_8/i0[10] ), .ZN(
        \SB1_1_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_8/Component_Function_4/N4  ( .A1(\SB1_1_8/i1[9] ), .A2(
        \SB1_1_8/i1_5 ), .A3(\SB1_1_8/i0_4 ), .ZN(
        \SB1_1_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_8/Component_Function_4/N2  ( .A1(\SB1_1_8/i3[0] ), .A2(
        \SB1_1_8/i0_0 ), .A3(\SB1_1_8/i1_7 ), .ZN(
        \SB1_1_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_4/N1  ( .A1(\SB1_1_8/i0[9] ), .A2(
        \SB1_1_8/i0_0 ), .A3(\SB1_1_8/i0[8] ), .ZN(
        \SB1_1_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_2/N4  ( .A1(\SB1_1_9/i1_5 ), .A2(
        \SB1_1_9/i0_0 ), .A3(\SB1_1_9/i0_4 ), .ZN(
        \SB1_1_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_9/Component_Function_2/N2  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i0[10] ), .A3(\SB1_1_9/i0[6] ), .ZN(
        \SB1_1_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_9/Component_Function_2/N1  ( .A1(\SB1_1_9/i1_5 ), .A2(
        \SB1_1_9/i0[10] ), .A3(\SB1_1_9/i1[9] ), .ZN(
        \SB1_1_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_3/N4  ( .A1(\SB1_1_9/i1_5 ), .A2(
        \SB1_1_9/i0[8] ), .A3(\SB1_1_9/i3[0] ), .ZN(
        \SB1_1_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_9/Component_Function_3/N1  ( .A1(\SB1_1_9/i1[9] ), .A2(
        \SB1_1_9/i0_3 ), .A3(\SB1_1_9/i0[6] ), .ZN(
        \SB1_1_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N4  ( .A1(\SB1_1_9/i1[9] ), .A2(
        \SB1_1_9/i1_5 ), .A3(\SB1_1_9/i0_4 ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N2  ( .A1(\SB1_1_9/i3[0] ), .A2(
        \SB1_1_9/i0_0 ), .A3(\SB1_1_9/i1_7 ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N1  ( .A1(\SB1_1_9/i0[9] ), .A2(
        \SB1_1_9/i0_0 ), .A3(\SB1_1_9/i0[8] ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_2/N3  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i0[8] ), .A3(\SB1_1_10/i0[9] ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_10/Component_Function_2/N2  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i0[10] ), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_10/Component_Function_2/N1  ( .A1(\SB1_1_10/i1_5 ), .A2(
        \SB1_1_10/i0[10] ), .A3(\SB1_1_10/i1[9] ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_3/N4  ( .A1(\SB1_1_10/i1_5 ), .A2(
        \SB1_1_10/i0[8] ), .A3(\SB1_1_10/i3[0] ), .ZN(
        \SB1_1_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_3/N1  ( .A1(\SB1_1_10/i1[9] ), .A2(
        n826), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_4/N4  ( .A1(\SB1_1_10/i1[9] ), .A2(
        \SB1_1_10/i1_5 ), .A3(\SB1_1_10/i0_4 ), .ZN(
        \SB1_1_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_4/N2  ( .A1(\SB1_1_10/i3[0] ), .A2(
        \SB1_1_10/i0_0 ), .A3(\SB1_1_10/i1_7 ), .ZN(
        \SB1_1_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_10/Component_Function_4/N1  ( .A1(\SB1_1_10/i0[9] ), .A2(
        \SB1_1_10/i0_0 ), .A3(\SB1_1_10/i0[8] ), .ZN(
        \SB1_1_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_2/N3  ( .A1(\SB1_1_11/i0_3 ), .A2(
        \SB1_1_11/i0[8] ), .A3(\SB1_1_11/i0[9] ), .ZN(
        \SB1_1_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_11/Component_Function_2/N2  ( .A1(n2141), .A2(
        \SB1_1_11/i0[10] ), .A3(\SB1_1_11/i0[6] ), .ZN(
        \SB1_1_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_11/Component_Function_2/N1  ( .A1(\SB1_1_11/i1_5 ), .A2(
        \SB1_1_11/i0[10] ), .A3(\SB1_1_11/i1[9] ), .ZN(
        \SB1_1_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_3/N4  ( .A1(\SB1_1_11/i1_5 ), .A2(
        \SB1_1_11/i0[8] ), .A3(\SB1_1_11/i3[0] ), .ZN(
        \SB1_1_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_11/Component_Function_3/N1  ( .A1(\SB1_1_11/i1[9] ), .A2(
        n2141), .A3(\SB1_1_11/i0[6] ), .ZN(
        \SB1_1_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_4/N4  ( .A1(\SB1_1_11/i1[9] ), .A2(
        \SB1_1_11/i1_5 ), .A3(\SB1_1_11/i0_4 ), .ZN(
        \SB1_1_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_11/Component_Function_4/N2  ( .A1(\SB1_1_11/i3[0] ), .A2(
        \SB1_1_11/i0_0 ), .A3(\SB1_1_11/i1_7 ), .ZN(
        \SB1_1_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_11/Component_Function_4/N1  ( .A1(\SB1_1_11/i0[9] ), .A2(
        \SB1_1_11/i0_0 ), .A3(\SB1_1_11/i0[8] ), .ZN(
        \SB1_1_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_2/N3  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i0[8] ), .A3(\SB1_1_12/i0[9] ), .ZN(
        \SB1_1_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_12/Component_Function_2/N2  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i0[10] ), .A3(\SB1_1_12/i0[6] ), .ZN(
        \SB1_1_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_2/N1  ( .A1(\SB1_1_12/i1_5 ), .A2(
        \SB1_1_12/i0[10] ), .A3(\SB1_1_12/i1[9] ), .ZN(
        \SB1_1_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_3/N4  ( .A1(\SB1_1_12/i1_5 ), .A2(
        \SB1_1_12/i0[8] ), .A3(\SB1_1_12/i3[0] ), .ZN(
        \SB1_1_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_12/Component_Function_3/N3  ( .A1(\SB1_1_12/i1[9] ), .A2(
        \SB1_1_12/i1_7 ), .A3(\SB1_1_12/i0[10] ), .ZN(
        \SB1_1_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_12/Component_Function_3/N1  ( .A1(\SB1_1_12/i1[9] ), .A2(
        \SB1_1_12/i0_3 ), .A3(\SB1_1_12/i0[6] ), .ZN(
        \SB1_1_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_4/N4  ( .A1(\SB1_1_12/i1[9] ), .A2(
        \SB1_1_12/i1_5 ), .A3(\SB1_1_12/i0_4 ), .ZN(
        \SB1_1_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_12/Component_Function_4/N2  ( .A1(\SB1_1_12/i3[0] ), .A2(
        \SB1_1_12/i0_0 ), .A3(\SB1_1_12/i1_7 ), .ZN(
        \SB1_1_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_4/N1  ( .A1(\SB1_1_12/i0[9] ), .A2(
        \SB1_1_12/i0_0 ), .A3(\SB1_1_12/i0[8] ), .ZN(
        \SB1_1_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_2/N2  ( .A1(\SB1_1_13/i0_3 ), .A2(
        \SB1_1_13/i0[10] ), .A3(\SB1_1_13/i0[6] ), .ZN(
        \SB1_1_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_13/Component_Function_2/N1  ( .A1(\SB1_1_13/i1_5 ), .A2(
        \SB1_1_13/i0[10] ), .A3(\SB1_1_13/i1[9] ), .ZN(
        \SB1_1_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_3/N4  ( .A1(\SB1_1_13/i1_5 ), .A2(
        \SB1_1_13/i0[8] ), .A3(\SB1_1_13/i3[0] ), .ZN(
        \SB1_1_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_13/Component_Function_3/N3  ( .A1(\SB1_1_13/i1[9] ), .A2(
        \SB1_1_13/i1_7 ), .A3(\SB1_1_13/i0[10] ), .ZN(
        \SB1_1_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_13/Component_Function_3/N1  ( .A1(\SB1_1_13/i1[9] ), .A2(
        \SB1_1_13/i0_3 ), .A3(\SB1_1_13/i0[6] ), .ZN(
        \SB1_1_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_4/N4  ( .A1(\SB1_1_13/i1[9] ), .A2(
        \SB1_1_13/i1_5 ), .A3(\SB1_1_13/i0_4 ), .ZN(
        \SB1_1_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_13/Component_Function_4/N2  ( .A1(\SB1_1_13/i3[0] ), .A2(
        \SB1_1_13/i0_0 ), .A3(\SB1_1_13/i1_7 ), .ZN(
        \SB1_1_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_13/Component_Function_4/N1  ( .A1(\SB1_1_13/i0[9] ), .A2(
        \SB1_1_13/i0_0 ), .A3(\SB1_1_13/i0[8] ), .ZN(
        \SB1_1_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_2/N4  ( .A1(\SB1_1_14/i1_5 ), .A2(
        \SB1_1_14/i0_0 ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_14/Component_Function_2/N2  ( .A1(\SB1_1_14/i0_3 ), .A2(
        \SB1_1_14/i0[10] ), .A3(\SB1_1_14/i0[6] ), .ZN(
        \SB1_1_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_14/Component_Function_2/N1  ( .A1(\SB1_1_14/i1_5 ), .A2(
        \SB1_1_14/i0[10] ), .A3(\SB1_1_14/i1[9] ), .ZN(
        \SB1_1_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_3/N3  ( .A1(\SB1_1_14/i1[9] ), .A2(
        \SB1_1_14/i1_7 ), .A3(\SB1_1_14/i0[10] ), .ZN(
        \SB1_1_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_14/Component_Function_3/N1  ( .A1(\SB1_1_14/i1[9] ), .A2(
        \SB1_1_14/i0_3 ), .A3(\SB1_1_14/i0[6] ), .ZN(
        \SB1_1_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_4/N4  ( .A1(\SB1_1_14/i1[9] ), .A2(
        \SB1_1_14/i1_5 ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_14/Component_Function_4/N2  ( .A1(\SB1_1_14/i3[0] ), .A2(
        \SB1_1_14/i0_0 ), .A3(\SB1_1_14/i1_7 ), .ZN(
        \SB1_1_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_14/Component_Function_4/N1  ( .A1(\SB1_1_14/i0[9] ), .A2(
        \SB1_1_14/i0_0 ), .A3(\SB1_1_14/i0[8] ), .ZN(
        \SB1_1_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_2/N4  ( .A1(\SB1_1_15/i1_5 ), .A2(
        \SB1_1_15/i0_0 ), .A3(\SB1_1_15/i0_4 ), .ZN(
        \SB1_1_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_15/Component_Function_2/N2  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i0[10] ), .A3(\SB1_1_15/i0[6] ), .ZN(
        \SB1_1_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_15/Component_Function_2/N1  ( .A1(\SB1_1_15/i1_5 ), .A2(
        \SB1_1_15/i0[10] ), .A3(\SB1_1_15/i1[9] ), .ZN(
        \SB1_1_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_3/N4  ( .A1(\SB1_1_15/i1_5 ), .A2(
        \SB1_1_15/i0[8] ), .A3(\SB1_1_15/i3[0] ), .ZN(
        \SB1_1_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_15/Component_Function_3/N1  ( .A1(\SB1_1_15/i1[9] ), .A2(
        \SB1_1_15/i0_3 ), .A3(\SB1_1_15/i0[6] ), .ZN(
        \SB1_1_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N4  ( .A1(\SB1_1_15/i1[9] ), .A2(
        \SB1_1_15/i1_5 ), .A3(\SB1_1_15/i0_4 ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N2  ( .A1(\SB1_1_15/i3[0] ), .A2(
        \SB1_1_15/i0_0 ), .A3(\SB1_1_15/i1_7 ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N1  ( .A1(\SB1_1_15/i0[9] ), .A2(
        \SB1_1_15/i0_0 ), .A3(\SB1_1_15/i0[8] ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_2/N2  ( .A1(\SB1_1_16/i0_3 ), .A2(
        \SB1_1_16/i0[10] ), .A3(\SB1_1_16/i0[6] ), .ZN(
        \SB1_1_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_16/Component_Function_2/N1  ( .A1(\SB1_1_16/i1_5 ), .A2(
        \SB1_1_16/i0[10] ), .A3(\SB1_1_16/i1[9] ), .ZN(
        \SB1_1_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_3/N4  ( .A1(\SB1_1_16/i1_5 ), .A2(
        \SB1_1_16/i0[8] ), .A3(\SB1_1_16/i3[0] ), .ZN(
        \SB1_1_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_16/Component_Function_3/N1  ( .A1(\SB1_1_16/i1[9] ), .A2(
        \SB1_1_16/i0_3 ), .A3(\SB1_1_16/i0[6] ), .ZN(
        \SB1_1_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_4/N2  ( .A1(\SB1_1_16/i3[0] ), .A2(
        \SB1_1_16/i0_0 ), .A3(\SB1_1_16/i1_7 ), .ZN(
        \SB1_1_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_16/Component_Function_4/N1  ( .A1(\SB1_1_16/i0[9] ), .A2(
        \SB1_1_16/i0_0 ), .A3(\SB1_1_16/i0[8] ), .ZN(
        \SB1_1_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_2/N2  ( .A1(n789), .A2(
        \SB1_1_17/i0[10] ), .A3(\SB1_1_17/i0[6] ), .ZN(
        \SB1_1_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_17/Component_Function_2/N1  ( .A1(\SB1_1_17/i1_5 ), .A2(
        \SB1_1_17/i0[10] ), .A3(\SB1_1_17/i1[9] ), .ZN(
        \SB1_1_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_3/N4  ( .A1(\SB1_1_17/i1_5 ), .A2(
        \SB1_1_17/i0[8] ), .A3(\SB1_1_17/i3[0] ), .ZN(
        \SB1_1_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_17/Component_Function_3/N3  ( .A1(\SB1_1_17/i1[9] ), .A2(
        \SB1_1_17/i1_7 ), .A3(\SB1_1_17/i0[10] ), .ZN(
        \SB1_1_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_17/Component_Function_3/N1  ( .A1(\SB1_1_17/i1[9] ), .A2(
        n789), .A3(\SB1_1_17/i0[6] ), .ZN(
        \SB1_1_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_4/N4  ( .A1(\SB1_1_17/i1[9] ), .A2(
        \SB1_1_17/i1_5 ), .A3(\SB1_1_17/i0_4 ), .ZN(
        \SB1_1_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_17/Component_Function_4/N2  ( .A1(\SB1_1_17/i3[0] ), .A2(
        \SB1_1_17/i0_0 ), .A3(\SB1_1_17/i1_7 ), .ZN(
        \SB1_1_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_17/Component_Function_4/N1  ( .A1(\SB1_1_17/i0[9] ), .A2(
        \SB1_1_17/i0_0 ), .A3(\SB1_1_17/i0[8] ), .ZN(
        \SB1_1_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_2/N2  ( .A1(\SB1_1_18/i0_3 ), .A2(
        \SB1_1_18/i0[10] ), .A3(\SB1_1_18/i0[6] ), .ZN(
        \SB1_1_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_18/Component_Function_2/N1  ( .A1(\SB1_1_18/i1_5 ), .A2(
        \SB1_1_18/i0[10] ), .A3(\SB1_1_18/i1[9] ), .ZN(
        \SB1_1_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_3/N4  ( .A1(\SB1_1_18/i1_5 ), .A2(
        \SB1_1_18/i0[8] ), .A3(\SB1_1_18/i3[0] ), .ZN(
        \SB1_1_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_18/Component_Function_3/N3  ( .A1(\SB1_1_18/i1[9] ), .A2(
        \SB1_1_18/i1_7 ), .A3(\SB1_1_18/i0[10] ), .ZN(
        \SB1_1_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_18/Component_Function_3/N1  ( .A1(\SB1_1_18/i1[9] ), .A2(
        \SB1_1_18/i0_3 ), .A3(\SB1_1_18/i0[6] ), .ZN(
        \SB1_1_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_4/N1  ( .A1(\SB1_1_18/i0[9] ), .A2(
        \SB1_1_18/i0_0 ), .A3(\SB1_1_18/i0[8] ), .ZN(
        \SB1_1_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_2/N2  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i0[10] ), .A3(\SB1_1_19/i0[6] ), .ZN(
        \SB1_1_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_19/Component_Function_2/N1  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0[10] ), .A3(\SB1_1_19/i1[9] ), .ZN(
        \SB1_1_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_3/N4  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0[8] ), .A3(\SB1_1_19/i3[0] ), .ZN(
        \SB1_1_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_3/N1  ( .A1(\SB1_1_19/i1[9] ), .A2(
        \SB1_1_19/i0_3 ), .A3(\SB1_1_19/i0[6] ), .ZN(
        \SB1_1_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_4/N4  ( .A1(\SB1_1_19/i1[9] ), .A2(
        \SB1_1_19/i1_5 ), .A3(\SB1_1_19/i0_4 ), .ZN(
        \SB1_1_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_4/N2  ( .A1(\SB1_1_19/i3[0] ), .A2(
        \SB1_1_19/i0_0 ), .A3(\SB1_1_19/i1_7 ), .ZN(
        \SB1_1_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_19/Component_Function_4/N1  ( .A1(\SB1_1_19/i0[9] ), .A2(
        \SB1_1_19/i0_0 ), .A3(\SB1_1_19/i0[8] ), .ZN(
        \SB1_1_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_2/N4  ( .A1(\SB1_1_20/i1_5 ), .A2(
        \SB1_1_20/i0_0 ), .A3(\SB1_1_20/i0_4 ), .ZN(
        \SB1_1_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_20/Component_Function_2/N3  ( .A1(\SB1_1_20/i0_3 ), .A2(
        \SB1_1_20/i0[8] ), .A3(\SB1_1_20/i0[9] ), .ZN(
        \SB1_1_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_20/Component_Function_2/N2  ( .A1(\SB1_1_20/i0_3 ), .A2(
        \SB1_1_20/i0[10] ), .A3(\SB1_1_20/i0[6] ), .ZN(
        \SB1_1_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_20/Component_Function_2/N1  ( .A1(\SB1_1_20/i1_5 ), .A2(
        \SB1_1_20/i0[10] ), .A3(\SB1_1_20/i1[9] ), .ZN(
        \SB1_1_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_3/N3  ( .A1(\SB1_1_20/i1[9] ), .A2(
        \SB1_1_20/i1_7 ), .A3(\SB1_1_20/i0[10] ), .ZN(
        \SB1_1_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_20/Component_Function_3/N1  ( .A1(\SB1_1_20/i1[9] ), .A2(
        \SB1_1_20/i0_3 ), .A3(\SB1_1_20/i0[6] ), .ZN(
        \SB1_1_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_4/N4  ( .A1(\SB1_1_20/i1[9] ), .A2(
        \SB1_1_20/i1_5 ), .A3(\SB1_1_20/i0_4 ), .ZN(
        \SB1_1_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_20/Component_Function_4/N2  ( .A1(\SB1_1_20/i3[0] ), .A2(
        \SB1_1_20/i0_0 ), .A3(\SB1_1_20/i1_7 ), .ZN(
        \SB1_1_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_20/Component_Function_4/N1  ( .A1(\SB1_1_20/i0[9] ), .A2(
        \SB1_1_20/i0_0 ), .A3(\SB1_1_20/i0[8] ), .ZN(
        \SB1_1_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_2/N4  ( .A1(\SB1_1_21/i1_5 ), .A2(
        \SB1_1_21/i0_0 ), .A3(\SB1_1_21/i0_4 ), .ZN(
        \SB1_1_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_2/N2  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i0[10] ), .A3(\SB1_1_21/i0[6] ), .ZN(
        \SB1_1_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_21/Component_Function_2/N1  ( .A1(\SB1_1_21/i1_5 ), .A2(
        \SB1_1_21/i0[10] ), .A3(\SB1_1_21/i1[9] ), .ZN(
        \SB1_1_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_3/N4  ( .A1(\SB1_1_21/i1_5 ), .A2(
        \SB1_1_21/i0[8] ), .A3(\SB1_1_21/i3[0] ), .ZN(
        \SB1_1_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_3/N1  ( .A1(\SB1_1_21/i1[9] ), .A2(
        \SB1_1_21/i0_3 ), .A3(\SB1_1_21/i0[6] ), .ZN(
        \SB1_1_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_4/N4  ( .A1(\SB1_1_21/i1[9] ), .A2(
        \SB1_1_21/i1_5 ), .A3(\SB1_1_21/i0_4 ), .ZN(
        \SB1_1_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_4/N2  ( .A1(\SB1_1_21/i3[0] ), .A2(
        \SB1_1_21/i0_0 ), .A3(\SB1_1_21/i1_7 ), .ZN(
        \SB1_1_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_21/Component_Function_4/N1  ( .A1(\SB1_1_21/i0[9] ), .A2(
        \SB1_1_21/i0_0 ), .A3(\SB1_1_21/i0[8] ), .ZN(
        \SB1_1_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_2/N2  ( .A1(\SB1_1_22/i0_3 ), .A2(
        \SB1_1_22/i0[10] ), .A3(\SB1_1_22/i0[6] ), .ZN(
        \SB1_1_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_22/Component_Function_2/N1  ( .A1(\SB1_1_22/i1_5 ), .A2(
        \SB1_1_22/i0[10] ), .A3(\SB1_1_22/i1[9] ), .ZN(
        \SB1_1_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_3/N4  ( .A1(\SB1_1_22/i1_5 ), .A2(
        \SB1_1_22/i0[8] ), .A3(\SB1_1_22/i3[0] ), .ZN(
        \SB1_1_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_22/Component_Function_3/N1  ( .A1(\SB1_1_22/i1[9] ), .A2(
        \SB1_1_22/i0_3 ), .A3(\SB1_1_22/i0[6] ), .ZN(
        \SB1_1_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_4/N4  ( .A1(\SB1_1_22/i1[9] ), .A2(
        \SB1_1_22/i1_5 ), .A3(\SB1_1_22/i0_4 ), .ZN(
        \SB1_1_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_22/Component_Function_4/N2  ( .A1(\SB1_1_22/i3[0] ), .A2(
        \SB1_1_22/i0_0 ), .A3(\SB1_1_22/i1_7 ), .ZN(
        \SB1_1_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_22/Component_Function_4/N1  ( .A1(\SB1_1_22/i0[9] ), .A2(
        \SB1_1_22/i0_0 ), .A3(\SB1_1_22/i0[8] ), .ZN(
        \SB1_1_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_2/N2  ( .A1(\SB1_1_23/i0_3 ), .A2(
        \SB1_1_23/i0[10] ), .A3(\SB1_1_23/i0[6] ), .ZN(
        \SB1_1_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_23/Component_Function_2/N1  ( .A1(\SB1_1_23/i1_5 ), .A2(
        \SB1_1_23/i0[10] ), .A3(\SB1_1_23/i1[9] ), .ZN(
        \SB1_1_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_3/N4  ( .A1(\SB1_1_23/i1_5 ), .A2(
        \SB1_1_23/i0[8] ), .A3(\SB1_1_23/i3[0] ), .ZN(
        \SB1_1_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_23/Component_Function_3/N1  ( .A1(\SB1_1_23/i1[9] ), .A2(
        \SB1_1_23/i0_3 ), .A3(\SB1_1_23/i0[6] ), .ZN(
        \SB1_1_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_4/N2  ( .A1(\SB1_1_23/i3[0] ), .A2(
        \SB1_1_23/i0_0 ), .A3(\SB1_1_23/i1_7 ), .ZN(
        \SB1_1_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_23/Component_Function_4/N1  ( .A1(\SB1_1_23/i0[9] ), .A2(
        \SB1_1_23/i0_0 ), .A3(\SB1_1_23/i0[8] ), .ZN(
        \SB1_1_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_2/N2  ( .A1(\SB1_1_24/i0_3 ), .A2(
        \SB1_1_24/i0[10] ), .A3(\SB1_1_24/i0[6] ), .ZN(
        \SB1_1_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_2/N1  ( .A1(\SB1_1_24/i1_5 ), .A2(
        \SB1_1_24/i0[10] ), .A3(\SB1_1_24/i1[9] ), .ZN(
        \SB1_1_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_3/N4  ( .A1(\SB1_1_24/i1_5 ), .A2(
        \SB1_1_24/i0[8] ), .A3(\SB1_1_24/i3[0] ), .ZN(
        \SB1_1_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_24/Component_Function_3/N3  ( .A1(\SB1_1_24/i1[9] ), .A2(
        \SB1_1_24/i1_7 ), .A3(\SB1_1_24/i0[10] ), .ZN(
        \SB1_1_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_24/Component_Function_3/N1  ( .A1(\SB1_1_24/i1[9] ), .A2(
        \SB1_1_24/i0_3 ), .A3(\SB1_1_24/i0[6] ), .ZN(
        \SB1_1_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N4  ( .A1(\SB1_1_24/i1[9] ), .A2(
        \SB1_1_24/i1_5 ), .A3(\SB1_1_24/i0_4 ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N3  ( .A1(\SB1_1_24/i0[9] ), .A2(
        \SB1_1_24/i0[10] ), .A3(\SB1_1_24/i0_3 ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N2  ( .A1(\SB1_1_24/i3[0] ), .A2(
        \SB1_1_24/i0_0 ), .A3(\SB1_1_24/i1_7 ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N1  ( .A1(\SB1_1_24/i0[9] ), .A2(
        \SB1_1_24/i0_0 ), .A3(\SB1_1_24/i0[8] ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_2/N2  ( .A1(\SB1_1_25/i0_3 ), .A2(
        \SB1_1_25/i0[10] ), .A3(\SB1_1_25/i0[6] ), .ZN(
        \SB1_1_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_25/Component_Function_2/N1  ( .A1(\SB1_1_25/i1_5 ), .A2(
        \SB1_1_25/i0[10] ), .A3(\SB1_1_25/i1[9] ), .ZN(
        \SB1_1_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_3/N4  ( .A1(\SB1_1_25/i1_5 ), .A2(
        \SB1_1_25/i0[8] ), .A3(\SB1_1_25/i3[0] ), .ZN(
        \SB1_1_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_3/N1  ( .A1(\SB1_1_25/i1[9] ), .A2(
        \SB1_1_25/i0_3 ), .A3(\SB1_1_25/i0[6] ), .ZN(
        \SB1_1_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N4  ( .A1(\SB1_1_25/i1[9] ), .A2(
        \SB1_1_25/i1_5 ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N2  ( .A1(\SB1_1_25/i3[0] ), .A2(
        \SB1_1_25/i0_0 ), .A3(\SB1_1_25/i1_7 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N1  ( .A1(\SB1_1_25/i0[9] ), .A2(
        \SB1_1_25/i0_0 ), .A3(\SB1_1_25/i0[8] ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_2/N4  ( .A1(\SB1_1_26/i1_5 ), .A2(
        \SB1_1_26/i0_0 ), .A3(\SB1_1_26/i0_4 ), .ZN(
        \SB1_1_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_26/Component_Function_2/N2  ( .A1(\SB1_1_26/i0_3 ), .A2(
        \SB1_1_26/i0[10] ), .A3(\SB1_1_26/i0[6] ), .ZN(
        \SB1_1_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_26/Component_Function_2/N1  ( .A1(\SB1_1_26/i1_5 ), .A2(
        \SB1_1_26/i0[10] ), .A3(\SB1_1_26/i1[9] ), .ZN(
        \SB1_1_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_3/N4  ( .A1(\SB1_1_26/i1_5 ), .A2(
        \SB1_1_26/i0[8] ), .A3(\SB1_1_26/i3[0] ), .ZN(
        \SB1_1_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_26/Component_Function_3/N3  ( .A1(\SB1_1_26/i1[9] ), .A2(
        \SB1_1_26/i1_7 ), .A3(\SB1_1_26/i0[10] ), .ZN(
        \SB1_1_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_26/Component_Function_3/N1  ( .A1(\SB1_1_26/i1[9] ), .A2(
        \SB1_1_26/i0_3 ), .A3(\SB1_1_26/i0[6] ), .ZN(
        \SB1_1_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N4  ( .A1(\SB1_1_26/i1[9] ), .A2(
        \SB1_1_26/i1_5 ), .A3(\SB1_1_26/i0_4 ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N2  ( .A1(\SB1_1_26/i3[0] ), .A2(
        \SB1_1_26/i0_0 ), .A3(\SB1_1_26/i1_7 ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N1  ( .A1(\SB1_1_26/i0[9] ), .A2(
        \SB1_1_26/i0_0 ), .A3(\SB1_1_26/i0[8] ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_2/N2  ( .A1(\SB1_1_27/i0_3 ), .A2(
        \SB1_1_27/i0[10] ), .A3(\SB1_1_27/i0[6] ), .ZN(
        \SB1_1_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_27/Component_Function_2/N1  ( .A1(\SB1_1_27/i1_5 ), .A2(
        \SB1_1_27/i0[10] ), .A3(\SB1_1_27/i1[9] ), .ZN(
        \SB1_1_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_3/N4  ( .A1(\SB1_1_27/i1_5 ), .A2(
        \SB1_1_27/i0[8] ), .A3(\SB1_1_27/i3[0] ), .ZN(
        \SB1_1_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_3/N3  ( .A1(\SB1_1_27/i1[9] ), .A2(
        \SB1_1_27/i1_7 ), .A3(\SB1_1_27/i0[10] ), .ZN(
        \SB1_1_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_27/Component_Function_3/N1  ( .A1(\SB1_1_27/i1[9] ), .A2(
        \SB1_1_27/i0_3 ), .A3(\SB1_1_27/i0[6] ), .ZN(
        \SB1_1_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_4/N4  ( .A1(\SB1_1_27/i1[9] ), .A2(
        \SB1_1_27/i1_5 ), .A3(\SB1_1_27/i0_4 ), .ZN(
        \SB1_1_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_4/N2  ( .A1(\SB1_1_27/i3[0] ), .A2(
        \SB1_1_27/i0_0 ), .A3(\SB1_1_27/i1_7 ), .ZN(
        \SB1_1_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_27/Component_Function_4/N1  ( .A1(\SB1_1_27/i0[9] ), .A2(
        \SB1_1_27/i0_0 ), .A3(\SB1_1_27/i0[8] ), .ZN(
        \SB1_1_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_2/N2  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i0[10] ), .A3(\SB1_1_28/i0[6] ), .ZN(
        \SB1_1_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_28/Component_Function_2/N1  ( .A1(\SB1_1_28/i1_5 ), .A2(
        \SB1_1_28/i0[10] ), .A3(\SB1_1_28/i1[9] ), .ZN(
        \SB1_1_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_3/N4  ( .A1(\SB1_1_28/i1_5 ), .A2(
        \SB1_1_28/i0[8] ), .A3(\SB1_1_28/i3[0] ), .ZN(
        \SB1_1_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_3/N3  ( .A1(\SB1_1_28/i1[9] ), .A2(
        \SB1_1_28/i1_7 ), .A3(\SB1_1_28/i0[10] ), .ZN(
        \SB1_1_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_28/Component_Function_3/N1  ( .A1(\SB1_1_28/i1[9] ), .A2(
        \SB1_1_28/i0_3 ), .A3(\SB1_1_28/i0[6] ), .ZN(
        \SB1_1_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_4/N4  ( .A1(\SB1_1_28/i1[9] ), .A2(
        \SB1_1_28/i1_5 ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_4/N2  ( .A1(\SB1_1_28/i3[0] ), .A2(
        \SB1_1_28/i0_0 ), .A3(\SB1_1_28/i1_7 ), .ZN(
        \SB1_1_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_28/Component_Function_4/N1  ( .A1(\SB1_1_28/i0[9] ), .A2(
        \SB1_1_28/i0_0 ), .A3(\SB1_1_28/i0[8] ), .ZN(
        \SB1_1_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_2/N2  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i0[10] ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_29/Component_Function_2/N1  ( .A1(\SB1_1_29/i1_5 ), .A2(
        \SB1_1_29/i0[10] ), .A3(\SB1_1_29/i1[9] ), .ZN(
        \SB1_1_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_3/N4  ( .A1(\SB1_1_29/i1_5 ), .A2(
        \SB1_1_29/i0[8] ), .A3(\SB1_1_29/i3[0] ), .ZN(
        \SB1_1_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_29/Component_Function_3/N1  ( .A1(\SB1_1_29/i1[9] ), .A2(
        \SB1_1_29/i0_3 ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_4/N4  ( .A1(\SB1_1_29/i1[9] ), .A2(
        \SB1_1_29/i1_5 ), .A3(\SB1_1_29/i0_4 ), .ZN(
        \SB1_1_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_29/Component_Function_4/N2  ( .A1(\SB1_1_29/i3[0] ), .A2(
        \SB1_1_29/i0_0 ), .A3(\SB1_1_29/i1_7 ), .ZN(
        \SB1_1_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_29/Component_Function_4/N1  ( .A1(\SB1_1_29/i0[9] ), .A2(
        \SB1_1_29/i0_0 ), .A3(\SB1_1_29/i0[8] ), .ZN(
        \SB1_1_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_2/N2  ( .A1(\SB1_1_30/i0_3 ), .A2(
        \SB1_1_30/i0[10] ), .A3(\SB1_1_30/i0[6] ), .ZN(
        \SB1_1_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_30/Component_Function_2/N1  ( .A1(\SB1_1_30/i1_5 ), .A2(
        \SB1_1_30/i0[10] ), .A3(\SB1_1_30/i1[9] ), .ZN(
        \SB1_1_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_3/N4  ( .A1(\SB1_1_30/i1_5 ), .A2(
        \SB1_1_30/i0[8] ), .A3(\SB1_1_30/i3[0] ), .ZN(
        \SB1_1_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_30/Component_Function_3/N1  ( .A1(\SB1_1_30/i1[9] ), .A2(
        \SB1_1_30/i0_3 ), .A3(\SB1_1_30/i0[6] ), .ZN(
        \SB1_1_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_4/N4  ( .A1(\SB1_1_30/i1[9] ), .A2(
        \SB1_1_30/i1_5 ), .A3(\SB1_1_30/i0_4 ), .ZN(
        \SB1_1_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_30/Component_Function_4/N2  ( .A1(\SB1_1_30/i3[0] ), .A2(
        \SB1_1_30/i0_0 ), .A3(\SB1_1_30/i1_7 ), .ZN(
        \SB1_1_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_30/Component_Function_4/N1  ( .A1(\SB1_1_30/i0[9] ), .A2(
        \SB1_1_30/i0_0 ), .A3(\SB1_1_30/i0[8] ), .ZN(
        \SB1_1_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_2/N2  ( .A1(\SB1_1_31/i0_3 ), .A2(
        \SB1_1_31/i0[10] ), .A3(\SB1_1_31/i0[6] ), .ZN(
        \SB1_1_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_31/Component_Function_2/N1  ( .A1(\SB1_1_31/i1_5 ), .A2(
        \SB1_1_31/i0[10] ), .A3(\SB1_1_31/i1[9] ), .ZN(
        \SB1_1_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_3/N4  ( .A1(\SB1_1_31/i1_5 ), .A2(
        \SB1_1_31/i0[8] ), .A3(\SB1_1_31/i3[0] ), .ZN(
        \SB1_1_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_31/Component_Function_3/N1  ( .A1(\SB1_1_31/i1[9] ), .A2(
        \SB1_1_31/i0_3 ), .A3(\SB1_1_31/i0[6] ), .ZN(
        \SB1_1_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_4/N2  ( .A1(\SB1_1_31/i3[0] ), .A2(
        \SB1_1_31/i0_0 ), .A3(\SB1_1_31/i1_7 ), .ZN(
        \SB1_1_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_31/Component_Function_4/N1  ( .A1(\SB1_1_31/i0[9] ), .A2(
        \SB1_1_31/i0_0 ), .A3(\SB1_1_31/i0[8] ), .ZN(
        \SB1_1_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_0/Component_Function_2/N2  ( .A1(\SB2_1_0/i0_3 ), .A2(
        \SB2_1_0/i0[10] ), .A3(\SB2_1_0/i0[6] ), .ZN(
        \SB2_1_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_0/Component_Function_3/N3  ( .A1(\SB2_1_0/i1[9] ), .A2(
        \SB2_1_0/i1_7 ), .A3(\SB2_1_0/i0[10] ), .ZN(
        \SB2_1_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_0/Component_Function_3/N2  ( .A1(\SB2_1_0/i0_3 ), .A2(
        \SB2_1_0/i0_0 ), .A3(\SB2_1_0/i0_4 ), .ZN(
        \SB2_1_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_0/Component_Function_4/N4  ( .A1(\SB2_1_0/i1[9] ), .A2(
        \SB2_1_0/i1_5 ), .A3(\SB2_1_0/i0_4 ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_0/Component_Function_4/N3  ( .A1(\SB2_1_0/i0[9] ), .A2(
        \SB2_1_0/i0[10] ), .A3(\SB2_1_0/i0_3 ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_0/Component_Function_4/N2  ( .A1(\SB2_1_0/i3[0] ), .A2(
        \SB2_1_0/i0_0 ), .A3(\SB2_1_0/i1_7 ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_0/Component_Function_4/N1  ( .A1(\SB2_1_0/i0[9] ), .A2(
        \SB2_1_0/i0_0 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_2/N4  ( .A1(\SB2_1_1/i1_5 ), .A2(
        \SB2_1_1/i0_0 ), .A3(\SB2_1_1/i0_4 ), .ZN(
        \SB2_1_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_1/Component_Function_2/N2  ( .A1(\SB2_1_1/i0_3 ), .A2(
        \SB2_1_1/i0[10] ), .A3(\SB2_1_1/i0[6] ), .ZN(
        \SB2_1_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_2/N1  ( .A1(\SB2_1_1/i1_5 ), .A2(
        \SB2_1_1/i0[10] ), .A3(\SB2_1_1/i1[9] ), .ZN(
        \SB2_1_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_3/N3  ( .A1(\SB2_1_1/i1[9] ), .A2(
        \SB2_1_1/i1_7 ), .A3(\SB2_1_1/i0[10] ), .ZN(
        \SB2_1_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_1/Component_Function_3/N2  ( .A1(\SB2_1_1/i0_0 ), .A2(
        \SB2_1_1/i0_3 ), .A3(\SB2_1_1/i0_4 ), .ZN(
        \SB2_1_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_3/N1  ( .A1(\SB2_1_1/i1[9] ), .A2(
        \SB2_1_1/i0_3 ), .A3(\SB2_1_1/i0[6] ), .ZN(
        \SB2_1_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N4  ( .A1(\SB2_1_1/i1[9] ), .A2(
        \SB2_1_1/i1_5 ), .A3(\SB2_1_1/i0_4 ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N2  ( .A1(\SB2_1_1/i3[0] ), .A2(
        \SB2_1_1/i0_0 ), .A3(\SB2_1_1/i1_7 ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N1  ( .A1(\SB2_1_1/i0[9] ), .A2(
        \SB2_1_1/i0_0 ), .A3(\SB2_1_1/i0[8] ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_2/N2  ( .A1(\SB2_1_2/i0_3 ), .A2(
        \SB2_1_2/i0[10] ), .A3(\SB2_1_2/i0[6] ), .ZN(
        \SB2_1_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_2/Component_Function_2/N1  ( .A1(\SB2_1_2/i1_5 ), .A2(
        \SB2_1_2/i0[10] ), .A3(\SB2_1_2/i1[9] ), .ZN(
        \SB2_1_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_3/N2  ( .A1(\SB2_1_2/i0_0 ), .A2(
        \SB2_1_2/i0_3 ), .A3(\SB2_1_2/i0_4 ), .ZN(
        \SB2_1_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_2/Component_Function_3/N1  ( .A1(\SB2_1_2/i1[9] ), .A2(
        \SB2_1_2/i0_3 ), .A3(\SB2_1_2/i0[6] ), .ZN(
        \SB2_1_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N4  ( .A1(\SB2_1_2/i1[9] ), .A2(
        \SB2_1_2/i1_5 ), .A3(\SB2_1_2/i0_4 ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N2  ( .A1(\SB2_1_2/i3[0] ), .A2(
        \SB2_1_2/i0_0 ), .A3(\SB2_1_2/i1_7 ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N1  ( .A1(\SB2_1_2/i0[9] ), .A2(
        \SB2_1_2/i0_0 ), .A3(\SB2_1_2/i0[8] ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_2/N2  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i0[10] ), .A3(\SB2_1_3/i0[6] ), .ZN(
        \SB2_1_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_3/Component_Function_2/N1  ( .A1(\SB2_1_3/i1_5 ), .A2(
        \SB2_1_3/i0[10] ), .A3(\SB2_1_3/i1[9] ), .ZN(
        \SB2_1_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_4/N3  ( .A1(\SB2_1_3/i0[9] ), .A2(
        \SB2_1_3/i0[10] ), .A3(\SB2_1_3/i0_3 ), .ZN(
        \SB2_1_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_3/Component_Function_4/N1  ( .A1(\SB2_1_3/i0[9] ), .A2(
        \SB2_1_3/i0_0 ), .A3(\SB2_1_3/i0[8] ), .ZN(
        \SB2_1_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_2/N4  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB2_1_4/i0_0 ), .A3(\SB2_1_4/i0_4 ), .ZN(
        \SB2_1_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_2/N2  ( .A1(\SB2_1_4/i0_3 ), .A2(
        \SB2_1_4/i0[10] ), .A3(\SB2_1_4/i0[6] ), .ZN(
        \SB2_1_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_4/Component_Function_2/N1  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB2_1_4/i0[10] ), .A3(\SB2_1_4/i1[9] ), .ZN(
        \SB2_1_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_3/N3  ( .A1(\SB2_1_4/i1[9] ), .A2(
        \SB2_1_4/i1_7 ), .A3(\SB2_1_4/i0[10] ), .ZN(
        \SB2_1_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_3/N1  ( .A1(\SB2_1_4/i1[9] ), .A2(
        \SB2_1_4/i0_3 ), .A3(\SB2_1_4/i0[6] ), .ZN(
        \SB2_1_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N4  ( .A1(\SB2_1_4/i1[9] ), .A2(
        \SB2_1_4/i1_5 ), .A3(\SB2_1_4/i0_4 ), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N3  ( .A1(\SB2_1_4/i0[9] ), .A2(
        \SB2_1_4/i0[10] ), .A3(\SB2_1_4/i0_3 ), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N2  ( .A1(\SB2_1_4/i3[0] ), .A2(
        \SB2_1_4/i0_0 ), .A3(\SB2_1_4/i1_7 ), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N1  ( .A1(\SB2_1_4/i0[9] ), .A2(
        \SB2_1_4/i0_0 ), .A3(\SB2_1_4/i0[8] ), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_2/N3  ( .A1(\SB2_1_5/i0_3 ), .A2(
        \SB2_1_5/i0[8] ), .A3(\SB2_1_5/i0[9] ), .ZN(
        \SB2_1_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_5/Component_Function_2/N2  ( .A1(\SB2_1_5/i0_3 ), .A2(
        \SB2_1_5/i0[10] ), .A3(\SB2_1_5/i0[6] ), .ZN(
        \SB2_1_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_5/Component_Function_3/N3  ( .A1(\SB2_1_5/i1[9] ), .A2(
        \SB2_1_5/i1_7 ), .A3(\SB2_1_5/i0[10] ), .ZN(
        \SB2_1_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_5/Component_Function_3/N1  ( .A1(\SB2_1_5/i1[9] ), .A2(
        \SB2_1_5/i0_3 ), .A3(\SB2_1_5/i0[6] ), .ZN(
        \SB2_1_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_4/N4  ( .A1(\SB2_1_5/i1[9] ), .A2(
        \SB2_1_5/i1_5 ), .A3(\SB2_1_5/i0_4 ), .ZN(
        \SB2_1_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_5/Component_Function_4/N2  ( .A1(\SB2_1_5/i3[0] ), .A2(
        \SB2_1_5/i0_0 ), .A3(\SB2_1_5/i1_7 ), .ZN(
        \SB2_1_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_5/Component_Function_4/N1  ( .A1(\SB2_1_5/i0[9] ), .A2(
        \SB2_1_5/i0_0 ), .A3(\SB2_1_5/i0[8] ), .ZN(
        \SB2_1_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_2/N2  ( .A1(\SB2_1_6/i0_3 ), .A2(
        \SB2_1_6/i0[10] ), .A3(\SB2_1_6/i0[6] ), .ZN(
        \SB2_1_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_6/Component_Function_2/N1  ( .A1(\SB2_1_6/i1_5 ), .A2(
        \SB2_1_6/i0[10] ), .A3(\SB2_1_6/i1[9] ), .ZN(
        \SB2_1_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_3/N2  ( .A1(\SB2_1_6/i0_0 ), .A2(
        \SB2_1_6/i0_3 ), .A3(\SB2_1_6/i0_4 ), .ZN(
        \SB2_1_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_6/Component_Function_3/N1  ( .A1(\SB2_1_6/i1[9] ), .A2(
        \SB2_1_6/i0_3 ), .A3(\SB2_1_6/i0[6] ), .ZN(
        \SB2_1_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N4  ( .A1(\SB2_1_6/i1[9] ), .A2(
        \SB2_1_6/i1_5 ), .A3(\SB2_1_6/i0_4 ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N2  ( .A1(\SB2_1_6/i3[0] ), .A2(
        \SB2_1_6/i0_0 ), .A3(\SB2_1_6/i1_7 ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N1  ( .A1(\SB2_1_6/i0[9] ), .A2(
        \SB2_1_6/i0_0 ), .A3(\SB2_1_6/i0[8] ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_2/N2  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i0[10] ), .A3(\SB2_1_7/i0[6] ), .ZN(
        \SB2_1_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_7/Component_Function_2/N1  ( .A1(\SB2_1_7/i1_5 ), .A2(
        \SB2_1_7/i0[10] ), .A3(\SB2_1_7/i1[9] ), .ZN(
        \SB2_1_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_3/N2  ( .A1(\SB2_1_7/i0_0 ), .A2(
        \SB2_1_7/i0_3 ), .A3(\SB2_1_7/i0_4 ), .ZN(
        \SB2_1_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_7/Component_Function_3/N1  ( .A1(\SB2_1_7/i1[9] ), .A2(
        \SB2_1_7/i0_3 ), .A3(\SB2_1_7/i0[6] ), .ZN(
        \SB2_1_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_4/N4  ( .A1(\SB2_1_7/i1[9] ), .A2(
        \SB2_1_7/i1_5 ), .A3(\SB2_1_7/i0_4 ), .ZN(
        \SB2_1_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_7/Component_Function_4/N1  ( .A1(\SB2_1_7/i0[9] ), .A2(
        \SB2_1_7/i0_0 ), .A3(\SB2_1_7/i0[8] ), .ZN(
        \SB2_1_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_2/N2  ( .A1(\SB2_1_8/i0_3 ), .A2(
        \SB2_1_8/i0[10] ), .A3(\SB2_1_8/i0[6] ), .ZN(
        \SB2_1_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_8/Component_Function_2/N1  ( .A1(\SB2_1_8/i1_5 ), .A2(
        \SB2_1_8/i0[10] ), .A3(\SB2_1_8/i1[9] ), .ZN(
        \SB2_1_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_3/N3  ( .A1(\SB2_1_8/i1[9] ), .A2(
        \SB2_1_8/i1_7 ), .A3(\SB2_1_8/i0[10] ), .ZN(
        \SB2_1_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_8/Component_Function_3/N1  ( .A1(\SB2_1_8/i1[9] ), .A2(
        \SB2_1_8/i0_3 ), .A3(\SB2_1_8/i0[6] ), .ZN(
        \SB2_1_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_4/N4  ( .A1(\SB2_1_8/i1[9] ), .A2(
        \SB2_1_8/i1_5 ), .A3(\SB2_1_8/i0_4 ), .ZN(
        \SB2_1_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_9/Component_Function_2/N3  ( .A1(\SB2_1_9/i0_3 ), .A2(
        \SB2_1_9/i0[8] ), .A3(\SB2_1_9/i0[9] ), .ZN(
        \SB2_1_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_9/Component_Function_2/N2  ( .A1(\SB2_1_9/i0_3 ), .A2(
        \SB2_1_9/i0[10] ), .A3(\SB2_1_9/i0[6] ), .ZN(
        \SB2_1_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_9/Component_Function_3/N3  ( .A1(\SB2_1_9/i1[9] ), .A2(
        \SB2_1_9/i1_7 ), .A3(\SB2_1_9/i0[10] ), .ZN(
        \SB2_1_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_9/Component_Function_3/N1  ( .A1(\SB2_1_9/i1[9] ), .A2(
        \SB2_1_9/i0_3 ), .A3(\SB2_1_9/i0[6] ), .ZN(
        \SB2_1_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_9/Component_Function_4/N4  ( .A1(\SB2_1_9/i1[9] ), .A2(
        \SB2_1_9/i1_5 ), .A3(\SB2_1_9/i0_4 ), .ZN(
        \SB2_1_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_9/Component_Function_4/N2  ( .A1(\SB2_1_9/i3[0] ), .A2(
        \SB2_1_9/i0_0 ), .A3(\SB2_1_9/i1_7 ), .ZN(
        \SB2_1_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_9/Component_Function_4/N1  ( .A1(\SB2_1_9/i0[9] ), .A2(
        \SB2_1_9/i0_0 ), .A3(\SB2_1_9/i0[8] ), .ZN(
        \SB2_1_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_10/Component_Function_2/N4  ( .A1(\SB2_1_10/i1_5 ), .A2(
        \SB2_1_10/i0_0 ), .A3(\SB2_1_10/i0_4 ), .ZN(
        \SB2_1_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_10/Component_Function_2/N2  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i0[10] ), .A3(\SB2_1_10/i0[6] ), .ZN(
        \SB2_1_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_10/Component_Function_3/N1  ( .A1(\SB2_1_10/i1[9] ), .A2(
        \SB2_1_10/i0_3 ), .A3(\SB2_1_10/i0[6] ), .ZN(
        \SB2_1_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_10/Component_Function_4/N4  ( .A1(\SB2_1_10/i1[9] ), .A2(
        \SB2_1_10/i1_5 ), .A3(\SB2_1_10/i0_4 ), .ZN(
        \SB2_1_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_10/Component_Function_4/N3  ( .A1(\SB2_1_10/i0[9] ), .A2(
        \SB2_1_10/i0[10] ), .A3(\SB2_1_10/i0_3 ), .ZN(
        \SB2_1_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_10/Component_Function_4/N2  ( .A1(\SB2_1_10/i3[0] ), .A2(
        \SB2_1_10/i0_0 ), .A3(\SB2_1_10/i1_7 ), .ZN(
        \SB2_1_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_10/Component_Function_4/N1  ( .A1(\SB2_1_10/i0[9] ), .A2(
        \SB2_1_10/i0_0 ), .A3(\SB2_1_10/i0[8] ), .ZN(
        \SB2_1_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_2/N2  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i0[10] ), .A3(\SB2_1_11/i0[6] ), .ZN(
        \SB2_1_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_11/Component_Function_2/N1  ( .A1(\SB2_1_11/i1_5 ), .A2(
        \SB2_1_11/i0[10] ), .A3(\SB2_1_11/i1[9] ), .ZN(
        \SB2_1_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_3/N3  ( .A1(\SB2_1_11/i1[9] ), .A2(
        \SB2_1_11/i1_7 ), .A3(\SB2_1_11/i0[10] ), .ZN(
        \SB2_1_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_11/Component_Function_3/N1  ( .A1(\SB2_1_11/i1[9] ), .A2(
        \SB2_1_11/i0_3 ), .A3(\SB2_1_11/i0[6] ), .ZN(
        \SB2_1_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_4/N2  ( .A1(\SB2_1_11/i3[0] ), .A2(
        \SB2_1_11/i0_0 ), .A3(\SB2_1_11/i1_7 ), .ZN(
        \SB2_1_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_11/Component_Function_4/N1  ( .A1(\SB2_1_11/i0[9] ), .A2(
        \SB2_1_11/i0_0 ), .A3(\SB2_1_11/i0[8] ), .ZN(
        \SB2_1_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_2/N4  ( .A1(\SB2_1_12/i1_5 ), .A2(
        \SB2_1_12/i0_0 ), .A3(\SB2_1_12/i0_4 ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_12/Component_Function_2/N2  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i0[10] ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_12/Component_Function_2/N1  ( .A1(\SB2_1_12/i1_5 ), .A2(
        \SB2_1_12/i0[10] ), .A3(\SB2_1_12/i1[9] ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_3/N3  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i1_7 ), .A3(\SB2_1_12/i0[10] ), .ZN(
        \SB2_1_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_12/Component_Function_3/N2  ( .A1(\SB2_1_12/i0_0 ), .A2(
        \SB2_1_12/i0_3 ), .A3(\SB2_1_12/i0_4 ), .ZN(
        \SB2_1_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_12/Component_Function_3/N1  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i0_3 ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N4  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i1_5 ), .A3(\SB2_1_12/i0_4 ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N2  ( .A1(\SB2_1_12/i3[0] ), .A2(
        \SB2_1_12/i0_0 ), .A3(\SB2_1_12/i1_7 ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N1  ( .A1(\SB2_1_12/i0[9] ), .A2(
        \SB2_1_12/i0_0 ), .A3(\SB2_1_12/i0[8] ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_2/N4  ( .A1(\SB2_1_13/i1_5 ), .A2(
        \SB2_1_13/i0_0 ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_13/Component_Function_2/N2  ( .A1(\SB2_1_13/i0_3 ), .A2(
        \SB2_1_13/i0[10] ), .A3(\SB2_1_13/i0[6] ), .ZN(
        \SB2_1_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_13/Component_Function_2/N1  ( .A1(\SB2_1_13/i1_5 ), .A2(
        \SB2_1_13/i0[10] ), .A3(\SB2_1_13/i1[9] ), .ZN(
        \SB2_1_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_3/N1  ( .A1(\SB2_1_13/i1[9] ), .A2(
        \SB2_1_13/i0_3 ), .A3(\SB2_1_13/i0[6] ), .ZN(
        \SB2_1_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N4  ( .A1(\SB2_1_13/i1[9] ), .A2(
        \SB2_1_13/i1_5 ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N3  ( .A1(\SB2_1_13/i0[9] ), .A2(
        \SB2_1_13/i0[10] ), .A3(\SB2_1_13/i0_3 ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N2  ( .A1(\SB2_1_13/i3[0] ), .A2(
        \SB2_1_13/i0_0 ), .A3(\SB2_1_13/i1_7 ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N1  ( .A1(\SB2_1_13/i0[9] ), .A2(
        \SB2_1_13/i0_0 ), .A3(\SB2_1_13/i0[8] ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_2/N2  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i0[10] ), .A3(\SB2_1_14/i0[6] ), .ZN(
        \SB2_1_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_14/Component_Function_3/N4  ( .A1(\SB2_1_14/i1_5 ), .A2(
        \SB2_1_14/i0[8] ), .A3(\SB2_1_14/i3[0] ), .ZN(
        \SB2_1_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_14/Component_Function_3/N3  ( .A1(\SB2_1_14/i1[9] ), .A2(
        \SB2_1_14/i1_7 ), .A3(\SB2_1_14/i0[10] ), .ZN(
        \SB2_1_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_14/Component_Function_3/N2  ( .A1(\SB2_1_14/i0_0 ), .A2(
        \SB2_1_14/i0_3 ), .A3(\SB2_1_14/i0_4 ), .ZN(
        \SB2_1_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_14/Component_Function_3/N1  ( .A1(\SB2_1_14/i1[9] ), .A2(
        \SB2_1_14/i0_3 ), .A3(\SB2_1_14/i0[6] ), .ZN(
        \SB2_1_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_4/N3  ( .A1(\SB2_1_14/i0[9] ), .A2(
        \SB2_1_14/i0[10] ), .A3(\SB2_1_14/i0_3 ), .ZN(
        \SB2_1_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_14/Component_Function_4/N2  ( .A1(\SB2_1_14/i3[0] ), .A2(
        \SB2_1_14/i0_0 ), .A3(\SB2_1_14/i1_7 ), .ZN(
        \SB2_1_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_14/Component_Function_4/N1  ( .A1(\SB2_1_14/i0[9] ), .A2(
        \SB2_1_14/i0_0 ), .A3(\SB2_1_14/i0[8] ), .ZN(
        \SB2_1_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_15/Component_Function_2/N4  ( .A1(\SB2_1_15/i1_5 ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i0_4 ), .ZN(
        \SB2_1_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_15/Component_Function_2/N2  ( .A1(\SB2_1_15/i0_3 ), .A2(
        \SB2_1_15/i0[10] ), .A3(\SB2_1_15/i0[6] ), .ZN(
        \SB2_1_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_15/Component_Function_3/N3  ( .A1(\SB2_1_15/i1[9] ), .A2(
        \SB2_1_15/i1_7 ), .A3(\SB2_1_15/i0[10] ), .ZN(
        \SB2_1_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_15/Component_Function_3/N1  ( .A1(\SB2_1_15/i1[9] ), .A2(
        \SB2_1_15/i0_3 ), .A3(\SB2_1_15/i0[6] ), .ZN(
        \SB2_1_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_15/Component_Function_4/N3  ( .A1(\SB2_1_15/i0[9] ), .A2(
        \SB2_1_15/i0[10] ), .A3(\SB2_1_15/i0_3 ), .ZN(
        \SB2_1_15/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_15/Component_Function_4/N2  ( .A1(\SB2_1_15/i3[0] ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i1_7 ), .ZN(
        \SB2_1_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_15/Component_Function_4/N1  ( .A1(\SB2_1_15/i0[9] ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i0[8] ), .ZN(
        \SB2_1_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_16/Component_Function_2/N4  ( .A1(\SB2_1_16/i1_5 ), .A2(
        \SB2_1_16/i0_0 ), .A3(\SB2_1_16/i0_4 ), .ZN(
        \SB2_1_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_16/Component_Function_2/N2  ( .A1(\SB2_1_16/i0_3 ), .A2(
        \SB2_1_16/i0[10] ), .A3(\SB2_1_16/i0[6] ), .ZN(
        \SB2_1_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_16/Component_Function_3/N2  ( .A1(\SB2_1_16/i0_0 ), .A2(
        \SB2_1_16/i0_3 ), .A3(\SB2_1_16/i0_4 ), .ZN(
        \SB2_1_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N4  ( .A1(\SB2_1_16/i1[9] ), .A2(
        \SB2_1_16/i1_5 ), .A3(\SB2_1_16/i0_4 ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N3  ( .A1(\SB2_1_16/i0[9] ), .A2(
        \SB2_1_16/i0[10] ), .A3(\SB2_1_16/i0_3 ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N2  ( .A1(\SB2_1_16/i3[0] ), .A2(
        \SB2_1_16/i0_0 ), .A3(\SB2_1_16/i1_7 ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N1  ( .A1(\SB2_1_16/i0[9] ), .A2(
        \SB2_1_16/i0_0 ), .A3(\SB2_1_16/i0[8] ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_2/N2  ( .A1(\SB2_1_17/i0_3 ), .A2(
        \SB2_1_17/i0[10] ), .A3(\SB2_1_17/i0[6] ), .ZN(
        \SB2_1_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_17/Component_Function_2/N1  ( .A1(\SB2_1_17/i1_5 ), .A2(
        \SB2_1_17/i0[10] ), .A3(\SB2_1_17/i1[9] ), .ZN(
        \SB2_1_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_3/N1  ( .A1(\SB2_1_17/i1[9] ), .A2(
        \SB2_1_17/i0_3 ), .A3(\SB2_1_17/i0[6] ), .ZN(
        \SB2_1_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N4  ( .A1(\SB2_1_17/i1[9] ), .A2(
        \SB2_1_17/i1_5 ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N3  ( .A1(\SB2_1_17/i0[9] ), .A2(
        \SB2_1_17/i0[10] ), .A3(\SB2_1_17/i0_3 ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N2  ( .A1(\SB2_1_17/i3[0] ), .A2(
        \SB2_1_17/i0_0 ), .A3(\SB2_1_17/i1_7 ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N1  ( .A1(\SB2_1_17/i0[9] ), .A2(
        \SB2_1_17/i0_0 ), .A3(\SB2_1_17/i0[8] ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_2/N2  ( .A1(\SB2_1_18/i0_3 ), .A2(
        \SB2_1_18/i0[10] ), .A3(\SB2_1_18/i0[6] ), .ZN(
        \SB2_1_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_18/Component_Function_2/N1  ( .A1(\SB2_1_18/i1_5 ), .A2(
        \SB2_1_18/i0[10] ), .A3(\SB2_1_18/i1[9] ), .ZN(
        \SB2_1_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_3/N4  ( .A1(\SB2_1_18/i1_5 ), .A2(
        \SB2_1_18/i0[8] ), .A3(\SB2_1_18/i3[0] ), .ZN(
        \SB2_1_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_18/Component_Function_3/N1  ( .A1(\SB2_1_18/i1[9] ), .A2(
        \SB2_1_18/i0_3 ), .A3(\SB2_1_18/i0[6] ), .ZN(
        \SB2_1_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_4/N4  ( .A1(\SB2_1_18/i1[9] ), .A2(
        \SB2_1_18/i1_5 ), .A3(\SB2_1_18/i0_4 ), .ZN(
        \SB2_1_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_18/Component_Function_4/N3  ( .A1(\SB2_1_18/i0[9] ), .A2(
        \SB2_1_18/i0[10] ), .A3(\SB2_1_18/i0_3 ), .ZN(
        \SB2_1_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_18/Component_Function_4/N2  ( .A1(\SB2_1_18/i3[0] ), .A2(
        \SB2_1_18/i0_0 ), .A3(\SB2_1_18/i1_7 ), .ZN(
        \SB2_1_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_18/Component_Function_4/N1  ( .A1(\SB2_1_18/i0[9] ), .A2(
        \SB2_1_18/i0_0 ), .A3(\SB2_1_18/i0[8] ), .ZN(
        \SB2_1_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_19/Component_Function_2/N3  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i0[8] ), .A3(\SB2_1_19/i0[9] ), .ZN(
        \SB2_1_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_19/Component_Function_2/N2  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i0[10] ), .A3(\SB2_1_19/i0[6] ), .ZN(
        \SB2_1_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_19/Component_Function_3/N3  ( .A1(\SB2_1_19/i1[9] ), .A2(
        \SB2_1_19/i1_7 ), .A3(\SB2_1_19/i0[10] ), .ZN(
        \SB2_1_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_19/Component_Function_3/N2  ( .A1(\SB2_1_19/i0_0 ), .A2(
        \SB2_1_19/i0_3 ), .A3(\SB2_1_19/i0_4 ), .ZN(
        \SB2_1_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_19/Component_Function_4/N4  ( .A1(\SB2_1_19/i1[9] ), .A2(
        \SB2_1_19/i1_5 ), .A3(\SB2_1_19/i0_4 ), .ZN(
        \SB2_1_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_19/Component_Function_4/N1  ( .A1(\SB2_1_19/i0[9] ), .A2(
        \SB2_1_19/i0_0 ), .A3(\SB2_1_19/i0[8] ), .ZN(
        \SB2_1_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_20/Component_Function_2/N3  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i0[8] ), .A3(\SB2_1_20/i0[9] ), .ZN(
        \SB2_1_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_20/Component_Function_2/N2  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i0[10] ), .A3(\SB2_1_20/i0[6] ), .ZN(
        \SB2_1_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_20/Component_Function_3/N3  ( .A1(\SB2_1_20/i1[9] ), .A2(
        \SB2_1_20/i1_7 ), .A3(\SB2_1_20/i0[10] ), .ZN(
        \SB2_1_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_20/Component_Function_3/N2  ( .A1(\SB2_1_20/i0_0 ), .A2(
        \SB2_1_20/i0_3 ), .A3(\SB2_1_20/i0_4 ), .ZN(
        \SB2_1_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_20/Component_Function_4/N3  ( .A1(\SB2_1_20/i0[9] ), .A2(
        \SB2_1_20/i0[10] ), .A3(\SB2_1_20/i0_3 ), .ZN(
        \SB2_1_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_20/Component_Function_4/N2  ( .A1(\SB2_1_20/i3[0] ), .A2(
        \SB2_1_20/i0_0 ), .A3(\SB2_1_20/i1_7 ), .ZN(
        \SB2_1_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_20/Component_Function_4/N1  ( .A1(\SB2_1_20/i0[9] ), .A2(
        \SB2_1_20/i0_0 ), .A3(\SB2_1_20/i0[8] ), .ZN(
        \SB2_1_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_21/Component_Function_2/N4  ( .A1(\SB2_1_21/i1_5 ), .A2(
        \SB2_1_21/i0_0 ), .A3(\SB2_1_21/i0_4 ), .ZN(
        \SB2_1_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_21/Component_Function_2/N2  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i0[10] ), .A3(\SB2_1_21/i0[6] ), .ZN(
        \SB2_1_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_21/Component_Function_2/N1  ( .A1(\SB2_1_21/i1_5 ), .A2(
        \SB2_1_21/i0[10] ), .A3(\SB2_1_21/i1[9] ), .ZN(
        \SB2_1_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_21/Component_Function_3/N1  ( .A1(\SB2_1_21/i1[9] ), .A2(
        \SB2_1_21/i0_3 ), .A3(\SB2_1_21/i0[6] ), .ZN(
        \SB2_1_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_21/Component_Function_4/N4  ( .A1(\SB2_1_21/i1[9] ), .A2(
        \SB2_1_21/i1_5 ), .A3(\SB2_1_21/i0_4 ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_21/Component_Function_4/N2  ( .A1(\SB2_1_21/i3[0] ), .A2(
        \SB2_1_21/i0_0 ), .A3(\SB2_1_21/i1_7 ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_21/Component_Function_4/N1  ( .A1(\SB2_1_21/i0[9] ), .A2(
        \SB2_1_21/i0_0 ), .A3(\SB2_1_21/i0[8] ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_2/N3  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i0[8] ), .A3(\SB2_1_22/i0[9] ), .ZN(
        \SB2_1_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_22/Component_Function_2/N2  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i0[10] ), .A3(\SB2_1_22/i0[6] ), .ZN(
        \SB2_1_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_22/Component_Function_2/N1  ( .A1(\SB2_1_22/i1_5 ), .A2(
        \SB2_1_22/i0[10] ), .A3(\SB2_1_22/i1[9] ), .ZN(
        \SB2_1_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_3/N3  ( .A1(\SB2_1_22/i1[9] ), .A2(
        \SB2_1_22/i1_7 ), .A3(\SB2_1_22/i0[10] ), .ZN(
        \SB2_1_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_22/Component_Function_3/N1  ( .A1(\SB2_1_22/i1[9] ), .A2(
        \SB2_1_22/i0_3 ), .A3(\SB2_1_22/i0[6] ), .ZN(
        \SB2_1_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_4/N4  ( .A1(\SB2_1_22/i1[9] ), .A2(
        \SB2_1_22/i1_5 ), .A3(\SB2_1_22/i0_4 ), .ZN(
        \SB2_1_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_22/Component_Function_4/N2  ( .A1(\SB2_1_22/i3[0] ), .A2(
        \SB2_1_22/i0_0 ), .A3(\SB2_1_22/i1_7 ), .ZN(
        \SB2_1_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_22/Component_Function_4/N1  ( .A1(\SB2_1_22/i0[9] ), .A2(
        \SB2_1_22/i0_0 ), .A3(\SB2_1_22/i0[8] ), .ZN(
        \SB2_1_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_2/N4  ( .A1(\SB2_1_23/i1_5 ), .A2(
        \SB2_1_23/i0_0 ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_23/Component_Function_2/N2  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i0[10] ), .A3(\SB2_1_23/i0[6] ), .ZN(
        \SB2_1_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_23/Component_Function_2/N1  ( .A1(\SB2_1_23/i1_5 ), .A2(
        \SB2_1_23/i0[10] ), .A3(\SB2_1_23/i1[9] ), .ZN(
        \SB2_1_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_3/N3  ( .A1(\SB2_1_23/i1[9] ), .A2(
        \SB2_1_23/i1_7 ), .A3(\SB2_1_23/i0[10] ), .ZN(
        \SB2_1_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_23/Component_Function_3/N2  ( .A1(\SB2_1_23/i0_0 ), .A2(
        \SB2_1_23/i0_3 ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_23/Component_Function_3/N1  ( .A1(\SB2_1_23/i1[9] ), .A2(
        \SB2_1_23/i0_3 ), .A3(\SB2_1_23/i0[6] ), .ZN(
        \SB2_1_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N4  ( .A1(\SB2_1_23/i1[9] ), .A2(
        \SB2_1_23/i1_5 ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N3  ( .A1(\SB2_1_23/i0[9] ), .A2(
        \SB2_1_23/i0[10] ), .A3(\SB2_1_23/i0_3 ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N2  ( .A1(\SB2_1_23/i3[0] ), .A2(
        \SB2_1_23/i0_0 ), .A3(\SB2_1_23/i1_7 ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N1  ( .A1(\SB2_1_23/i0[9] ), .A2(
        \SB2_1_23/i0_0 ), .A3(\SB2_1_23/i0[8] ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_2/N3  ( .A1(\SB2_1_24/i0_3 ), .A2(
        \SB2_1_24/i0[8] ), .A3(\SB2_1_24/i0[9] ), .ZN(
        \SB2_1_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_24/Component_Function_2/N2  ( .A1(\SB2_1_24/i0_3 ), .A2(
        \SB2_1_24/i0[10] ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_24/Component_Function_3/N1  ( .A1(\SB2_1_24/i1[9] ), .A2(
        \SB2_1_24/i0_3 ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_4/N4  ( .A1(\SB2_1_24/i1[9] ), .A2(
        \SB2_1_24/i1_5 ), .A3(\SB2_1_24/i0_4 ), .ZN(
        \SB2_1_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_24/Component_Function_4/N2  ( .A1(\SB2_1_24/i3[0] ), .A2(
        \SB2_1_24/i0_0 ), .A3(\SB2_1_24/i1_7 ), .ZN(
        \SB2_1_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_24/Component_Function_4/N1  ( .A1(\SB2_1_24/i0[9] ), .A2(
        \SB2_1_24/i0_0 ), .A3(\SB2_1_24/i0[8] ), .ZN(
        \SB2_1_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_2/N4  ( .A1(\SB2_1_25/i1_5 ), .A2(
        \SB2_1_25/i0_0 ), .A3(\SB2_1_25/i0_4 ), .ZN(
        \SB2_1_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_25/Component_Function_2/N3  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i0[8] ), .A3(\SB2_1_25/i0[9] ), .ZN(
        \SB2_1_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_25/Component_Function_2/N2  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i0[10] ), .A3(\SB2_1_25/i0[6] ), .ZN(
        \SB2_1_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_25/Component_Function_2/N1  ( .A1(\SB2_1_25/i1_5 ), .A2(
        \SB2_1_25/i0[10] ), .A3(\SB2_1_25/i1[9] ), .ZN(
        \SB2_1_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_3/N3  ( .A1(\SB2_1_25/i1[9] ), .A2(
        \SB2_1_25/i1_7 ), .A3(\SB2_1_25/i0[10] ), .ZN(
        \SB2_1_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_25/Component_Function_3/N1  ( .A1(\SB2_1_25/i1[9] ), .A2(
        \SB2_1_25/i0_3 ), .A3(\SB2_1_25/i0[6] ), .ZN(
        \SB2_1_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N4  ( .A1(\SB2_1_25/i1[9] ), .A2(
        \SB2_1_25/i1_5 ), .A3(\SB2_1_25/i0_4 ), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N2  ( .A1(\SB2_1_25/i3[0] ), .A2(
        \SB2_1_25/i0_0 ), .A3(\SB2_1_25/i1_7 ), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N1  ( .A1(\SB2_1_25/i0[9] ), .A2(
        \SB2_1_25/i0_0 ), .A3(\SB2_1_25/i0[8] ), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_2/N4  ( .A1(\SB2_1_26/i1_5 ), .A2(
        \SB2_1_26/i0_0 ), .A3(\SB2_1_26/i0_4 ), .ZN(
        \SB2_1_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_26/Component_Function_2/N3  ( .A1(\SB2_1_26/i0_3 ), .A2(
        \SB2_1_26/i0[8] ), .A3(\SB2_1_26/i0[9] ), .ZN(
        \SB2_1_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_26/Component_Function_3/N3  ( .A1(\SB2_1_26/i1[9] ), .A2(
        \SB2_1_26/i1_7 ), .A3(\SB2_1_26/i0[10] ), .ZN(
        \SB2_1_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_26/Component_Function_3/N2  ( .A1(\SB2_1_26/i0_0 ), .A2(
        \SB2_1_26/i0_3 ), .A3(\SB2_1_26/i0_4 ), .ZN(
        \SB2_1_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N4  ( .A1(\SB2_1_26/i1[9] ), .A2(
        \SB2_1_26/i1_5 ), .A3(\SB2_1_26/i0_4 ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N3  ( .A1(\SB2_1_26/i0[9] ), .A2(
        \SB2_1_26/i0[10] ), .A3(\SB2_1_26/i0_3 ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N2  ( .A1(\SB2_1_26/i3[0] ), .A2(
        \SB2_1_26/i0_0 ), .A3(\SB2_1_26/i1_7 ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N1  ( .A1(\SB2_1_26/i0[9] ), .A2(
        \SB2_1_26/i0_0 ), .A3(\SB2_1_26/i0[8] ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_2/N4  ( .A1(\SB2_1_27/i1_5 ), .A2(
        \SB2_1_27/i0_0 ), .A3(\SB2_1_27/i0_4 ), .ZN(
        \SB2_1_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_27/Component_Function_2/N2  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i0[10] ), .A3(\SB2_1_27/i0[6] ), .ZN(
        \SB2_1_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_27/Component_Function_2/N1  ( .A1(\SB2_1_27/i1_5 ), .A2(
        \SB2_1_27/i0[10] ), .A3(\SB2_1_27/i1[9] ), .ZN(
        \SB2_1_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_3/N3  ( .A1(\SB2_1_27/i1[9] ), .A2(
        \SB2_1_27/i1_7 ), .A3(\SB2_1_27/i0[10] ), .ZN(
        \SB2_1_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_27/Component_Function_3/N1  ( .A1(\SB2_1_27/i1[9] ), .A2(
        \SB2_1_27/i0_3 ), .A3(\SB2_1_27/i0[6] ), .ZN(
        \SB2_1_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_4/N4  ( .A1(\SB2_1_27/i1[9] ), .A2(
        \SB2_1_27/i1_5 ), .A3(\SB2_1_27/i0_4 ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_27/Component_Function_4/N2  ( .A1(\SB2_1_27/i3[0] ), .A2(
        \SB2_1_27/i0_0 ), .A3(\SB2_1_27/i1_7 ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_27/Component_Function_4/N1  ( .A1(\SB2_1_27/i0[9] ), .A2(
        \SB2_1_27/i0_0 ), .A3(\SB2_1_27/i0[8] ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_2/N4  ( .A1(\SB2_1_28/i1_5 ), .A2(
        \SB2_1_28/i0_0 ), .A3(\SB2_1_28/i0_4 ), .ZN(
        \SB2_1_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_28/Component_Function_2/N2  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i0[10] ), .A3(\SB2_1_28/i0[6] ), .ZN(
        \SB2_1_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_2/N1  ( .A1(\SB2_1_28/i1_5 ), .A2(
        \SB2_1_28/i0[10] ), .A3(\SB2_1_28/i1[9] ), .ZN(
        \SB2_1_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_3/N3  ( .A1(\SB2_1_28/i1[9] ), .A2(
        \SB2_1_28/i1_7 ), .A3(\SB2_1_28/i0[10] ), .ZN(
        \SB2_1_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_28/Component_Function_3/N2  ( .A1(\SB2_1_28/i0_0 ), .A2(
        \SB2_1_28/i0_3 ), .A3(\SB2_1_28/i0_4 ), .ZN(
        \SB2_1_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_3/N1  ( .A1(\SB2_1_28/i1[9] ), .A2(
        \SB2_1_28/i0_3 ), .A3(\SB2_1_28/i0[6] ), .ZN(
        \SB2_1_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N4  ( .A1(\SB2_1_28/i1[9] ), .A2(
        \SB2_1_28/i1_5 ), .A3(\SB2_1_28/i0_4 ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N2  ( .A1(\SB2_1_28/i3[0] ), .A2(
        \SB2_1_28/i0_0 ), .A3(\SB2_1_28/i1_7 ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N1  ( .A1(\SB2_1_28/i0[9] ), .A2(
        \SB2_1_28/i0_0 ), .A3(\SB2_1_28/i0[8] ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_2/N2  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i0[10] ), .A3(\SB2_1_29/i0[6] ), .ZN(
        \SB2_1_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_29/Component_Function_3/N3  ( .A1(\SB2_1_29/i1[9] ), .A2(
        \SB2_1_29/i1_7 ), .A3(\SB2_1_29/i0[10] ), .ZN(
        \SB2_1_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_29/Component_Function_3/N1  ( .A1(\SB2_1_29/i1[9] ), .A2(
        \SB2_1_29/i0_3 ), .A3(\SB2_1_29/i0[6] ), .ZN(
        \SB2_1_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N3  ( .A1(\SB2_1_29/i0[9] ), .A2(
        \SB2_1_29/i0[10] ), .A3(\SB2_1_29/i0_3 ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N2  ( .A1(\SB2_1_29/i3[0] ), .A2(
        \SB2_1_29/i0_0 ), .A3(\SB2_1_29/i1_7 ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N1  ( .A1(\SB2_1_29/i0[9] ), .A2(
        \SB2_1_29/i0_0 ), .A3(\SB2_1_29/i0[8] ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_2/N1  ( .A1(\SB2_1_30/i1_5 ), .A2(
        \SB2_1_30/i0[10] ), .A3(\SB2_1_30/i1[9] ), .ZN(
        \SB2_1_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_3/N3  ( .A1(\SB2_1_30/i1[9] ), .A2(
        \SB2_1_30/i1_7 ), .A3(\SB2_1_30/i0[10] ), .ZN(
        \SB2_1_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_30/Component_Function_3/N1  ( .A1(\SB2_1_30/i1[9] ), .A2(
        \SB2_1_30/i0_3 ), .A3(\SB2_1_30/i0[6] ), .ZN(
        \SB2_1_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N4  ( .A1(\SB2_1_30/i1[9] ), .A2(
        \SB2_1_30/i1_5 ), .A3(\SB2_1_30/i0_4 ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N2  ( .A1(\SB2_1_30/i3[0] ), .A2(
        \SB2_1_30/i0_0 ), .A3(\SB2_1_30/i1_7 ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N1  ( .A1(\SB2_1_30/i0[9] ), .A2(
        \SB2_1_30/i0_0 ), .A3(\SB2_1_30/i0[8] ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_2/N1  ( .A1(\SB2_1_31/i1_5 ), .A2(
        \SB2_1_31/i0[10] ), .A3(\SB2_1_31/i1[9] ), .ZN(
        \SB2_1_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_3/N3  ( .A1(\SB2_1_31/i1[9] ), .A2(
        \SB2_1_31/i1_7 ), .A3(\SB2_1_31/i0[10] ), .ZN(
        \SB2_1_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_31/Component_Function_3/N1  ( .A1(\SB2_1_31/i1[9] ), .A2(
        \SB2_1_31/i0_3 ), .A3(\SB2_1_31/i0[6] ), .ZN(
        \SB2_1_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_4/N4  ( .A1(\SB2_1_31/i1[9] ), .A2(
        \SB2_1_31/i1_5 ), .A3(\SB2_1_31/i0_4 ), .ZN(
        \SB2_1_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_31/Component_Function_4/N2  ( .A1(\SB2_1_31/i3[0] ), .A2(
        \SB2_1_31/i0_0 ), .A3(\SB2_1_31/i1_7 ), .ZN(
        \SB2_1_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_31/Component_Function_4/N1  ( .A1(\SB2_1_31/i0[9] ), .A2(
        \SB2_1_31/i0_0 ), .A3(\SB2_1_31/i0[8] ), .ZN(
        \SB2_1_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_2/N2  ( .A1(\SB1_2_0/i0_3 ), .A2(
        \SB1_2_0/i0[10] ), .A3(\SB1_2_0/i0[6] ), .ZN(
        \SB1_2_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_2/N1  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[10] ), .A3(\SB1_2_0/i1[9] ), .ZN(
        \SB1_2_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_3/N4  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[8] ), .A3(\SB1_2_0/i3[0] ), .ZN(
        \SB1_2_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_0/Component_Function_3/N1  ( .A1(\SB1_2_0/i1[9] ), .A2(
        \SB1_2_0/i0_3 ), .A3(\SB1_2_0/i0[6] ), .ZN(
        \SB1_2_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_4/N2  ( .A1(\SB1_2_0/i3[0] ), .A2(
        \SB1_2_0/i0_0 ), .A3(\SB1_2_0/i1_7 ), .ZN(
        \SB1_2_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_4/N1  ( .A1(\SB1_2_0/i0[9] ), .A2(
        \SB1_2_0/i0_0 ), .A3(\SB1_2_0/i0[8] ), .ZN(
        \SB1_2_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_2/N2  ( .A1(\SB1_2_1/i0_3 ), .A2(
        \SB1_2_1/i0[10] ), .A3(\SB1_2_1/i0[6] ), .ZN(
        \SB1_2_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_1/Component_Function_2/N1  ( .A1(\SB1_2_1/i1_5 ), .A2(
        \SB1_2_1/i0[10] ), .A3(\SB1_2_1/i1[9] ), .ZN(
        \SB1_2_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_4/N4  ( .A1(\SB1_2_1/i1[9] ), .A2(
        \SB1_2_1/i1_5 ), .A3(\SB1_2_1/i0_4 ), .ZN(
        \SB1_2_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_1/Component_Function_4/N2  ( .A1(\SB1_2_1/i3[0] ), .A2(
        \SB1_2_1/i0_0 ), .A3(\SB1_2_1/i1_7 ), .ZN(
        \SB1_2_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_1/Component_Function_4/N1  ( .A1(\SB1_2_1/i0[9] ), .A2(
        \SB1_2_1/i0_0 ), .A3(\SB1_2_1/i0[8] ), .ZN(
        \SB1_2_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_2/N2  ( .A1(\SB1_2_2/i0_3 ), .A2(
        \SB1_2_2/i0[10] ), .A3(\SB1_2_2/i0[6] ), .ZN(
        \SB1_2_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_2/Component_Function_2/N1  ( .A1(\SB1_2_2/i1_5 ), .A2(
        \SB1_2_2/i0[10] ), .A3(\SB1_2_2/i1[9] ), .ZN(
        \SB1_2_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_3/N4  ( .A1(\SB1_2_2/i1_5 ), .A2(
        \SB1_2_2/i0[8] ), .A3(\SB1_2_2/i3[0] ), .ZN(
        \SB1_2_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_3/N3  ( .A1(\SB1_2_2/i1[9] ), .A2(
        \SB1_2_2/i1_7 ), .A3(\SB1_2_2/i0[10] ), .ZN(
        \SB1_2_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_2/Component_Function_3/N1  ( .A1(\SB1_2_2/i1[9] ), .A2(n1648), .A3(\SB1_2_2/i0[6] ), .ZN(\SB1_2_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_4/N4  ( .A1(\SB1_2_2/i1[9] ), .A2(
        \SB1_2_2/i1_5 ), .A3(\SB1_2_2/i0_4 ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_4/N2  ( .A1(\SB1_2_2/i3[0] ), .A2(
        \SB1_2_2/i0_0 ), .A3(\SB1_2_2/i1_7 ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_2/Component_Function_4/N1  ( .A1(\SB1_2_2/i0[9] ), .A2(
        \SB1_2_2/i0_0 ), .A3(\SB1_2_2/i0[8] ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_2/N2  ( .A1(\SB1_2_3/i0_3 ), .A2(
        \SB1_2_3/i0[10] ), .A3(\SB1_2_3/i0[6] ), .ZN(
        \SB1_2_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_3/Component_Function_2/N1  ( .A1(\SB1_2_3/i1_5 ), .A2(
        \SB1_2_3/i0[10] ), .A3(\SB1_2_3/i1[9] ), .ZN(
        \SB1_2_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_3/N4  ( .A1(\SB1_2_3/i1_5 ), .A2(
        \SB1_2_3/i0[8] ), .A3(\SB1_2_3/i3[0] ), .ZN(
        \SB1_2_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_3/Component_Function_3/N1  ( .A1(\SB1_2_3/i1[9] ), .A2(
        \SB1_2_3/i0_3 ), .A3(\SB1_2_3/i0[6] ), .ZN(
        \SB1_2_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_4/N4  ( .A1(\SB1_2_3/i1[9] ), .A2(
        \SB1_2_3/i1_5 ), .A3(\SB1_2_3/i0_4 ), .ZN(
        \SB1_2_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_3/Component_Function_4/N2  ( .A1(\SB1_2_3/i3[0] ), .A2(
        \SB1_2_3/i0_0 ), .A3(\SB1_2_3/i1_7 ), .ZN(
        \SB1_2_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_3/Component_Function_4/N1  ( .A1(\SB1_2_3/i0[9] ), .A2(
        \SB1_2_3/i0_0 ), .A3(\SB1_2_3/i0[8] ), .ZN(
        \SB1_2_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_2/N3  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i0[8] ), .A3(\SB1_2_4/i0[9] ), .ZN(
        \SB1_2_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_4/Component_Function_2/N2  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i0[10] ), .A3(\SB1_2_4/i0[6] ), .ZN(
        \SB1_2_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_4/Component_Function_2/N1  ( .A1(\SB1_2_4/i1_5 ), .A2(
        \SB1_2_4/i0[10] ), .A3(\SB1_2_4/i1[9] ), .ZN(
        \SB1_2_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_3/N4  ( .A1(\SB1_2_4/i1_5 ), .A2(
        \SB1_2_4/i0[8] ), .A3(\SB1_2_4/i3[0] ), .ZN(
        \SB1_2_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_4/Component_Function_3/N3  ( .A1(\SB1_2_4/i1[9] ), .A2(
        \SB1_2_4/i1_7 ), .A3(\SB1_2_4/i0[10] ), .ZN(
        \SB1_2_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_4/Component_Function_3/N1  ( .A1(\SB1_2_4/i1[9] ), .A2(
        \SB1_2_4/i0_3 ), .A3(\SB1_2_4/i0[6] ), .ZN(
        \SB1_2_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_4/N4  ( .A1(\SB1_2_4/i1[9] ), .A2(
        \SB1_2_4/i1_5 ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_4/Component_Function_4/N2  ( .A1(\SB1_2_4/i3[0] ), .A2(
        \SB1_2_4/i0_0 ), .A3(\SB1_2_4/i1_7 ), .ZN(
        \SB1_2_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_4/Component_Function_4/N1  ( .A1(\SB1_2_4/i0[9] ), .A2(
        \SB1_2_4/i0_0 ), .A3(\SB1_2_4/i0[8] ), .ZN(
        \SB1_2_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_2/N2  ( .A1(\SB1_2_5/i0_3 ), .A2(
        \SB1_2_5/i0[10] ), .A3(\SB1_2_5/i0[6] ), .ZN(
        \SB1_2_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_5/Component_Function_2/N1  ( .A1(\SB1_2_5/i1_5 ), .A2(
        \SB1_2_5/i0[10] ), .A3(\SB1_2_5/i1[9] ), .ZN(
        \SB1_2_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_3/N4  ( .A1(\SB1_2_5/i1_5 ), .A2(
        \SB1_2_5/i0[8] ), .A3(\SB1_2_5/i3[0] ), .ZN(
        \SB1_2_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_5/Component_Function_3/N3  ( .A1(\SB1_2_5/i1[9] ), .A2(
        \SB1_2_5/i1_7 ), .A3(\SB1_2_5/i0[10] ), .ZN(
        \SB1_2_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_5/Component_Function_3/N1  ( .A1(\SB1_2_5/i1[9] ), .A2(
        \SB1_2_5/i0_3 ), .A3(\SB1_2_5/i0[6] ), .ZN(
        \SB1_2_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_4/N4  ( .A1(\SB1_2_5/i1[9] ), .A2(
        \SB1_2_5/i1_5 ), .A3(\SB1_2_5/i0_4 ), .ZN(
        \SB1_2_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_5/Component_Function_4/N2  ( .A1(\SB1_2_5/i3[0] ), .A2(
        \SB1_2_5/i0_0 ), .A3(\SB1_2_5/i1_7 ), .ZN(
        \SB1_2_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_5/Component_Function_4/N1  ( .A1(\SB1_2_5/i0[9] ), .A2(
        \SB1_2_5/i0_0 ), .A3(\SB1_2_5/i0[8] ), .ZN(
        \SB1_2_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_2/N2  ( .A1(\SB1_2_6/i0_3 ), .A2(
        \SB1_2_6/i0[10] ), .A3(\SB1_2_6/i0[6] ), .ZN(
        \SB1_2_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_6/Component_Function_2/N1  ( .A1(\SB1_2_6/i1_5 ), .A2(
        \SB1_2_6/i0[10] ), .A3(\SB1_2_6/i1[9] ), .ZN(
        \SB1_2_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_3/N4  ( .A1(\SB1_2_6/i1_5 ), .A2(
        \SB1_2_6/i0[8] ), .A3(\SB1_2_6/i3[0] ), .ZN(
        \SB1_2_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_6/Component_Function_3/N3  ( .A1(\SB1_2_6/i1[9] ), .A2(
        \RI1[2][151] ), .A3(\SB1_2_6/i0[10] ), .ZN(
        \SB1_2_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_6/Component_Function_3/N1  ( .A1(\SB1_2_6/i1[9] ), .A2(
        \SB1_2_6/i0_3 ), .A3(\SB1_2_6/i0[6] ), .ZN(
        \SB1_2_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_4/N4  ( .A1(\SB1_2_6/i1[9] ), .A2(
        \SB1_2_6/i1_5 ), .A3(\SB1_2_6/i0_4 ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_6/Component_Function_4/N2  ( .A1(\SB1_2_6/i3[0] ), .A2(
        \SB1_2_6/i0_0 ), .A3(\SB1_2_6/i1_7 ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_6/Component_Function_4/N1  ( .A1(\SB1_2_6/i0[9] ), .A2(
        \SB1_2_6/i0_0 ), .A3(\SB1_2_6/i0[8] ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_2/N2  ( .A1(\SB1_2_7/i0_3 ), .A2(
        \SB1_2_7/i0[10] ), .A3(\SB1_2_7/i0[6] ), .ZN(
        \SB1_2_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_7/Component_Function_2/N1  ( .A1(\SB1_2_7/i1_5 ), .A2(
        \SB1_2_7/i0[10] ), .A3(\SB1_2_7/i1[9] ), .ZN(
        \SB1_2_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_3/N4  ( .A1(\SB1_2_7/i1_5 ), .A2(
        \SB1_2_7/i0[8] ), .A3(\SB1_2_7/i3[0] ), .ZN(
        \SB1_2_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_7/Component_Function_3/N3  ( .A1(\SB1_2_7/i1[9] ), .A2(
        \SB1_2_7/i1_7 ), .A3(\SB1_2_7/i0[10] ), .ZN(
        \SB1_2_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_7/Component_Function_3/N1  ( .A1(\SB1_2_7/i1[9] ), .A2(
        \SB1_2_7/i0_3 ), .A3(\SB1_2_7/i0[6] ), .ZN(
        \SB1_2_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N4  ( .A1(\SB1_2_7/i1[9] ), .A2(
        \SB1_2_7/i1_5 ), .A3(\SB1_2_7/i0_4 ), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N2  ( .A1(\SB1_2_7/i3[0] ), .A2(
        \SB1_2_7/i0_0 ), .A3(\SB1_2_7/i1_7 ), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N1  ( .A1(\SB1_2_7/i0[9] ), .A2(
        \SB1_2_7/i0_0 ), .A3(\SB1_2_7/i0[8] ), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_2/N2  ( .A1(\SB1_2_8/i0_3 ), .A2(
        \SB1_2_8/i0[10] ), .A3(\SB1_2_8/i0[6] ), .ZN(
        \SB1_2_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_8/Component_Function_2/N1  ( .A1(\SB1_2_8/i1_5 ), .A2(
        \SB1_2_8/i0[10] ), .A3(\SB1_2_8/i1[9] ), .ZN(
        \SB1_2_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_3/N4  ( .A1(\SB1_2_8/i1_5 ), .A2(
        \SB1_2_8/i0[8] ), .A3(\SB1_2_8/i3[0] ), .ZN(
        \SB1_2_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_8/Component_Function_3/N3  ( .A1(\SB1_2_8/i1[9] ), .A2(
        \SB1_2_8/i1_7 ), .A3(\SB1_2_8/i0[10] ), .ZN(
        \SB1_2_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_8/Component_Function_3/N1  ( .A1(\SB1_2_8/i1[9] ), .A2(
        \SB1_2_8/i0_3 ), .A3(\SB1_2_8/i0[6] ), .ZN(
        \SB1_2_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_4/N4  ( .A1(\SB1_2_8/i1[9] ), .A2(
        \SB1_2_8/i1_5 ), .A3(\SB1_2_8/i0_4 ), .ZN(
        \SB1_2_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_8/Component_Function_4/N2  ( .A1(\SB1_2_8/i3[0] ), .A2(
        \SB1_2_8/i0_0 ), .A3(\SB1_2_8/i1_7 ), .ZN(
        \SB1_2_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_8/Component_Function_4/N1  ( .A1(\SB1_2_8/i0[9] ), .A2(
        \SB1_2_8/i0_0 ), .A3(\SB1_2_8/i0[8] ), .ZN(
        \SB1_2_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_2/N2  ( .A1(n1657), .A2(
        \SB1_2_9/i0[10] ), .A3(\SB1_2_9/i0[6] ), .ZN(
        \SB1_2_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_9/Component_Function_2/N1  ( .A1(\SB1_2_9/i1_5 ), .A2(
        \SB1_2_9/i0[10] ), .A3(\SB1_2_9/i1[9] ), .ZN(
        \SB1_2_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_3/N4  ( .A1(\SB1_2_9/i1_5 ), .A2(
        \SB1_2_9/i0[8] ), .A3(\SB1_2_9/i3[0] ), .ZN(
        \SB1_2_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_9/Component_Function_3/N1  ( .A1(\SB1_2_9/i1[9] ), .A2(n1657), .A3(\SB1_2_9/i0[6] ), .ZN(\SB1_2_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_4/N4  ( .A1(\SB1_2_9/i1[9] ), .A2(
        \SB1_2_9/i1_5 ), .A3(\SB1_2_9/i0_4 ), .ZN(
        \SB1_2_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_9/Component_Function_4/N2  ( .A1(\SB1_2_9/i3[0] ), .A2(
        \SB1_2_9/i0_0 ), .A3(\SB1_2_9/i1_7 ), .ZN(
        \SB1_2_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_9/Component_Function_4/N1  ( .A1(\SB1_2_9/i0[9] ), .A2(
        \SB1_2_9/i0_0 ), .A3(\SB1_2_9/i0[8] ), .ZN(
        \SB1_2_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_2/N2  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i0[10] ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_10/Component_Function_2/N1  ( .A1(\SB1_2_10/i1_5 ), .A2(
        \SB1_2_10/i0[10] ), .A3(\SB1_2_10/i1[9] ), .ZN(
        \SB1_2_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_3/N4  ( .A1(\SB1_2_10/i1_5 ), .A2(
        \SB1_2_10/i0[8] ), .A3(\SB1_2_10/i3[0] ), .ZN(
        \SB1_2_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_10/Component_Function_3/N1  ( .A1(\SB1_2_10/i1[9] ), .A2(
        \SB1_2_10/i0_3 ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_4/N4  ( .A1(\SB1_2_10/i1[9] ), .A2(
        \SB1_2_10/i1_5 ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_10/Component_Function_4/N2  ( .A1(\SB1_2_10/i3[0] ), .A2(
        \SB1_2_10/i0_0 ), .A3(\SB1_2_10/i1_7 ), .ZN(
        \SB1_2_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_10/Component_Function_4/N1  ( .A1(\SB1_2_10/i0[9] ), .A2(
        \SB1_2_10/i0_0 ), .A3(\SB1_2_10/i0[8] ), .ZN(
        \SB1_2_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_2/N2  ( .A1(\SB1_2_11/i0_3 ), .A2(
        \SB1_2_11/i0[10] ), .A3(\SB1_2_11/i0[6] ), .ZN(
        \SB1_2_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_11/Component_Function_2/N1  ( .A1(\SB1_2_11/i1_5 ), .A2(
        \SB1_2_11/i0[10] ), .A3(\SB1_2_11/i1[9] ), .ZN(
        \SB1_2_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_3/N4  ( .A1(\SB1_2_11/i1_5 ), .A2(
        \SB1_2_11/i0[8] ), .A3(\SB1_2_11/i3[0] ), .ZN(
        \SB1_2_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_11/Component_Function_3/N1  ( .A1(\SB1_2_11/i1[9] ), .A2(
        \SB1_2_11/i0_3 ), .A3(\SB1_2_11/i0[6] ), .ZN(
        \SB1_2_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_4/N4  ( .A1(\SB1_2_11/i1[9] ), .A2(
        \SB1_2_11/i1_5 ), .A3(\SB1_2_11/i0_4 ), .ZN(
        \SB1_2_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_11/Component_Function_4/N2  ( .A1(\SB1_2_11/i3[0] ), .A2(
        \SB1_2_11/i0_0 ), .A3(\SB1_2_11/i1_7 ), .ZN(
        \SB1_2_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_11/Component_Function_4/N1  ( .A1(\SB1_2_11/i0[9] ), .A2(
        \SB1_2_11/i0_0 ), .A3(\SB1_2_11/i0[8] ), .ZN(
        \SB1_2_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_2/N2  ( .A1(\SB1_2_12/i0[10] ), .A2(
        \SB1_2_12/i0_3 ), .A3(\SB1_2_12/i0[6] ), .ZN(
        \SB1_2_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_12/Component_Function_2/N1  ( .A1(\SB1_2_12/i1_5 ), .A2(
        \SB1_2_12/i0[10] ), .A3(\SB1_2_12/i1[9] ), .ZN(
        \SB1_2_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_3/N1  ( .A1(\SB1_2_12/i1[9] ), .A2(
        \SB1_2_12/i0_3 ), .A3(\SB1_2_12/i0[6] ), .ZN(
        \SB1_2_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_4/N4  ( .A1(\SB1_2_12/i1[9] ), .A2(
        \SB1_2_12/i1_5 ), .A3(\SB1_2_12/i0_4 ), .ZN(
        \SB1_2_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_12/Component_Function_4/N2  ( .A1(\SB1_2_12/i3[0] ), .A2(
        \SB1_2_12/i0_0 ), .A3(\SB1_2_12/i1_7 ), .ZN(
        \SB1_2_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_12/Component_Function_4/N1  ( .A1(\SB1_2_12/i0[9] ), .A2(
        \SB1_2_12/i0_0 ), .A3(\SB1_2_12/i0[8] ), .ZN(
        \SB1_2_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_2/N2  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i0[10] ), .A3(\SB1_2_13/i0[6] ), .ZN(
        \SB1_2_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_13/Component_Function_2/N1  ( .A1(\SB1_2_13/i1_5 ), .A2(
        \SB1_2_13/i0[10] ), .A3(\SB1_2_13/i1[9] ), .ZN(
        \SB1_2_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_3/N4  ( .A1(\SB1_2_13/i1_5 ), .A2(
        \SB1_2_13/i0[8] ), .A3(\SB1_2_13/i3[0] ), .ZN(
        \SB1_2_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_13/Component_Function_3/N3  ( .A1(\SB1_2_13/i1[9] ), .A2(
        \SB1_2_13/i1_7 ), .A3(\SB1_2_13/i0[10] ), .ZN(
        \SB1_2_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_13/Component_Function_3/N1  ( .A1(\SB1_2_13/i1[9] ), .A2(
        \SB1_2_13/i0_3 ), .A3(\SB1_2_13/i0[6] ), .ZN(
        \SB1_2_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_4/N4  ( .A1(\SB1_2_13/i1[9] ), .A2(
        \SB1_2_13/i1_5 ), .A3(\SB1_2_13/i0_4 ), .ZN(
        \SB1_2_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_13/Component_Function_4/N2  ( .A1(\SB1_2_13/i3[0] ), .A2(
        \SB1_2_13/i0_0 ), .A3(\SB1_2_13/i1_7 ), .ZN(
        \SB1_2_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_13/Component_Function_4/N1  ( .A1(\SB1_2_13/i0[9] ), .A2(
        \SB1_2_13/i0_0 ), .A3(\SB1_2_13/i0[8] ), .ZN(
        \SB1_2_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_2/N2  ( .A1(\SB1_2_14/i0_3 ), .A2(
        \SB1_2_14/i0[10] ), .A3(\SB1_2_14/i0[6] ), .ZN(
        \SB1_2_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_14/Component_Function_2/N1  ( .A1(\SB1_2_14/i1_5 ), .A2(
        \SB1_2_14/i0[10] ), .A3(\SB1_2_14/i1[9] ), .ZN(
        \SB1_2_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_3/N4  ( .A1(\SB1_2_14/i1_5 ), .A2(
        \SB1_2_14/i0[8] ), .A3(\SB1_2_14/i3[0] ), .ZN(
        \SB1_2_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_14/Component_Function_3/N1  ( .A1(\SB1_2_14/i1[9] ), .A2(
        \SB1_2_14/i0_3 ), .A3(\SB1_2_14/i0[6] ), .ZN(
        \SB1_2_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N4  ( .A1(\SB1_2_14/i1[9] ), .A2(
        \SB1_2_14/i1_5 ), .A3(\SB1_2_14/i0_4 ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N2  ( .A1(\SB1_2_14/i3[0] ), .A2(
        \SB1_2_14/i0_0 ), .A3(\SB1_2_14/i1_7 ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N1  ( .A1(\SB1_2_14/i0[9] ), .A2(
        \SB1_2_14/i0_0 ), .A3(\SB1_2_14/i0[8] ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_2/N2  ( .A1(\SB1_2_15/i0_3 ), .A2(
        \SB1_2_15/i0[10] ), .A3(\SB1_2_15/i0[6] ), .ZN(
        \SB1_2_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_15/Component_Function_2/N1  ( .A1(\SB1_2_15/i1_5 ), .A2(
        \SB1_2_15/i0[10] ), .A3(\SB1_2_15/i1[9] ), .ZN(
        \SB1_2_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_3/N4  ( .A1(\SB1_2_15/i1_5 ), .A2(
        \SB1_2_15/i0[8] ), .A3(\SB1_2_15/i3[0] ), .ZN(
        \SB1_2_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_15/Component_Function_3/N1  ( .A1(\SB1_2_15/i1[9] ), .A2(
        \SB1_2_15/i0_3 ), .A3(\SB1_2_15/i0[6] ), .ZN(
        \SB1_2_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_4/N4  ( .A1(\SB1_2_15/i1[9] ), .A2(
        \SB1_2_15/i1_5 ), .A3(\SB1_2_15/i0_4 ), .ZN(
        \SB1_2_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_15/Component_Function_4/N2  ( .A1(\SB1_2_15/i3[0] ), .A2(
        \SB1_2_15/i0_0 ), .A3(\SB1_2_15/i1_7 ), .ZN(
        \SB1_2_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_15/Component_Function_4/N1  ( .A1(\SB1_2_15/i0[9] ), .A2(
        \SB1_2_15/i0_0 ), .A3(\SB1_2_15/i0[8] ), .ZN(
        \SB1_2_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_2/N3  ( .A1(\SB1_2_16/i0_3 ), .A2(
        \SB1_2_16/i0[8] ), .A3(\SB1_2_16/i0[9] ), .ZN(
        \SB1_2_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_16/Component_Function_2/N2  ( .A1(\SB1_2_16/i0_3 ), .A2(
        \SB1_2_16/i0[10] ), .A3(\SB1_2_16/i0[6] ), .ZN(
        \SB1_2_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_16/Component_Function_2/N1  ( .A1(\SB1_2_16/i1_5 ), .A2(
        \SB1_2_16/i0[10] ), .A3(\SB1_2_16/i1[9] ), .ZN(
        \SB1_2_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_3/N4  ( .A1(\SB1_2_16/i1_5 ), .A2(
        \SB1_2_16/i0[8] ), .A3(\SB1_2_16/i3[0] ), .ZN(
        \SB1_2_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_16/Component_Function_3/N3  ( .A1(\SB1_2_16/i1[9] ), .A2(
        \SB1_2_16/i1_7 ), .A3(\SB1_2_16/i0[10] ), .ZN(
        \SB1_2_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_16/Component_Function_3/N1  ( .A1(\SB1_2_16/i1[9] ), .A2(
        \SB1_2_16/i0_3 ), .A3(\SB1_2_16/i0[6] ), .ZN(
        \SB1_2_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_4/N2  ( .A1(\SB1_2_16/i3[0] ), .A2(
        \SB1_2_16/i0_0 ), .A3(\SB1_2_16/i1_7 ), .ZN(
        \SB1_2_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_16/Component_Function_4/N1  ( .A1(\SB1_2_16/i0[9] ), .A2(
        \SB1_2_16/i0_0 ), .A3(\SB1_2_16/i0[8] ), .ZN(
        \SB1_2_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_2/N2  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i0[10] ), .A3(\SB1_2_17/i0[6] ), .ZN(
        \SB1_2_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_17/Component_Function_2/N1  ( .A1(\SB1_2_17/i1_5 ), .A2(
        \SB1_2_17/i0[10] ), .A3(\SB1_2_17/i1[9] ), .ZN(
        \SB1_2_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_3/N3  ( .A1(\SB1_2_17/i1[9] ), .A2(
        \SB1_2_17/i1_7 ), .A3(\SB1_2_17/i0[10] ), .ZN(
        \SB1_2_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_17/Component_Function_3/N1  ( .A1(\SB1_2_17/i1[9] ), .A2(
        \SB1_2_17/i0_3 ), .A3(\SB1_2_17/i0[6] ), .ZN(
        \SB1_2_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_4/N2  ( .A1(\SB1_2_17/i3[0] ), .A2(
        \SB1_2_17/i0_0 ), .A3(\SB1_2_17/i1_7 ), .ZN(
        \SB1_2_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_17/Component_Function_4/N1  ( .A1(\SB1_2_17/i0[9] ), .A2(
        \SB1_2_17/i0_0 ), .A3(\SB1_2_17/i0[8] ), .ZN(
        \SB1_2_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_2/N2  ( .A1(\SB1_2_18/i0_3 ), .A2(
        \SB1_2_18/i0[10] ), .A3(\SB1_2_18/i0[6] ), .ZN(
        \SB1_2_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_18/Component_Function_2/N1  ( .A1(\SB1_2_18/i1_5 ), .A2(
        \SB1_2_18/i0[10] ), .A3(\SB1_2_18/i1[9] ), .ZN(
        \SB1_2_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_3/N4  ( .A1(\SB1_2_18/i1_5 ), .A2(
        \SB1_2_18/i0[8] ), .A3(\SB1_2_18/i3[0] ), .ZN(
        \SB1_2_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_18/Component_Function_3/N1  ( .A1(\SB1_2_18/i1[9] ), .A2(
        \SB1_2_18/i0_3 ), .A3(\SB1_2_18/i0[6] ), .ZN(
        \SB1_2_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_4/N4  ( .A1(\SB1_2_18/i1[9] ), .A2(
        \SB1_2_18/i1_5 ), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_18/Component_Function_4/N2  ( .A1(\SB1_2_18/i3[0] ), .A2(
        \SB1_2_18/i0_0 ), .A3(\SB1_2_18/i1_7 ), .ZN(
        \SB1_2_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_18/Component_Function_4/N1  ( .A1(\SB1_2_18/i0[9] ), .A2(
        \SB1_2_18/i0_0 ), .A3(\SB1_2_18/i0[8] ), .ZN(
        \SB1_2_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_2/N2  ( .A1(n1649), .A2(
        \SB1_2_19/i0[10] ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_19/Component_Function_2/N1  ( .A1(\SB1_2_19/i1_5 ), .A2(
        \SB1_2_19/i0[10] ), .A3(\SB1_2_19/i1[9] ), .ZN(
        \SB1_2_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_3/N4  ( .A1(\SB1_2_19/i1_5 ), .A2(
        \SB1_2_19/i0[8] ), .A3(\SB1_2_19/i3[0] ), .ZN(
        \SB1_2_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_3/N3  ( .A1(\SB1_2_19/i1[9] ), .A2(
        \SB1_2_19/i1_7 ), .A3(\SB1_2_19/i0[10] ), .ZN(
        \SB1_2_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_19/Component_Function_3/N1  ( .A1(\SB1_2_19/i1[9] ), .A2(
        n1649), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_4/N4  ( .A1(\SB1_2_19/i1[9] ), .A2(
        \SB1_2_19/i1_5 ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_4/N2  ( .A1(\SB1_2_19/i3[0] ), .A2(
        \SB1_2_19/i0_0 ), .A3(\SB1_2_19/i1_7 ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_19/Component_Function_4/N1  ( .A1(\SB1_2_19/i0[9] ), .A2(
        \SB1_2_19/i0_0 ), .A3(\SB1_2_19/i0[8] ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_2/N2  ( .A1(\SB1_2_20/i0_3 ), .A2(
        \SB1_2_20/i0[10] ), .A3(\SB1_2_20/i0[6] ), .ZN(
        \SB1_2_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_20/Component_Function_2/N1  ( .A1(\SB1_2_20/i1_5 ), .A2(
        \SB1_2_20/i0[10] ), .A3(\SB1_2_20/i1[9] ), .ZN(
        \SB1_2_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_3/N4  ( .A1(\SB1_2_20/i1_5 ), .A2(
        \SB1_2_20/i0[8] ), .A3(\SB1_2_20/i3[0] ), .ZN(
        \SB1_2_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_3/N1  ( .A1(\SB1_2_20/i1[9] ), .A2(
        n1644), .A3(\SB1_2_20/i0[6] ), .ZN(
        \SB1_2_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N4  ( .A1(\SB1_2_20/i1[9] ), .A2(
        \SB1_2_20/i1_5 ), .A3(\SB1_2_20/i0_4 ), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N2  ( .A1(\SB1_2_20/i3[0] ), .A2(
        \SB1_2_20/i0_0 ), .A3(\SB1_2_20/i1_7 ), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N1  ( .A1(\SB1_2_20/i0[9] ), .A2(
        \SB1_2_20/i0_0 ), .A3(\SB1_2_20/i0[8] ), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_2/N2  ( .A1(\SB1_2_21/i0_3 ), .A2(
        \SB1_2_21/i0[10] ), .A3(\SB1_2_21/i0[6] ), .ZN(
        \SB1_2_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_21/Component_Function_2/N1  ( .A1(\SB1_2_21/i1_5 ), .A2(
        \SB1_2_21/i0[10] ), .A3(\SB1_2_21/i1[9] ), .ZN(
        \SB1_2_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_3/N4  ( .A1(\SB1_2_21/i1_5 ), .A2(
        \SB1_2_21/i0[8] ), .A3(\SB1_2_21/i3[0] ), .ZN(
        \SB1_2_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_21/Component_Function_3/N1  ( .A1(\SB1_2_21/i1[9] ), .A2(
        \SB1_2_21/i0_3 ), .A3(\SB1_2_21/i0[6] ), .ZN(
        \SB1_2_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_4/N4  ( .A1(\SB1_2_21/i1[9] ), .A2(
        \SB1_2_21/i1_5 ), .A3(\SB1_2_21/i0_4 ), .ZN(
        \SB1_2_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_21/Component_Function_4/N2  ( .A1(\SB1_2_21/i3[0] ), .A2(
        \SB1_2_21/i0_0 ), .A3(\SB1_2_21/i1_7 ), .ZN(
        \SB1_2_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_21/Component_Function_4/N1  ( .A1(\SB1_2_21/i0[9] ), .A2(
        \SB1_2_21/i0_0 ), .A3(\SB1_2_21/i0[8] ), .ZN(
        \SB1_2_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_2/N2  ( .A1(\SB1_2_22/i0_3 ), .A2(
        \SB1_2_22/i0[10] ), .A3(\SB1_2_22/i0[6] ), .ZN(
        \SB1_2_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_22/Component_Function_2/N1  ( .A1(\SB1_2_22/i1_5 ), .A2(
        \SB1_2_22/i0[10] ), .A3(\SB1_2_22/i1[9] ), .ZN(
        \SB1_2_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_3/N4  ( .A1(\SB1_2_22/i1_5 ), .A2(
        \SB1_2_22/i0[8] ), .A3(\SB1_2_22/i3[0] ), .ZN(
        \SB1_2_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_22/Component_Function_3/N1  ( .A1(\SB1_2_22/i1[9] ), .A2(
        \SB1_2_22/i0_3 ), .A3(\SB1_2_22/i0[6] ), .ZN(
        \SB1_2_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_4/N4  ( .A1(\SB1_2_22/i1[9] ), .A2(
        \SB1_2_22/i1_5 ), .A3(\SB1_2_22/i0_4 ), .ZN(
        \SB1_2_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_22/Component_Function_4/N2  ( .A1(\SB1_2_22/i3[0] ), .A2(
        \SB1_2_22/i0_0 ), .A3(\SB1_2_22/i1_7 ), .ZN(
        \SB1_2_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_22/Component_Function_4/N1  ( .A1(\SB1_2_22/i0[9] ), .A2(
        \SB1_2_22/i0_0 ), .A3(\SB1_2_22/i0[8] ), .ZN(
        \SB1_2_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_2/N2  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_2/N1  ( .A1(\SB1_2_23/i1_5 ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i1[9] ), .ZN(
        \SB1_2_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_3/N4  ( .A1(\SB1_2_23/i1_5 ), .A2(
        \SB1_2_23/i0[8] ), .A3(\SB1_2_23/i3[0] ), .ZN(
        \SB1_2_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_23/Component_Function_3/N1  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i0_3 ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N4  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i1_5 ), .A3(\SB1_2_23/i0_4 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N2  ( .A1(\SB1_2_23/i3[0] ), .A2(
        \SB1_2_23/i0_0 ), .A3(\SB1_2_23/i1_7 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N1  ( .A1(\SB1_2_23/i0[9] ), .A2(
        \SB1_2_23/i0_0 ), .A3(\SB1_2_23/i0[8] ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_2/N2  ( .A1(\SB1_2_24/i0_3 ), .A2(
        \SB1_2_24/i0[10] ), .A3(\SB1_2_24/i0[6] ), .ZN(
        \SB1_2_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_24/Component_Function_2/N1  ( .A1(\SB1_2_24/i1_5 ), .A2(
        \SB1_2_24/i0[10] ), .A3(\SB1_2_24/i1[9] ), .ZN(
        \SB1_2_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_3/N4  ( .A1(\SB1_2_24/i1_5 ), .A2(
        \SB1_2_24/i0[8] ), .A3(\SB1_2_24/i3[0] ), .ZN(
        \SB1_2_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_24/Component_Function_3/N2  ( .A1(\SB1_2_24/i0_0 ), .A2(
        \SB1_2_24/i0_3 ), .A3(\SB1_2_24/i0_4 ), .ZN(
        \SB1_2_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_24/Component_Function_3/N1  ( .A1(\SB1_2_24/i1[9] ), .A2(
        \SB1_2_24/i0_3 ), .A3(\SB1_2_24/i0[6] ), .ZN(
        \SB1_2_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_4/N4  ( .A1(\SB1_2_24/i1[9] ), .A2(
        \SB1_2_24/i1_5 ), .A3(\SB1_2_24/i0_4 ), .ZN(
        \SB1_2_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_24/Component_Function_4/N2  ( .A1(\SB1_2_24/i3[0] ), .A2(
        \SB1_2_24/i0_0 ), .A3(\SB1_2_24/i1_7 ), .ZN(
        \SB1_2_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_24/Component_Function_4/N1  ( .A1(\SB1_2_24/i0[9] ), .A2(
        \SB1_2_24/i0_0 ), .A3(\SB1_2_24/i0[8] ), .ZN(
        \SB1_2_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_2/N2  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i0[10] ), .A3(\SB1_2_25/i0[6] ), .ZN(
        \SB1_2_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_25/Component_Function_2/N1  ( .A1(\SB1_2_25/i1_5 ), .A2(
        \SB1_2_25/i0[10] ), .A3(\SB1_2_25/i1[9] ), .ZN(
        \SB1_2_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_3/N4  ( .A1(\SB1_2_25/i1_5 ), .A2(
        \SB1_2_25/i0[8] ), .A3(\SB1_2_25/i3[0] ), .ZN(
        \SB1_2_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_3/N3  ( .A1(\SB1_2_25/i1[9] ), .A2(
        \SB1_2_25/i1_7 ), .A3(\SB1_2_25/i0[10] ), .ZN(
        \SB1_2_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_3/N1  ( .A1(\SB1_2_25/i1[9] ), .A2(
        \SB1_2_25/i0_3 ), .A3(\SB1_2_25/i0[6] ), .ZN(
        \SB1_2_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_4/N4  ( .A1(\SB1_2_25/i1[9] ), .A2(
        \SB1_2_25/i1_5 ), .A3(\SB1_2_25/i0_4 ), .ZN(
        \SB1_2_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_4/N2  ( .A1(\SB1_2_25/i3[0] ), .A2(
        \SB1_2_25/i0_0 ), .A3(\SB1_2_25/i1_7 ), .ZN(
        \SB1_2_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_25/Component_Function_4/N1  ( .A1(\SB1_2_25/i0[9] ), .A2(
        \SB1_2_25/i0_0 ), .A3(\SB1_2_25/i0[8] ), .ZN(
        \SB1_2_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_2/N2  ( .A1(\SB1_2_26/i0_3 ), .A2(
        \SB1_2_26/i0[10] ), .A3(\SB1_2_26/i0[6] ), .ZN(
        \SB1_2_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_26/Component_Function_2/N1  ( .A1(\SB1_2_26/i1_5 ), .A2(
        \SB1_2_26/i0[10] ), .A3(\SB1_2_26/i1[9] ), .ZN(
        \SB1_2_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_3/N4  ( .A1(\SB1_2_26/i1_5 ), .A2(
        \SB1_2_26/i0[8] ), .A3(\SB1_2_26/i3[0] ), .ZN(
        \SB1_2_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_26/Component_Function_3/N3  ( .A1(\SB1_2_26/i1[9] ), .A2(
        \SB1_2_26/i1_7 ), .A3(\SB1_2_26/i0[10] ), .ZN(
        \SB1_2_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_26/Component_Function_3/N1  ( .A1(\SB1_2_26/i1[9] ), .A2(
        \SB1_2_26/i0_3 ), .A3(\SB1_2_26/i0[6] ), .ZN(
        \SB1_2_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_4/N4  ( .A1(\SB1_2_26/i1[9] ), .A2(
        \SB1_2_26/i1_5 ), .A3(\SB1_2_26/i0_4 ), .ZN(
        \SB1_2_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_26/Component_Function_4/N2  ( .A1(\SB1_2_26/i3[0] ), .A2(
        \SB1_2_26/i0_0 ), .A3(\SB1_2_26/i1_7 ), .ZN(
        \SB1_2_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_26/Component_Function_4/N1  ( .A1(\SB1_2_26/i0[9] ), .A2(
        \SB1_2_26/i0_0 ), .A3(\SB1_2_26/i0[8] ), .ZN(
        \SB1_2_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_2/N2  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i0[10] ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_27/Component_Function_2/N1  ( .A1(\SB1_2_27/i1_5 ), .A2(
        \SB1_2_27/i0[10] ), .A3(\SB1_2_27/i1[9] ), .ZN(
        \SB1_2_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_3/N4  ( .A1(\SB1_2_27/i1_5 ), .A2(
        \SB1_2_27/i0[8] ), .A3(\SB1_2_27/i3[0] ), .ZN(
        \SB1_2_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_3/N3  ( .A1(\SB1_2_27/i1[9] ), .A2(
        \SB1_2_27/i1_7 ), .A3(\SB1_2_27/i0[10] ), .ZN(
        \SB1_2_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_27/Component_Function_3/N1  ( .A1(\SB1_2_27/i1[9] ), .A2(
        \SB1_2_27/i0_3 ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_4/N4  ( .A1(\SB1_2_27/i1[9] ), .A2(
        \SB1_2_27/i1_5 ), .A3(\SB1_2_27/i0_4 ), .ZN(
        \SB1_2_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_4/N2  ( .A1(\SB1_2_27/i3[0] ), .A2(
        \SB1_2_27/i0_0 ), .A3(\SB1_2_27/i1_7 ), .ZN(
        \SB1_2_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_27/Component_Function_4/N1  ( .A1(\SB1_2_27/i0[9] ), .A2(
        \SB1_2_27/i0_0 ), .A3(\SB1_2_27/i0[8] ), .ZN(
        \SB1_2_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_2/N2  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i0[10] ), .A3(\SB1_2_28/i0[6] ), .ZN(
        \SB1_2_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_28/Component_Function_2/N1  ( .A1(\SB1_2_28/i1_5 ), .A2(
        \SB1_2_28/i0[10] ), .A3(\SB1_2_28/i1[9] ), .ZN(
        \SB1_2_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_3/N4  ( .A1(\SB1_2_28/i1_5 ), .A2(
        \SB1_2_28/i0[8] ), .A3(\SB1_2_28/i3[0] ), .ZN(
        \SB1_2_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_3/N1  ( .A1(\SB1_2_28/i1[9] ), .A2(
        \SB1_2_28/i0_3 ), .A3(\SB1_2_28/i0[6] ), .ZN(
        \SB1_2_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_4/N4  ( .A1(\SB1_2_28/i1[9] ), .A2(
        \SB1_2_28/i1_5 ), .A3(\SB1_2_28/i0_4 ), .ZN(
        \SB1_2_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_4/N1  ( .A1(\SB1_2_28/i0[9] ), .A2(
        \SB1_2_28/i0_0 ), .A3(\SB1_2_28/i0[8] ), .ZN(
        \SB1_2_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_2/N2  ( .A1(\SB1_2_29/i0_3 ), .A2(
        \SB1_2_29/i0[10] ), .A3(\SB1_2_29/i0[6] ), .ZN(
        \SB1_2_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_29/Component_Function_2/N1  ( .A1(\SB1_2_29/i1_5 ), .A2(
        \SB1_2_29/i0[10] ), .A3(\SB1_2_29/i1[9] ), .ZN(
        \SB1_2_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_3/N4  ( .A1(\SB1_2_29/i1_5 ), .A2(
        \SB1_2_29/i0[8] ), .A3(\SB1_2_29/i3[0] ), .ZN(
        \SB1_2_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_29/Component_Function_3/N1  ( .A1(\SB1_2_29/i1[9] ), .A2(
        n814), .A3(\SB1_2_29/i0[6] ), .ZN(
        \SB1_2_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_4/N4  ( .A1(\SB1_2_29/i1[9] ), .A2(
        \SB1_2_29/i1_5 ), .A3(\SB1_2_29/i0_4 ), .ZN(
        \SB1_2_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_29/Component_Function_4/N2  ( .A1(\SB1_2_29/i3[0] ), .A2(
        \SB1_2_29/i0_0 ), .A3(\SB1_2_29/i1_7 ), .ZN(
        \SB1_2_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_29/Component_Function_4/N1  ( .A1(\SB1_2_29/i0[9] ), .A2(
        \SB1_2_29/i0_0 ), .A3(\SB1_2_29/i0[8] ), .ZN(
        \SB1_2_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_2/N2  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i0[10] ), .A3(\SB1_2_30/i0[6] ), .ZN(
        \SB1_2_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_30/Component_Function_2/N1  ( .A1(\SB1_2_30/i1_5 ), .A2(
        \SB1_2_30/i0[10] ), .A3(\SB1_2_30/i1[9] ), .ZN(
        \SB1_2_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_3/N4  ( .A1(\SB1_2_30/i1_5 ), .A2(
        \SB1_2_30/i0[8] ), .A3(\SB1_2_30/i3[0] ), .ZN(
        \SB1_2_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_30/Component_Function_3/N1  ( .A1(\SB1_2_30/i1[9] ), .A2(
        \SB1_2_30/i0_3 ), .A3(\SB1_2_30/i0[6] ), .ZN(
        \SB1_2_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_4/N4  ( .A1(\SB1_2_30/i1[9] ), .A2(
        \SB1_2_30/i1_5 ), .A3(\SB1_2_30/i0_4 ), .ZN(
        \SB1_2_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_30/Component_Function_4/N2  ( .A1(\SB1_2_30/i3[0] ), .A2(
        \SB1_2_30/i0_0 ), .A3(\SB1_2_30/i1_7 ), .ZN(
        \SB1_2_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_30/Component_Function_4/N1  ( .A1(\SB1_2_30/i0[9] ), .A2(
        \SB1_2_30/i0_0 ), .A3(\SB1_2_30/i0[8] ), .ZN(
        \SB1_2_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_2/N4  ( .A1(\SB1_2_31/i1_5 ), .A2(
        \SB1_2_31/i0_0 ), .A3(\SB1_2_31/i0_4 ), .ZN(
        \SB1_2_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_31/Component_Function_2/N2  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i0[10] ), .A3(\SB1_2_31/i0[6] ), .ZN(
        \SB1_2_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_31/Component_Function_2/N1  ( .A1(\SB1_2_31/i1_5 ), .A2(
        \SB1_2_31/i0[10] ), .A3(\SB1_2_31/i1[9] ), .ZN(
        \SB1_2_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_4/N4  ( .A1(\SB1_2_31/i1[9] ), .A2(
        \SB1_2_31/i1_5 ), .A3(\SB1_2_31/i0_4 ), .ZN(
        \SB1_2_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_31/Component_Function_4/N2  ( .A1(\SB1_2_31/i3[0] ), .A2(
        \SB1_2_31/i0_0 ), .A3(\SB1_2_31/i1_7 ), .ZN(
        \SB1_2_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_31/Component_Function_4/N1  ( .A1(\SB1_2_31/i0[9] ), .A2(
        \SB1_2_31/i0_0 ), .A3(\SB1_2_31/i0[8] ), .ZN(
        \SB1_2_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_2/N3  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i0[8] ), .A3(\SB2_2_0/i0[9] ), .ZN(
        \SB2_2_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_0/Component_Function_2/N2  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i0[10] ), .A3(\SB2_2_0/i0[6] ), .ZN(
        \SB2_2_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_0/Component_Function_3/N3  ( .A1(\SB2_2_0/i1[9] ), .A2(
        \SB2_2_0/i1_7 ), .A3(\SB2_2_0/i0[10] ), .ZN(
        \SB2_2_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_0/Component_Function_3/N1  ( .A1(\SB2_2_0/i1[9] ), .A2(
        \SB2_2_0/i0_3 ), .A3(\SB2_2_0/i0[6] ), .ZN(
        \SB2_2_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_4/N4  ( .A1(\SB2_2_0/i1[9] ), .A2(
        \SB2_2_0/i1_5 ), .A3(\SB2_2_0/i0_4 ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_0/Component_Function_4/N2  ( .A1(\SB2_2_0/i3[0] ), .A2(
        \SB2_2_0/i0_0 ), .A3(\SB2_2_0/i1_7 ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_0/Component_Function_4/N1  ( .A1(\SB2_2_0/i0[9] ), .A2(
        \SB2_2_0/i0_0 ), .A3(\SB2_2_0/i0[8] ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_2/N1  ( .A1(\SB2_2_1/i1_5 ), .A2(
        \SB2_2_1/i0[10] ), .A3(\SB2_2_1/i1[9] ), .ZN(
        \SB2_2_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_3/N3  ( .A1(\SB2_2_1/i1[9] ), .A2(
        \SB2_2_1/i1_7 ), .A3(\SB2_2_1/i0[10] ), .ZN(
        \SB2_2_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_1/Component_Function_3/N2  ( .A1(\SB2_2_1/i0_0 ), .A2(
        \SB2_2_1/i0_3 ), .A3(\SB2_2_1/i0_4 ), .ZN(
        \SB2_2_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_1/Component_Function_4/N3  ( .A1(\SB2_2_1/i0[9] ), .A2(
        \SB2_2_1/i0[10] ), .A3(\SB2_2_1/i0_3 ), .ZN(
        \SB2_2_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_1/Component_Function_4/N2  ( .A1(\SB2_2_1/i3[0] ), .A2(
        \SB2_2_1/i0_0 ), .A3(\SB2_2_1/i1_7 ), .ZN(
        \SB2_2_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_1/Component_Function_4/N1  ( .A1(\SB2_2_1/i0[9] ), .A2(
        \SB2_2_1/i0_0 ), .A3(\SB2_2_1/i0[8] ), .ZN(
        \SB2_2_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_2/N2  ( .A1(\SB2_2_2/i0_3 ), .A2(
        \SB2_2_2/i0[10] ), .A3(\SB2_2_2/i0[6] ), .ZN(
        \SB2_2_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_2/Component_Function_2/N1  ( .A1(\SB2_2_2/i1_5 ), .A2(
        \SB2_2_2/i0[10] ), .A3(\SB2_2_2/i1[9] ), .ZN(
        \SB2_2_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_3/N3  ( .A1(\SB2_2_2/i1[9] ), .A2(
        \SB2_2_2/i1_7 ), .A3(\SB2_2_2/i0[10] ), .ZN(
        \SB2_2_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_2/Component_Function_3/N2  ( .A1(\SB2_2_2/i0_0 ), .A2(
        \SB2_2_2/i0_3 ), .A3(\SB2_2_2/i0_4 ), .ZN(
        \SB2_2_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_2/Component_Function_4/N3  ( .A1(\SB2_2_2/i0[9] ), .A2(
        \SB2_2_2/i0[10] ), .A3(\SB2_2_2/i0_3 ), .ZN(
        \SB2_2_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_2/Component_Function_4/N1  ( .A1(\SB2_2_2/i0[9] ), .A2(
        \SB2_2_2/i0_0 ), .A3(\SB2_2_2/i0[8] ), .ZN(
        \SB2_2_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_3/Component_Function_2/N4  ( .A1(\SB2_2_3/i1_5 ), .A2(
        \SB2_2_3/i0_0 ), .A3(\SB2_2_3/i0_4 ), .ZN(
        \SB2_2_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_3/Component_Function_2/N2  ( .A1(\SB2_2_3/i0_3 ), .A2(
        \SB2_2_3/i0[10] ), .A3(\SB2_2_3/i0[6] ), .ZN(
        \SB2_2_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_3/Component_Function_2/N1  ( .A1(\SB2_2_3/i1_5 ), .A2(
        \SB2_2_3/i0[10] ), .A3(\SB2_2_3/i1[9] ), .ZN(
        \SB2_2_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_3/Component_Function_3/N3  ( .A1(\SB2_2_3/i1[9] ), .A2(
        \SB2_2_3/i1_7 ), .A3(\SB2_2_3/i0[10] ), .ZN(
        \SB2_2_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_3/Component_Function_3/N2  ( .A1(\SB2_2_3/i0_0 ), .A2(
        \SB2_2_3/i0_3 ), .A3(\SB2_2_3/i0_4 ), .ZN(
        \SB2_2_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_3/Component_Function_3/N1  ( .A1(\SB2_2_3/i1[9] ), .A2(
        \SB2_2_3/i0_3 ), .A3(\SB2_2_3/i0[6] ), .ZN(
        \SB2_2_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_3/Component_Function_4/N4  ( .A1(\SB2_2_3/i1[9] ), .A2(
        \SB2_2_3/i1_5 ), .A3(\SB2_2_3/i0_4 ), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_3/Component_Function_4/N2  ( .A1(\SB2_2_3/i3[0] ), .A2(
        \SB2_2_3/i0_0 ), .A3(\SB2_2_3/i1_7 ), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_3/Component_Function_4/N1  ( .A1(\SB2_2_3/i0[9] ), .A2(
        \SB2_2_3/i0_0 ), .A3(\SB2_2_3/i0[8] ), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_2/N4  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0_0 ), .A3(\SB2_2_4/i0_4 ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_4/Component_Function_2/N2  ( .A1(\SB2_2_4/i0_3 ), .A2(
        \SB2_2_4/i0[10] ), .A3(\SB2_2_4/i0[6] ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_4/Component_Function_2/N1  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0[10] ), .A3(\SB2_2_4/i1[9] ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_3/N3  ( .A1(\SB2_2_4/i1[9] ), .A2(
        \SB2_2_4/i1_7 ), .A3(\SB2_2_4/i0[10] ), .ZN(
        \SB2_2_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_4/Component_Function_3/N1  ( .A1(\SB2_2_4/i1[9] ), .A2(
        \SB2_2_4/i0_3 ), .A3(\SB2_2_4/i0[6] ), .ZN(
        \SB2_2_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_4/N4  ( .A1(\SB2_2_4/i1[9] ), .A2(
        \SB2_2_4/i1_5 ), .A3(\SB2_2_4/i0_4 ), .ZN(
        \SB2_2_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_4/Component_Function_4/N2  ( .A1(\SB2_2_4/i3[0] ), .A2(
        \SB2_2_4/i0_0 ), .A3(\SB2_2_4/i1_7 ), .ZN(
        \SB2_2_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_4/Component_Function_4/N1  ( .A1(\SB2_2_4/i0[9] ), .A2(
        \SB2_2_4/i0_0 ), .A3(\SB2_2_4/i0[8] ), .ZN(
        \SB2_2_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_2/N2  ( .A1(\SB2_2_5/i0_3 ), .A2(
        \SB2_2_5/i0[10] ), .A3(\SB2_2_5/i0[6] ), .ZN(
        \SB2_2_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_5/Component_Function_2/N1  ( .A1(\SB2_2_5/i1_5 ), .A2(
        \SB2_2_5/i0[10] ), .A3(\SB2_2_5/i1[9] ), .ZN(
        \SB2_2_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_3/N3  ( .A1(\SB2_2_5/i1[9] ), .A2(
        \SB2_2_5/i1_7 ), .A3(\SB2_2_5/i0[10] ), .ZN(
        \SB2_2_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_5/Component_Function_3/N1  ( .A1(\SB2_2_5/i1[9] ), .A2(
        \SB2_2_5/i0_3 ), .A3(\SB2_2_5/i0[6] ), .ZN(
        \SB2_2_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_4/N3  ( .A1(\SB2_2_5/i0[9] ), .A2(
        \SB2_2_5/i0[10] ), .A3(\SB2_2_5/i0_3 ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_5/Component_Function_4/N2  ( .A1(\SB2_2_5/i3[0] ), .A2(
        \SB2_2_5/i0_0 ), .A3(\SB2_2_5/i1_7 ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_5/Component_Function_4/N1  ( .A1(\SB2_2_5/i0[9] ), .A2(
        \SB2_2_5/i0_0 ), .A3(\SB2_2_5/i0[8] ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_2/N2  ( .A1(\SB2_2_6/i0_3 ), .A2(
        \SB2_2_6/i0[10] ), .A3(\SB2_2_6/i0[6] ), .ZN(
        \SB2_2_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_6/Component_Function_3/N3  ( .A1(\SB2_2_6/i1[9] ), .A2(
        \SB2_2_6/i1_7 ), .A3(\SB2_2_6/i0[10] ), .ZN(
        \SB2_2_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_6/Component_Function_3/N2  ( .A1(\SB2_2_6/i0_0 ), .A2(
        \SB2_2_6/i0_3 ), .A3(\SB2_2_6/i0_4 ), .ZN(
        \SB2_2_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_6/Component_Function_3/N1  ( .A1(\SB2_2_6/i1[9] ), .A2(
        \SB2_2_6/i0_3 ), .A3(\SB2_2_6/i0[6] ), .ZN(
        \SB2_2_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_4/N3  ( .A1(\SB2_2_6/i0[9] ), .A2(
        \SB2_2_6/i0[10] ), .A3(\SB2_2_6/i0_3 ), .ZN(
        \SB2_2_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_6/Component_Function_4/N2  ( .A1(\SB2_2_6/i3[0] ), .A2(
        \SB2_2_6/i0_0 ), .A3(\SB2_2_6/i1_7 ), .ZN(
        \SB2_2_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_6/Component_Function_4/N1  ( .A1(\SB2_2_6/i0[9] ), .A2(
        \SB2_2_6/i0_0 ), .A3(\SB2_2_6/i0[8] ), .ZN(
        \SB2_2_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_7/Component_Function_2/N2  ( .A1(\SB2_2_7/i0_3 ), .A2(
        \SB2_2_7/i0[10] ), .A3(\SB2_2_7/i0[6] ), .ZN(
        \SB2_2_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_7/Component_Function_2/N1  ( .A1(\SB2_2_7/i1_5 ), .A2(
        \SB2_2_7/i0[10] ), .A3(\SB2_2_7/i1[9] ), .ZN(
        \SB2_2_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_7/Component_Function_3/N3  ( .A1(\SB2_2_7/i1[9] ), .A2(
        \SB2_2_7/i1_7 ), .A3(\SB2_2_7/i0[10] ), .ZN(
        \SB2_2_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_7/Component_Function_4/N4  ( .A1(\SB2_2_7/i1[9] ), .A2(
        \SB2_2_7/i1_5 ), .A3(\SB2_2_7/i0_4 ), .ZN(
        \SB2_2_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_7/Component_Function_4/N2  ( .A1(\SB2_2_7/i3[0] ), .A2(
        \SB2_2_7/i0_0 ), .A3(\SB2_2_7/i1_7 ), .ZN(
        \SB2_2_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_7/Component_Function_4/N1  ( .A1(\SB2_2_7/i0[9] ), .A2(
        \SB2_2_7/i0_0 ), .A3(\SB2_2_7/i0[8] ), .ZN(
        \SB2_2_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_8/Component_Function_2/N2  ( .A1(\SB2_2_8/i0_3 ), .A2(
        \SB2_2_8/i0[10] ), .A3(\SB2_2_8/i0[6] ), .ZN(
        \SB2_2_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_8/Component_Function_3/N2  ( .A1(\SB2_2_8/i0_0 ), .A2(
        \SB2_2_8/i0_3 ), .A3(\SB2_2_8/i0_4 ), .ZN(
        \SB2_2_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_8/Component_Function_4/N3  ( .A1(\SB2_2_8/i0[9] ), .A2(
        \SB2_2_8/i0[10] ), .A3(\SB2_2_8/i0_3 ), .ZN(
        \SB2_2_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_8/Component_Function_4/N2  ( .A1(\SB2_2_8/i3[0] ), .A2(
        \SB2_2_8/i0_0 ), .A3(\SB2_2_8/i1_7 ), .ZN(
        \SB2_2_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_8/Component_Function_4/N1  ( .A1(\SB2_2_8/i0[9] ), .A2(
        \SB2_2_8/i0_0 ), .A3(\SB2_2_8/i0[8] ), .ZN(
        \SB2_2_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_2/N2  ( .A1(\SB2_2_9/i0_3 ), .A2(
        \SB2_2_9/i0[10] ), .A3(\SB2_2_9/i0[6] ), .ZN(
        \SB2_2_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_9/Component_Function_3/N4  ( .A1(\SB2_2_9/i1_5 ), .A2(
        \SB2_2_9/i0[8] ), .A3(\SB2_2_9/i3[0] ), .ZN(
        \SB2_2_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_9/Component_Function_3/N3  ( .A1(\SB2_2_9/i1[9] ), .A2(
        \SB2_2_9/i1_7 ), .A3(\SB2_2_9/i0[10] ), .ZN(
        \SB2_2_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_9/Component_Function_3/N1  ( .A1(\SB2_2_9/i0_3 ), .A2(
        \SB2_2_9/i1[9] ), .A3(\SB2_2_9/i0[6] ), .ZN(
        \SB2_2_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_4/N2  ( .A1(\SB2_2_9/i3[0] ), .A2(
        \SB2_2_9/i0_0 ), .A3(\SB2_2_9/i1_7 ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_9/Component_Function_4/N1  ( .A1(\SB2_2_9/i0[9] ), .A2(
        \SB2_2_9/i0_0 ), .A3(\SB2_2_9/i0[8] ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_10/Component_Function_2/N2  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i0[10] ), .A3(\SB2_2_10/i0[6] ), .ZN(
        \SB2_2_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_10/Component_Function_3/N3  ( .A1(\SB2_2_10/i1[9] ), .A2(
        \SB2_2_10/i1_7 ), .A3(\SB2_2_10/i0[10] ), .ZN(
        \SB2_2_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_10/Component_Function_3/N2  ( .A1(\SB2_2_10/i0_0 ), .A2(
        \SB2_2_10/i0_3 ), .A3(\SB2_2_10/i0_4 ), .ZN(
        \SB2_2_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_10/Component_Function_4/N3  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i0[10] ), .A3(\SB2_2_10/i0[9] ), .ZN(
        \SB2_2_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_10/Component_Function_4/N1  ( .A1(\SB2_2_10/i0[9] ), .A2(
        \SB2_2_10/i0_0 ), .A3(\SB2_2_10/i0[8] ), .ZN(
        \SB2_2_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_2/N2  ( .A1(\SB2_2_11/i0_3 ), .A2(
        \SB2_2_11/i0[10] ), .A3(\SB2_2_11/i0[6] ), .ZN(
        \SB2_2_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_11/Component_Function_2/N1  ( .A1(\SB2_2_11/i1_5 ), .A2(
        \SB2_2_11/i0[10] ), .A3(\SB2_2_11/i1[9] ), .ZN(
        \SB2_2_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_3/N3  ( .A1(\SB2_2_11/i1[9] ), .A2(
        \SB2_2_11/i1_7 ), .A3(\SB2_2_11/i0[10] ), .ZN(
        \SB2_2_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_11/Component_Function_3/N2  ( .A1(\SB2_2_11/i0_0 ), .A2(
        \SB2_2_11/i0_3 ), .A3(\SB2_2_11/i0_4 ), .ZN(
        \SB2_2_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N3  ( .A1(\SB2_2_11/i0[9] ), .A2(
        \SB2_2_11/i0[10] ), .A3(\SB2_2_11/i0_3 ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N2  ( .A1(\SB2_2_11/i3[0] ), .A2(
        \SB2_2_11/i0_0 ), .A3(\SB2_2_11/i1_7 ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N1  ( .A1(\SB2_2_11/i0[9] ), .A2(
        \SB2_2_11/i0_0 ), .A3(\SB2_2_11/i0[8] ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_2/N2  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i0[10] ), .A3(\SB2_2_12/i0[6] ), .ZN(
        \SB2_2_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_12/Component_Function_3/N3  ( .A1(\SB2_2_12/i1[9] ), .A2(
        \SB2_2_12/i1_7 ), .A3(\SB2_2_12/i0[10] ), .ZN(
        \SB2_2_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_12/Component_Function_3/N1  ( .A1(\SB2_2_12/i1[9] ), .A2(
        \SB2_2_12/i0_3 ), .A3(\SB2_2_12/i0[6] ), .ZN(
        \SB2_2_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_4/N2  ( .A1(\SB2_2_12/i3[0] ), .A2(
        \SB2_2_12/i0_0 ), .A3(\SB2_2_12/i1_7 ), .ZN(
        \SB2_2_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_12/Component_Function_4/N1  ( .A1(\SB2_2_12/i0[8] ), .A2(
        \SB2_2_12/i0_0 ), .A3(\SB2_2_12/i0[9] ), .ZN(
        \SB2_2_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_2/N4  ( .A1(\SB2_2_13/i1_5 ), .A2(
        \SB2_2_13/i0_0 ), .A3(\SB2_2_13/i0_4 ), .ZN(
        \SB2_2_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_13/Component_Function_2/N2  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i0[10] ), .A3(\SB2_2_13/i0[6] ), .ZN(
        \SB2_2_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_13/Component_Function_2/N1  ( .A1(\SB2_2_13/i1_5 ), .A2(
        \SB2_2_13/i0[10] ), .A3(\SB2_2_13/i1[9] ), .ZN(
        \SB2_2_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_3/N4  ( .A1(\SB2_2_13/i1_5 ), .A2(
        \SB2_2_13/i0[8] ), .A3(\SB2_2_13/i3[0] ), .ZN(
        \SB2_2_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_13/Component_Function_3/N3  ( .A1(\SB2_2_13/i1[9] ), .A2(
        \SB2_2_13/i1_7 ), .A3(\SB2_2_13/i0[10] ), .ZN(
        \SB2_2_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_13/Component_Function_3/N1  ( .A1(\SB2_2_13/i1[9] ), .A2(
        \SB2_2_13/i0_3 ), .A3(\SB2_2_13/i0[6] ), .ZN(
        \SB2_2_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_4/N4  ( .A1(\SB2_2_13/i1[9] ), .A2(
        \SB2_2_13/i1_5 ), .A3(\SB2_2_13/i0_4 ), .ZN(
        \SB2_2_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_13/Component_Function_4/N1  ( .A1(\SB2_2_13/i0[9] ), .A2(
        \SB2_2_13/i0_0 ), .A3(\SB2_2_13/i0[8] ), .ZN(
        \SB2_2_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_2/N2  ( .A1(\SB2_2_14/i0_3 ), .A2(
        \SB2_2_14/i0[10] ), .A3(\SB2_2_14/i0[6] ), .ZN(
        \SB2_2_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_14/Component_Function_2/N1  ( .A1(\SB2_2_14/i1_5 ), .A2(
        \SB2_2_14/i0[10] ), .A3(\SB2_2_14/i1[9] ), .ZN(
        \SB2_2_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_3/N3  ( .A1(\SB2_2_14/i1[9] ), .A2(
        \SB2_2_14/i1_7 ), .A3(\SB2_2_14/i0[10] ), .ZN(
        \SB2_2_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_14/Component_Function_3/N1  ( .A1(\SB2_2_14/i1[9] ), .A2(
        \SB2_2_14/i0_3 ), .A3(\SB2_2_14/i0[6] ), .ZN(
        \SB2_2_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_4/N3  ( .A1(\SB2_2_14/i0[9] ), .A2(
        \SB2_2_14/i0[10] ), .A3(\SB2_2_14/i0_3 ), .ZN(
        \SB2_2_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_14/Component_Function_4/N2  ( .A1(\SB2_2_14/i3[0] ), .A2(
        \SB2_2_14/i0_0 ), .A3(\SB2_2_14/i1_7 ), .ZN(
        \SB2_2_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_14/Component_Function_4/N1  ( .A1(\SB2_2_14/i0[9] ), .A2(
        \SB2_2_14/i0_0 ), .A3(\SB2_2_14/i0[8] ), .ZN(
        \SB2_2_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_15/Component_Function_2/N2  ( .A1(\SB2_2_15/i0_3 ), .A2(
        \SB2_2_15/i0[10] ), .A3(\SB2_2_15/i0[6] ), .ZN(
        \SB2_2_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_15/Component_Function_3/N3  ( .A1(\SB2_2_15/i1[9] ), .A2(
        \SB2_2_15/i1_7 ), .A3(\SB2_2_15/i0[10] ), .ZN(
        \SB2_2_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_15/Component_Function_3/N2  ( .A1(\SB2_2_15/i0_0 ), .A2(
        \SB2_2_15/i0_3 ), .A3(\SB2_2_15/i0_4 ), .ZN(
        \SB2_2_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_15/Component_Function_3/N1  ( .A1(\SB2_2_15/i1[9] ), .A2(
        \SB2_2_15/i0_3 ), .A3(\SB2_2_15/i0[6] ), .ZN(
        \SB2_2_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_15/Component_Function_4/N2  ( .A1(\SB2_2_15/i3[0] ), .A2(
        \SB2_2_15/i0_0 ), .A3(\SB2_2_15/i1_7 ), .ZN(
        \SB2_2_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_15/Component_Function_4/N1  ( .A1(\SB2_2_15/i0[9] ), .A2(
        \SB2_2_15/i0_0 ), .A3(\SB2_2_15/i0[8] ), .ZN(
        \SB2_2_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_2/N4  ( .A1(\SB2_2_16/i1_5 ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i0_4 ), .ZN(
        \SB2_2_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_16/Component_Function_2/N2  ( .A1(\SB2_2_16/i0_3 ), .A2(
        \SB2_2_16/i0[10] ), .A3(\SB2_2_16/i0[6] ), .ZN(
        \SB2_2_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_16/Component_Function_2/N1  ( .A1(\SB2_2_16/i1_5 ), .A2(
        \SB2_2_16/i0[10] ), .A3(\SB2_2_16/i1[9] ), .ZN(
        \SB2_2_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_3/N3  ( .A1(\SB2_2_16/i1[9] ), .A2(
        \SB2_2_16/i1_7 ), .A3(\SB2_2_16/i0[10] ), .ZN(
        \SB2_2_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_16/Component_Function_3/N1  ( .A1(\SB2_2_16/i1[9] ), .A2(
        \SB2_2_16/i0_3 ), .A3(\SB2_2_16/i0[6] ), .ZN(
        \SB2_2_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N4  ( .A1(\SB2_2_16/i1[9] ), .A2(
        \SB2_2_16/i1_5 ), .A3(\SB2_2_16/i0_4 ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N2  ( .A1(\SB2_2_16/i3[0] ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i1_7 ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N1  ( .A1(\SB2_2_16/i0[9] ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i0[8] ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_2/N2  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i0[10] ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_17/Component_Function_2/N1  ( .A1(\SB2_2_17/i1_5 ), .A2(
        \SB2_2_17/i0[10] ), .A3(\SB2_2_17/i1[9] ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_3/N3  ( .A1(\SB2_2_17/i1[9] ), .A2(
        \SB2_2_17/i1_7 ), .A3(\SB2_2_17/i0[10] ), .ZN(
        \SB2_2_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_17/Component_Function_3/N2  ( .A1(\SB2_2_17/i0_0 ), .A2(
        \SB2_2_17/i0_3 ), .A3(\SB2_2_17/i0_4 ), .ZN(
        \SB2_2_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_17/Component_Function_3/N1  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i1[9] ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_4/N3  ( .A1(\SB2_2_17/i0[9] ), .A2(
        \SB2_2_17/i0[10] ), .A3(\SB2_2_17/i0_3 ), .ZN(
        \SB2_2_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_17/Component_Function_4/N2  ( .A1(\SB2_2_17/i3[0] ), .A2(
        \SB2_2_17/i0_0 ), .A3(\SB2_2_17/i1_7 ), .ZN(
        \SB2_2_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_17/Component_Function_4/N1  ( .A1(\SB2_2_17/i0[9] ), .A2(
        \SB2_2_17/i0_0 ), .A3(\SB2_2_17/i0[8] ), .ZN(
        \SB2_2_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_2/N3  ( .A1(\SB2_2_18/i0_3 ), .A2(
        \SB2_2_18/i0[8] ), .A3(\SB2_2_18/i0[9] ), .ZN(
        \SB2_2_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_18/Component_Function_2/N2  ( .A1(\SB2_2_18/i0_3 ), .A2(
        \SB2_2_18/i0[10] ), .A3(\SB2_2_18/i0[6] ), .ZN(
        \SB2_2_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_18/Component_Function_2/N1  ( .A1(\SB2_2_18/i1_5 ), .A2(
        \SB2_2_18/i0[10] ), .A3(\SB2_2_18/i1[9] ), .ZN(
        \SB2_2_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_3/N3  ( .A1(\SB2_2_18/i1[9] ), .A2(
        \SB2_2_18/i1_7 ), .A3(\SB2_2_18/i0[10] ), .ZN(
        \SB2_2_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_18/Component_Function_3/N2  ( .A1(\SB2_2_18/i0_0 ), .A2(
        \SB2_2_18/i0_3 ), .A3(\SB2_2_18/i0_4 ), .ZN(
        \SB2_2_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_18/Component_Function_4/N3  ( .A1(\SB2_2_18/i0[9] ), .A2(
        \SB2_2_18/i0[10] ), .A3(\SB2_2_18/i0_3 ), .ZN(
        \SB2_2_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_18/Component_Function_4/N2  ( .A1(\SB2_2_18/i3[0] ), .A2(
        \SB2_2_18/i0_0 ), .A3(\SB2_2_18/i1_7 ), .ZN(
        \SB2_2_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_18/Component_Function_4/N1  ( .A1(\SB2_2_18/i0[9] ), .A2(
        \SB2_2_18/i0_0 ), .A3(\SB2_2_18/i0[8] ), .ZN(
        \SB2_2_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_2/N4  ( .A1(\SB2_2_19/i1_5 ), .A2(
        \SB2_2_19/i0_0 ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_19/Component_Function_2/N2  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i0[10] ), .A3(\SB2_2_19/i0[6] ), .ZN(
        \SB2_2_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_19/Component_Function_2/N1  ( .A1(\SB2_2_19/i1_5 ), .A2(
        \SB2_2_19/i0[10] ), .A3(\SB2_2_19/i1[9] ), .ZN(
        \SB2_2_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_3/N3  ( .A1(\SB2_2_19/i1[9] ), .A2(
        \SB2_2_19/i1_7 ), .A3(\SB2_2_19/i0[10] ), .ZN(
        \SB2_2_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_19/Component_Function_3/N1  ( .A1(\SB2_2_19/i1[9] ), .A2(
        \SB2_2_19/i0_3 ), .A3(\SB2_2_19/i0[6] ), .ZN(
        \SB2_2_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_4/N4  ( .A1(\SB2_2_19/i1[9] ), .A2(
        \SB2_2_19/i1_5 ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_19/Component_Function_4/N2  ( .A1(\SB2_2_19/i3[0] ), .A2(
        \SB2_2_19/i0_0 ), .A3(\SB2_2_19/i1_7 ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_19/Component_Function_4/N1  ( .A1(\SB2_2_19/i0[9] ), .A2(
        \SB2_2_19/i0_0 ), .A3(\SB2_2_19/i0[8] ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_2/N2  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i0[10] ), .A3(\SB2_2_20/i0[6] ), .ZN(
        \SB2_2_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_2/N1  ( .A1(\SB2_2_20/i1_5 ), .A2(
        \SB2_2_20/i0[10] ), .A3(\SB2_2_20/i1[9] ), .ZN(
        \SB2_2_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_3/N3  ( .A1(\SB2_2_20/i1[9] ), .A2(
        \SB2_2_20/i1_7 ), .A3(\SB2_2_20/i0[10] ), .ZN(
        \SB2_2_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_20/Component_Function_3/N1  ( .A1(\SB2_2_20/i1[9] ), .A2(
        \SB2_2_20/i0_3 ), .A3(\SB2_2_20/i0[6] ), .ZN(
        \SB2_2_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N4  ( .A1(\SB2_2_20/i1[9] ), .A2(
        \SB2_2_20/i1_5 ), .A3(\SB2_2_20/i0_4 ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N2  ( .A1(\SB2_2_20/i3[0] ), .A2(
        \SB2_2_20/i0_0 ), .A3(\SB2_2_20/i1_7 ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N1  ( .A1(\SB2_2_20/i0[9] ), .A2(
        \SB2_2_20/i0_0 ), .A3(\SB2_2_20/i0[8] ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_2/N2  ( .A1(\SB2_2_21/i0_3 ), .A2(
        \SB2_2_21/i0[10] ), .A3(\SB2_2_21/i0[6] ), .ZN(
        \SB2_2_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_21/Component_Function_3/N3  ( .A1(\SB2_2_21/i1[9] ), .A2(
        \SB2_2_21/i1_7 ), .A3(\SB2_2_21/i0[10] ), .ZN(
        \SB2_2_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_21/Component_Function_3/N2  ( .A1(\SB2_2_21/i0_0 ), .A2(
        \SB2_2_21/i0_3 ), .A3(\SB2_2_21/i0_4 ), .ZN(
        \SB2_2_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_21/Component_Function_3/N1  ( .A1(\SB2_2_21/i1[9] ), .A2(
        \SB2_2_21/i0_3 ), .A3(\SB2_2_21/i0[6] ), .ZN(
        \SB2_2_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_4/N3  ( .A1(\SB2_2_21/i0[9] ), .A2(
        \SB2_2_21/i0[10] ), .A3(\SB2_2_21/i0_3 ), .ZN(
        \SB2_2_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_21/Component_Function_4/N2  ( .A1(\SB2_2_21/i3[0] ), .A2(
        \SB2_2_21/i0_0 ), .A3(\SB2_2_21/i1_7 ), .ZN(
        \SB2_2_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_21/Component_Function_4/N1  ( .A1(\SB2_2_21/i0[9] ), .A2(
        \SB2_2_21/i0_0 ), .A3(\SB2_2_21/i0[8] ), .ZN(
        \SB2_2_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_22/Component_Function_2/N4  ( .A1(\SB2_2_22/i1_5 ), .A2(
        \SB2_2_22/i0_0 ), .A3(\SB2_2_22/i0_4 ), .ZN(
        \SB2_2_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_22/Component_Function_2/N2  ( .A1(\SB2_2_22/i0_3 ), .A2(
        \SB2_2_22/i0[10] ), .A3(\SB2_2_22/i0[6] ), .ZN(
        \SB2_2_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_22/Component_Function_2/N1  ( .A1(\SB2_2_22/i1_5 ), .A2(
        \SB2_2_22/i0[10] ), .A3(\SB2_2_22/i1[9] ), .ZN(
        \SB2_2_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_22/Component_Function_3/N3  ( .A1(\SB2_2_22/i1[9] ), .A2(
        \SB2_2_22/i1_7 ), .A3(\SB2_2_22/i0[10] ), .ZN(
        \SB2_2_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_22/Component_Function_3/N1  ( .A1(\SB2_2_22/i1[9] ), .A2(
        \SB2_2_22/i0_3 ), .A3(\SB2_2_22/i0[6] ), .ZN(
        \SB2_2_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_22/Component_Function_4/N4  ( .A1(\SB2_2_22/i1[9] ), .A2(
        \SB2_2_22/i1_5 ), .A3(\SB2_2_22/i0_4 ), .ZN(
        \SB2_2_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_22/Component_Function_4/N2  ( .A1(\SB2_2_22/i3[0] ), .A2(
        \SB2_2_22/i0_0 ), .A3(\SB2_2_22/i1_7 ), .ZN(
        \SB2_2_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_22/Component_Function_4/N1  ( .A1(\SB2_2_22/i0[9] ), .A2(
        \SB2_2_22/i0_0 ), .A3(\SB2_2_22/i0[8] ), .ZN(
        \SB2_2_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_23/Component_Function_2/N4  ( .A1(\SB2_2_23/i1_5 ), .A2(
        \SB2_2_23/i0_0 ), .A3(\RI3[2][52] ), .ZN(
        \SB2_2_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_23/Component_Function_2/N2  ( .A1(\SB2_2_23/i0_3 ), .A2(
        \SB2_2_23/i0[10] ), .A3(\SB2_2_23/i0[6] ), .ZN(
        \SB2_2_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_23/Component_Function_3/N3  ( .A1(\SB2_2_23/i1[9] ), .A2(
        \SB2_2_23/i1_7 ), .A3(\SB2_2_23/i0[10] ), .ZN(
        \SB2_2_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_23/Component_Function_3/N2  ( .A1(\SB2_2_23/i0_0 ), .A2(
        \SB2_2_23/i0_3 ), .A3(\SB2_2_23/i0_4 ), .ZN(
        \SB2_2_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_23/Component_Function_4/N3  ( .A1(\SB2_2_23/i0[9] ), .A2(
        \SB2_2_23/i0[10] ), .A3(\SB2_2_23/i0_3 ), .ZN(
        \SB2_2_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_23/Component_Function_4/N2  ( .A1(\SB2_2_23/i3[0] ), .A2(
        \SB2_2_23/i0_0 ), .A3(\SB2_2_23/i1_7 ), .ZN(
        \SB2_2_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_23/Component_Function_4/N1  ( .A1(\RI3[2][48] ), .A2(
        \SB2_2_23/i0_0 ), .A3(\SB2_2_23/i0[8] ), .ZN(
        \SB2_2_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_2/N3  ( .A1(\SB2_2_24/i0_3 ), .A2(
        \SB2_2_24/i0[8] ), .A3(\SB2_2_24/i0[9] ), .ZN(
        \SB2_2_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_24/Component_Function_2/N2  ( .A1(\SB2_2_24/i0_3 ), .A2(
        \SB2_2_24/i0[10] ), .A3(\SB2_2_24/i0[6] ), .ZN(
        \SB2_2_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_24/Component_Function_3/N3  ( .A1(\SB2_2_24/i1[9] ), .A2(
        \SB2_2_24/i1_7 ), .A3(\SB2_2_24/i0[10] ), .ZN(
        \SB2_2_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_24/Component_Function_3/N2  ( .A1(\SB2_2_24/i0_0 ), .A2(
        \SB2_2_24/i0_3 ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_24/Component_Function_3/N1  ( .A1(\SB2_2_24/i1[9] ), .A2(
        \SB2_2_24/i0_3 ), .A3(\SB2_2_24/i0[6] ), .ZN(
        \SB2_2_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N4  ( .A1(\SB2_2_24/i1[9] ), .A2(
        \SB2_2_24/i1_5 ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N2  ( .A1(\SB2_2_24/i3[0] ), .A2(
        \SB2_2_24/i0_0 ), .A3(\SB2_2_24/i1_7 ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N1  ( .A1(\SB2_2_24/i0[9] ), .A2(
        \SB2_2_24/i0_0 ), .A3(\SB2_2_24/i0[8] ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_2/N2  ( .A1(\SB2_2_25/i0_3 ), .A2(
        \SB2_2_25/i0[10] ), .A3(\SB2_2_25/i0[6] ), .ZN(
        \SB2_2_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_25/Component_Function_2/N1  ( .A1(\SB2_2_25/i1_5 ), .A2(
        \SB2_2_25/i0[10] ), .A3(\SB2_2_25/i1[9] ), .ZN(
        \SB2_2_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_3/N3  ( .A1(\SB2_2_25/i1[9] ), .A2(
        \SB2_2_25/i1_7 ), .A3(\SB2_2_25/i0[10] ), .ZN(
        \SB2_2_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_25/Component_Function_3/N2  ( .A1(\SB2_2_25/i0_0 ), .A2(
        \SB2_2_25/i0_3 ), .A3(\SB2_2_25/i0_4 ), .ZN(
        \SB2_2_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_25/Component_Function_3/N1  ( .A1(\SB2_2_25/i1[9] ), .A2(
        \SB2_2_25/i0_3 ), .A3(\SB2_2_25/i0[6] ), .ZN(
        \SB2_2_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N3  ( .A1(\SB2_2_25/i0[9] ), .A2(
        \SB2_2_25/i0[10] ), .A3(\SB2_2_25/i0_3 ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N2  ( .A1(\SB2_2_25/i3[0] ), .A2(
        \SB2_2_25/i0_0 ), .A3(\SB2_2_25/i1_7 ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N1  ( .A1(\SB2_2_25/i0[9] ), .A2(
        \SB2_2_25/i0_0 ), .A3(\SB2_2_25/i0[8] ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_2/N2  ( .A1(\SB2_2_26/i0_3 ), .A2(
        \SB2_2_26/i0[10] ), .A3(\SB2_2_26/i0[6] ), .ZN(
        \SB2_2_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_26/Component_Function_3/N3  ( .A1(\SB2_2_26/i1[9] ), .A2(
        \SB2_2_26/i1_7 ), .A3(\SB2_2_26/i0[10] ), .ZN(
        \SB2_2_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_26/Component_Function_3/N2  ( .A1(\SB2_2_26/i0_0 ), .A2(
        \SB2_2_26/i0_3 ), .A3(\SB2_2_26/i0_4 ), .ZN(
        \SB2_2_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_26/Component_Function_4/N3  ( .A1(\SB2_2_26/i0[9] ), .A2(
        \SB2_2_26/i0[10] ), .A3(\SB2_2_26/i0_3 ), .ZN(
        \SB2_2_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_26/Component_Function_4/N2  ( .A1(\SB2_2_26/i3[0] ), .A2(
        \SB2_2_26/i0_0 ), .A3(\SB2_2_26/i1_7 ), .ZN(
        \SB2_2_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_26/Component_Function_4/N1  ( .A1(\SB2_2_26/i0[9] ), .A2(
        \SB2_2_26/i0_0 ), .A3(\SB2_2_26/i0[8] ), .ZN(
        \SB2_2_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_27/Component_Function_3/N3  ( .A1(\SB2_2_27/i1[9] ), .A2(
        \SB2_2_27/i1_7 ), .A3(\SB2_2_27/i0[10] ), .ZN(
        \SB2_2_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_27/Component_Function_3/N2  ( .A1(\SB2_2_27/i0_0 ), .A2(
        \SB2_2_27/i0_3 ), .A3(\SB2_2_27/i0_4 ), .ZN(
        \SB2_2_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_27/Component_Function_4/N3  ( .A1(\SB2_2_27/i0[9] ), .A2(
        \SB2_2_27/i0[10] ), .A3(\SB2_2_27/i0_3 ), .ZN(
        \SB2_2_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_27/Component_Function_4/N2  ( .A1(\SB2_2_27/i3[0] ), .A2(
        \SB2_2_27/i0_0 ), .A3(\SB2_2_27/i1_7 ), .ZN(
        \SB2_2_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_27/Component_Function_4/N1  ( .A1(\SB2_2_27/i0[9] ), .A2(
        \SB2_2_27/i0_0 ), .A3(\SB2_2_27/i0[8] ), .ZN(
        \SB2_2_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_2/N1  ( .A1(\SB2_2_28/i1_5 ), .A2(
        \SB2_2_28/i0[10] ), .A3(\SB2_2_28/i1[9] ), .ZN(
        \SB2_2_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_3/N3  ( .A1(\SB2_2_28/i1[9] ), .A2(
        \SB2_2_28/i1_7 ), .A3(\SB2_2_28/i0[10] ), .ZN(
        \SB2_2_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_28/Component_Function_3/N1  ( .A1(\SB2_2_28/i1[9] ), .A2(
        \SB2_2_28/i0_3 ), .A3(\SB2_2_28/i0[6] ), .ZN(
        \SB2_2_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_4/N4  ( .A1(\SB2_2_28/i1[9] ), .A2(
        \SB2_2_28/i1_5 ), .A3(\SB2_2_28/i0_4 ), .ZN(
        \SB2_2_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_28/Component_Function_4/N1  ( .A1(\SB2_2_28/i0[9] ), .A2(
        \SB2_2_28/i0_0 ), .A3(\SB2_2_28/i0[8] ), .ZN(
        \SB2_2_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_2/N2  ( .A1(\SB2_2_29/i0_3 ), .A2(
        \SB2_2_29/i0[10] ), .A3(\SB2_2_29/i0[6] ), .ZN(
        \SB2_2_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_29/Component_Function_2/N1  ( .A1(\SB2_2_29/i1_5 ), .A2(
        \SB2_2_29/i0[10] ), .A3(\SB2_2_29/i1[9] ), .ZN(
        \SB2_2_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_3/N4  ( .A1(\SB2_2_29/i1_5 ), .A2(
        \SB2_2_29/i0[8] ), .A3(\SB2_2_29/i3[0] ), .ZN(
        \SB2_2_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_29/Component_Function_3/N2  ( .A1(\SB2_2_29/i0_0 ), .A2(
        \SB2_2_29/i0_3 ), .A3(\SB2_2_29/i0_4 ), .ZN(
        \SB2_2_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_29/Component_Function_3/N1  ( .A1(\SB2_2_29/i1[9] ), .A2(
        \SB2_2_29/i0_3 ), .A3(\SB2_2_29/i0[6] ), .ZN(
        \SB2_2_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_4/N2  ( .A1(\SB2_2_29/i3[0] ), .A2(
        \SB2_2_29/i0_0 ), .A3(\SB2_2_29/i1_7 ), .ZN(
        \SB2_2_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_29/Component_Function_4/N1  ( .A1(\SB2_2_29/i0[9] ), .A2(
        \SB2_2_29/i0_0 ), .A3(\SB2_2_29/i0[8] ), .ZN(
        \SB2_2_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_2/N4  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0_0 ), .A3(\SB2_2_30/i0_4 ), .ZN(
        \SB2_2_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_30/Component_Function_2/N2  ( .A1(\SB2_2_30/i0_3 ), .A2(
        \SB2_2_30/i0[10] ), .A3(\SB2_2_30/i0[6] ), .ZN(
        \SB2_2_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_30/Component_Function_2/N1  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0[10] ), .A3(n2118), .ZN(
        \SB2_2_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_3/N3  ( .A1(n2118), .A2(
        \SB2_2_30/i1_7 ), .A3(\SB2_2_30/i0[10] ), .ZN(
        \SB2_2_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_30/Component_Function_3/N1  ( .A1(n2118), .A2(
        \SB2_2_30/i0_3 ), .A3(\SB2_2_30/i0[6] ), .ZN(
        \SB2_2_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N4  ( .A1(n2118), .A2(
        \SB2_2_30/i1_5 ), .A3(\SB2_2_30/i0_4 ), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N2  ( .A1(\SB2_2_30/i3[0] ), .A2(
        \SB2_2_30/i0_0 ), .A3(\SB2_2_30/i1_7 ), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N1  ( .A1(\SB2_2_30/i0[9] ), .A2(
        \SB2_2_30/i0_0 ), .A3(\SB2_2_30/i0[8] ), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_31/Component_Function_2/N2  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i0[10] ), .A3(\SB2_2_31/i0[6] ), .ZN(
        \SB2_2_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_31/Component_Function_2/N1  ( .A1(\SB2_2_31/i1_5 ), .A2(
        \SB2_2_31/i0[10] ), .A3(\SB2_2_31/i1[9] ), .ZN(
        \SB2_2_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_31/Component_Function_3/N3  ( .A1(\SB2_2_31/i1[9] ), .A2(
        \SB2_2_31/i1_7 ), .A3(\SB2_2_31/i0[10] ), .ZN(
        \SB2_2_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_31/Component_Function_3/N2  ( .A1(\SB2_2_31/i0_0 ), .A2(
        \SB2_2_31/i0_3 ), .A3(\SB2_2_31/i0_4 ), .ZN(
        \SB2_2_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_31/Component_Function_3/N1  ( .A1(\SB2_2_31/i1[9] ), .A2(
        \SB2_2_31/i0_3 ), .A3(\SB2_2_31/i0[6] ), .ZN(
        \SB2_2_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N4  ( .A1(\SB2_2_31/i1[9] ), .A2(
        \SB2_2_31/i1_5 ), .A3(\SB2_2_31/i0_4 ), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N2  ( .A1(\SB2_2_31/i3[0] ), .A2(
        \SB2_2_31/i0_0 ), .A3(\SB2_2_31/i1_7 ), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N1  ( .A1(\SB2_2_31/i0[9] ), .A2(
        \SB2_2_31/i0_0 ), .A3(\SB2_2_31/i0[8] ), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_2/N2  ( .A1(n809), .A2(\SB1_3_0/i0[10] ), .A3(\SB1_3_0/i0[6] ), .ZN(\SB1_3_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_0/Component_Function_2/N1  ( .A1(\SB1_3_0/i1_5 ), .A2(
        \SB1_3_0/i0[10] ), .A3(\SB1_3_0/i1[9] ), .ZN(
        \SB1_3_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_3/N4  ( .A1(\SB1_3_0/i1_5 ), .A2(
        \SB1_3_0/i0[8] ), .A3(\SB1_3_0/i3[0] ), .ZN(
        \SB1_3_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_0/Component_Function_3/N3  ( .A1(\SB1_3_0/i0[10] ), .A2(
        \SB1_3_0/i1_7 ), .A3(\SB1_3_0/i1[9] ), .ZN(
        \SB1_3_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_0/Component_Function_3/N2  ( .A1(\SB1_3_0/i0_0 ), .A2(n809), 
        .A3(\SB1_3_0/i0_4 ), .ZN(\SB1_3_0/Component_Function_3/NAND4_in[1] )
         );
  NAND3_X1 \SB1_3_0/Component_Function_3/N1  ( .A1(\SB1_3_0/i1[9] ), .A2(n809), 
        .A3(\SB1_3_0/i0[6] ), .ZN(\SB1_3_0/Component_Function_3/NAND4_in[0] )
         );
  NAND3_X1 \SB1_3_0/Component_Function_4/N4  ( .A1(\SB1_3_0/i1[9] ), .A2(
        \SB1_3_0/i1_5 ), .A3(\SB1_3_0/i0_4 ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N3  ( .A1(\SB1_3_0/i0[9] ), .A2(
        \SB1_3_0/i0[10] ), .A3(n809), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N2  ( .A1(\SB1_3_0/i3[0] ), .A2(
        \SB1_3_0/i0_0 ), .A3(\SB1_3_0/i1_7 ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N1  ( .A1(\SB1_3_0/i0[9] ), .A2(
        \SB1_3_0/i0_0 ), .A3(\SB1_3_0/i0[8] ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_2/N2  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i0[10] ), .A3(\SB1_3_1/i0[6] ), .ZN(
        \SB1_3_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_1/Component_Function_2/N1  ( .A1(\SB1_3_1/i1_5 ), .A2(
        \SB1_3_1/i0[10] ), .A3(\SB1_3_1/i1[9] ), .ZN(
        \SB1_3_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_3/N4  ( .A1(\SB1_3_1/i1_5 ), .A2(
        \SB1_3_1/i0[8] ), .A3(\SB1_3_1/i3[0] ), .ZN(
        \SB1_3_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_1/Component_Function_3/N2  ( .A1(\SB1_3_1/i0_0 ), .A2(
        \SB1_3_1/i0_3 ), .A3(\SB1_3_1/i0_4 ), .ZN(
        \SB1_3_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_1/Component_Function_3/N1  ( .A1(\SB1_3_1/i1[9] ), .A2(
        \SB1_3_1/i0_3 ), .A3(\SB1_3_1/i0[6] ), .ZN(
        \SB1_3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_4/N4  ( .A1(\SB1_3_1/i1[9] ), .A2(
        \SB1_3_1/i1_5 ), .A3(\SB1_3_1/i0_4 ), .ZN(
        \SB1_3_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_1/Component_Function_4/N2  ( .A1(\SB1_3_1/i3[0] ), .A2(
        \SB1_3_1/i0_0 ), .A3(\SB1_3_1/i1_7 ), .ZN(
        \SB1_3_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_1/Component_Function_4/N1  ( .A1(\SB1_3_1/i0[9] ), .A2(
        \SB1_3_1/i0_0 ), .A3(\SB1_3_1/i0[8] ), .ZN(
        \SB1_3_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_2/N2  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i0[10] ), .A3(\SB1_3_2/i0[6] ), .ZN(
        \SB1_3_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_3/N4  ( .A1(\SB1_3_2/i1_5 ), .A2(
        \SB1_3_2/i0[8] ), .A3(\SB1_3_2/i3[0] ), .ZN(
        \SB1_3_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_2/Component_Function_3/N2  ( .A1(\SB1_3_2/i0_4 ), .A2(
        \SB1_3_2/i0_3 ), .A3(\SB1_3_2/i0_0 ), .ZN(
        \SB1_3_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_3/N1  ( .A1(\SB1_3_2/i1[9] ), .A2(
        \SB1_3_2/i0_3 ), .A3(\SB1_3_2/i0[6] ), .ZN(
        \SB1_3_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_4/N4  ( .A1(\SB1_3_2/i1[9] ), .A2(
        \SB1_3_2/i1_5 ), .A3(\SB1_3_2/i0_4 ), .ZN(
        \SB1_3_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_2/Component_Function_4/N2  ( .A1(\SB1_3_2/i3[0] ), .A2(
        \SB1_3_2/i0_0 ), .A3(\SB1_3_2/i1_7 ), .ZN(
        \SB1_3_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_4/N1  ( .A1(\SB1_3_2/i0[9] ), .A2(
        \SB1_3_2/i0_0 ), .A3(\SB1_3_2/i0[8] ), .ZN(
        \SB1_3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_2/N3  ( .A1(\SB1_3_3/i0_3 ), .A2(
        \SB1_3_3/i0[8] ), .A3(\SB1_3_3/i0[9] ), .ZN(
        \SB1_3_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_3/Component_Function_2/N2  ( .A1(\SB1_3_3/i0_3 ), .A2(
        \SB1_3_3/i0[10] ), .A3(\SB1_3_3/i0[6] ), .ZN(
        \SB1_3_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_3/N4  ( .A1(\SB1_3_3/i1_5 ), .A2(
        \SB1_3_3/i0[8] ), .A3(\SB1_3_3/i3[0] ), .ZN(
        \SB1_3_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_3/Component_Function_3/N3  ( .A1(\SB1_3_3/i1[9] ), .A2(
        \SB1_3_3/i1_7 ), .A3(\SB1_3_3/i0[10] ), .ZN(
        \SB1_3_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_3/Component_Function_3/N2  ( .A1(\SB1_3_3/i0_0 ), .A2(
        \SB1_3_3/i0_3 ), .A3(\SB1_3_3/i0_4 ), .ZN(
        \SB1_3_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_3/N1  ( .A1(\SB1_3_3/i1[9] ), .A2(
        \SB1_3_3/i0_3 ), .A3(\SB1_3_3/i0[6] ), .ZN(
        \SB1_3_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N4  ( .A1(\SB1_3_3/i1[9] ), .A2(
        \SB1_3_3/i1_5 ), .A3(\SB1_3_3/i0_4 ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N2  ( .A1(\SB1_3_3/i3[0] ), .A2(
        \SB1_3_3/i0_0 ), .A3(\SB1_3_3/i1_7 ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N1  ( .A1(\SB1_3_3/i0[9] ), .A2(
        \SB1_3_3/i0_0 ), .A3(\SB1_3_3/i0[8] ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_2/N2  ( .A1(\SB1_3_4/i0_3 ), .A2(
        \SB1_3_4/i0[10] ), .A3(\SB1_3_4/i0[6] ), .ZN(
        \SB1_3_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_4/Component_Function_2/N1  ( .A1(\SB1_3_4/i1_5 ), .A2(
        \SB1_3_4/i0[10] ), .A3(\SB1_3_4/i1[9] ), .ZN(
        \SB1_3_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_3/N4  ( .A1(\SB1_3_4/i1_5 ), .A2(
        \SB1_3_4/i0[8] ), .A3(\SB1_3_4/i3[0] ), .ZN(
        \SB1_3_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_4/Component_Function_3/N3  ( .A1(\SB1_3_4/i1[9] ), .A2(
        \SB1_3_4/i1_7 ), .A3(\SB1_3_4/i0[10] ), .ZN(
        \SB1_3_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_4/Component_Function_3/N2  ( .A1(\SB1_3_4/i0_0 ), .A2(
        \SB1_3_4/i0_3 ), .A3(\SB1_3_4/i0_4 ), .ZN(
        \SB1_3_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_4/Component_Function_3/N1  ( .A1(\SB1_3_4/i1[9] ), .A2(
        \SB1_3_4/i0_3 ), .A3(\SB1_3_4/i0[6] ), .ZN(
        \SB1_3_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_4/N4  ( .A1(\SB1_3_4/i1[9] ), .A2(
        \SB1_3_4/i1_5 ), .A3(\SB1_3_4/i0_4 ), .ZN(
        \SB1_3_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_4/Component_Function_4/N2  ( .A1(\SB1_3_4/i3[0] ), .A2(
        \SB1_3_4/i0_0 ), .A3(\SB1_3_4/i1_7 ), .ZN(
        \SB1_3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_4/Component_Function_4/N1  ( .A1(\SB1_3_4/i0[9] ), .A2(
        \SB1_3_4/i0_0 ), .A3(\SB1_3_4/i0[8] ), .ZN(
        \SB1_3_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_2/N2  ( .A1(\SB1_3_5/i0_3 ), .A2(
        \SB1_3_5/i0[10] ), .A3(\SB1_3_5/i0[6] ), .ZN(
        \SB1_3_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_5/Component_Function_2/N1  ( .A1(\SB1_3_5/i1_5 ), .A2(
        \SB1_3_5/i0[10] ), .A3(\SB1_3_5/i1[9] ), .ZN(
        \SB1_3_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_3/N4  ( .A1(\SB1_3_5/i1_5 ), .A2(
        \SB1_3_5/i0[8] ), .A3(\SB1_3_5/i3[0] ), .ZN(
        \SB1_3_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_5/Component_Function_3/N3  ( .A1(\SB1_3_5/i0[10] ), .A2(
        \SB1_3_5/i1_7 ), .A3(\SB1_3_5/i1[9] ), .ZN(
        \SB1_3_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_5/Component_Function_3/N1  ( .A1(\SB1_3_5/i1[9] ), .A2(
        \SB1_3_5/i0_3 ), .A3(\SB1_3_5/i0[6] ), .ZN(
        \SB1_3_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N4  ( .A1(\SB1_3_5/i1[9] ), .A2(
        \SB1_3_5/i1_5 ), .A3(\SB1_3_5/i0_4 ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N2  ( .A1(\SB1_3_5/i3[0] ), .A2(
        \SB1_3_5/i0_0 ), .A3(\SB1_3_5/i1_7 ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N1  ( .A1(\SB1_3_5/i0[9] ), .A2(
        \SB1_3_5/i0_0 ), .A3(\SB1_3_5/i0[8] ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_2/N2  ( .A1(\SB1_3_6/i0_3 ), .A2(
        \SB1_3_6/i0[10] ), .A3(\SB1_3_6/i0[6] ), .ZN(
        \SB1_3_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_6/Component_Function_2/N1  ( .A1(\SB1_3_6/i1_5 ), .A2(
        \SB1_3_6/i0[10] ), .A3(\SB1_3_6/i1[9] ), .ZN(
        \SB1_3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_3/N4  ( .A1(\SB1_3_6/i1_5 ), .A2(
        \SB1_3_6/i0[8] ), .A3(\SB1_3_6/i3[0] ), .ZN(
        \SB1_3_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_6/Component_Function_3/N2  ( .A1(\SB1_3_6/i0_0 ), .A2(
        \SB1_3_6/i0_3 ), .A3(\SB1_3_6/i0_4 ), .ZN(
        \SB1_3_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_6/Component_Function_3/N1  ( .A1(\SB1_3_6/i1[9] ), .A2(
        \SB1_3_6/i0_3 ), .A3(\SB1_3_6/i0[6] ), .ZN(
        \SB1_3_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_4/N4  ( .A1(\SB1_3_6/i1[9] ), .A2(
        \SB1_3_6/i1_5 ), .A3(\SB1_3_6/i0_4 ), .ZN(
        \SB1_3_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_6/Component_Function_4/N3  ( .A1(\SB1_3_6/i0[9] ), .A2(
        \SB1_3_6/i0[10] ), .A3(\SB1_3_6/i0_3 ), .ZN(
        \SB1_3_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_6/Component_Function_4/N2  ( .A1(\SB1_3_6/i3[0] ), .A2(
        \SB1_3_6/i0_0 ), .A3(\SB1_3_6/i1_7 ), .ZN(
        \SB1_3_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_6/Component_Function_4/N1  ( .A1(\SB1_3_6/i0[9] ), .A2(
        \SB1_3_6/i0_0 ), .A3(\SB1_3_6/i0[8] ), .ZN(
        \SB1_3_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_2/N2  ( .A1(\SB1_3_7/i0_3 ), .A2(
        \SB1_3_7/i0[10] ), .A3(\SB1_3_7/i0[6] ), .ZN(
        \SB1_3_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_7/Component_Function_2/N1  ( .A1(\SB1_3_7/i1_5 ), .A2(
        \SB1_3_7/i0[10] ), .A3(\SB1_3_7/i1[9] ), .ZN(
        \SB1_3_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_3/N4  ( .A1(\SB1_3_7/i1_5 ), .A2(
        \SB1_3_7/i0[8] ), .A3(\SB1_3_7/i3[0] ), .ZN(
        \SB1_3_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_7/Component_Function_3/N1  ( .A1(\SB1_3_7/i1[9] ), .A2(
        \SB1_3_7/i0_3 ), .A3(\SB1_3_7/i0[6] ), .ZN(
        \SB1_3_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_4/N4  ( .A1(\SB1_3_7/i1[9] ), .A2(
        \SB1_3_7/i1_5 ), .A3(\SB1_3_7/i0_4 ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_7/Component_Function_4/N3  ( .A1(\SB1_3_7/i0[9] ), .A2(
        \SB1_3_7/i0[10] ), .A3(\SB1_3_7/i0_3 ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_7/Component_Function_4/N2  ( .A1(\SB1_3_7/i3[0] ), .A2(
        \SB1_3_7/i0_0 ), .A3(\SB1_3_7/i1_7 ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_7/Component_Function_4/N1  ( .A1(\SB1_3_7/i0[9] ), .A2(
        \SB1_3_7/i0_0 ), .A3(\SB1_3_7/i0[8] ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_2/N2  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i0[10] ), .A3(\SB1_3_8/i0[6] ), .ZN(
        \SB1_3_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_8/Component_Function_2/N1  ( .A1(\SB1_3_8/i1_5 ), .A2(
        \SB1_3_8/i0[10] ), .A3(\SB1_3_8/i1[9] ), .ZN(
        \SB1_3_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_3/N4  ( .A1(\SB1_3_8/i1_5 ), .A2(
        \SB1_3_8/i0[8] ), .A3(\SB1_3_8/i3[0] ), .ZN(
        \SB1_3_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_8/Component_Function_3/N3  ( .A1(\SB1_3_8/i1[9] ), .A2(
        \SB1_3_8/i1_7 ), .A3(\SB1_3_8/i0[10] ), .ZN(
        \SB1_3_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_8/Component_Function_3/N2  ( .A1(\SB1_3_8/i0_0 ), .A2(
        \SB1_3_8/i0_3 ), .A3(\SB1_3_8/i0_4 ), .ZN(
        \SB1_3_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_8/Component_Function_3/N1  ( .A1(\SB1_3_8/i1[9] ), .A2(
        \SB1_3_8/i0_3 ), .A3(\SB1_3_8/i0[6] ), .ZN(
        \SB1_3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_4/N4  ( .A1(\SB1_3_8/i1[9] ), .A2(
        \SB1_3_8/i1_5 ), .A3(\SB1_3_8/i0_4 ), .ZN(
        \SB1_3_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_8/Component_Function_4/N2  ( .A1(\SB1_3_8/i3[0] ), .A2(
        \SB1_3_8/i0_0 ), .A3(\SB1_3_8/i1_7 ), .ZN(
        \SB1_3_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_8/Component_Function_4/N1  ( .A1(\SB1_3_8/i0[9] ), .A2(
        \SB1_3_8/i0_0 ), .A3(\SB1_3_8/i0[8] ), .ZN(
        \SB1_3_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_2/N2  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i0[10] ), .A3(\SB1_3_9/i0[6] ), .ZN(
        \SB1_3_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_9/Component_Function_2/N1  ( .A1(\SB1_3_9/i1_5 ), .A2(
        \SB1_3_9/i0[10] ), .A3(\SB1_3_9/i1[9] ), .ZN(
        \SB1_3_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_3/N3  ( .A1(\SB1_3_9/i1[9] ), .A2(
        \SB1_3_9/i1_7 ), .A3(\SB1_3_9/i0[10] ), .ZN(
        \SB1_3_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_9/Component_Function_3/N2  ( .A1(\SB1_3_9/i0_0 ), .A2(
        \SB1_3_9/i0_3 ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N4  ( .A1(\SB1_3_9/i1[9] ), .A2(
        \SB1_3_9/i1_5 ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N3  ( .A1(\SB1_3_9/i0[9] ), .A2(
        \SB1_3_9/i0[10] ), .A3(\SB1_3_9/i0_3 ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N2  ( .A1(\SB1_3_9/i3[0] ), .A2(
        \SB1_3_9/i0_0 ), .A3(\SB1_3_9/i1_7 ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N1  ( .A1(\SB1_3_9/i0[9] ), .A2(
        \SB1_3_9/i0_0 ), .A3(\SB1_3_9/i0[8] ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_2/N3  ( .A1(\SB1_3_10/i0_3 ), .A2(
        \SB1_3_10/i0[8] ), .A3(\SB1_3_10/i0[9] ), .ZN(
        \SB1_3_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_10/Component_Function_2/N1  ( .A1(\SB1_3_10/i1_5 ), .A2(
        \SB1_3_10/i0[10] ), .A3(\SB1_3_10/i1[9] ), .ZN(
        \SB1_3_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_3/N4  ( .A1(\SB1_3_10/i1_5 ), .A2(
        \SB1_3_10/i0[8] ), .A3(\SB1_3_10/i3[0] ), .ZN(
        \SB1_3_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_10/Component_Function_3/N1  ( .A1(\SB1_3_10/i1[9] ), .A2(
        \SB1_3_10/i0_3 ), .A3(\SB1_3_10/i0[6] ), .ZN(
        \SB1_3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_4/N4  ( .A1(\SB1_3_10/i1[9] ), .A2(
        \SB1_3_10/i1_5 ), .A3(\SB1_3_10/i0_4 ), .ZN(
        \SB1_3_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_10/Component_Function_4/N2  ( .A1(\SB1_3_10/i3[0] ), .A2(
        \SB1_3_10/i0_0 ), .A3(\SB1_3_10/i1_7 ), .ZN(
        \SB1_3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_10/Component_Function_4/N1  ( .A1(\SB1_3_10/i0[9] ), .A2(
        \SB1_3_10/i0_0 ), .A3(\SB1_3_10/i0[8] ), .ZN(
        \SB1_3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_2/N2  ( .A1(n831), .A2(
        \SB1_3_11/i0[10] ), .A3(\SB1_3_11/i0[6] ), .ZN(
        \SB1_3_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_11/Component_Function_2/N1  ( .A1(\SB1_3_11/i1_5 ), .A2(
        \SB1_3_11/i0[10] ), .A3(\SB1_3_11/i1[9] ), .ZN(
        \SB1_3_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_3/N3  ( .A1(\SB1_3_11/i1[9] ), .A2(
        \SB1_3_11/i1_7 ), .A3(\SB1_3_11/i0[10] ), .ZN(
        \SB1_3_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_11/Component_Function_3/N2  ( .A1(\SB1_3_11/i0_0 ), .A2(
        \SB1_3_11/i0_3 ), .A3(\SB1_3_11/i0_4 ), .ZN(
        \SB1_3_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_11/Component_Function_3/N1  ( .A1(\SB1_3_11/i1[9] ), .A2(
        n831), .A3(\SB1_3_11/i0[6] ), .ZN(
        \SB1_3_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_4/N4  ( .A1(\SB1_3_11/i1[9] ), .A2(
        \SB1_3_11/i1_5 ), .A3(\SB1_3_11/i0_4 ), .ZN(
        \SB1_3_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_11/Component_Function_4/N2  ( .A1(\SB1_3_11/i3[0] ), .A2(
        \SB1_3_11/i0_0 ), .A3(\SB1_3_11/i1_7 ), .ZN(
        \SB1_3_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_11/Component_Function_4/N1  ( .A1(\SB1_3_11/i0[9] ), .A2(
        \SB1_3_11/i0_0 ), .A3(\SB1_3_11/i0[8] ), .ZN(
        \SB1_3_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_12/Component_Function_2/N2  ( .A1(\SB1_3_12/i0_3 ), .A2(
        \SB1_3_12/i0[10] ), .A3(\SB1_3_12/i0[6] ), .ZN(
        \SB1_3_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_12/Component_Function_2/N1  ( .A1(\SB1_3_12/i1_5 ), .A2(
        \SB1_3_12/i0[10] ), .A3(\SB1_3_12/i1[9] ), .ZN(
        \SB1_3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_12/Component_Function_3/N3  ( .A1(\SB1_3_12/i1[9] ), .A2(
        \SB1_3_12/i1_7 ), .A3(\SB1_3_12/i0[10] ), .ZN(
        \SB1_3_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_12/Component_Function_3/N2  ( .A1(\SB1_3_12/i0_0 ), .A2(
        \SB1_3_12/i0_3 ), .A3(\SB1_3_12/i0_4 ), .ZN(
        \SB1_3_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_12/Component_Function_4/N4  ( .A1(\SB1_3_12/i1[9] ), .A2(
        \SB1_3_12/i1_5 ), .A3(\SB1_3_12/i0_4 ), .ZN(
        \SB1_3_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_12/Component_Function_4/N3  ( .A1(\SB1_3_12/i0[9] ), .A2(
        \SB1_3_12/i0[10] ), .A3(\SB1_3_12/i0_3 ), .ZN(
        \SB1_3_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_12/Component_Function_4/N2  ( .A1(\SB1_3_12/i3[0] ), .A2(
        \SB1_3_12/i0_0 ), .A3(\SB1_3_12/i1_7 ), .ZN(
        \SB1_3_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_12/Component_Function_4/N1  ( .A1(\SB1_3_12/i0[9] ), .A2(
        \SB1_3_12/i0_0 ), .A3(\SB1_3_12/i0[8] ), .ZN(
        \SB1_3_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_2/N2  ( .A1(\SB1_3_13/i0_3 ), .A2(
        \SB1_3_13/i0[10] ), .A3(\SB1_3_13/i0[6] ), .ZN(
        \SB1_3_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_13/Component_Function_2/N1  ( .A1(\SB1_3_13/i1_5 ), .A2(
        \SB1_3_13/i0[10] ), .A3(\SB1_3_13/i1[9] ), .ZN(
        \SB1_3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_3/N4  ( .A1(\SB1_3_13/i1_5 ), .A2(
        \SB1_3_13/i0[8] ), .A3(\SB1_3_13/i3[0] ), .ZN(
        \SB1_3_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_13/Component_Function_3/N3  ( .A1(\SB1_3_13/i1[9] ), .A2(
        \SB1_3_13/i1_7 ), .A3(\SB1_3_13/i0[10] ), .ZN(
        \SB1_3_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_3/N1  ( .A1(\SB1_3_13/i1[9] ), .A2(
        \SB1_3_13/i0_3 ), .A3(\SB1_3_13/i0[6] ), .ZN(
        \SB1_3_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_4/N4  ( .A1(\SB1_3_13/i1[9] ), .A2(
        \SB1_3_13/i1_5 ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_13/Component_Function_4/N2  ( .A1(\SB1_3_13/i3[0] ), .A2(
        \SB1_3_13/i0_0 ), .A3(\SB1_3_13/i1_7 ), .ZN(
        \SB1_3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_13/Component_Function_4/N1  ( .A1(\SB1_3_13/i0[9] ), .A2(
        \SB1_3_13/i0_0 ), .A3(\SB1_3_13/i0[8] ), .ZN(
        \SB1_3_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_2/N4  ( .A1(\SB1_3_14/i1_5 ), .A2(
        \SB1_3_14/i0_0 ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_2/N2  ( .A1(\SB1_3_14/i0_3 ), .A2(
        \SB1_3_14/i0[10] ), .A3(\SB1_3_14/i0[6] ), .ZN(
        \SB1_3_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_14/Component_Function_2/N1  ( .A1(\SB1_3_14/i1_5 ), .A2(
        \SB1_3_14/i0[10] ), .A3(\SB1_3_14/i1[9] ), .ZN(
        \SB1_3_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_3/N4  ( .A1(\SB1_3_14/i1_5 ), .A2(
        \SB1_3_14/i0[8] ), .A3(\SB1_3_14/i3[0] ), .ZN(
        \SB1_3_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_3/N3  ( .A1(\SB1_3_14/i1[9] ), .A2(
        \SB1_3_14/i1_7 ), .A3(\SB1_3_14/i0[10] ), .ZN(
        \SB1_3_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_14/Component_Function_3/N1  ( .A1(\SB1_3_14/i1[9] ), .A2(
        \SB1_3_14/i0_3 ), .A3(\SB1_3_14/i0[6] ), .ZN(
        \SB1_3_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_4/N4  ( .A1(\SB1_3_14/i1[9] ), .A2(
        \SB1_3_14/i1_5 ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_4/N2  ( .A1(\SB1_3_14/i3[0] ), .A2(
        \SB1_3_14/i0_0 ), .A3(\SB1_3_14/i1_7 ), .ZN(
        \SB1_3_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_14/Component_Function_4/N1  ( .A1(\SB1_3_14/i0[9] ), .A2(
        \SB1_3_14/i0_0 ), .A3(\SB1_3_14/i0[8] ), .ZN(
        \SB1_3_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_2/N3  ( .A1(\SB1_3_15/i0_3 ), .A2(
        \SB1_3_15/i0[8] ), .A3(\SB1_3_15/i0[9] ), .ZN(
        \SB1_3_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_15/Component_Function_2/N2  ( .A1(n1647), .A2(
        \SB1_3_15/i0[10] ), .A3(\SB1_3_15/i0[6] ), .ZN(
        \SB1_3_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_15/Component_Function_3/N4  ( .A1(\SB1_3_15/i1_5 ), .A2(
        \SB1_3_15/i0[8] ), .A3(\SB1_3_15/i3[0] ), .ZN(
        \SB1_3_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_15/Component_Function_3/N2  ( .A1(\SB1_3_15/i0_0 ), .A2(
        \SB1_3_15/i0_3 ), .A3(\SB1_3_15/i0_4 ), .ZN(
        \SB1_3_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_15/Component_Function_3/N1  ( .A1(\SB1_3_15/i1[9] ), .A2(
        n1647), .A3(\SB1_3_15/i0[6] ), .ZN(
        \SB1_3_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_4/N4  ( .A1(\SB1_3_15/i1[9] ), .A2(
        \SB1_3_15/i1_5 ), .A3(\SB1_3_15/i0_4 ), .ZN(
        \SB1_3_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_15/Component_Function_4/N2  ( .A1(\SB1_3_15/i3[0] ), .A2(
        \SB1_3_15/i0_0 ), .A3(\SB1_3_15/i1_7 ), .ZN(
        \SB1_3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_15/Component_Function_4/N1  ( .A1(\SB1_3_15/i0[9] ), .A2(
        \SB1_3_15/i0_0 ), .A3(\SB1_3_15/i0[8] ), .ZN(
        \SB1_3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_2/N2  ( .A1(\SB1_3_16/i0_3 ), .A2(
        \SB1_3_16/i0[10] ), .A3(\SB1_3_16/i0[6] ), .ZN(
        \SB1_3_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_16/Component_Function_2/N1  ( .A1(\SB1_3_16/i1_5 ), .A2(
        \SB1_3_16/i0[10] ), .A3(\SB1_3_16/i1[9] ), .ZN(
        \SB1_3_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_3/N4  ( .A1(\SB1_3_16/i1_5 ), .A2(
        \SB1_3_16/i0[8] ), .A3(\SB1_3_16/i3[0] ), .ZN(
        \SB1_3_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_3/N3  ( .A1(\SB1_3_16/i1[9] ), .A2(
        \SB1_3_16/i1_7 ), .A3(\SB1_3_16/i0[10] ), .ZN(
        \SB1_3_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_16/Component_Function_3/N2  ( .A1(\SB1_3_16/i0_0 ), .A2(
        \SB1_3_16/i0_3 ), .A3(\SB1_3_16/i0_4 ), .ZN(
        \SB1_3_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_16/Component_Function_3/N1  ( .A1(\SB1_3_16/i1[9] ), .A2(
        \SB1_3_16/i0_3 ), .A3(\SB1_3_16/i0[6] ), .ZN(
        \SB1_3_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_4/N4  ( .A1(\SB1_3_16/i1[9] ), .A2(
        \SB1_3_16/i1_5 ), .A3(\SB1_3_16/i0_4 ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_4/N3  ( .A1(\SB1_3_16/i0[9] ), .A2(
        \SB1_3_16/i0[10] ), .A3(\SB1_3_16/i0_3 ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_16/Component_Function_4/N2  ( .A1(\SB1_3_16/i3[0] ), .A2(
        \SB1_3_16/i0_0 ), .A3(\SB1_3_16/i1_7 ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_16/Component_Function_4/N1  ( .A1(\SB1_3_16/i0[9] ), .A2(
        \SB1_3_16/i0_0 ), .A3(\SB1_3_16/i0[8] ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_17/Component_Function_2/N2  ( .A1(\SB1_3_17/i0_3 ), .A2(
        \SB1_3_17/i0[10] ), .A3(\SB1_3_17/i0[6] ), .ZN(
        \SB1_3_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_17/Component_Function_2/N1  ( .A1(\SB1_3_17/i1_5 ), .A2(
        \SB1_3_17/i0[10] ), .A3(\SB1_3_17/i1[9] ), .ZN(
        \SB1_3_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_17/Component_Function_3/N4  ( .A1(\SB1_3_17/i1_5 ), .A2(
        \SB1_3_17/i0[8] ), .A3(\SB1_3_17/i3[0] ), .ZN(
        \SB1_3_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_17/Component_Function_3/N2  ( .A1(\SB1_3_17/i0_0 ), .A2(
        \SB1_3_17/i0_3 ), .A3(\SB1_3_17/i0_4 ), .ZN(
        \SB1_3_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_17/Component_Function_3/N1  ( .A1(\SB1_3_17/i1[9] ), .A2(
        \SB1_3_17/i0_3 ), .A3(\SB1_3_17/i0[6] ), .ZN(
        \SB1_3_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_17/Component_Function_4/N4  ( .A1(\SB1_3_17/i1[9] ), .A2(
        \SB1_3_17/i1_5 ), .A3(\SB1_3_17/i0_4 ), .ZN(
        \SB1_3_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_17/Component_Function_4/N2  ( .A1(\SB1_3_17/i3[0] ), .A2(
        \SB1_3_17/i0_0 ), .A3(\SB1_3_17/i1_7 ), .ZN(
        \SB1_3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_17/Component_Function_4/N1  ( .A1(\SB1_3_17/i0[9] ), .A2(
        \SB1_3_17/i0_0 ), .A3(\SB1_3_17/i0[8] ), .ZN(
        \SB1_3_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_2/N3  ( .A1(\SB1_3_18/i0_3 ), .A2(
        \SB1_3_18/i0[8] ), .A3(\SB1_3_18/i0[9] ), .ZN(
        \SB1_3_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_18/Component_Function_2/N2  ( .A1(\SB1_3_18/i0_3 ), .A2(
        \SB1_3_18/i0[10] ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_3/N4  ( .A1(\SB1_3_18/i1_5 ), .A2(
        \SB1_3_18/i0[8] ), .A3(\SB1_3_18/i3[0] ), .ZN(
        \SB1_3_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_18/Component_Function_3/N2  ( .A1(\SB1_3_18/i0_0 ), .A2(
        \SB1_3_18/i0_3 ), .A3(\SB1_3_18/i0_4 ), .ZN(
        \SB1_3_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_3/N1  ( .A1(\SB1_3_18/i1[9] ), .A2(
        \SB1_3_18/i0_3 ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_4/N4  ( .A1(\SB1_3_18/i1[9] ), .A2(
        \SB1_3_18/i1_5 ), .A3(\SB1_3_18/i0_4 ), .ZN(
        \SB1_3_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_18/Component_Function_4/N2  ( .A1(\SB1_3_18/i3[0] ), .A2(
        \SB1_3_18/i0_0 ), .A3(\SB1_3_18/i1_7 ), .ZN(
        \SB1_3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_4/N1  ( .A1(\SB1_3_18/i0[9] ), .A2(
        \SB1_3_18/i0_0 ), .A3(\SB1_3_18/i0[8] ), .ZN(
        \SB1_3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_2/N2  ( .A1(\SB1_3_19/i0_3 ), .A2(
        \SB1_3_19/i0[10] ), .A3(\SB1_3_19/i0[6] ), .ZN(
        \SB1_3_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_19/Component_Function_2/N1  ( .A1(\SB1_3_19/i1_5 ), .A2(
        \SB1_3_19/i0[10] ), .A3(\SB1_3_19/i1[9] ), .ZN(
        \SB1_3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_3/N3  ( .A1(\SB1_3_19/i1[9] ), .A2(
        \SB1_3_19/i0[10] ), .A3(\SB1_3_19/i1_7 ), .ZN(
        \SB1_3_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_19/Component_Function_3/N2  ( .A1(\SB1_3_19/i0_0 ), .A2(
        \SB1_3_19/i0_3 ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N3  ( .A1(\SB1_3_19/i0[9] ), .A2(
        \SB1_3_19/i0[10] ), .A3(\SB1_3_19/i0_3 ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N2  ( .A1(\SB1_3_19/i3[0] ), .A2(
        \SB1_3_19/i0_0 ), .A3(\SB1_3_19/i1_7 ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N1  ( .A1(\SB1_3_19/i0[9] ), .A2(
        \SB1_3_19/i0_0 ), .A3(\SB1_3_19/i0[8] ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_2/N2  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i0[10] ), .A3(\SB1_3_20/i0[6] ), .ZN(
        \SB1_3_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_20/Component_Function_2/N1  ( .A1(\SB1_3_20/i1_5 ), .A2(
        \SB1_3_20/i0[10] ), .A3(\SB1_3_20/i1[9] ), .ZN(
        \SB1_3_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_3/N4  ( .A1(\SB1_3_20/i1_5 ), .A2(
        \SB1_3_20/i0[8] ), .A3(\SB1_3_20/i3[0] ), .ZN(
        \SB1_3_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_20/Component_Function_3/N1  ( .A1(\SB1_3_20/i1[9] ), .A2(
        \SB1_3_20/i0_3 ), .A3(\SB1_3_20/i0[6] ), .ZN(
        \SB1_3_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_4/N4  ( .A1(\SB1_3_20/i1[9] ), .A2(
        \SB1_3_20/i1_5 ), .A3(\SB1_3_20/i0_4 ), .ZN(
        \SB1_3_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_20/Component_Function_4/N3  ( .A1(\SB1_3_20/i0[9] ), .A2(
        \SB1_3_20/i0[10] ), .A3(\SB1_3_20/i0_3 ), .ZN(
        \SB1_3_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_20/Component_Function_4/N2  ( .A1(\SB1_3_20/i3[0] ), .A2(
        \SB1_3_20/i0_0 ), .A3(\SB1_3_20/i1_7 ), .ZN(
        \SB1_3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_20/Component_Function_4/N1  ( .A1(\SB1_3_20/i0[9] ), .A2(
        \SB1_3_20/i0_0 ), .A3(\SB1_3_20/i0[8] ), .ZN(
        \SB1_3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_2/N2  ( .A1(\SB1_3_21/i0_3 ), .A2(
        \SB1_3_21/i0[10] ), .A3(\SB1_3_21/i0[6] ), .ZN(
        \SB1_3_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_21/Component_Function_2/N1  ( .A1(\SB1_3_21/i0[10] ), .A2(
        \SB1_3_21/i1_5 ), .A3(\SB1_3_21/i1[9] ), .ZN(
        \SB1_3_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_3/N4  ( .A1(\SB1_3_21/i1_5 ), .A2(
        \SB1_3_21/i0[8] ), .A3(\SB1_3_21/i3[0] ), .ZN(
        \SB1_3_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_21/Component_Function_3/N1  ( .A1(\SB1_3_21/i1[9] ), .A2(
        \SB1_3_21/i0_3 ), .A3(\SB1_3_21/i0[6] ), .ZN(
        \SB1_3_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_4/N2  ( .A1(\SB1_3_21/i3[0] ), .A2(
        \SB1_3_21/i0_0 ), .A3(\SB1_3_21/i1_7 ), .ZN(
        \SB1_3_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_21/Component_Function_4/N1  ( .A1(\SB1_3_21/i0[9] ), .A2(
        \SB1_3_21/i0_0 ), .A3(\SB1_3_21/i0[8] ), .ZN(
        \SB1_3_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_2/N2  ( .A1(\SB1_3_22/i0_3 ), .A2(
        \SB1_3_22/i0[10] ), .A3(\SB1_3_22/i0[6] ), .ZN(
        \SB1_3_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_22/Component_Function_2/N1  ( .A1(\SB1_3_22/i1_5 ), .A2(
        \SB1_3_22/i0[10] ), .A3(\SB1_3_22/i1[9] ), .ZN(
        \SB1_3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_3/N4  ( .A1(\SB1_3_22/i1_5 ), .A2(
        \SB1_3_22/i0[8] ), .A3(\SB1_3_22/i3[0] ), .ZN(
        \SB1_3_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_22/Component_Function_3/N3  ( .A1(\SB1_3_22/i1[9] ), .A2(
        \SB1_3_22/i1_7 ), .A3(\SB1_3_22/i0[10] ), .ZN(
        \SB1_3_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_22/Component_Function_3/N2  ( .A1(\SB1_3_22/i0_0 ), .A2(
        \SB1_3_22/i0_3 ), .A3(\SB1_3_22/i0_4 ), .ZN(
        \SB1_3_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_22/Component_Function_3/N1  ( .A1(\SB1_3_22/i1[9] ), .A2(
        \SB1_3_22/i0_3 ), .A3(\SB1_3_22/i0[6] ), .ZN(
        \SB1_3_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_4/N2  ( .A1(\SB1_3_22/i3[0] ), .A2(
        \SB1_3_22/i0_0 ), .A3(\SB1_3_22/i1_7 ), .ZN(
        \SB1_3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_22/Component_Function_4/N1  ( .A1(\SB1_3_22/i0[9] ), .A2(
        \SB1_3_22/i0_0 ), .A3(\SB1_3_22/i0[8] ), .ZN(
        \SB1_3_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_2/N3  ( .A1(\SB1_3_23/i0_3 ), .A2(
        \SB1_3_23/i0[8] ), .A3(\SB1_3_23/i0[9] ), .ZN(
        \SB1_3_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_23/Component_Function_2/N2  ( .A1(\SB1_3_23/i0_3 ), .A2(
        \SB1_3_23/i0[10] ), .A3(\SB1_3_23/i0[6] ), .ZN(
        \SB1_3_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_23/Component_Function_2/N1  ( .A1(\SB1_3_23/i1_5 ), .A2(
        \SB1_3_23/i0[10] ), .A3(\SB1_3_23/i1[9] ), .ZN(
        \SB1_3_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_3/N4  ( .A1(\SB1_3_23/i1_5 ), .A2(
        \SB1_3_23/i0[8] ), .A3(\SB1_3_23/i3[0] ), .ZN(
        \SB1_3_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_23/Component_Function_3/N2  ( .A1(\SB1_3_23/i0_0 ), .A2(
        \SB1_3_23/i0_3 ), .A3(\SB1_3_23/i0_4 ), .ZN(
        \SB1_3_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_23/Component_Function_3/N1  ( .A1(\SB1_3_23/i1[9] ), .A2(
        \SB1_3_23/i0_3 ), .A3(\SB1_3_23/i0[6] ), .ZN(
        \SB1_3_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_4/N2  ( .A1(\SB1_3_23/i3[0] ), .A2(
        \SB1_3_23/i0_0 ), .A3(\SB1_3_23/i1_7 ), .ZN(
        \SB1_3_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_24/Component_Function_2/N3  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i0[8] ), .A3(\SB1_3_24/i0[9] ), .ZN(
        \SB1_3_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_24/Component_Function_2/N2  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i0[10] ), .A3(\SB1_3_24/i0[6] ), .ZN(
        \SB1_3_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_24/Component_Function_2/N1  ( .A1(\SB1_3_24/i1_5 ), .A2(
        \SB1_3_24/i0[10] ), .A3(\SB1_3_24/i1[9] ), .ZN(
        \SB1_3_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_3/N4  ( .A1(\SB1_3_24/i1_5 ), .A2(
        \SB1_3_24/i0[8] ), .A3(\SB1_3_24/i3[0] ), .ZN(
        \SB1_3_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_3/N2  ( .A1(\SB1_3_24/i0_0 ), .A2(
        \SB1_3_24/i0_3 ), .A3(\SB1_3_24/i0_4 ), .ZN(
        \SB1_3_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_24/Component_Function_3/N1  ( .A1(\SB1_3_24/i1[9] ), .A2(
        \SB1_3_24/i0_3 ), .A3(\SB1_3_24/i0[6] ), .ZN(
        \SB1_3_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_4/N4  ( .A1(\SB1_3_24/i1[9] ), .A2(
        \SB1_3_24/i1_5 ), .A3(\SB1_3_24/i0_4 ), .ZN(
        \SB1_3_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_4/N2  ( .A1(\SB1_3_24/i3[0] ), .A2(
        \SB1_3_24/i0_0 ), .A3(\SB1_3_24/i1_7 ), .ZN(
        \SB1_3_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_24/Component_Function_4/N1  ( .A1(\SB1_3_24/i0[9] ), .A2(
        \SB1_3_24/i0_0 ), .A3(\SB1_3_24/i0[8] ), .ZN(
        \SB1_3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_2/N2  ( .A1(n804), .A2(
        \SB1_3_25/i0[10] ), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_25/Component_Function_2/N1  ( .A1(\SB1_3_25/i1_5 ), .A2(
        \SB1_3_25/i0[10] ), .A3(\SB1_3_25/i1[9] ), .ZN(
        \SB1_3_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_3/N4  ( .A1(\SB1_3_25/i1_5 ), .A2(
        \SB1_3_25/i0[8] ), .A3(\SB1_3_25/i3[0] ), .ZN(
        \SB1_3_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_25/Component_Function_3/N3  ( .A1(\SB1_3_25/i1[9] ), .A2(
        \SB1_3_25/i1_7 ), .A3(\SB1_3_25/i0[10] ), .ZN(
        \SB1_3_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_25/Component_Function_3/N1  ( .A1(\SB1_3_25/i1[9] ), .A2(
        n804), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_4/N4  ( .A1(\SB1_3_25/i1[9] ), .A2(
        \SB1_3_25/i1_5 ), .A3(\SB1_3_25/i0_4 ), .ZN(
        \SB1_3_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_25/Component_Function_4/N2  ( .A1(\SB1_3_25/i3[0] ), .A2(
        \SB1_3_25/i0_0 ), .A3(\SB1_3_25/i1_7 ), .ZN(
        \SB1_3_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_25/Component_Function_4/N1  ( .A1(\SB1_3_25/i0[9] ), .A2(
        \SB1_3_25/i0_0 ), .A3(\SB1_3_25/i0[8] ), .ZN(
        \SB1_3_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_2/N2  ( .A1(\SB1_3_26/i0_3 ), .A2(
        \SB1_3_26/i0[10] ), .A3(\SB1_3_26/i0[6] ), .ZN(
        \SB1_3_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_26/Component_Function_3/N4  ( .A1(\SB1_3_26/i1_5 ), .A2(
        \SB1_3_26/i0[8] ), .A3(\SB1_3_26/i3[0] ), .ZN(
        \SB1_3_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_26/Component_Function_3/N2  ( .A1(\SB1_3_26/i0_0 ), .A2(
        \SB1_3_26/i0_3 ), .A3(\SB1_3_26/i0_4 ), .ZN(
        \SB1_3_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_26/Component_Function_3/N1  ( .A1(\SB1_3_26/i1[9] ), .A2(
        \SB1_3_26/i0_3 ), .A3(\SB1_3_26/i0[6] ), .ZN(
        \SB1_3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_4/N2  ( .A1(\SB1_3_26/i3[0] ), .A2(
        \SB1_3_26/i0_0 ), .A3(\SB1_3_26/i1_7 ), .ZN(
        \SB1_3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_26/Component_Function_4/N1  ( .A1(\SB1_3_26/i0[9] ), .A2(
        \SB1_3_26/i0_0 ), .A3(\SB1_3_26/i0[8] ), .ZN(
        \SB1_3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_2/N2  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i0[10] ), .A3(\SB1_3_27/i0[6] ), .ZN(
        \SB1_3_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_27/Component_Function_2/N1  ( .A1(\SB1_3_27/i1_5 ), .A2(
        \SB1_3_27/i0[10] ), .A3(\SB1_3_27/i1[9] ), .ZN(
        \SB1_3_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_3/N4  ( .A1(\SB1_3_27/i1_5 ), .A2(
        \SB1_3_27/i0[8] ), .A3(\SB1_3_27/i3[0] ), .ZN(
        \SB1_3_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_27/Component_Function_3/N3  ( .A1(\SB1_3_27/i0[10] ), .A2(
        \SB1_3_27/i1_7 ), .A3(\SB1_3_27/i1[9] ), .ZN(
        \SB1_3_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_27/Component_Function_3/N2  ( .A1(\SB1_3_27/i0_0 ), .A2(
        \SB1_3_27/i0_3 ), .A3(\SB1_3_27/i0_4 ), .ZN(
        \SB1_3_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_27/Component_Function_3/N1  ( .A1(\SB1_3_27/i1[9] ), .A2(
        \SB1_3_27/i0_3 ), .A3(\SB1_3_27/i0[6] ), .ZN(
        \SB1_3_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_4/N3  ( .A1(\SB1_3_27/i0[9] ), .A2(
        \SB1_3_27/i0[10] ), .A3(\SB1_3_27/i0_3 ), .ZN(
        \SB1_3_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_27/Component_Function_4/N2  ( .A1(\SB1_3_27/i3[0] ), .A2(
        \SB1_3_27/i0_0 ), .A3(\SB1_3_27/i1_7 ), .ZN(
        \SB1_3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_27/Component_Function_4/N1  ( .A1(\SB1_3_27/i0[9] ), .A2(
        \SB1_3_27/i0_0 ), .A3(\SB1_3_27/i0[8] ), .ZN(
        \SB1_3_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_2/N2  ( .A1(\SB1_3_28/i0_3 ), .A2(
        \SB1_3_28/i0[10] ), .A3(\SB1_3_28/i0[6] ), .ZN(
        \SB1_3_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_28/Component_Function_2/N1  ( .A1(\SB1_3_28/i1_5 ), .A2(
        \SB1_3_28/i0[10] ), .A3(\SB1_3_28/i1[9] ), .ZN(
        \SB1_3_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_3/N4  ( .A1(\SB1_3_28/i1_5 ), .A2(
        \SB1_3_28/i0[8] ), .A3(\SB1_3_28/i3[0] ), .ZN(
        \SB1_3_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_28/Component_Function_3/N3  ( .A1(\SB1_3_28/i1[9] ), .A2(
        \SB1_3_28/i1_7 ), .A3(\SB1_3_28/i0[10] ), .ZN(
        \SB1_3_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_28/Component_Function_3/N2  ( .A1(\SB1_3_28/i0_0 ), .A2(
        \SB1_3_28/i0_3 ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_28/Component_Function_3/N1  ( .A1(\SB1_3_28/i1[9] ), .A2(
        \SB1_3_28/i0_3 ), .A3(\SB1_3_28/i0[6] ), .ZN(
        \SB1_3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N4  ( .A1(\SB1_3_28/i1[9] ), .A2(
        \SB1_3_28/i1_5 ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N3  ( .A1(\SB1_3_28/i0[9] ), .A2(
        \SB1_3_28/i0[10] ), .A3(\SB1_3_28/i0_3 ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N2  ( .A1(\SB1_3_28/i3[0] ), .A2(
        \SB1_3_28/i0_0 ), .A3(\SB1_3_28/i1_7 ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N1  ( .A1(\SB1_3_28/i0[9] ), .A2(
        \SB1_3_28/i0_0 ), .A3(\SB1_3_28/i0[8] ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_2/N1  ( .A1(\SB1_3_29/i1_5 ), .A2(
        \SB1_3_29/i0[10] ), .A3(\SB1_3_29/i1[9] ), .ZN(
        \SB1_3_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_3/N4  ( .A1(\SB1_3_29/i1_5 ), .A2(
        \SB1_3_29/i0[8] ), .A3(\SB1_3_29/i3[0] ), .ZN(
        \SB1_3_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_29/Component_Function_3/N2  ( .A1(\SB1_3_29/i0_0 ), .A2(
        \SB1_3_29/i0_3 ), .A3(\SB1_3_29/i0_4 ), .ZN(
        \SB1_3_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_29/Component_Function_3/N1  ( .A1(\SB1_3_29/i1[9] ), .A2(
        \SB1_3_29/i0_3 ), .A3(\SB1_3_29/i0[6] ), .ZN(
        \SB1_3_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_4/N2  ( .A1(\SB1_3_29/i3[0] ), .A2(
        \SB1_3_29/i0_0 ), .A3(\SB1_3_29/i1_7 ), .ZN(
        \SB1_3_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_29/Component_Function_4/N1  ( .A1(\SB1_3_29/i0[9] ), .A2(
        \SB1_3_29/i0_0 ), .A3(\SB1_3_29/i0[8] ), .ZN(
        \SB1_3_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_2/N2  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i0[10] ), .A3(\SB1_3_30/i0[6] ), .ZN(
        \SB1_3_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_30/Component_Function_2/N1  ( .A1(\SB1_3_30/i1_5 ), .A2(
        \SB1_3_30/i0[10] ), .A3(\SB1_3_30/i1[9] ), .ZN(
        \SB1_3_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_3/N3  ( .A1(\SB1_3_30/i1[9] ), .A2(
        \SB1_3_30/i1_7 ), .A3(\SB1_3_30/i0[10] ), .ZN(
        \SB1_3_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_30/Component_Function_3/N2  ( .A1(\SB1_3_30/i0_0 ), .A2(
        \SB1_3_30/i0_3 ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_30/Component_Function_3/N1  ( .A1(\SB1_3_30/i1[9] ), .A2(
        \SB1_3_30/i0_3 ), .A3(\SB1_3_30/i0[6] ), .ZN(
        \SB1_3_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_4/N4  ( .A1(\SB1_3_30/i1[9] ), .A2(
        \SB1_3_30/i1_5 ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_30/Component_Function_4/N2  ( .A1(\SB1_3_30/i3[0] ), .A2(
        \SB1_3_30/i0_0 ), .A3(\SB1_3_30/i1_7 ), .ZN(
        \SB1_3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_30/Component_Function_4/N1  ( .A1(\SB1_3_30/i0[9] ), .A2(
        \SB1_3_30/i0_0 ), .A3(\SB1_3_30/i0[8] ), .ZN(
        \SB1_3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_31/Component_Function_2/N2  ( .A1(\SB1_3_31/i0_3 ), .A2(
        \SB1_3_31/i0[10] ), .A3(\SB1_3_31/i0[6] ), .ZN(
        \SB1_3_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_31/Component_Function_2/N1  ( .A1(\SB1_3_31/i1_5 ), .A2(
        \SB1_3_31/i0[10] ), .A3(\SB1_3_31/i1[9] ), .ZN(
        \SB1_3_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_31/Component_Function_3/N4  ( .A1(\SB1_3_31/i1_5 ), .A2(
        \SB1_3_31/i0[8] ), .A3(\SB1_3_31/i3[0] ), .ZN(
        \SB1_3_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_31/Component_Function_3/N2  ( .A1(\SB1_3_31/i0_0 ), .A2(
        \SB1_3_31/i0_3 ), .A3(\SB1_3_31/i0_4 ), .ZN(
        \SB1_3_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_31/Component_Function_3/N1  ( .A1(\SB1_3_31/i1[9] ), .A2(
        \SB1_3_31/i0_3 ), .A3(\SB1_3_31/i0[6] ), .ZN(
        \SB1_3_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_31/Component_Function_4/N4  ( .A1(\SB1_3_31/i1[9] ), .A2(
        \SB1_3_31/i1_5 ), .A3(\SB1_3_31/i0_4 ), .ZN(
        \SB1_3_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_31/Component_Function_4/N2  ( .A1(\SB1_3_31/i3[0] ), .A2(
        \SB1_3_31/i0_0 ), .A3(\SB1_3_31/i1_7 ), .ZN(
        \SB1_3_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_31/Component_Function_4/N1  ( .A1(\SB1_3_31/i0[9] ), .A2(
        \SB1_3_31/i0_0 ), .A3(\SB1_3_31/i0[8] ), .ZN(
        \SB1_3_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_2/N3  ( .A1(\SB2_3_0/i0_3 ), .A2(
        \SB2_3_0/i0[8] ), .A3(\SB2_3_0/i0[9] ), .ZN(
        \SB2_3_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_0/Component_Function_2/N2  ( .A1(\SB2_3_0/i0_3 ), .A2(
        \SB2_3_0/i0[10] ), .A3(\SB2_3_0/i0[6] ), .ZN(
        \SB2_3_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_0/Component_Function_2/N1  ( .A1(\SB2_3_0/i1_5 ), .A2(
        \SB2_3_0/i0[10] ), .A3(\SB2_3_0/i1[9] ), .ZN(
        \SB2_3_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_3/N4  ( .A1(\SB2_3_0/i1_5 ), .A2(
        \SB2_3_0/i0[8] ), .A3(\SB2_3_0/i3[0] ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_0/Component_Function_3/N3  ( .A1(\SB2_3_0/i1[9] ), .A2(
        \SB2_3_0/i1_7 ), .A3(\SB2_3_0/i0[10] ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_0/Component_Function_3/N2  ( .A1(\SB2_3_0/i0_0 ), .A2(
        \SB2_3_0/i0_3 ), .A3(\SB2_3_0/i0_4 ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_0/Component_Function_3/N1  ( .A1(\SB2_3_0/i1[9] ), .A2(
        \SB2_3_0/i0_3 ), .A3(\SB2_3_0/i0[6] ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_4/N4  ( .A1(\SB2_3_0/i1[9] ), .A2(
        \SB2_3_0/i1_5 ), .A3(\SB2_3_0/i0_4 ), .ZN(
        \SB2_3_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_0/Component_Function_4/N3  ( .A1(\SB2_3_0/i0[9] ), .A2(
        \SB2_3_0/i0[10] ), .A3(\SB2_3_0/i0_3 ), .ZN(
        \SB2_3_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_0/Component_Function_4/N2  ( .A1(\SB2_3_0/i3[0] ), .A2(
        \SB2_3_0/i0_0 ), .A3(\SB2_3_0/i1_7 ), .ZN(
        \SB2_3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_0/Component_Function_4/N1  ( .A1(\SB2_3_0/i0[9] ), .A2(
        \SB2_3_0/i0_0 ), .A3(\SB2_3_0/i0[8] ), .ZN(
        \SB2_3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_2/N3  ( .A1(\SB2_3_1/i0_3 ), .A2(
        \SB2_3_1/i0[8] ), .A3(\SB2_3_1/i0[9] ), .ZN(
        \SB2_3_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_1/Component_Function_2/N2  ( .A1(\SB2_3_1/i0_3 ), .A2(
        \SB2_3_1/i0[10] ), .A3(n1637), .ZN(
        \SB2_3_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_1/Component_Function_2/N1  ( .A1(\SB2_3_1/i1_5 ), .A2(
        \SB2_3_1/i0[10] ), .A3(\SB2_3_1/i1[9] ), .ZN(
        \SB2_3_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_3/N3  ( .A1(\SB2_3_1/i1[9] ), .A2(
        \SB2_3_1/i1_7 ), .A3(\SB2_3_1/i0[10] ), .ZN(
        \SB2_3_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_1/Component_Function_3/N2  ( .A1(\SB2_3_1/i0_0 ), .A2(
        \SB2_3_1/i0_3 ), .A3(\SB2_3_1/i0_4 ), .ZN(
        \SB2_3_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_1/Component_Function_3/N1  ( .A1(\SB2_3_1/i1[9] ), .A2(
        \SB2_3_1/i0_3 ), .A3(n1637), .ZN(
        \SB2_3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_4/N3  ( .A1(\SB2_3_1/i0[9] ), .A2(
        \SB2_3_1/i0[10] ), .A3(\SB2_3_1/i0_3 ), .ZN(
        \SB2_3_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_1/Component_Function_4/N2  ( .A1(\SB2_3_1/i3[0] ), .A2(
        \SB2_3_1/i0_0 ), .A3(\SB2_3_1/i1_7 ), .ZN(
        \SB2_3_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_1/Component_Function_4/N1  ( .A1(\SB2_3_1/i0[9] ), .A2(
        \SB2_3_1/i0_0 ), .A3(\SB2_3_1/i0[8] ), .ZN(
        \SB2_3_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_2/N2  ( .A1(\SB2_3_2/i0_3 ), .A2(
        \SB2_3_2/i0[10] ), .A3(\SB2_3_2/i0[6] ), .ZN(
        \SB2_3_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_2/Component_Function_2/N1  ( .A1(\SB2_3_2/i1_5 ), .A2(
        \SB2_3_2/i0[10] ), .A3(\SB2_3_2/i1[9] ), .ZN(
        \SB2_3_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_3/N4  ( .A1(\SB2_3_2/i1_5 ), .A2(
        \SB2_3_2/i0[8] ), .A3(\SB2_3_2/i3[0] ), .ZN(
        \SB2_3_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_2/Component_Function_3/N2  ( .A1(\SB2_3_2/i0_0 ), .A2(
        \SB2_3_2/i0_3 ), .A3(\SB2_3_2/i0_4 ), .ZN(
        \SB2_3_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_2/Component_Function_3/N1  ( .A1(\SB2_3_2/i1[9] ), .A2(
        \SB2_3_2/i0_3 ), .A3(\SB2_3_2/i0[6] ), .ZN(
        \SB2_3_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_4/N4  ( .A1(\SB2_3_2/i1[9] ), .A2(
        \SB2_3_2/i1_5 ), .A3(\SB2_3_2/i0_4 ), .ZN(
        \SB2_3_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_2/Component_Function_4/N3  ( .A1(\SB2_3_2/i0[9] ), .A2(
        \SB2_3_2/i0[10] ), .A3(\SB2_3_2/i0_3 ), .ZN(
        \SB2_3_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_2/Component_Function_4/N2  ( .A1(\SB2_3_2/i3[0] ), .A2(
        \SB2_3_2/i0_0 ), .A3(\SB2_3_2/i1_7 ), .ZN(
        \SB2_3_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_2/Component_Function_4/N1  ( .A1(\SB2_3_2/i0[9] ), .A2(
        \SB2_3_2/i0_0 ), .A3(\SB2_3_2/i0[8] ), .ZN(
        \SB2_3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_2/N4  ( .A1(\SB2_3_3/i1_5 ), .A2(
        \SB2_3_3/i0_0 ), .A3(\SB2_3_3/i0_4 ), .ZN(
        \SB2_3_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_2/N3  ( .A1(\SB2_3_3/i0_3 ), .A2(
        \SB2_3_3/i0[8] ), .A3(\SB2_3_3/i0[9] ), .ZN(
        \SB2_3_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_3/Component_Function_2/N2  ( .A1(\SB2_3_3/i0_3 ), .A2(
        \SB2_3_3/i0[10] ), .A3(\SB2_3_3/i0[6] ), .ZN(
        \SB2_3_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_3/Component_Function_2/N1  ( .A1(\SB2_3_3/i1_5 ), .A2(
        \SB2_3_3/i0[10] ), .A3(\SB2_3_3/i1[9] ), .ZN(
        \SB2_3_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_3/N4  ( .A1(\SB2_3_3/i1_5 ), .A2(
        \SB2_3_3/i0[8] ), .A3(\SB2_3_3/i3[0] ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_3/N3  ( .A1(\SB2_3_3/i1[9] ), .A2(
        \SB2_3_3/i1_7 ), .A3(\SB2_3_3/i0[10] ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_3/Component_Function_3/N2  ( .A1(\SB2_3_3/i0_0 ), .A2(
        \SB2_3_3/i0_3 ), .A3(\SB2_3_3/i0_4 ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_3/Component_Function_3/N1  ( .A1(\SB2_3_3/i1[9] ), .A2(
        \SB2_3_3/i0_3 ), .A3(\SB2_3_3/i0[6] ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_4/N4  ( .A1(\SB2_3_3/i1[9] ), .A2(
        \SB2_3_3/i1_5 ), .A3(\SB2_3_3/i0_4 ), .ZN(
        \SB2_3_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_4/N1  ( .A1(\SB2_3_3/i0[9] ), .A2(
        \SB2_3_3/i0_0 ), .A3(\SB2_3_3/i0[8] ), .ZN(
        \SB2_3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_2/N4  ( .A1(\SB2_3_4/i1_5 ), .A2(
        \SB2_3_4/i0_0 ), .A3(\SB2_3_4/i0_4 ), .ZN(
        \SB2_3_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_2/N3  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i0[8] ), .A3(n2133), .ZN(
        \SB2_3_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_4/Component_Function_2/N2  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i0[10] ), .A3(\SB2_3_4/i0[6] ), .ZN(
        \SB2_3_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_3/N3  ( .A1(\SB2_3_4/i1[9] ), .A2(
        \SB2_3_4/i1_7 ), .A3(\SB2_3_4/i0[10] ), .ZN(
        \SB2_3_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_4/Component_Function_3/N2  ( .A1(\SB2_3_4/i0_0 ), .A2(
        \SB2_3_4/i0_3 ), .A3(\SB2_3_4/i0_4 ), .ZN(
        \SB2_3_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_3/N1  ( .A1(\SB2_3_4/i1[9] ), .A2(
        \SB2_3_4/i0_3 ), .A3(\SB2_3_4/i0[6] ), .ZN(
        \SB2_3_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N4  ( .A1(\SB2_3_4/i1[9] ), .A2(
        \SB2_3_4/i1_5 ), .A3(\SB2_3_4/i0_4 ), .ZN(
        \SB2_3_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N2  ( .A1(\SB2_3_4/i3[0] ), .A2(
        \SB2_3_4/i0_0 ), .A3(\SB2_3_4/i1_7 ), .ZN(
        \SB2_3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N1  ( .A1(n2133), .A2(\SB2_3_4/i0_0 ), 
        .A3(\SB2_3_4/i0[8] ), .ZN(\SB2_3_4/Component_Function_4/NAND4_in[0] )
         );
  NAND3_X1 \SB2_3_5/Component_Function_2/N3  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i0[8] ), .A3(n2110), .ZN(
        \SB2_3_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_5/Component_Function_2/N2  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i0[10] ), .A3(\SB2_3_5/i0[6] ), .ZN(
        \SB2_3_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_5/Component_Function_2/N1  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[10] ), .A3(\SB2_3_5/i1[9] ), .ZN(
        \SB2_3_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_3/N4  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[8] ), .A3(\SB2_3_5/i3[0] ), .ZN(
        \SB2_3_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_5/Component_Function_3/N3  ( .A1(\SB2_3_5/i1[9] ), .A2(
        \SB2_3_5/i1_7 ), .A3(\SB2_3_5/i0[10] ), .ZN(
        \SB2_3_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_5/Component_Function_3/N2  ( .A1(\SB2_3_5/i0_0 ), .A2(
        \SB2_3_5/i0_3 ), .A3(\SB2_3_5/i0_4 ), .ZN(
        \SB2_3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_5/Component_Function_3/N1  ( .A1(\SB2_3_5/i1[9] ), .A2(
        \SB2_3_5/i0_3 ), .A3(\SB2_3_5/i0[6] ), .ZN(
        \SB2_3_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_4/N4  ( .A1(\SB2_3_5/i1[9] ), .A2(
        \SB2_3_5/i1_5 ), .A3(\SB2_3_5/i0_4 ), .ZN(
        \SB2_3_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_5/Component_Function_4/N3  ( .A1(n2110), .A2(
        \SB2_3_5/i0[10] ), .A3(\SB2_3_5/i0_3 ), .ZN(
        \SB2_3_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_5/Component_Function_4/N2  ( .A1(\SB2_3_5/i3[0] ), .A2(
        \SB2_3_5/i0_0 ), .A3(\SB2_3_5/i1_7 ), .ZN(
        \SB2_3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_5/Component_Function_4/N1  ( .A1(n2110), .A2(\SB2_3_5/i0_0 ), 
        .A3(\SB2_3_5/i0[8] ), .ZN(\SB2_3_5/Component_Function_4/NAND4_in[0] )
         );
  NAND3_X1 \SB2_3_6/Component_Function_2/N2  ( .A1(\SB2_3_6/i0_3 ), .A2(
        \SB2_3_6/i0[10] ), .A3(n2143), .ZN(
        \SB2_3_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_6/Component_Function_2/N1  ( .A1(\SB2_3_6/i1_5 ), .A2(
        \SB2_3_6/i0[10] ), .A3(\SB2_3_6/i1[9] ), .ZN(
        \SB2_3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_3/N3  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \SB2_3_6/i1_7 ), .A3(\SB2_3_6/i0[10] ), .ZN(
        \SB2_3_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_6/Component_Function_3/N2  ( .A1(\SB2_3_6/i0_0 ), .A2(
        \SB2_3_6/i0_3 ), .A3(\RI3[3][154] ), .ZN(
        \SB2_3_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_6/Component_Function_3/N1  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \SB2_3_6/i0_3 ), .A3(n2143), .ZN(
        \SB2_3_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_4/N4  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \SB2_3_6/i1_5 ), .A3(\RI3[3][154] ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_6/Component_Function_4/N3  ( .A1(\SB2_3_6/i0[9] ), .A2(
        \SB2_3_6/i0[10] ), .A3(\SB2_3_6/i0_3 ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_6/Component_Function_4/N2  ( .A1(\SB2_3_6/i3[0] ), .A2(
        \SB2_3_6/i0_0 ), .A3(\SB2_3_6/i1_7 ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_6/Component_Function_4/N1  ( .A1(\SB2_3_6/i0[9] ), .A2(
        \SB2_3_6/i0_0 ), .A3(\SB2_3_6/i0[8] ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_2/N4  ( .A1(\SB2_3_7/i1_5 ), .A2(
        \SB2_3_7/i0_0 ), .A3(\SB2_3_7/i0_4 ), .ZN(
        \SB2_3_7/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_7/Component_Function_2/N3  ( .A1(\SB2_3_7/i0_3 ), .A2(
        \SB2_3_7/i0[8] ), .A3(\SB2_3_7/i0[9] ), .ZN(
        \SB2_3_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_7/Component_Function_2/N2  ( .A1(\SB2_3_7/i0_3 ), .A2(
        \SB2_3_7/i0[10] ), .A3(\SB2_3_7/i0[6] ), .ZN(
        \SB2_3_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_7/Component_Function_2/N1  ( .A1(\SB2_3_7/i1_5 ), .A2(
        \SB2_3_7/i0[10] ), .A3(\SB2_3_7/i1[9] ), .ZN(
        \SB2_3_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_3/N4  ( .A1(\SB2_3_7/i1_5 ), .A2(
        \SB2_3_7/i0[8] ), .A3(\SB2_3_7/i3[0] ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_7/Component_Function_3/N3  ( .A1(\SB2_3_7/i1[9] ), .A2(
        \SB2_3_7/i1_7 ), .A3(\SB2_3_7/i0[10] ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_7/Component_Function_3/N2  ( .A1(\SB2_3_7/i0_0 ), .A2(
        \SB2_3_7/i0_3 ), .A3(\SB2_3_7/i0_4 ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_7/Component_Function_3/N1  ( .A1(\SB2_3_7/i1[9] ), .A2(
        \SB2_3_7/i0_3 ), .A3(\SB2_3_7/i0[6] ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_4/N4  ( .A1(\SB2_3_7/i1[9] ), .A2(
        \SB2_3_7/i1_5 ), .A3(\SB2_3_7/i0_4 ), .ZN(
        \SB2_3_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_7/Component_Function_4/N3  ( .A1(\SB2_3_7/i0_3 ), .A2(
        \SB2_3_7/i0[10] ), .A3(\SB2_3_7/i0[9] ), .ZN(
        \SB2_3_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_7/Component_Function_4/N1  ( .A1(\SB2_3_7/i0[9] ), .A2(
        \SB2_3_7/i0_0 ), .A3(\SB2_3_7/i0[8] ), .ZN(
        \SB2_3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_2/N4  ( .A1(\SB2_3_8/i1_5 ), .A2(
        \SB2_3_8/i0_0 ), .A3(\SB2_3_8/i0_4 ), .ZN(
        \SB2_3_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_2/N2  ( .A1(\SB2_3_8/i0_3 ), .A2(
        \SB2_3_8/i0[10] ), .A3(\SB2_3_8/i0[6] ), .ZN(
        \SB2_3_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_8/Component_Function_2/N1  ( .A1(\SB2_3_8/i1_5 ), .A2(
        \SB2_3_8/i0[10] ), .A3(\SB2_3_8/i1[9] ), .ZN(
        \SB2_3_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_3/N4  ( .A1(\SB2_3_8/i1_5 ), .A2(
        \SB2_3_8/i0[8] ), .A3(\SB2_3_8/i3[0] ), .ZN(
        \SB2_3_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_3/N3  ( .A1(\SB2_3_8/i1[9] ), .A2(
        \SB2_3_8/i1_7 ), .A3(\SB2_3_8/i0[10] ), .ZN(
        \SB2_3_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_8/Component_Function_3/N2  ( .A1(\SB2_3_8/i0_0 ), .A2(
        \SB2_3_8/i0_3 ), .A3(\SB2_3_8/i0_4 ), .ZN(
        \SB2_3_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_8/Component_Function_3/N1  ( .A1(\SB2_3_8/i1[9] ), .A2(
        \SB2_3_8/i0_3 ), .A3(\SB2_3_8/i0[6] ), .ZN(
        \SB2_3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_4/N4  ( .A1(\SB2_3_8/i1[9] ), .A2(
        \SB2_3_8/i1_5 ), .A3(\SB2_3_8/i0_4 ), .ZN(
        \SB2_3_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_4/N3  ( .A1(n1639), .A2(
        \SB2_3_8/i0[10] ), .A3(\SB2_3_8/i0_3 ), .ZN(
        \SB2_3_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_8/Component_Function_4/N2  ( .A1(\SB2_3_8/i3[0] ), .A2(
        \SB2_3_8/i0_0 ), .A3(\SB2_3_8/i1_7 ), .ZN(
        \SB2_3_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_8/Component_Function_4/N1  ( .A1(n1639), .A2(\SB2_3_8/i0_0 ), 
        .A3(\SB2_3_8/i0[8] ), .ZN(\SB2_3_8/Component_Function_4/NAND4_in[0] )
         );
  NAND3_X1 \SB2_3_9/Component_Function_2/N4  ( .A1(\SB2_3_9/i1_5 ), .A2(
        \SB2_3_9/i0_0 ), .A3(\SB2_3_9/i0_4 ), .ZN(
        \SB2_3_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_9/Component_Function_2/N3  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i0[8] ), .A3(n546), .ZN(
        \SB2_3_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_9/Component_Function_2/N2  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i0[10] ), .A3(\SB2_3_9/i0[6] ), .ZN(
        \SB2_3_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_9/Component_Function_2/N1  ( .A1(\SB2_3_9/i1_5 ), .A2(
        \SB2_3_9/i0[10] ), .A3(\SB2_3_9/i1[9] ), .ZN(
        \SB2_3_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_3/N3  ( .A1(\SB2_3_9/i1[9] ), .A2(
        \SB2_3_9/i1_7 ), .A3(\SB2_3_9/i0[10] ), .ZN(
        \SB2_3_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_9/Component_Function_3/N2  ( .A1(\SB2_3_9/i0_0 ), .A2(
        \SB2_3_9/i0_3 ), .A3(\SB2_3_9/i0_4 ), .ZN(
        \SB2_3_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_9/Component_Function_3/N1  ( .A1(\SB2_3_9/i1[9] ), .A2(
        \SB2_3_9/i0_3 ), .A3(\SB2_3_9/i0[6] ), .ZN(
        \SB2_3_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_4/N4  ( .A1(\SB2_3_9/i1[9] ), .A2(
        \SB2_3_9/i1_5 ), .A3(\SB2_3_9/i0_4 ), .ZN(
        \SB2_3_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_9/Component_Function_4/N3  ( .A1(n546), .A2(\SB2_3_9/i0[10] ), .A3(\SB2_3_9/i0_3 ), .ZN(\SB2_3_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_9/Component_Function_4/N1  ( .A1(n546), .A2(\SB2_3_9/i0_0 ), 
        .A3(\SB2_3_9/i0[8] ), .ZN(\SB2_3_9/Component_Function_4/NAND4_in[0] )
         );
  NAND3_X1 \SB2_3_10/Component_Function_2/N4  ( .A1(\SB2_3_10/i1_5 ), .A2(
        \SB2_3_10/i0_0 ), .A3(\SB2_3_10/i0_4 ), .ZN(
        \SB2_3_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_10/Component_Function_2/N3  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i0[8] ), .A3(\SB2_3_10/i0[9] ), .ZN(
        \SB2_3_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_10/Component_Function_2/N2  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i0[10] ), .A3(\SB2_3_10/i0[6] ), .ZN(
        \SB2_3_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_10/Component_Function_2/N1  ( .A1(\SB2_3_10/i1_5 ), .A2(
        \SB2_3_10/i0[10] ), .A3(\SB2_3_10/i1[9] ), .ZN(
        \SB2_3_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_3/N4  ( .A1(\SB2_3_10/i1_5 ), .A2(
        \SB2_3_10/i0[8] ), .A3(\SB2_3_10/i3[0] ), .ZN(
        \SB2_3_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_10/Component_Function_3/N3  ( .A1(\SB2_3_10/i1[9] ), .A2(
        \SB2_3_10/i1_7 ), .A3(\SB2_3_10/i0[10] ), .ZN(
        \SB2_3_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_10/Component_Function_3/N1  ( .A1(\SB2_3_10/i1[9] ), .A2(
        \SB2_3_10/i0_3 ), .A3(\SB2_3_10/i0[6] ), .ZN(
        \SB2_3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N3  ( .A1(\SB2_3_10/i0[9] ), .A2(
        \SB2_3_10/i0[10] ), .A3(\SB2_3_10/i0_3 ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N2  ( .A1(\SB2_3_10/i3[0] ), .A2(
        \SB2_3_10/i0_0 ), .A3(\SB2_3_10/i1_7 ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N1  ( .A1(\SB2_3_10/i0[9] ), .A2(
        \SB2_3_10/i0_0 ), .A3(\SB2_3_10/i0[8] ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_2/N4  ( .A1(\SB2_3_11/i1_5 ), .A2(
        \SB2_3_11/i0_0 ), .A3(\RI3[3][124] ), .ZN(
        \SB2_3_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_2/N3  ( .A1(\SB2_3_11/i0_3 ), .A2(
        \SB2_3_11/i0[8] ), .A3(\SB2_3_11/i0[9] ), .ZN(
        \SB2_3_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_11/Component_Function_2/N2  ( .A1(\SB2_3_11/i0_3 ), .A2(
        \SB2_3_11/i0[10] ), .A3(\SB2_3_11/i0[6] ), .ZN(
        \SB2_3_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_11/Component_Function_3/N4  ( .A1(\SB2_3_11/i1_5 ), .A2(
        \SB2_3_11/i0[8] ), .A3(\SB2_3_11/i3[0] ), .ZN(
        \SB2_3_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_3/N3  ( .A1(\SB2_3_11/i1[9] ), .A2(
        \SB2_3_11/i1_7 ), .A3(\SB2_3_11/i0[10] ), .ZN(
        \SB2_3_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_11/Component_Function_3/N2  ( .A1(\SB2_3_11/i0_0 ), .A2(
        \SB2_3_11/i0_3 ), .A3(\RI3[3][124] ), .ZN(
        \SB2_3_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_11/Component_Function_3/N1  ( .A1(\SB2_3_11/i1[9] ), .A2(
        \SB2_3_11/i0_3 ), .A3(\SB2_3_11/i0[6] ), .ZN(
        \SB2_3_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N4  ( .A1(\SB2_3_11/i1[9] ), .A2(
        \SB2_3_11/i1_5 ), .A3(\RI3[3][124] ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N3  ( .A1(\SB2_3_11/i0[9] ), .A2(
        \SB2_3_11/i0[10] ), .A3(\SB2_3_11/i0_3 ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N2  ( .A1(\SB2_3_11/i3[0] ), .A2(
        \SB2_3_11/i0_0 ), .A3(\SB2_3_11/i1_7 ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N1  ( .A1(\SB2_3_11/i0[9] ), .A2(
        \SB2_3_11/i0_0 ), .A3(\SB2_3_11/i0[8] ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_2/N4  ( .A1(\SB2_3_12/i1_5 ), .A2(
        \SB2_3_12/i0_0 ), .A3(\SB2_3_12/i0_4 ), .ZN(
        \SB2_3_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_2/N2  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i0[10] ), .A3(\SB2_3_12/i0[6] ), .ZN(
        \SB2_3_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_12/Component_Function_2/N1  ( .A1(\SB2_3_12/i1_5 ), .A2(
        \SB2_3_12/i0[10] ), .A3(\SB2_3_12/i1[9] ), .ZN(
        \SB2_3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_3/N4  ( .A1(\SB2_3_12/i1_5 ), .A2(
        \SB2_3_12/i0[8] ), .A3(\SB2_3_12/i3[0] ), .ZN(
        \SB2_3_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_3/N2  ( .A1(\SB2_3_12/i0_0 ), .A2(
        \SB2_3_12/i0_3 ), .A3(\SB2_3_12/i0_4 ), .ZN(
        \SB2_3_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_12/Component_Function_3/N1  ( .A1(\SB2_3_12/i1[9] ), .A2(
        \SB2_3_12/i0_3 ), .A3(\SB2_3_12/i0[6] ), .ZN(
        \SB2_3_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N4  ( .A1(\SB2_3_12/i1[9] ), .A2(
        \SB2_3_12/i1_5 ), .A3(\SB2_3_12/i0_4 ), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N3  ( .A1(\SB2_3_12/i0[9] ), .A2(
        \SB2_3_12/i0[10] ), .A3(\SB2_3_12/i0_3 ), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N1  ( .A1(\SB2_3_12/i0[9] ), .A2(
        \SB2_3_12/i0_0 ), .A3(\SB2_3_12/i0[8] ), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_2/N3  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i0[8] ), .A3(n2107), .ZN(
        \SB2_3_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_2/N2  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i0[10] ), .A3(\SB2_3_13/i0[6] ), .ZN(
        \SB2_3_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_13/Component_Function_2/N1  ( .A1(\SB2_3_13/i1_5 ), .A2(
        \SB2_3_13/i0[10] ), .A3(\SB2_3_13/i1[9] ), .ZN(
        \SB2_3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_3/N3  ( .A1(\SB2_3_13/i1[9] ), .A2(
        \SB2_3_13/i1_7 ), .A3(\SB2_3_13/i0[10] ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_3/N2  ( .A1(\SB2_3_13/i0_0 ), .A2(
        \SB2_3_13/i0_3 ), .A3(\SB2_3_13/i0_4 ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_13/Component_Function_3/N1  ( .A1(\SB2_3_13/i1[9] ), .A2(
        \SB2_3_13/i0_3 ), .A3(\SB2_3_13/i0[6] ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_4/N4  ( .A1(\SB2_3_13/i1[9] ), .A2(
        \SB2_3_13/i1_5 ), .A3(\SB2_3_13/i0_4 ), .ZN(
        \SB2_3_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_13/Component_Function_4/N2  ( .A1(\SB2_3_13/i3[0] ), .A2(
        \SB2_3_13/i0_0 ), .A3(\SB2_3_13/i1_7 ), .ZN(
        \SB2_3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_13/Component_Function_4/N1  ( .A1(n2107), .A2(
        \SB2_3_13/i0_0 ), .A3(\SB2_3_13/i0[8] ), .ZN(
        \SB2_3_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_2/N4  ( .A1(\SB2_3_14/i1_5 ), .A2(
        \SB2_3_14/i0_0 ), .A3(n1945), .ZN(
        \SB2_3_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_2/N3  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i0[8] ), .A3(\SB2_3_14/i0[9] ), .ZN(
        \SB2_3_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_14/Component_Function_2/N2  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i0[10] ), .A3(\SB2_3_14/i0[6] ), .ZN(
        \SB2_3_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_2/N1  ( .A1(\SB2_3_14/i1_5 ), .A2(
        \SB2_3_14/i0[10] ), .A3(\SB2_3_14/i1[9] ), .ZN(
        \SB2_3_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_3/N4  ( .A1(\SB2_3_14/i1_5 ), .A2(
        \SB2_3_14/i0[8] ), .A3(\SB2_3_14/i3[0] ), .ZN(
        \SB2_3_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_3/N3  ( .A1(\SB2_3_14/i1[9] ), .A2(
        \SB2_3_14/i1_7 ), .A3(\SB2_3_14/i0[10] ), .ZN(
        \SB2_3_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_14/Component_Function_3/N2  ( .A1(\SB2_3_14/i0_0 ), .A2(
        \SB2_3_14/i0_3 ), .A3(n1945), .ZN(
        \SB2_3_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_3/N1  ( .A1(\SB2_3_14/i1[9] ), .A2(
        \SB2_3_14/i0_3 ), .A3(\SB2_3_14/i0[6] ), .ZN(
        \SB2_3_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N4  ( .A1(\SB2_3_14/i1[9] ), .A2(
        \SB2_3_14/i1_5 ), .A3(n1945), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N3  ( .A1(\SB2_3_14/i0[9] ), .A2(
        \SB2_3_14/i0[10] ), .A3(\SB2_3_14/i0_3 ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N2  ( .A1(\SB2_3_14/i3[0] ), .A2(
        \SB2_3_14/i0_0 ), .A3(\SB2_3_14/i1_7 ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N1  ( .A1(\RI3[3][102] ), .A2(
        \SB2_3_14/i0_0 ), .A3(\SB2_3_14/i0[8] ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_2/N3  ( .A1(\SB2_3_15/i0_3 ), .A2(
        \SB2_3_15/i0[8] ), .A3(\SB2_3_15/i0[9] ), .ZN(
        \SB2_3_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_15/Component_Function_2/N2  ( .A1(\SB2_3_15/i0_3 ), .A2(
        \SB2_3_15/i0[10] ), .A3(n2097), .ZN(
        \SB2_3_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_15/Component_Function_2/N1  ( .A1(\SB2_3_15/i1_5 ), .A2(
        \SB2_3_15/i0[10] ), .A3(\SB2_3_15/i1[9] ), .ZN(
        \SB2_3_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_3/N3  ( .A1(\SB2_3_15/i1[9] ), .A2(
        n1965), .A3(\SB2_3_15/i0[10] ), .ZN(
        \SB2_3_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_15/Component_Function_3/N2  ( .A1(\SB2_3_15/i0_0 ), .A2(
        \SB2_3_15/i0_3 ), .A3(\SB2_3_15/i0_4 ), .ZN(
        \SB2_3_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_15/Component_Function_3/N1  ( .A1(\SB2_3_15/i1[9] ), .A2(
        \SB2_3_15/i0_3 ), .A3(n2097), .ZN(
        \SB2_3_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N4  ( .A1(\SB2_3_15/i1[9] ), .A2(
        \SB2_3_15/i1_5 ), .A3(\SB2_3_15/i0_4 ), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N2  ( .A1(\SB2_3_15/i3[0] ), .A2(
        \SB2_3_15/i0_0 ), .A3(n1965), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N1  ( .A1(\SB2_3_15/i0[9] ), .A2(
        \SB2_3_15/i0_0 ), .A3(\SB2_3_15/i0[8] ), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_2/N2  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i0[10] ), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_16/Component_Function_2/N1  ( .A1(\SB2_3_16/i1_5 ), .A2(
        \SB2_3_16/i0[10] ), .A3(\SB2_3_16/i1[9] ), .ZN(
        \SB2_3_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_3/N3  ( .A1(\SB2_3_16/i1[9] ), .A2(
        \SB2_3_16/i1_7 ), .A3(\SB2_3_16/i0[10] ), .ZN(
        \SB2_3_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_16/Component_Function_3/N2  ( .A1(\SB2_3_16/i0_0 ), .A2(
        \SB2_3_16/i0_3 ), .A3(\RI3[3][94] ), .ZN(
        \SB2_3_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_16/Component_Function_3/N1  ( .A1(\SB2_3_16/i1[9] ), .A2(
        \SB2_3_16/i0_3 ), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_4/N4  ( .A1(\SB2_3_16/i1[9] ), .A2(
        \SB2_3_16/i1_5 ), .A3(\RI3[3][94] ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_16/Component_Function_4/N3  ( .A1(n2114), .A2(
        \SB2_3_16/i0[10] ), .A3(\SB2_3_16/i0_3 ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_16/Component_Function_4/N2  ( .A1(\SB2_3_16/i3[0] ), .A2(
        \SB2_3_16/i0_0 ), .A3(\SB2_3_16/i1_7 ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_16/Component_Function_4/N1  ( .A1(n2114), .A2(
        \SB2_3_16/i0_0 ), .A3(\SB2_3_16/i0[8] ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_17/Component_Function_2/N4  ( .A1(\SB2_3_17/i1_5 ), .A2(
        \SB2_3_17/i0_0 ), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_2/N3  ( .A1(\SB2_3_17/i0_3 ), .A2(
        \SB2_3_17/i0[8] ), .A3(\SB2_3_17/i0[9] ), .ZN(
        \SB2_3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_17/Component_Function_2/N2  ( .A1(\SB2_3_17/i0_3 ), .A2(
        \SB2_3_17/i0[10] ), .A3(\SB2_3_17/i0[6] ), .ZN(
        \SB2_3_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_17/Component_Function_3/N4  ( .A1(\SB2_3_17/i1_5 ), .A2(
        \SB2_3_17/i0[8] ), .A3(\SB2_3_17/i3[0] ), .ZN(
        \SB2_3_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_3/N3  ( .A1(\SB2_3_17/i1[9] ), .A2(
        \SB2_3_17/i1_7 ), .A3(\SB2_3_17/i0[10] ), .ZN(
        \SB2_3_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_17/Component_Function_3/N2  ( .A1(\SB2_3_17/i0_0 ), .A2(
        \SB2_3_17/i0_3 ), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_17/Component_Function_3/N1  ( .A1(\SB2_3_17/i1[9] ), .A2(
        \SB2_3_17/i0_3 ), .A3(\SB2_3_17/i0[6] ), .ZN(
        \SB2_3_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_17/Component_Function_4/N4  ( .A1(\SB2_3_17/i1[9] ), .A2(
        \SB2_3_17/i1_5 ), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_4/N3  ( .A1(\SB2_3_17/i0[9] ), .A2(
        \SB2_3_17/i0[10] ), .A3(\SB2_3_17/i0_3 ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_17/Component_Function_4/N2  ( .A1(\SB2_3_17/i3[0] ), .A2(
        \SB2_3_17/i0_0 ), .A3(\SB2_3_17/i1_7 ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_17/Component_Function_4/N1  ( .A1(\SB2_3_17/i0[9] ), .A2(
        \SB2_3_17/i0_0 ), .A3(\SB2_3_17/i0[8] ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_2/N3  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i0[8] ), .A3(\SB2_3_18/i0[9] ), .ZN(
        \SB2_3_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_18/Component_Function_2/N2  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i0[10] ), .A3(\SB2_3_18/i0[6] ), .ZN(
        \SB2_3_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_18/Component_Function_2/N1  ( .A1(\SB2_3_18/i1_5 ), .A2(
        \SB2_3_18/i0[10] ), .A3(\SB2_3_18/i1[9] ), .ZN(
        \SB2_3_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_3/N3  ( .A1(\SB2_3_18/i1[9] ), .A2(
        \SB2_3_18/i1_7 ), .A3(\SB2_3_18/i0[10] ), .ZN(
        \SB2_3_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_18/Component_Function_3/N1  ( .A1(\SB2_3_18/i1[9] ), .A2(
        \SB2_3_18/i0_3 ), .A3(\SB2_3_18/i0[6] ), .ZN(
        \SB2_3_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N4  ( .A1(\SB2_3_18/i1[9] ), .A2(
        \SB2_3_18/i1_5 ), .A3(\SB2_3_18/i0_4 ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N2  ( .A1(\SB2_3_18/i3[0] ), .A2(
        \SB2_3_18/i0_0 ), .A3(\SB2_3_18/i1_7 ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N1  ( .A1(\SB2_3_18/i0[9] ), .A2(
        \SB2_3_18/i0_0 ), .A3(\SB2_3_18/i0[8] ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_2/N4  ( .A1(\SB2_3_19/i1_5 ), .A2(
        \SB2_3_19/i0_0 ), .A3(\SB2_3_19/i0_4 ), .ZN(
        \SB2_3_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_19/Component_Function_2/N3  ( .A1(\SB2_3_19/i0_3 ), .A2(
        \SB2_3_19/i0[8] ), .A3(n1623), .ZN(
        \SB2_3_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_19/Component_Function_2/N2  ( .A1(\SB2_3_19/i0_3 ), .A2(
        \SB2_3_19/i0[10] ), .A3(\SB2_3_19/i0[6] ), .ZN(
        \SB2_3_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_19/Component_Function_2/N1  ( .A1(\SB2_3_19/i1_5 ), .A2(
        \SB2_3_19/i0[10] ), .A3(\SB2_3_19/i1[9] ), .ZN(
        \SB2_3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_3/N4  ( .A1(\SB2_3_19/i1_5 ), .A2(
        \SB2_3_19/i0[8] ), .A3(\SB2_3_19/i3[0] ), .ZN(
        \SB2_3_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_19/Component_Function_3/N3  ( .A1(\SB2_3_19/i1[9] ), .A2(
        \SB2_3_19/i1_7 ), .A3(\SB2_3_19/i0[10] ), .ZN(
        \SB2_3_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_19/Component_Function_3/N2  ( .A1(\SB2_3_19/i0_0 ), .A2(
        \SB2_3_19/i0_3 ), .A3(\SB2_3_19/i0_4 ), .ZN(
        \SB2_3_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_19/Component_Function_3/N1  ( .A1(\SB2_3_19/i1[9] ), .A2(
        \SB2_3_19/i0_3 ), .A3(\SB2_3_19/i0[6] ), .ZN(
        \SB2_3_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_4/N4  ( .A1(\SB2_3_19/i1[9] ), .A2(
        \SB2_3_19/i1_5 ), .A3(\SB2_3_19/i0_4 ), .ZN(
        \SB2_3_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_19/Component_Function_4/N1  ( .A1(n1623), .A2(
        \SB2_3_19/i0_0 ), .A3(\SB2_3_19/i0[8] ), .ZN(
        \SB2_3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_2/N4  ( .A1(\SB2_3_20/i1_5 ), .A2(
        \SB2_3_20/i0_0 ), .A3(\SB2_3_20/i0_4 ), .ZN(
        \SB2_3_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_2/N2  ( .A1(\SB2_3_20/i0_3 ), .A2(
        \SB2_3_20/i0[10] ), .A3(\SB2_3_20/i0[6] ), .ZN(
        \SB2_3_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_20/Component_Function_2/N1  ( .A1(\SB2_3_20/i1_5 ), .A2(
        \SB2_3_20/i0[10] ), .A3(\SB2_3_20/i1[9] ), .ZN(
        \SB2_3_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_3/N4  ( .A1(\SB2_3_20/i1_5 ), .A2(
        \SB2_3_20/i0[8] ), .A3(\SB2_3_20/i3[0] ), .ZN(
        \SB2_3_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_3/N3  ( .A1(\SB2_3_20/i0[10] ), .A2(
        \SB2_3_20/i1_7 ), .A3(\SB2_3_20/i1[9] ), .ZN(
        \SB2_3_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_20/Component_Function_3/N2  ( .A1(\SB2_3_20/i0_0 ), .A2(
        \SB2_3_20/i0_3 ), .A3(\SB2_3_20/i0_4 ), .ZN(
        \SB2_3_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_20/Component_Function_4/N4  ( .A1(\SB2_3_20/i1[9] ), .A2(
        \SB2_3_20/i1_5 ), .A3(\SB2_3_20/i0_4 ), .ZN(
        \SB2_3_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_4/N3  ( .A1(\SB2_3_20/i0[9] ), .A2(
        \SB2_3_20/i0[10] ), .A3(\SB2_3_20/i0_3 ), .ZN(
        \SB2_3_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_20/Component_Function_4/N2  ( .A1(\SB2_3_20/i3[0] ), .A2(
        \SB2_3_20/i0_0 ), .A3(\SB2_3_20/i1_7 ), .ZN(
        \SB2_3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_20/Component_Function_4/N1  ( .A1(\SB2_3_20/i0[9] ), .A2(
        \SB2_3_20/i0_0 ), .A3(\SB2_3_20/i0[8] ), .ZN(
        \SB2_3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_2/N2  ( .A1(\SB2_3_21/i0_3 ), .A2(
        \SB2_3_21/i0[10] ), .A3(\SB2_3_21/i0[6] ), .ZN(
        \SB2_3_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_21/Component_Function_2/N1  ( .A1(\SB2_3_21/i1_5 ), .A2(
        \SB2_3_21/i0[10] ), .A3(\SB2_3_21/i1[9] ), .ZN(
        \SB2_3_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_3/N3  ( .A1(\SB2_3_21/i1[9] ), .A2(
        \SB2_3_21/i1_7 ), .A3(\SB2_3_21/i0[10] ), .ZN(
        \SB2_3_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_21/Component_Function_3/N2  ( .A1(\SB2_3_21/i0_0 ), .A2(
        \SB2_3_21/i0_3 ), .A3(\RI3[3][64] ), .ZN(
        \SB2_3_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_21/Component_Function_4/N3  ( .A1(\SB2_3_21/i0[9] ), .A2(
        \SB2_3_21/i0[10] ), .A3(\SB2_3_21/i0_3 ), .ZN(
        \SB2_3_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_21/Component_Function_4/N1  ( .A1(\SB2_3_21/i0[9] ), .A2(
        \SB2_3_21/i0_0 ), .A3(\SB2_3_21/i0[8] ), .ZN(
        \SB2_3_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_2/N4  ( .A1(\SB2_3_22/i1_5 ), .A2(
        \SB2_3_22/i0_0 ), .A3(\SB2_3_22/i0_4 ), .ZN(
        \SB2_3_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_22/Component_Function_2/N3  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i0[8] ), .A3(\SB2_3_22/i0[9] ), .ZN(
        \SB2_3_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_22/Component_Function_2/N2  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i0[10] ), .A3(\SB2_3_22/i0[6] ), .ZN(
        \SB2_3_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_22/Component_Function_2/N1  ( .A1(\SB2_3_22/i1_5 ), .A2(
        \SB2_3_22/i0[10] ), .A3(\SB2_3_22/i1[9] ), .ZN(
        \SB2_3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_3/N3  ( .A1(\SB2_3_22/i1[9] ), .A2(
        \SB2_3_22/i1_7 ), .A3(\SB2_3_22/i0[10] ), .ZN(
        \SB2_3_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_22/Component_Function_3/N2  ( .A1(\SB2_3_22/i0_0 ), .A2(
        \SB2_3_22/i0_3 ), .A3(\SB2_3_22/i0_4 ), .ZN(
        \SB2_3_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_22/Component_Function_3/N1  ( .A1(\SB2_3_22/i1[9] ), .A2(
        \SB2_3_22/i0_3 ), .A3(\SB2_3_22/i0[6] ), .ZN(
        \SB2_3_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_4/N4  ( .A1(\SB2_3_22/i1[9] ), .A2(
        \SB2_3_22/i1_5 ), .A3(\SB2_3_22/i0_4 ), .ZN(
        \SB2_3_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_22/Component_Function_4/N3  ( .A1(\SB2_3_22/i0[9] ), .A2(
        \SB2_3_22/i0[10] ), .A3(\SB2_3_22/i0_3 ), .ZN(
        \SB2_3_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_22/Component_Function_4/N2  ( .A1(\SB2_3_22/i3[0] ), .A2(
        \SB2_3_22/i0_0 ), .A3(\SB2_3_22/i1_7 ), .ZN(
        \SB2_3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_22/Component_Function_4/N1  ( .A1(\SB2_3_22/i0[9] ), .A2(
        \SB2_3_22/i0_0 ), .A3(\SB2_3_22/i0[8] ), .ZN(
        \SB2_3_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_2/N4  ( .A1(\SB2_3_23/i1_5 ), .A2(
        \SB2_3_23/i0_0 ), .A3(\SB2_3_23/i0_4 ), .ZN(
        \SB2_3_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_23/Component_Function_2/N2  ( .A1(\SB2_3_23/i0_3 ), .A2(
        \SB2_3_23/i0[10] ), .A3(\SB2_3_23/i0[6] ), .ZN(
        \SB2_3_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_23/Component_Function_2/N1  ( .A1(\SB2_3_23/i1_5 ), .A2(
        \SB2_3_23/i0[10] ), .A3(\SB2_3_23/i1[9] ), .ZN(
        \SB2_3_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_3/N3  ( .A1(\SB2_3_23/i1[9] ), .A2(
        \SB2_3_23/i1_7 ), .A3(\SB2_3_23/i0[10] ), .ZN(
        \SB2_3_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_23/Component_Function_3/N2  ( .A1(\SB2_3_23/i0_0 ), .A2(
        \SB2_3_23/i0_3 ), .A3(\SB2_3_23/i0_4 ), .ZN(
        \SB2_3_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_23/Component_Function_3/N1  ( .A1(\SB2_3_23/i1[9] ), .A2(
        \SB2_3_23/i0_3 ), .A3(\SB2_3_23/i0[6] ), .ZN(
        \SB2_3_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N4  ( .A1(\SB2_3_23/i1[9] ), .A2(
        \SB2_3_23/i1_5 ), .A3(\SB2_3_23/i0_4 ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N3  ( .A1(\SB2_3_23/i0[9] ), .A2(
        \SB2_3_23/i0[10] ), .A3(\SB2_3_23/i0_3 ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N2  ( .A1(\SB2_3_23/i3[0] ), .A2(
        \SB2_3_23/i0_0 ), .A3(\SB2_3_23/i1_7 ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N1  ( .A1(\SB2_3_23/i0[9] ), .A2(
        \SB2_3_23/i0_0 ), .A3(\SB2_3_23/i0[8] ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_24/Component_Function_2/N4  ( .A1(\SB2_3_24/i1_5 ), .A2(
        \SB2_3_24/i0_0 ), .A3(\SB2_3_24/i0_4 ), .ZN(
        \SB2_3_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_2/N3  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB2_3_24/i0[8] ), .A3(\SB2_3_24/i0[9] ), .ZN(
        \SB2_3_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_24/Component_Function_2/N2  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB2_3_24/i0[10] ), .A3(\SB2_3_24/i0[6] ), .ZN(
        \SB2_3_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_3/N4  ( .A1(\SB2_3_24/i1_5 ), .A2(
        \SB2_3_24/i0[8] ), .A3(\SB2_3_24/i3[0] ), .ZN(
        \SB2_3_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_3/N3  ( .A1(\SB2_3_24/i1[9] ), .A2(
        \SB2_3_24/i1_7 ), .A3(\SB2_3_24/i0[10] ), .ZN(
        \SB2_3_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_24/Component_Function_3/N2  ( .A1(\SB2_3_24/i0_0 ), .A2(
        \SB2_3_24/i0_3 ), .A3(\SB2_3_24/i0_4 ), .ZN(
        \SB2_3_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_3/N1  ( .A1(\SB2_3_24/i1[9] ), .A2(
        \SB2_3_24/i0_3 ), .A3(\SB2_3_24/i0[6] ), .ZN(
        \SB2_3_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N4  ( .A1(\SB2_3_24/i1[9] ), .A2(
        \SB2_3_24/i1_5 ), .A3(\SB2_3_24/i0_4 ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N3  ( .A1(\SB2_3_24/i0[9] ), .A2(
        \SB2_3_24/i0[10] ), .A3(\SB2_3_24/i0_3 ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N2  ( .A1(\SB2_3_24/i3[0] ), .A2(
        \SB2_3_24/i0_0 ), .A3(\SB2_3_24/i1_7 ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N1  ( .A1(\SB2_3_24/i0[9] ), .A2(
        \SB2_3_24/i0_0 ), .A3(\SB2_3_24/i0[8] ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_25/Component_Function_2/N4  ( .A1(\SB2_3_25/i1_5 ), .A2(
        \SB2_3_25/i0_0 ), .A3(\SB2_3_25/i0_4 ), .ZN(
        \SB2_3_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_25/Component_Function_2/N3  ( .A1(\SB2_3_25/i0_3 ), .A2(
        \SB2_3_25/i0[8] ), .A3(\SB2_3_25/i0[9] ), .ZN(
        \SB2_3_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_25/Component_Function_2/N2  ( .A1(\SB2_3_25/i0_3 ), .A2(
        \SB2_3_25/i0[10] ), .A3(\SB2_3_25/i0[6] ), .ZN(
        \SB2_3_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_25/Component_Function_3/N4  ( .A1(\SB2_3_25/i1_5 ), .A2(
        \SB2_3_25/i0[8] ), .A3(\SB2_3_25/i3[0] ), .ZN(
        \SB2_3_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_25/Component_Function_3/N3  ( .A1(\SB2_3_25/i1[9] ), .A2(
        \SB2_3_25/i1_7 ), .A3(\SB2_3_25/i0[10] ), .ZN(
        \SB2_3_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_25/Component_Function_3/N2  ( .A1(\SB2_3_25/i0_0 ), .A2(
        \SB2_3_25/i0_3 ), .A3(\SB2_3_25/i0_4 ), .ZN(
        \SB2_3_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_25/Component_Function_3/N1  ( .A1(\SB2_3_25/i1[9] ), .A2(
        \SB2_3_25/i0[6] ), .A3(\SB2_3_25/i0_3 ), .ZN(
        \SB2_3_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_25/Component_Function_4/N4  ( .A1(\SB2_3_25/i0_4 ), .A2(
        \SB2_3_25/i1_5 ), .A3(\SB2_3_25/i1[9] ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_25/Component_Function_4/N3  ( .A1(\SB2_3_25/i0[9] ), .A2(
        \SB2_3_25/i0[10] ), .A3(\SB2_3_25/i0_3 ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_25/Component_Function_4/N2  ( .A1(\SB2_3_25/i3[0] ), .A2(
        \SB2_3_25/i0_0 ), .A3(\SB2_3_25/i1_7 ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_25/Component_Function_4/N1  ( .A1(\SB2_3_25/i0[9] ), .A2(
        \SB2_3_25/i0_0 ), .A3(\SB2_3_25/i0[8] ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_2/N4  ( .A1(\SB2_3_26/i1_5 ), .A2(
        \SB2_3_26/i0_0 ), .A3(\SB2_3_26/i0_4 ), .ZN(
        \SB2_3_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_26/Component_Function_2/N3  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i0[8] ), .A3(\SB2_3_26/i0[9] ), .ZN(
        \SB2_3_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_26/Component_Function_2/N2  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i0[10] ), .A3(\SB2_3_26/i0[6] ), .ZN(
        \SB2_3_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_26/Component_Function_2/N1  ( .A1(\SB2_3_26/i1_5 ), .A2(
        \SB2_3_26/i0[10] ), .A3(\SB2_3_26/i1[9] ), .ZN(
        \SB2_3_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_3/N4  ( .A1(\SB2_3_26/i1_5 ), .A2(
        \SB2_3_26/i0[8] ), .A3(\SB2_3_26/i3[0] ), .ZN(
        \SB2_3_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_26/Component_Function_3/N3  ( .A1(\SB2_3_26/i1[9] ), .A2(
        \SB2_3_26/i1_7 ), .A3(\SB2_3_26/i0[10] ), .ZN(
        \SB2_3_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_26/Component_Function_3/N2  ( .A1(\SB2_3_26/i0_0 ), .A2(
        \SB2_3_26/i0_3 ), .A3(\SB2_3_26/i0_4 ), .ZN(
        \SB2_3_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_26/Component_Function_3/N1  ( .A1(\SB2_3_26/i1[9] ), .A2(
        \SB2_3_26/i0_3 ), .A3(\SB2_3_26/i0[6] ), .ZN(
        \SB2_3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N4  ( .A1(\SB2_3_26/i1[9] ), .A2(
        \SB2_3_26/i1_5 ), .A3(\SB2_3_26/i0_4 ), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N2  ( .A1(\SB2_3_26/i3[0] ), .A2(
        \SB2_3_26/i0_0 ), .A3(\SB2_3_26/i1_7 ), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N1  ( .A1(\SB2_3_26/i0[9] ), .A2(
        \SB2_3_26/i0_0 ), .A3(\SB2_3_26/i0[8] ), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_2/N4  ( .A1(n1630), .A2(
        \SB2_3_27/i0_0 ), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_27/Component_Function_2/N2  ( .A1(\SB2_3_27/i0_3 ), .A2(
        \SB2_3_27/i0[10] ), .A3(\SB2_3_27/i0[6] ), .ZN(
        \SB2_3_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_27/Component_Function_2/N1  ( .A1(n1630), .A2(
        \SB2_3_27/i0[10] ), .A3(\SB2_3_27/i1[9] ), .ZN(
        \SB2_3_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_3/N3  ( .A1(\SB2_3_27/i1[9] ), .A2(
        \SB2_3_27/i1_7 ), .A3(\SB2_3_27/i0[10] ), .ZN(
        \SB2_3_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_27/Component_Function_3/N2  ( .A1(\SB2_3_27/i0_0 ), .A2(
        \SB2_3_27/i0_3 ), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_27/Component_Function_3/N1  ( .A1(\SB2_3_27/i1[9] ), .A2(
        \SB2_3_27/i0_3 ), .A3(\SB2_3_27/i0[6] ), .ZN(
        \SB2_3_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N4  ( .A1(\SB2_3_27/i1[9] ), .A2(
        n1630), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N3  ( .A1(\SB2_3_27/i0[9] ), .A2(
        \SB2_3_27/i0[10] ), .A3(\SB2_3_27/i0_3 ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N2  ( .A1(\SB2_3_27/i3[0] ), .A2(
        \SB2_3_27/i0_0 ), .A3(\SB2_3_27/i1_7 ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N1  ( .A1(\SB2_3_27/i0[9] ), .A2(
        \SB2_3_27/i0_0 ), .A3(\SB2_3_27/i0[8] ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_2/N4  ( .A1(\SB2_3_28/i1_5 ), .A2(
        \SB2_3_28/i0_0 ), .A3(\SB2_3_28/i0_4 ), .ZN(
        \SB2_3_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_28/Component_Function_2/N3  ( .A1(\SB2_3_28/i0_3 ), .A2(
        \SB2_3_28/i0[8] ), .A3(\SB2_3_28/i0[9] ), .ZN(
        \SB2_3_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_28/Component_Function_2/N2  ( .A1(\SB2_3_28/i0_3 ), .A2(
        \SB2_3_28/i0[10] ), .A3(\SB2_3_28/i0[6] ), .ZN(
        \SB2_3_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_28/Component_Function_3/N3  ( .A1(\SB2_3_28/i1[9] ), .A2(
        \SB2_3_28/i1_7 ), .A3(\SB2_3_28/i0[10] ), .ZN(
        \SB2_3_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_28/Component_Function_3/N2  ( .A1(\SB2_3_28/i0_0 ), .A2(
        \SB2_3_28/i0_3 ), .A3(\SB2_3_28/i0_4 ), .ZN(
        \SB2_3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_28/Component_Function_3/N1  ( .A1(\SB2_3_28/i1[9] ), .A2(
        \SB2_3_28/i0_3 ), .A3(\SB2_3_28/i0[6] ), .ZN(
        \SB2_3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_4/N4  ( .A1(\SB2_3_28/i1[9] ), .A2(
        \SB2_3_28/i1_5 ), .A3(\SB2_3_28/i0_4 ), .ZN(
        \SB2_3_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_28/Component_Function_4/N3  ( .A1(\SB2_3_28/i0[9] ), .A2(
        \SB2_3_28/i0[10] ), .A3(\SB2_3_28/i0_3 ), .ZN(
        \SB2_3_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_28/Component_Function_4/N2  ( .A1(\SB2_3_28/i3[0] ), .A2(
        \SB2_3_28/i0_0 ), .A3(\SB2_3_28/i1_7 ), .ZN(
        \SB2_3_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_28/Component_Function_4/N1  ( .A1(\SB2_3_28/i0[9] ), .A2(
        \SB2_3_28/i0_0 ), .A3(\SB2_3_28/i0[8] ), .ZN(
        \SB2_3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_29/Component_Function_2/N4  ( .A1(\SB2_3_29/i1_5 ), .A2(
        \SB2_3_29/i0_0 ), .A3(\SB2_3_29/i0_4 ), .ZN(
        \SB2_3_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_29/Component_Function_2/N3  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i0[8] ), .A3(\SB2_3_29/i0[9] ), .ZN(
        \SB2_3_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_29/Component_Function_2/N2  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i0[10] ), .A3(n2115), .ZN(
        \SB2_3_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_29/Component_Function_3/N4  ( .A1(\SB2_3_29/i1_5 ), .A2(
        \SB2_3_29/i0[8] ), .A3(\SB2_3_29/i3[0] ), .ZN(
        \SB2_3_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_29/Component_Function_3/N3  ( .A1(\SB2_3_29/i1[9] ), .A2(
        \SB2_3_29/i1_7 ), .A3(\SB2_3_29/i0[10] ), .ZN(
        \SB2_3_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_29/Component_Function_3/N2  ( .A1(\SB2_3_29/i0_0 ), .A2(
        \SB2_3_29/i0_3 ), .A3(\SB2_3_29/i0_4 ), .ZN(
        \SB2_3_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_29/Component_Function_3/N1  ( .A1(\SB2_3_29/i1[9] ), .A2(
        \SB2_3_29/i0_3 ), .A3(n2115), .ZN(
        \SB2_3_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_29/Component_Function_4/N4  ( .A1(\SB2_3_29/i1[9] ), .A2(
        \SB2_3_29/i1_5 ), .A3(\SB2_3_29/i0_4 ), .ZN(
        \SB2_3_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_29/Component_Function_4/N3  ( .A1(\SB2_3_29/i0[9] ), .A2(
        \SB2_3_29/i0[10] ), .A3(\SB2_3_29/i0_3 ), .ZN(
        \SB2_3_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_29/Component_Function_4/N2  ( .A1(\SB2_3_29/i3[0] ), .A2(
        \SB2_3_29/i0_0 ), .A3(\SB2_3_29/i1_7 ), .ZN(
        \SB2_3_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_29/Component_Function_4/N1  ( .A1(\SB2_3_29/i0[9] ), .A2(
        \SB2_3_29/i0_0 ), .A3(\SB2_3_29/i0[8] ), .ZN(
        \SB2_3_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_2/N4  ( .A1(\SB2_3_30/i1_5 ), .A2(
        \SB2_3_30/i0_0 ), .A3(\SB2_3_30/i0_4 ), .ZN(
        \SB2_3_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_30/Component_Function_2/N2  ( .A1(\SB2_3_30/i0_3 ), .A2(
        \SB2_3_30/i0[10] ), .A3(\SB2_3_30/i0[6] ), .ZN(
        \SB2_3_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_30/Component_Function_2/N1  ( .A1(\SB2_3_30/i1_5 ), .A2(
        \SB2_3_30/i0[10] ), .A3(\SB2_3_30/i1[9] ), .ZN(
        \SB2_3_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_3/N4  ( .A1(\SB2_3_30/i1_5 ), .A2(
        \SB2_3_30/i0[8] ), .A3(\SB2_3_30/i3[0] ), .ZN(
        \SB2_3_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_30/Component_Function_3/N3  ( .A1(\SB2_3_30/i1[9] ), .A2(
        \SB2_3_30/i1_7 ), .A3(\SB2_3_30/i0[10] ), .ZN(
        \SB2_3_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_30/Component_Function_3/N2  ( .A1(\SB2_3_30/i0_0 ), .A2(
        \SB2_3_30/i0_3 ), .A3(\SB2_3_30/i0_4 ), .ZN(
        \SB2_3_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_30/Component_Function_3/N1  ( .A1(\SB2_3_30/i1[9] ), .A2(
        \SB2_3_30/i0_3 ), .A3(\SB2_3_30/i0[6] ), .ZN(
        \SB2_3_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N4  ( .A1(\SB2_3_30/i1[9] ), .A2(
        \SB2_3_30/i1_5 ), .A3(\SB2_3_30/i0_4 ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N3  ( .A1(\SB2_3_30/i0[9] ), .A2(
        \SB2_3_30/i0[10] ), .A3(\SB2_3_30/i0_3 ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N2  ( .A1(\SB2_3_30/i3[0] ), .A2(
        \SB2_3_30/i0_0 ), .A3(\SB2_3_30/i1_7 ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N1  ( .A1(\SB2_3_30/i0[9] ), .A2(
        \SB2_3_30/i0_0 ), .A3(\SB2_3_30/i0[8] ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_2/N3  ( .A1(\SB2_3_31/i0_3 ), .A2(
        \SB2_3_31/i0[8] ), .A3(\SB2_3_31/i0[9] ), .ZN(
        \SB2_3_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_31/Component_Function_2/N2  ( .A1(\SB2_3_31/i0_3 ), .A2(
        \SB2_3_31/i0[10] ), .A3(\SB2_3_31/i0[6] ), .ZN(
        \SB2_3_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_31/Component_Function_2/N1  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0[10] ), .A3(\SB2_3_31/i1[9] ), .ZN(
        \SB2_3_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_3/N3  ( .A1(\SB2_3_31/i1[9] ), .A2(
        \SB2_3_31/i1_7 ), .A3(\SB2_3_31/i0[10] ), .ZN(
        \SB2_3_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_31/Component_Function_3/N2  ( .A1(\SB2_3_31/i0_0 ), .A2(
        \SB2_3_31/i0_3 ), .A3(n1651), .ZN(
        \SB2_3_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_31/Component_Function_3/N1  ( .A1(\SB2_3_31/i1[9] ), .A2(
        \SB2_3_31/i0_3 ), .A3(\SB2_3_31/i0[6] ), .ZN(
        \SB2_3_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_4/N4  ( .A1(\SB2_3_31/i1[9] ), .A2(
        \SB2_3_31/i1_5 ), .A3(n1652), .ZN(
        \SB2_3_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_31/Component_Function_4/N3  ( .A1(\SB2_3_31/i0[9] ), .A2(
        \SB2_3_31/i0[10] ), .A3(\SB2_3_31/i0_3 ), .ZN(
        \SB2_3_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_31/Component_Function_4/N2  ( .A1(\SB2_3_31/i3[0] ), .A2(
        \SB2_3_31/i0_0 ), .A3(\SB2_3_31/i1_7 ), .ZN(
        \SB2_3_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_31/Component_Function_4/N1  ( .A1(\SB2_3_31/i0[9] ), .A2(
        \SB2_3_31/i0_0 ), .A3(\SB2_3_31/i0[8] ), .ZN(
        \SB2_3_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_2/N3  ( .A1(\SB3_0/i0_3 ), .A2(
        \SB3_0/i0[8] ), .A3(\SB3_0/i0[9] ), .ZN(
        \SB3_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_0/Component_Function_2/N2  ( .A1(\SB3_0/i0_3 ), .A2(
        \SB3_0/i0[10] ), .A3(\SB3_0/i0[6] ), .ZN(
        \SB3_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_0/Component_Function_2/N1  ( .A1(\SB3_0/i1_5 ), .A2(
        \SB3_0/i0[10] ), .A3(\SB3_0/i1[9] ), .ZN(
        \SB3_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_3/N3  ( .A1(\SB3_0/i1[9] ), .A2(
        \SB3_0/i1_7 ), .A3(\SB3_0/i0[10] ), .ZN(
        \SB3_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_0/Component_Function_3/N2  ( .A1(\SB3_0/i0_0 ), .A2(
        \SB3_0/i0_3 ), .A3(\SB3_0/i0_4 ), .ZN(
        \SB3_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_0/Component_Function_3/N1  ( .A1(\SB3_0/i1[9] ), .A2(
        \SB3_0/i0_3 ), .A3(\SB3_0/i0[6] ), .ZN(
        \SB3_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_4/N2  ( .A1(\SB3_0/i3[0] ), .A2(
        \SB3_0/i0_0 ), .A3(\SB3_0/i1_7 ), .ZN(
        \SB3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_0/Component_Function_4/N1  ( .A1(\SB3_0/i0[9] ), .A2(
        \SB3_0/i0_0 ), .A3(\SB3_0/i0[8] ), .ZN(
        \SB3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_2/N4  ( .A1(\SB3_1/i1_5 ), .A2(
        \SB3_1/i0_0 ), .A3(\SB3_1/i0_4 ), .ZN(
        \SB3_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_1/Component_Function_2/N3  ( .A1(n856), .A2(\SB3_1/i0[8] ), 
        .A3(\SB3_1/i0[9] ), .ZN(\SB3_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_1/Component_Function_2/N2  ( .A1(n856), .A2(\SB3_1/i0[10] ), 
        .A3(\SB3_1/i0[6] ), .ZN(\SB3_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_1/Component_Function_2/N1  ( .A1(\SB3_1/i1_5 ), .A2(
        \SB3_1/i0[10] ), .A3(\SB3_1/i1[9] ), .ZN(
        \SB3_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_3/N4  ( .A1(\SB3_1/i1_5 ), .A2(
        \SB3_1/i0[8] ), .A3(\SB3_1/i3[0] ), .ZN(
        \SB3_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_1/Component_Function_3/N3  ( .A1(\SB3_1/i1[9] ), .A2(
        \SB3_1/i1_7 ), .A3(\SB3_1/i0[10] ), .ZN(
        \SB3_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_1/Component_Function_3/N2  ( .A1(\SB3_1/i0_0 ), .A2(
        \SB3_1/i0_3 ), .A3(\SB3_1/i0_4 ), .ZN(
        \SB3_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_1/Component_Function_3/N1  ( .A1(\SB3_1/i1[9] ), .A2(n856), 
        .A3(\SB3_1/i0[6] ), .ZN(\SB3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_4/N4  ( .A1(\SB3_1/i1[9] ), .A2(
        \SB3_1/i1_5 ), .A3(\SB3_1/i0_4 ), .ZN(
        \SB3_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_1/Component_Function_4/N3  ( .A1(\SB3_1/i0[9] ), .A2(
        \SB3_1/i0[10] ), .A3(\SB3_1/i0_3 ), .ZN(
        \SB3_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_1/Component_Function_4/N2  ( .A1(\SB3_1/i3[0] ), .A2(
        \SB3_1/i0_0 ), .A3(\SB3_1/i1_7 ), .ZN(
        \SB3_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_1/Component_Function_4/N1  ( .A1(\SB3_1/i0[9] ), .A2(
        \SB3_1/i0_0 ), .A3(\SB3_1/i0[8] ), .ZN(
        \SB3_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_2/N3  ( .A1(\SB3_2/i0_3 ), .A2(
        \SB3_2/i0[8] ), .A3(\SB3_2/i0[9] ), .ZN(
        \SB3_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_2/Component_Function_2/N2  ( .A1(\SB3_2/i0_3 ), .A2(
        \SB3_2/i0[10] ), .A3(\SB3_2/i0[6] ), .ZN(
        \SB3_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_2/Component_Function_2/N1  ( .A1(\SB3_2/i1_5 ), .A2(
        \SB3_2/i0[10] ), .A3(\SB3_2/i1[9] ), .ZN(
        \SB3_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_3/N4  ( .A1(\SB3_2/i1_5 ), .A2(
        \SB3_2/i0[8] ), .A3(\SB3_2/i3[0] ), .ZN(
        \SB3_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_2/Component_Function_3/N3  ( .A1(\SB3_2/i1[9] ), .A2(
        \SB3_2/i1_7 ), .A3(\SB3_2/i0[10] ), .ZN(
        \SB3_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_2/Component_Function_3/N1  ( .A1(\SB3_2/i1[9] ), .A2(
        \SB3_2/i0_3 ), .A3(\SB3_2/i0[6] ), .ZN(
        \SB3_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_4/N2  ( .A1(\SB3_2/i3[0] ), .A2(
        \SB3_2/i0_0 ), .A3(\SB3_2/i1_7 ), .ZN(
        \SB3_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_2/Component_Function_4/N1  ( .A1(\SB3_2/i0[9] ), .A2(
        \SB3_2/i0_0 ), .A3(\SB3_2/i0[8] ), .ZN(
        \SB3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_2/N3  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i0[8] ), .A3(\SB3_3/i0[9] ), .ZN(
        \SB3_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_3/Component_Function_2/N2  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i0[10] ), .A3(\SB3_3/i0[6] ), .ZN(
        \SB3_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_3/Component_Function_2/N1  ( .A1(\SB3_3/i1_5 ), .A2(
        \SB3_3/i0[10] ), .A3(\SB3_3/i1[9] ), .ZN(
        \SB3_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_3/N4  ( .A1(\SB3_3/i1_5 ), .A2(
        \SB3_3/i0[8] ), .A3(\SB3_3/i3[0] ), .ZN(
        \SB3_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_3/Component_Function_3/N3  ( .A1(\SB3_3/i1[9] ), .A2(
        \SB3_3/i1_7 ), .A3(\SB3_3/i0[10] ), .ZN(
        \SB3_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_3/Component_Function_3/N2  ( .A1(\SB3_3/i0_0 ), .A2(
        \SB3_3/i0_3 ), .A3(\SB3_3/i0_4 ), .ZN(
        \SB3_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_3/Component_Function_3/N1  ( .A1(\SB3_3/i1[9] ), .A2(
        \SB3_3/i0_3 ), .A3(\SB3_3/i0[6] ), .ZN(
        \SB3_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N4  ( .A1(\SB3_3/i1[9] ), .A2(
        \SB3_3/i1_5 ), .A3(\SB3_3/i0_4 ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N2  ( .A1(\SB3_3/i3[0] ), .A2(
        \SB3_3/i0_0 ), .A3(\SB3_3/i1_7 ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N1  ( .A1(\SB3_3/i0[9] ), .A2(
        \SB3_3/i0_0 ), .A3(\SB3_3/i0[8] ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_2/N4  ( .A1(\SB3_4/i1_5 ), .A2(
        \SB3_4/i0_0 ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_2/N2  ( .A1(\SB3_4/i0_3 ), .A2(
        \SB3_4/i0[10] ), .A3(\SB3_4/i0[6] ), .ZN(
        \SB3_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_4/Component_Function_2/N1  ( .A1(\SB3_4/i1_5 ), .A2(
        \SB3_4/i0[10] ), .A3(\SB3_4/i1[9] ), .ZN(
        \SB3_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_3/N4  ( .A1(\SB3_4/i1_5 ), .A2(
        \SB3_4/i0[8] ), .A3(\SB3_4/i3[0] ), .ZN(
        \SB3_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_3/N3  ( .A1(\SB3_4/i1[9] ), .A2(
        \SB3_4/i1_7 ), .A3(\SB3_4/i0[10] ), .ZN(
        \SB3_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_4/Component_Function_3/N1  ( .A1(\SB3_4/i1[9] ), .A2(
        \SB3_4/i0_3 ), .A3(\SB3_4/i0[6] ), .ZN(
        \SB3_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N4  ( .A1(\SB3_4/i1[9] ), .A2(
        \SB3_4/i1_5 ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N2  ( .A1(\SB3_4/i3[0] ), .A2(
        \SB3_4/i0_0 ), .A3(\SB3_4/i1_7 ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N1  ( .A1(\SB3_4/i0[9] ), .A2(
        \SB3_4/i0_0 ), .A3(\SB3_4/i0[8] ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_2/N3  ( .A1(\SB3_5/i0_3 ), .A2(
        \SB3_5/i0[8] ), .A3(\SB3_5/i0[9] ), .ZN(
        \SB3_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_5/Component_Function_2/N2  ( .A1(\SB3_5/i0_3 ), .A2(
        \SB3_5/i0[10] ), .A3(\SB3_5/i0[6] ), .ZN(
        \SB3_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_5/Component_Function_2/N1  ( .A1(\SB3_5/i1_5 ), .A2(
        \SB3_5/i0[10] ), .A3(\SB3_5/i1[9] ), .ZN(
        \SB3_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_3/N3  ( .A1(\SB3_5/i1[9] ), .A2(
        \SB3_5/i1_7 ), .A3(\SB3_5/i0[10] ), .ZN(
        \SB3_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_5/Component_Function_3/N2  ( .A1(\SB3_5/i0_0 ), .A2(
        \SB3_5/i0_3 ), .A3(\SB3_5/i0_4 ), .ZN(
        \SB3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_5/Component_Function_3/N1  ( .A1(\SB3_5/i1[9] ), .A2(
        \SB3_5/i0_3 ), .A3(\SB3_5/i0[6] ), .ZN(
        \SB3_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_4/N4  ( .A1(\SB3_5/i1[9] ), .A2(
        \SB3_5/i1_5 ), .A3(\SB3_5/i0_4 ), .ZN(
        \SB3_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_5/Component_Function_4/N2  ( .A1(\SB3_5/i3[0] ), .A2(
        \SB3_5/i0_0 ), .A3(\SB3_5/i1_7 ), .ZN(
        \SB3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_5/Component_Function_4/N1  ( .A1(\SB3_5/i0[9] ), .A2(
        \SB3_5/i0_0 ), .A3(\SB3_5/i0[8] ), .ZN(
        \SB3_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_2/N4  ( .A1(\SB3_6/i1_5 ), .A2(
        \SB3_6/i0_0 ), .A3(\SB3_6/i0_4 ), .ZN(
        \SB3_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_2/N2  ( .A1(n833), .A2(\SB3_6/i0[10] ), 
        .A3(\SB3_6/i0[6] ), .ZN(\SB3_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_6/Component_Function_2/N1  ( .A1(\SB3_6/i1_5 ), .A2(
        \SB3_6/i0[10] ), .A3(\SB3_6/i1[9] ), .ZN(
        \SB3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_3/N4  ( .A1(\SB3_6/i1_5 ), .A2(
        \SB3_6/i0[8] ), .A3(\SB3_6/i3[0] ), .ZN(
        \SB3_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_3/N3  ( .A1(\SB3_6/i1[9] ), .A2(
        \SB3_6/i1_7 ), .A3(\SB3_6/i0[10] ), .ZN(
        \SB3_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_6/Component_Function_3/N2  ( .A1(\SB3_6/i0_0 ), .A2(
        \SB3_6/i0_3 ), .A3(\SB3_6/i0_4 ), .ZN(
        \SB3_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_6/Component_Function_3/N1  ( .A1(\SB3_6/i1[9] ), .A2(n833), 
        .A3(\SB3_6/i0[6] ), .ZN(\SB3_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_4/N4  ( .A1(\SB3_6/i1[9] ), .A2(
        \SB3_6/i1_5 ), .A3(\SB3_6/i0_4 ), .ZN(
        \SB3_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_4/N3  ( .A1(\SB3_6/i0[9] ), .A2(
        \SB3_6/i0[10] ), .A3(\SB3_6/i0_3 ), .ZN(
        \SB3_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_6/Component_Function_4/N2  ( .A1(\SB3_6/i3[0] ), .A2(
        \SB3_6/i0_0 ), .A3(\SB3_6/i1_7 ), .ZN(
        \SB3_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_6/Component_Function_4/N1  ( .A1(\SB3_6/i0[9] ), .A2(
        \SB3_6/i0_0 ), .A3(\SB3_6/i0[8] ), .ZN(
        \SB3_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_2/N3  ( .A1(\SB3_7/i0_3 ), .A2(n798), 
        .A3(\SB3_7/i0[9] ), .ZN(\SB3_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_7/Component_Function_2/N2  ( .A1(\SB3_7/i0[10] ), .A2(
        \SB3_7/i0_3 ), .A3(\SB3_7/i0[6] ), .ZN(
        \SB3_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_7/Component_Function_2/N1  ( .A1(\SB3_7/i1_5 ), .A2(
        \SB3_7/i0[10] ), .A3(\SB3_7/i1[9] ), .ZN(
        \SB3_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_3/N4  ( .A1(\SB3_7/i1_5 ), .A2(n798), 
        .A3(\SB3_7/i3[0] ), .ZN(\SB3_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_7/Component_Function_3/N2  ( .A1(\SB3_7/i0_0 ), .A2(
        \SB3_7/i0_3 ), .A3(\SB3_7/i0_4 ), .ZN(
        \SB3_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_7/Component_Function_3/N1  ( .A1(\SB3_7/i1[9] ), .A2(
        \SB3_7/i0_3 ), .A3(\SB3_7/i0[6] ), .ZN(
        \SB3_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_4/N4  ( .A1(\SB3_7/i1[9] ), .A2(
        \SB3_7/i1_5 ), .A3(\SB3_7/i0_4 ), .ZN(
        \SB3_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_7/Component_Function_4/N2  ( .A1(\SB3_7/i3[0] ), .A2(
        \SB3_7/i0_0 ), .A3(\SB3_7/i1_7 ), .ZN(
        \SB3_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_7/Component_Function_4/N1  ( .A1(\SB3_7/i0[9] ), .A2(
        \SB3_7/i0_0 ), .A3(n798), .ZN(\SB3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_2/N4  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0_0 ), .A3(\SB3_8/i0_4 ), .ZN(
        \SB3_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_2/N3  ( .A1(\SB3_8/i0_3 ), .A2(
        \SB3_8/i0[8] ), .A3(\SB3_8/i0[9] ), .ZN(
        \SB3_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_8/Component_Function_2/N2  ( .A1(\SB3_8/i0_3 ), .A2(
        \SB3_8/i0[10] ), .A3(\SB3_8/i0[6] ), .ZN(
        \SB3_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_8/Component_Function_2/N1  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[10] ), .A3(\SB3_8/i1[9] ), .ZN(
        \SB3_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_3/N4  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[8] ), .A3(\SB3_8/i3[0] ), .ZN(
        \SB3_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_3/N3  ( .A1(\SB3_8/i1[9] ), .A2(
        \SB3_8/i1_7 ), .A3(\SB3_8/i0[10] ), .ZN(
        \SB3_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_8/Component_Function_3/N2  ( .A1(\SB3_8/i0_0 ), .A2(
        \SB3_8/i0_3 ), .A3(\SB3_8/i0_4 ), .ZN(
        \SB3_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_8/Component_Function_3/N1  ( .A1(\SB3_8/i1[9] ), .A2(
        \SB3_8/i0_3 ), .A3(\SB3_8/i0[6] ), .ZN(
        \SB3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_4/N4  ( .A1(\SB3_8/i1[9] ), .A2(
        \SB3_8/i1_5 ), .A3(\SB3_8/i0_4 ), .ZN(
        \SB3_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_4/N2  ( .A1(\SB3_8/i3[0] ), .A2(
        \SB3_8/i0_0 ), .A3(\SB3_8/i1_7 ), .ZN(
        \SB3_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_8/Component_Function_4/N1  ( .A1(\SB3_8/i0[9] ), .A2(
        \SB3_8/i0_0 ), .A3(\SB3_8/i0[8] ), .ZN(
        \SB3_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_2/N3  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i0[8] ), .A3(\SB3_9/i0[9] ), .ZN(
        \SB3_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_9/Component_Function_2/N2  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i0[10] ), .A3(\SB3_9/i0[6] ), .ZN(
        \SB3_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_2/N1  ( .A1(\SB3_9/i1_5 ), .A2(
        \SB3_9/i0[10] ), .A3(\SB3_9/i1[9] ), .ZN(
        \SB3_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_3/N4  ( .A1(\SB3_9/i1_5 ), .A2(
        \SB3_9/i0[8] ), .A3(\SB3_9/i3[0] ), .ZN(
        \SB3_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_3/N3  ( .A1(\SB3_9/i1[9] ), .A2(
        \SB3_9/i1_7 ), .A3(\SB3_9/i0[10] ), .ZN(
        \SB3_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_9/Component_Function_3/N2  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i0_3 ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_3/N1  ( .A1(\SB3_9/i1[9] ), .A2(
        \SB3_9/i0_3 ), .A3(\SB3_9/i0[6] ), .ZN(
        \SB3_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N4  ( .A1(\SB3_9/i1[9] ), .A2(
        \SB3_9/i1_5 ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N2  ( .A1(\SB3_9/i3[0] ), .A2(
        \SB3_9/i0_0 ), .A3(\SB3_9/i1_7 ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N1  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i0[9] ), .A3(\SB3_9/i0[8] ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_2/N4  ( .A1(\SB3_10/i1_5 ), .A2(
        \SB3_10/i0_0 ), .A3(\SB3_10/i0_4 ), .ZN(
        \SB3_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_10/Component_Function_2/N3  ( .A1(n835), .A2(\SB3_10/i0[8] ), 
        .A3(\SB3_10/i0[9] ), .ZN(\SB3_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_10/Component_Function_2/N2  ( .A1(n835), .A2(\SB3_10/i0[10] ), 
        .A3(\SB3_10/i0[6] ), .ZN(\SB3_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_10/Component_Function_2/N1  ( .A1(\SB3_10/i1_5 ), .A2(
        \SB3_10/i0[10] ), .A3(\SB3_10/i1[9] ), .ZN(
        \SB3_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_3/N3  ( .A1(\SB3_10/i1[9] ), .A2(
        \SB3_10/i1_7 ), .A3(\SB3_10/i0[10] ), .ZN(
        \SB3_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_10/Component_Function_3/N2  ( .A1(\SB3_10/i0_0 ), .A2(
        \SB3_10/i0_3 ), .A3(\SB3_10/i0_4 ), .ZN(
        \SB3_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_10/Component_Function_3/N1  ( .A1(\SB3_10/i1[9] ), .A2(n835), 
        .A3(\SB3_10/i0[6] ), .ZN(\SB3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_4/N4  ( .A1(\SB3_10/i1[9] ), .A2(
        \SB3_10/i1_5 ), .A3(\SB3_10/i0_4 ), .ZN(
        \SB3_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_10/Component_Function_4/N2  ( .A1(\SB3_10/i3[0] ), .A2(
        \SB3_10/i0_0 ), .A3(\SB3_10/i1_7 ), .ZN(
        \SB3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_10/Component_Function_4/N1  ( .A1(\SB3_10/i0[9] ), .A2(
        \SB3_10/i0_0 ), .A3(\SB3_10/i0[8] ), .ZN(
        \SB3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_2/N4  ( .A1(\SB3_11/i1_5 ), .A2(
        \SB3_11/i0_0 ), .A3(\SB3_11/i0_4 ), .ZN(
        \SB3_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_11/Component_Function_2/N3  ( .A1(n840), .A2(\SB3_11/i0[8] ), 
        .A3(\SB3_11/i0[9] ), .ZN(\SB3_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_11/Component_Function_2/N2  ( .A1(n840), .A2(\SB3_11/i0[10] ), 
        .A3(\SB3_11/i0[6] ), .ZN(\SB3_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_11/Component_Function_2/N1  ( .A1(\SB3_11/i1_5 ), .A2(
        \SB3_11/i0[10] ), .A3(\SB3_11/i1[9] ), .ZN(
        \SB3_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_3/N3  ( .A1(\SB3_11/i1[9] ), .A2(
        \SB3_11/i1_7 ), .A3(\SB3_11/i0[10] ), .ZN(
        \SB3_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_11/Component_Function_3/N2  ( .A1(\SB3_11/i0_0 ), .A2(
        \SB3_11/i0_3 ), .A3(\SB3_11/i0_4 ), .ZN(
        \SB3_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_11/Component_Function_3/N1  ( .A1(\SB3_11/i1[9] ), .A2(n840), 
        .A3(\SB3_11/i0[6] ), .ZN(\SB3_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_4/N4  ( .A1(\SB3_11/i1[9] ), .A2(
        \SB3_11/i1_5 ), .A3(\SB3_11/i0_4 ), .ZN(
        \SB3_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_11/Component_Function_4/N3  ( .A1(\SB3_11/i0[9] ), .A2(
        \SB3_11/i0[10] ), .A3(\SB3_11/i0_3 ), .ZN(
        \SB3_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_11/Component_Function_4/N2  ( .A1(\SB3_11/i3[0] ), .A2(
        \SB3_11/i0_0 ), .A3(\SB3_11/i1_7 ), .ZN(
        \SB3_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_11/Component_Function_4/N1  ( .A1(\SB3_11/i0[9] ), .A2(
        \SB3_11/i0_0 ), .A3(\SB3_11/i0[8] ), .ZN(
        \SB3_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_2/N4  ( .A1(\SB3_12/i1_5 ), .A2(
        \SB3_12/i0_0 ), .A3(\SB3_12/i0_4 ), .ZN(
        \SB3_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_12/Component_Function_2/N2  ( .A1(\SB3_12/i0_3 ), .A2(
        \SB3_12/i0[10] ), .A3(\SB3_12/i0[6] ), .ZN(
        \SB3_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_12/Component_Function_2/N1  ( .A1(\SB3_12/i1_5 ), .A2(
        \SB3_12/i0[10] ), .A3(\SB3_12/i1[9] ), .ZN(
        \SB3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_3/N4  ( .A1(\SB3_12/i1_5 ), .A2(
        \SB3_12/i0[8] ), .A3(\SB3_12/i3[0] ), .ZN(
        \SB3_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_12/Component_Function_3/N3  ( .A1(\SB3_12/i1[9] ), .A2(
        \SB3_12/i1_7 ), .A3(\SB3_12/i0[10] ), .ZN(
        \SB3_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_12/Component_Function_3/N1  ( .A1(\SB3_12/i1[9] ), .A2(
        \SB3_12/i0_3 ), .A3(\SB3_12/i0[6] ), .ZN(
        \SB3_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_4/N4  ( .A1(\SB3_12/i1[9] ), .A2(
        \SB3_12/i1_5 ), .A3(\SB3_12/i0_4 ), .ZN(
        \SB3_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_12/Component_Function_4/N3  ( .A1(\SB3_12/i0_3 ), .A2(
        \SB3_12/i0[10] ), .A3(\SB3_12/i0[9] ), .ZN(
        \SB3_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_12/Component_Function_4/N2  ( .A1(\SB3_12/i3[0] ), .A2(
        \SB3_12/i0_0 ), .A3(\SB3_12/i1_7 ), .ZN(
        \SB3_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_12/Component_Function_4/N1  ( .A1(\SB3_12/i0[9] ), .A2(
        \SB3_12/i0_0 ), .A3(\SB3_12/i0[8] ), .ZN(
        \SB3_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_2/N4  ( .A1(\SB3_13/i1_5 ), .A2(
        \SB3_13/i0_0 ), .A3(\SB3_13/i0_4 ), .ZN(
        \SB3_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_2/N3  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i0[8] ), .A3(\SB3_13/i0[9] ), .ZN(
        \SB3_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_13/Component_Function_2/N2  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i0[10] ), .A3(\SB3_13/i0[6] ), .ZN(
        \SB3_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_13/Component_Function_2/N1  ( .A1(\SB3_13/i1_5 ), .A2(
        \SB3_13/i0[10] ), .A3(\SB3_13/i1[9] ), .ZN(
        \SB3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_3/N4  ( .A1(\SB3_13/i1_5 ), .A2(
        \SB3_13/i0[8] ), .A3(\SB3_13/i3[0] ), .ZN(
        \SB3_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_3/N2  ( .A1(\SB3_13/i0_0 ), .A2(
        \SB3_13/i0_3 ), .A3(\SB3_13/i0_4 ), .ZN(
        \SB3_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_13/Component_Function_3/N1  ( .A1(\SB3_13/i1[9] ), .A2(
        \SB3_13/i0_3 ), .A3(\SB3_13/i0[6] ), .ZN(
        \SB3_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_4/N4  ( .A1(\SB3_13/i1[9] ), .A2(
        \SB3_13/i1_5 ), .A3(\SB3_13/i0_4 ), .ZN(
        \SB3_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_4/N2  ( .A1(\SB3_13/i3[0] ), .A2(
        \SB3_13/i0_0 ), .A3(\SB3_13/i1_7 ), .ZN(
        \SB3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_13/Component_Function_4/N1  ( .A1(\SB3_13/i0[9] ), .A2(
        \SB3_13/i0_0 ), .A3(\SB3_13/i0[8] ), .ZN(
        \SB3_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_2/N3  ( .A1(\SB3_14/i0_3 ), .A2(
        \SB3_14/i0[8] ), .A3(\SB3_14/i0[9] ), .ZN(
        \SB3_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_2/N2  ( .A1(n860), .A2(\SB3_14/i0[10] ), 
        .A3(\SB3_14/i0[6] ), .ZN(\SB3_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_14/Component_Function_2/N1  ( .A1(\SB3_14/i1_5 ), .A2(
        \SB3_14/i0[10] ), .A3(\SB3_14/i1[9] ), .ZN(
        \SB3_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_3/N3  ( .A1(\SB3_14/i1[9] ), .A2(
        \SB3_14/i1_7 ), .A3(\SB3_14/i0[10] ), .ZN(
        \SB3_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_3/N2  ( .A1(\SB3_14/i0_0 ), .A2(
        \SB3_14/i0_3 ), .A3(\SB3_14/i0_4 ), .ZN(
        \SB3_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_14/Component_Function_3/N1  ( .A1(\SB3_14/i1[9] ), .A2(n860), 
        .A3(\SB3_14/i0[6] ), .ZN(\SB3_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N4  ( .A1(\SB3_14/i1[9] ), .A2(
        \SB3_14/i1_5 ), .A3(\SB3_14/i0_4 ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N3  ( .A1(\SB3_14/i0[9] ), .A2(
        \SB3_14/i0[10] ), .A3(\SB3_14/i0_3 ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N2  ( .A1(\SB3_14/i3[0] ), .A2(
        \SB3_14/i0_0 ), .A3(\SB3_14/i1_7 ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N1  ( .A1(\SB3_14/i0[9] ), .A2(
        \SB3_14/i0_0 ), .A3(\SB3_14/i0[8] ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_15/Component_Function_2/N3  ( .A1(\SB3_15/i0_3 ), .A2(
        \SB3_15/i0[8] ), .A3(\SB3_15/i0[9] ), .ZN(
        \SB3_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_2/N2  ( .A1(\SB3_15/i0[10] ), .A2(
        \SB3_15/i0_3 ), .A3(\SB3_15/i0[6] ), .ZN(
        \SB3_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_15/Component_Function_2/N1  ( .A1(\SB3_15/i1_5 ), .A2(
        \SB3_15/i0[10] ), .A3(\SB3_15/i1[9] ), .ZN(
        \SB3_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_15/Component_Function_3/N4  ( .A1(\SB3_15/i1_5 ), .A2(
        \SB3_15/i0[8] ), .A3(\SB3_15/i3[0] ), .ZN(
        \SB3_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_15/Component_Function_3/N3  ( .A1(\SB3_15/i1[9] ), .A2(
        \SB3_15/i1_7 ), .A3(\SB3_15/i0[10] ), .ZN(
        \SB3_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_3/N2  ( .A1(\SB3_15/i0_0 ), .A2(
        \SB3_15/i0_3 ), .A3(\SB3_15/i0_4 ), .ZN(
        \SB3_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_15/Component_Function_3/N1  ( .A1(\SB3_15/i1[9] ), .A2(
        \SB3_15/i0_3 ), .A3(\SB3_15/i0[6] ), .ZN(
        \SB3_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_15/Component_Function_4/N4  ( .A1(\SB3_15/i1[9] ), .A2(
        \SB3_15/i1_5 ), .A3(\SB3_15/i0_4 ), .ZN(
        \SB3_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_15/Component_Function_4/N3  ( .A1(\SB3_15/i0[9] ), .A2(
        \SB3_15/i0[10] ), .A3(\SB3_15/i0_3 ), .ZN(
        \SB3_15/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_4/N2  ( .A1(\SB3_15/i3[0] ), .A2(
        \SB3_15/i0_0 ), .A3(\SB3_15/i1_7 ), .ZN(
        \SB3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_15/Component_Function_4/N1  ( .A1(\SB3_15/i0[9] ), .A2(
        \SB3_15/i0_0 ), .A3(\SB3_15/i0[8] ), .ZN(
        \SB3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_2/N4  ( .A1(\SB3_16/i1_5 ), .A2(
        \SB3_16/i0_0 ), .A3(\SB3_16/i0_4 ), .ZN(
        \SB3_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_16/Component_Function_2/N3  ( .A1(\SB3_16/i0_3 ), .A2(
        \SB3_16/i0[8] ), .A3(\SB3_16/i0[9] ), .ZN(
        \SB3_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_16/Component_Function_2/N2  ( .A1(n876), .A2(\SB3_16/i0[10] ), 
        .A3(\SB3_16/i0[6] ), .ZN(\SB3_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_2/N1  ( .A1(\SB3_16/i1_5 ), .A2(
        \SB3_16/i0[10] ), .A3(\SB3_16/i1[9] ), .ZN(
        \SB3_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_3/N4  ( .A1(\SB3_16/i1_5 ), .A2(
        \SB3_16/i0[8] ), .A3(\SB3_16/i3[0] ), .ZN(
        \SB3_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_16/Component_Function_3/N3  ( .A1(\SB3_16/i1[9] ), .A2(
        \SB3_16/i1_7 ), .A3(\SB3_16/i0[10] ), .ZN(
        \SB3_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_16/Component_Function_3/N2  ( .A1(\SB3_16/i0_0 ), .A2(
        \SB3_16/i0_3 ), .A3(\SB3_16/i0_4 ), .ZN(
        \SB3_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_3/N1  ( .A1(\SB3_16/i1[9] ), .A2(n876), 
        .A3(\SB3_16/i0[6] ), .ZN(\SB3_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N4  ( .A1(\SB3_16/i1[9] ), .A2(
        \SB3_16/i1_5 ), .A3(\SB3_16/i0_4 ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N2  ( .A1(\SB3_16/i3[0] ), .A2(
        \SB3_16/i0_0 ), .A3(\SB3_16/i1_7 ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N1  ( .A1(\SB3_16/i0[9] ), .A2(
        \SB3_16/i0_0 ), .A3(\SB3_16/i0[8] ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_2/N4  ( .A1(\SB3_17/i1_5 ), .A2(
        \SB3_17/i0_0 ), .A3(\SB3_17/i0_4 ), .ZN(
        \SB3_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_17/Component_Function_2/N3  ( .A1(\SB3_17/i0_3 ), .A2(
        \SB3_17/i0[8] ), .A3(\SB3_17/i0[9] ), .ZN(
        \SB3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_17/Component_Function_2/N2  ( .A1(\SB3_17/i0_3 ), .A2(
        \SB3_17/i0[10] ), .A3(\SB3_17/i0[6] ), .ZN(
        \SB3_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_17/Component_Function_2/N1  ( .A1(\SB3_17/i1_5 ), .A2(
        \SB3_17/i0[10] ), .A3(\SB3_17/i1[9] ), .ZN(
        \SB3_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_3/N4  ( .A1(\SB3_17/i1_5 ), .A2(
        \SB3_17/i0[8] ), .A3(\SB3_17/i3[0] ), .ZN(
        \SB3_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_17/Component_Function_3/N3  ( .A1(\SB3_17/i1[9] ), .A2(
        \SB3_17/i1_7 ), .A3(\SB3_17/i0[10] ), .ZN(
        \SB3_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_17/Component_Function_3/N2  ( .A1(\SB3_17/i0_0 ), .A2(
        \SB3_17/i0_3 ), .A3(\SB3_17/i0_4 ), .ZN(
        \SB3_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_17/Component_Function_3/N1  ( .A1(\SB3_17/i1[9] ), .A2(n867), 
        .A3(\SB3_17/i0[6] ), .ZN(\SB3_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N4  ( .A1(\SB3_17/i1[9] ), .A2(
        \SB3_17/i1_5 ), .A3(\SB3_17/i0_4 ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N3  ( .A1(\SB3_17/i0[9] ), .A2(
        \SB3_17/i0[10] ), .A3(\SB3_17/i0_3 ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N2  ( .A1(\SB3_17/i3[0] ), .A2(
        \SB3_17/i0_0 ), .A3(\SB3_17/i1_7 ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N1  ( .A1(\SB3_17/i0[9] ), .A2(
        \SB3_17/i0_0 ), .A3(\SB3_17/i0[8] ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_18/Component_Function_2/N4  ( .A1(\SB3_18/i1_5 ), .A2(
        \SB3_18/i0_0 ), .A3(\SB3_18/i0_4 ), .ZN(
        \SB3_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_18/Component_Function_2/N3  ( .A1(n869), .A2(\SB3_18/i0[8] ), 
        .A3(\SB3_18/i0[9] ), .ZN(\SB3_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_2/N2  ( .A1(n869), .A2(\SB3_18/i0[10] ), 
        .A3(\SB3_18/i0[6] ), .ZN(\SB3_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_18/Component_Function_2/N1  ( .A1(\SB3_18/i1_5 ), .A2(
        \SB3_18/i0[10] ), .A3(\SB3_18/i1[9] ), .ZN(
        \SB3_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_18/Component_Function_3/N4  ( .A1(\SB3_18/i1_5 ), .A2(
        \SB3_18/i0[8] ), .A3(\SB3_18/i3[0] ), .ZN(
        \SB3_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_18/Component_Function_3/N3  ( .A1(\SB3_18/i1[9] ), .A2(
        \SB3_18/i1_7 ), .A3(\SB3_18/i0[10] ), .ZN(
        \SB3_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_3/N2  ( .A1(\SB3_18/i0_0 ), .A2(
        \SB3_18/i0_3 ), .A3(\SB3_18/i0_4 ), .ZN(
        \SB3_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_18/Component_Function_3/N1  ( .A1(\SB3_18/i1[9] ), .A2(n869), 
        .A3(\SB3_18/i0[6] ), .ZN(\SB3_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N4  ( .A1(\SB3_18/i1[9] ), .A2(
        \SB3_18/i1_5 ), .A3(\SB3_18/i0_4 ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N3  ( .A1(\SB3_18/i0[9] ), .A2(
        \SB3_18/i0[10] ), .A3(\SB3_18/i0_3 ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N2  ( .A1(\SB3_18/i3[0] ), .A2(
        \SB3_18/i0_0 ), .A3(\SB3_18/i1_7 ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N1  ( .A1(\SB3_18/i0[9] ), .A2(
        \SB3_18/i0_0 ), .A3(\SB3_18/i0[8] ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_2/N4  ( .A1(\SB3_19/i1_5 ), .A2(
        \SB3_19/i0_0 ), .A3(\SB3_19/i0_4 ), .ZN(
        \SB3_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_19/Component_Function_2/N2  ( .A1(\SB3_19/i0_3 ), .A2(
        \SB3_19/i0[10] ), .A3(\SB3_19/i0[6] ), .ZN(
        \SB3_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_19/Component_Function_2/N1  ( .A1(\SB3_19/i1_5 ), .A2(
        \SB3_19/i0[10] ), .A3(\SB3_19/i1[9] ), .ZN(
        \SB3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_3/N4  ( .A1(\SB3_19/i1_5 ), .A2(
        \SB3_19/i0[8] ), .A3(\SB3_19/i3[0] ), .ZN(
        \SB3_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_19/Component_Function_3/N3  ( .A1(\SB3_19/i1[9] ), .A2(
        \SB3_19/i1_7 ), .A3(\SB3_19/i0[10] ), .ZN(
        \SB3_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_19/Component_Function_3/N1  ( .A1(\SB3_19/i1[9] ), .A2(
        \SB3_19/i0_3 ), .A3(\SB3_19/i0[6] ), .ZN(
        \SB3_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N4  ( .A1(\SB3_19/i1[9] ), .A2(
        \SB3_19/i1_5 ), .A3(\SB3_19/i0_4 ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N2  ( .A1(\SB3_19/i3[0] ), .A2(
        \SB3_19/i0_0 ), .A3(\SB3_19/i1_7 ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N1  ( .A1(\SB3_19/i0[9] ), .A2(
        \SB3_19/i0_0 ), .A3(\SB3_19/i0[8] ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_2/N4  ( .A1(\SB3_20/i1_5 ), .A2(
        \SB3_20/i0_0 ), .A3(\SB3_20/i0_4 ), .ZN(
        \SB3_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_20/Component_Function_2/N3  ( .A1(n864), .A2(\SB3_20/i0[8] ), 
        .A3(\SB3_20/i0[9] ), .ZN(\SB3_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_20/Component_Function_2/N2  ( .A1(\SB3_20/i0_3 ), .A2(
        \SB3_20/i0[10] ), .A3(\SB3_20/i0[6] ), .ZN(
        \SB3_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_20/Component_Function_2/N1  ( .A1(\SB3_20/i1_5 ), .A2(
        \SB3_20/i0[10] ), .A3(\SB3_20/i1[9] ), .ZN(
        \SB3_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_3/N3  ( .A1(\SB3_20/i1[9] ), .A2(
        \SB3_20/i1_7 ), .A3(\SB3_20/i0[10] ), .ZN(
        \SB3_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_20/Component_Function_3/N2  ( .A1(\SB3_20/i0_0 ), .A2(
        \SB3_20/i0_3 ), .A3(\SB3_20/i0_4 ), .ZN(
        \SB3_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_20/Component_Function_3/N1  ( .A1(\SB3_20/i1[9] ), .A2(n864), 
        .A3(\SB3_20/i0[6] ), .ZN(\SB3_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_4/N4  ( .A1(\SB3_20/i1[9] ), .A2(
        \SB3_20/i1_5 ), .A3(\SB3_20/i0_4 ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_20/Component_Function_4/N3  ( .A1(\SB3_20/i0[9] ), .A2(
        \SB3_20/i0[10] ), .A3(\SB3_20/i0_3 ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_20/Component_Function_4/N2  ( .A1(\SB3_20/i3[0] ), .A2(
        \SB3_20/i0_0 ), .A3(\SB3_20/i1_7 ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_20/Component_Function_4/N1  ( .A1(\SB3_20/i0[9] ), .A2(
        \SB3_20/i0_0 ), .A3(\SB3_20/i0[8] ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_2/N4  ( .A1(\SB3_21/i1_5 ), .A2(
        \SB3_21/i0_0 ), .A3(\SB3_21/i0_4 ), .ZN(
        \SB3_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_21/Component_Function_2/N3  ( .A1(n843), .A2(\SB3_21/i0[8] ), 
        .A3(\SB3_21/i0[9] ), .ZN(\SB3_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_21/Component_Function_2/N2  ( .A1(n843), .A2(\SB3_21/i0[10] ), 
        .A3(\SB3_21/i0[6] ), .ZN(\SB3_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_21/Component_Function_2/N1  ( .A1(\SB3_21/i1_5 ), .A2(
        \SB3_21/i0[10] ), .A3(\SB3_21/i1[9] ), .ZN(
        \SB3_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_3/N4  ( .A1(\SB3_21/i1_5 ), .A2(
        \SB3_21/i0[8] ), .A3(\SB3_21/i3[0] ), .ZN(
        \SB3_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_21/Component_Function_3/N3  ( .A1(\SB3_21/i1[9] ), .A2(
        \SB3_21/i1_7 ), .A3(\SB3_21/i0[10] ), .ZN(
        \SB3_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_21/Component_Function_3/N2  ( .A1(\SB3_21/i0_0 ), .A2(n843), 
        .A3(\SB3_21/i0_4 ), .ZN(\SB3_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_21/Component_Function_3/N1  ( .A1(\SB3_21/i1[9] ), .A2(n843), 
        .A3(\SB3_21/i0[6] ), .ZN(\SB3_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_4/N4  ( .A1(\SB3_21/i1[9] ), .A2(
        \SB3_21/i1_5 ), .A3(\SB3_21/i0_4 ), .ZN(
        \SB3_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_21/Component_Function_4/N2  ( .A1(\SB3_21/i3[0] ), .A2(
        \SB3_21/i0_0 ), .A3(\SB3_21/i1_7 ), .ZN(
        \SB3_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_21/Component_Function_4/N1  ( .A1(\SB3_21/i0[9] ), .A2(
        \SB3_21/i0_0 ), .A3(\SB3_21/i0[8] ), .ZN(
        \SB3_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_2/N3  ( .A1(\SB3_22/i0_3 ), .A2(
        \SB3_22/i0[8] ), .A3(\SB3_22/i0[9] ), .ZN(
        \SB3_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_22/Component_Function_2/N2  ( .A1(\SB3_22/i0_3 ), .A2(
        \SB3_22/i0[10] ), .A3(\SB3_22/i0[6] ), .ZN(
        \SB3_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_22/Component_Function_2/N1  ( .A1(\SB3_22/i1_5 ), .A2(
        \SB3_22/i0[10] ), .A3(\SB3_22/i1[9] ), .ZN(
        \SB3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_3/N4  ( .A1(\SB3_22/i1_5 ), .A2(
        \SB3_22/i0[8] ), .A3(\SB3_22/i3[0] ), .ZN(
        \SB3_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_22/Component_Function_3/N3  ( .A1(\SB3_22/i1[9] ), .A2(
        \SB3_22/i1_7 ), .A3(\SB3_22/i0[10] ), .ZN(
        \SB3_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_22/Component_Function_3/N2  ( .A1(\SB3_22/i0_0 ), .A2(
        \SB3_22/i0_3 ), .A3(\SB3_22/i0_4 ), .ZN(
        \SB3_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_22/Component_Function_3/N1  ( .A1(\SB3_22/i1[9] ), .A2(
        \SB3_22/i0_3 ), .A3(\SB3_22/i0[6] ), .ZN(
        \SB3_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N4  ( .A1(\SB3_22/i1[9] ), .A2(
        \SB3_22/i1_5 ), .A3(\SB3_22/i0_4 ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N2  ( .A1(\SB3_22/i3[0] ), .A2(
        \SB3_22/i0_0 ), .A3(\SB3_22/i1_7 ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N1  ( .A1(\SB3_22/i0[9] ), .A2(
        \SB3_22/i0_0 ), .A3(\SB3_22/i0[8] ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_2/N4  ( .A1(\SB3_23/i1_5 ), .A2(
        \SB3_23/i0_0 ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_2/N3  ( .A1(\SB3_23/i0_3 ), .A2(
        \SB3_23/i0[8] ), .A3(\SB3_23/i0[9] ), .ZN(
        \SB3_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_23/Component_Function_2/N2  ( .A1(n847), .A2(\SB3_23/i0[10] ), 
        .A3(\SB3_23/i0[6] ), .ZN(\SB3_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_23/Component_Function_2/N1  ( .A1(\SB3_23/i1_5 ), .A2(
        \SB3_23/i0[10] ), .A3(\SB3_23/i1[9] ), .ZN(
        \SB3_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_3/N3  ( .A1(\SB3_23/i1[9] ), .A2(
        \SB3_23/i1_7 ), .A3(\SB3_23/i0[10] ), .ZN(
        \SB3_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_23/Component_Function_3/N2  ( .A1(\SB3_23/i0_0 ), .A2(
        \SB3_23/i0_3 ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_23/Component_Function_3/N1  ( .A1(\SB3_23/i1[9] ), .A2(n847), 
        .A3(\SB3_23/i0[6] ), .ZN(\SB3_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_4/N4  ( .A1(\SB3_23/i1[9] ), .A2(
        \SB3_23/i1_5 ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_4/N2  ( .A1(\SB3_23/i3[0] ), .A2(
        \SB3_23/i0_0 ), .A3(\SB3_23/i1_7 ), .ZN(
        \SB3_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_23/Component_Function_4/N1  ( .A1(\SB3_23/i0[9] ), .A2(
        \SB3_23/i0_0 ), .A3(\SB3_23/i0[8] ), .ZN(
        \SB3_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_2/N4  ( .A1(\SB3_24/i1_5 ), .A2(
        \SB3_24/i0_0 ), .A3(\SB3_24/i0_4 ), .ZN(
        \SB3_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_24/Component_Function_2/N3  ( .A1(\SB3_24/i0_3 ), .A2(
        \SB3_24/i0[8] ), .A3(\SB3_24/i0[9] ), .ZN(
        \SB3_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_24/Component_Function_2/N2  ( .A1(n872), .A2(\SB3_24/i0[10] ), 
        .A3(\SB3_24/i0[6] ), .ZN(\SB3_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_24/Component_Function_2/N1  ( .A1(\SB3_24/i1_5 ), .A2(
        \SB3_24/i0[10] ), .A3(\SB3_24/i1[9] ), .ZN(
        \SB3_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_3/N3  ( .A1(\SB3_24/i1[9] ), .A2(
        \SB3_24/i1_7 ), .A3(\SB3_24/i0[10] ), .ZN(
        \SB3_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_24/Component_Function_3/N2  ( .A1(\SB3_24/i0_0 ), .A2(
        \SB3_24/i0_3 ), .A3(\SB3_24/i0_4 ), .ZN(
        \SB3_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_24/Component_Function_4/N4  ( .A1(\SB3_24/i1[9] ), .A2(
        \SB3_24/i1_5 ), .A3(\SB3_24/i0_4 ), .ZN(
        \SB3_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_24/Component_Function_4/N3  ( .A1(\SB3_24/i0[9] ), .A2(
        \SB3_24/i0[10] ), .A3(\SB3_24/i0_3 ), .ZN(
        \SB3_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_24/Component_Function_4/N2  ( .A1(\SB3_24/i3[0] ), .A2(
        \SB3_24/i0_0 ), .A3(\SB3_24/i1_7 ), .ZN(
        \SB3_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_24/Component_Function_4/N1  ( .A1(\SB3_24/i0[9] ), .A2(
        \SB3_24/i0_0 ), .A3(\SB3_24/i0[8] ), .ZN(
        \SB3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_2/N4  ( .A1(\SB3_25/i1_5 ), .A2(
        \SB3_25/i0_0 ), .A3(\SB3_25/i0_4 ), .ZN(
        \SB3_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_25/Component_Function_2/N3  ( .A1(n845), .A2(\SB3_25/i0[8] ), 
        .A3(\SB3_25/i0[9] ), .ZN(\SB3_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_25/Component_Function_2/N2  ( .A1(n845), .A2(\SB3_25/i0[10] ), 
        .A3(\SB3_25/i0[6] ), .ZN(\SB3_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_25/Component_Function_2/N1  ( .A1(\SB3_25/i1_5 ), .A2(
        \SB3_25/i0[10] ), .A3(\SB3_25/i1[9] ), .ZN(
        \SB3_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_3/N4  ( .A1(\SB3_25/i1_5 ), .A2(
        \SB3_25/i0[8] ), .A3(\SB3_25/i3[0] ), .ZN(
        \SB3_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_25/Component_Function_3/N3  ( .A1(\SB3_25/i1[9] ), .A2(
        \SB3_25/i1_7 ), .A3(\SB3_25/i0[10] ), .ZN(
        \SB3_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_25/Component_Function_3/N2  ( .A1(\SB3_25/i0_0 ), .A2(
        \SB3_25/i0_3 ), .A3(\SB3_25/i0_4 ), .ZN(
        \SB3_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_25/Component_Function_3/N1  ( .A1(\SB3_25/i1[9] ), .A2(n845), 
        .A3(\SB3_25/i0[6] ), .ZN(\SB3_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_4/N4  ( .A1(\SB3_25/i1[9] ), .A2(
        \SB3_25/i1_5 ), .A3(\SB3_25/i0_4 ), .ZN(
        \SB3_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_25/Component_Function_4/N2  ( .A1(\SB3_25/i3[0] ), .A2(
        \SB3_25/i0_0 ), .A3(\SB3_25/i1_7 ), .ZN(
        \SB3_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_25/Component_Function_4/N1  ( .A1(\SB3_25/i0[9] ), .A2(
        \SB3_25/i0_0 ), .A3(\SB3_25/i0[8] ), .ZN(
        \SB3_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_2/N3  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i0[8] ), .A3(\SB3_26/i0[9] ), .ZN(
        \SB3_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_26/Component_Function_2/N2  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i0[10] ), .A3(\SB3_26/i0[6] ), .ZN(
        \SB3_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_2/N1  ( .A1(\SB3_26/i1_5 ), .A2(
        \SB3_26/i0[10] ), .A3(\SB3_26/i1[9] ), .ZN(
        \SB3_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_3/N4  ( .A1(\SB3_26/i1_5 ), .A2(
        \SB3_26/i0[8] ), .A3(\SB3_26/i3[0] ), .ZN(
        \SB3_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_26/Component_Function_3/N2  ( .A1(\SB3_26/i0_0 ), .A2(
        \SB3_26/i0_3 ), .A3(\SB3_26/i0_4 ), .ZN(
        \SB3_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_3/N1  ( .A1(\SB3_26/i1[9] ), .A2(
        \SB3_26/i0_3 ), .A3(\SB3_26/i0[6] ), .ZN(
        \SB3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N4  ( .A1(\SB3_26/i1[9] ), .A2(
        \SB3_26/i1_5 ), .A3(\SB3_26/i0_4 ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N3  ( .A1(\SB3_26/i0[9] ), .A2(
        \SB3_26/i0[10] ), .A3(\SB3_26/i0_3 ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N2  ( .A1(\SB3_26/i3[0] ), .A2(
        \SB3_26/i0_0 ), .A3(\SB3_26/i1_7 ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N1  ( .A1(\SB3_26/i0[9] ), .A2(
        \SB3_26/i0_0 ), .A3(\SB3_26/i0[8] ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_2/N3  ( .A1(\SB3_27/i0_3 ), .A2(
        \SB3_27/i0[8] ), .A3(\SB3_27/i0[9] ), .ZN(
        \SB3_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_27/Component_Function_2/N2  ( .A1(\SB3_27/i0_3 ), .A2(
        \SB3_27/i0[10] ), .A3(\SB3_27/i0[6] ), .ZN(
        \SB3_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_27/Component_Function_2/N1  ( .A1(\SB3_27/i1_5 ), .A2(
        \SB3_27/i0[10] ), .A3(\SB3_27/i1[9] ), .ZN(
        \SB3_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_3/N4  ( .A1(\SB3_27/i1_5 ), .A2(
        \SB3_27/i3[0] ), .A3(\SB3_27/i0[8] ), .ZN(
        \SB3_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_27/Component_Function_3/N3  ( .A1(\SB3_27/i1[9] ), .A2(
        \SB3_27/i1_7 ), .A3(\SB3_27/i0[10] ), .ZN(
        \SB3_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_27/Component_Function_3/N2  ( .A1(\SB3_27/i0_0 ), .A2(
        \SB3_27/i0_3 ), .A3(\SB3_27/i0_4 ), .ZN(
        \SB3_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_27/Component_Function_3/N1  ( .A1(\SB3_27/i1[9] ), .A2(n819), 
        .A3(\SB3_27/i0[6] ), .ZN(\SB3_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_4/N4  ( .A1(\SB3_27/i1[9] ), .A2(
        \SB3_27/i1_5 ), .A3(\SB3_27/i0_4 ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_27/Component_Function_4/N2  ( .A1(\SB3_27/i3[0] ), .A2(
        \SB3_27/i0_0 ), .A3(\SB3_27/i1_7 ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_27/Component_Function_4/N1  ( .A1(\SB3_27/i0[9] ), .A2(
        \SB3_27/i0_0 ), .A3(\SB3_27/i0[8] ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_2/N4  ( .A1(\SB3_28/i1_5 ), .A2(
        \SB3_28/i0_0 ), .A3(\SB3_28/i0_4 ), .ZN(
        \SB3_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_28/Component_Function_2/N3  ( .A1(\SB3_28/i0_3 ), .A2(
        \SB3_28/i0[8] ), .A3(\SB3_28/i0[9] ), .ZN(
        \SB3_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_2/N2  ( .A1(n865), .A2(\SB3_28/i0[10] ), 
        .A3(\SB3_28/i0[6] ), .ZN(\SB3_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_28/Component_Function_2/N1  ( .A1(\SB3_28/i1_5 ), .A2(
        \SB3_28/i0[10] ), .A3(\SB3_28/i1[9] ), .ZN(
        \SB3_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_3/N4  ( .A1(\SB3_28/i1_5 ), .A2(
        \SB3_28/i0[8] ), .A3(\SB3_28/i3[0] ), .ZN(
        \SB3_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_28/Component_Function_3/N2  ( .A1(\SB3_28/i0_0 ), .A2(n865), 
        .A3(\SB3_28/i0_4 ), .ZN(\SB3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_28/Component_Function_3/N1  ( .A1(\SB3_28/i1[9] ), .A2(n865), 
        .A3(\SB3_28/i0[6] ), .ZN(\SB3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N4  ( .A1(\SB3_28/i1[9] ), .A2(
        \SB3_28/i1_5 ), .A3(\SB3_28/i0_4 ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N3  ( .A1(\SB3_28/i0[9] ), .A2(
        \SB3_28/i0[10] ), .A3(\SB3_28/i0_3 ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N2  ( .A1(\SB3_28/i3[0] ), .A2(
        \SB3_28/i0_0 ), .A3(\SB3_28/i1_7 ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N1  ( .A1(\SB3_28/i0[9] ), .A2(
        \SB3_28/i0_0 ), .A3(\SB3_28/i0[8] ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_2/N2  ( .A1(n861), .A2(\SB3_29/i0[10] ), 
        .A3(\SB3_29/i0[6] ), .ZN(\SB3_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_29/Component_Function_2/N1  ( .A1(\SB3_29/i1_5 ), .A2(
        \SB3_29/i0[10] ), .A3(\SB3_29/i1[9] ), .ZN(
        \SB3_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_3/N3  ( .A1(\SB3_29/i1[9] ), .A2(
        \SB3_29/i1_7 ), .A3(\SB3_29/i0[10] ), .ZN(
        \SB3_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_3/N2  ( .A1(\SB3_29/i0_0 ), .A2(n861), 
        .A3(\SB3_29/i0_4 ), .ZN(\SB3_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_29/Component_Function_3/N1  ( .A1(\SB3_29/i1[9] ), .A2(n861), 
        .A3(\SB3_29/i0[6] ), .ZN(\SB3_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_4/N4  ( .A1(\SB3_29/i1[9] ), .A2(
        \SB3_29/i1_5 ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_29/Component_Function_4/N3  ( .A1(\SB3_29/i0[9] ), .A2(
        \SB3_29/i0[10] ), .A3(\SB3_29/i0_3 ), .ZN(
        \SB3_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_4/N2  ( .A1(\SB3_29/i3[0] ), .A2(
        \SB3_29/i0_0 ), .A3(\SB3_29/i1_7 ), .ZN(
        \SB3_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_29/Component_Function_4/N1  ( .A1(\SB3_29/i0[9] ), .A2(
        \SB3_29/i0_0 ), .A3(\SB3_29/i0[8] ), .ZN(
        \SB3_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_2/N3  ( .A1(\SB3_30/i0_3 ), .A2(
        \SB3_30/i0[8] ), .A3(\SB3_30/i0[9] ), .ZN(
        \SB3_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_30/Component_Function_2/N2  ( .A1(\SB3_30/i0[10] ), .A2(
        \SB3_30/i0_3 ), .A3(\SB3_30/i0[6] ), .ZN(
        \SB3_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_30/Component_Function_2/N1  ( .A1(\SB3_30/i1_5 ), .A2(
        \SB3_30/i0[10] ), .A3(\SB3_30/i1[9] ), .ZN(
        \SB3_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_3/N4  ( .A1(\SB3_30/i1_5 ), .A2(
        \SB3_30/i0[8] ), .A3(\SB3_30/i3[0] ), .ZN(
        \SB3_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_30/Component_Function_3/N2  ( .A1(\SB3_30/i0_0 ), .A2(
        \SB3_30/i0_3 ), .A3(\SB3_30/i0_4 ), .ZN(
        \SB3_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_30/Component_Function_3/N1  ( .A1(\SB3_30/i1[9] ), .A2(
        \SB3_30/i0_3 ), .A3(\SB3_30/i0[6] ), .ZN(
        \SB3_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_4/N4  ( .A1(\SB3_30/i1[9] ), .A2(
        \SB3_30/i1_5 ), .A3(\SB3_30/i0_4 ), .ZN(
        \SB3_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_30/Component_Function_4/N2  ( .A1(\SB3_30/i3[0] ), .A2(
        \SB3_30/i0_0 ), .A3(\SB3_30/i1_7 ), .ZN(
        \SB3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_30/Component_Function_4/N1  ( .A1(\SB3_30/i0[9] ), .A2(
        \SB3_30/i0_0 ), .A3(\SB3_30/i0[8] ), .ZN(
        \SB3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_2/N3  ( .A1(n1669), .A2(\SB3_31/i0[8] ), 
        .A3(\SB3_31/i0[9] ), .ZN(\SB3_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_31/Component_Function_2/N2  ( .A1(\SB3_31/i0_3 ), .A2(
        \SB3_31/i0[10] ), .A3(\SB3_31/i0[6] ), .ZN(
        \SB3_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_31/Component_Function_2/N1  ( .A1(\SB3_31/i1_5 ), .A2(
        \SB3_31/i0[10] ), .A3(\SB3_31/i1[9] ), .ZN(
        \SB3_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_3/N4  ( .A1(\SB3_31/i1_5 ), .A2(
        \SB3_31/i0[8] ), .A3(\SB3_31/i3[0] ), .ZN(
        \SB3_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_31/Component_Function_3/N2  ( .A1(\SB3_31/i0_0 ), .A2(
        \SB3_31/i0_3 ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_31/Component_Function_3/N1  ( .A1(n1669), .A2(\SB3_31/i1[9] ), 
        .A3(\SB3_31/i0[6] ), .ZN(\SB3_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_4/N4  ( .A1(\SB3_31/i1[9] ), .A2(
        \SB3_31/i1_5 ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_31/Component_Function_4/N2  ( .A1(\SB3_31/i3[0] ), .A2(
        \SB3_31/i0_0 ), .A3(\SB3_31/i1_7 ), .ZN(
        \SB3_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_31/Component_Function_4/N1  ( .A1(\SB3_31/i0[9] ), .A2(
        \SB3_31/i0_0 ), .A3(\SB3_31/i0[8] ), .ZN(
        \SB3_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_0/Component_Function_2/N4  ( .A1(\SB4_0/i1_5 ), .A2(
        \SB4_0/i0_0 ), .A3(\SB4_0/i0_4 ), .ZN(
        \SB4_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_0/Component_Function_2/N3  ( .A1(n1672), .A2(\SB4_0/i0[8] ), 
        .A3(\SB4_0/i0[9] ), .ZN(\SB4_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_0/Component_Function_2/N2  ( .A1(\SB4_0/i0_3 ), .A2(
        \SB4_0/i0[10] ), .A3(\SB4_0/i0[6] ), .ZN(
        \SB4_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_0/Component_Function_4/N4  ( .A1(\SB4_0/i1[9] ), .A2(
        \SB4_0/i1_5 ), .A3(\SB4_0/i0_4 ), .ZN(
        \SB4_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_0/Component_Function_4/N1  ( .A1(\SB4_0/i0[9] ), .A2(
        \SB4_0/i0_0 ), .A3(\SB4_0/i0[8] ), .ZN(
        \SB4_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_1/Component_Function_2/N4  ( .A1(\SB4_1/i1_5 ), .A2(
        \SB4_1/i0_0 ), .A3(\SB4_1/i0_4 ), .ZN(
        \SB4_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_1/Component_Function_2/N3  ( .A1(n857), .A2(\SB4_1/i0[8] ), 
        .A3(\SB4_1/i0[9] ), .ZN(\SB4_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_1/Component_Function_2/N2  ( .A1(\SB4_1/i0_3 ), .A2(
        \SB4_1/i0[10] ), .A3(\SB4_1/i0[6] ), .ZN(
        \SB4_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_1/Component_Function_3/N4  ( .A1(\SB4_1/i1_5 ), .A2(
        \SB4_1/i0[8] ), .A3(\SB4_1/i3[0] ), .ZN(
        \SB4_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_1/Component_Function_4/N4  ( .A1(\SB4_1/i1[9] ), .A2(
        \SB4_1/i1_5 ), .A3(\SB4_1/i0_4 ), .ZN(
        \SB4_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_2/Component_Function_2/N3  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i0[8] ), .A3(n785), .ZN(
        \SB4_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_2/Component_Function_2/N2  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i0[10] ), .A3(\SB4_2/i0[6] ), .ZN(
        \SB4_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_2/Component_Function_2/N1  ( .A1(\SB4_2/i1_5 ), .A2(
        \SB4_2/i0[10] ), .A3(\SB4_2/i1[9] ), .ZN(
        \SB4_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_3/N4  ( .A1(\SB4_2/i1_5 ), .A2(
        \SB4_2/i0[8] ), .A3(n556), .ZN(
        \SB4_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_3/Component_Function_2/N3  ( .A1(\SB4_3/i0_3 ), .A2(
        \SB4_3/i0[8] ), .A3(\SB4_3/i0[9] ), .ZN(
        \SB4_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_3/Component_Function_2/N2  ( .A1(n859), .A2(\SB4_3/i0[10] ), 
        .A3(\SB4_3/i0[6] ), .ZN(\SB4_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_3/Component_Function_3/N4  ( .A1(\SB4_3/i1_5 ), .A2(
        \SB4_3/i0[8] ), .A3(\SB4_3/i3[0] ), .ZN(
        \SB4_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_3/Component_Function_3/N3  ( .A1(\SB4_3/i1[9] ), .A2(
        \SB4_3/i1_7 ), .A3(\SB4_3/i0[10] ), .ZN(
        \SB4_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_3/Component_Function_4/N3  ( .A1(\SB4_3/i0[9] ), .A2(
        \SB4_3/i0[10] ), .A3(\SB4_3/i0_3 ), .ZN(
        \SB4_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_3/Component_Function_4/N2  ( .A1(\SB4_3/i3[0] ), .A2(
        \SB4_3/i0_0 ), .A3(\SB4_3/i1_7 ), .ZN(
        \SB4_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_3/Component_Function_4/N1  ( .A1(\SB4_3/i0[9] ), .A2(
        \SB4_3/i0_0 ), .A3(\SB4_3/i0[8] ), .ZN(
        \SB4_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_4/Component_Function_2/N3  ( .A1(n1667), .A2(\SB4_4/i0[8] ), 
        .A3(\SB4_4/i0[9] ), .ZN(\SB4_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_4/Component_Function_2/N2  ( .A1(\SB4_4/i0_3 ), .A2(
        \SB4_4/i0[10] ), .A3(\SB4_4/i0[6] ), .ZN(
        \SB4_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_4/Component_Function_2/N1  ( .A1(\SB4_4/i1_5 ), .A2(
        \SB4_4/i0[10] ), .A3(\SB4_4/i1[9] ), .ZN(
        \SB4_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_4/Component_Function_3/N4  ( .A1(\SB4_4/i1_5 ), .A2(
        \SB4_4/i0[8] ), .A3(\SB4_4/i3[0] ), .ZN(
        \SB4_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_4/Component_Function_4/N4  ( .A1(\SB4_4/i1[9] ), .A2(
        \SB4_4/i1_5 ), .A3(\SB4_4/i0_4 ), .ZN(
        \SB4_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_4/Component_Function_4/N3  ( .A1(\SB4_4/i0[9] ), .A2(
        \SB4_4/i0[10] ), .A3(\SB4_4/i0_3 ), .ZN(
        \SB4_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_4/Component_Function_4/N1  ( .A1(\SB4_4/i0[9] ), .A2(
        \SB4_4/i0_0 ), .A3(\SB4_4/i0[8] ), .ZN(
        \SB4_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_2/N3  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i0[8] ), .A3(\SB4_5/i0[9] ), .ZN(
        \SB4_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_5/Component_Function_2/N2  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i0[10] ), .A3(n810), .ZN(
        \SB4_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_5/Component_Function_4/N1  ( .A1(\SB4_5/i0[9] ), .A2(
        \SB4_5/i0_0 ), .A3(\SB4_5/i0[8] ), .ZN(
        \SB4_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_6/Component_Function_2/N4  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0_0 ), .A3(\SB4_6/i0_4 ), .ZN(
        \SB4_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_2/N3  ( .A1(n858), .A2(\SB4_6/i0[8] ), 
        .A3(\SB4_6/i0[9] ), .ZN(\SB4_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_6/Component_Function_2/N2  ( .A1(\SB4_6/i0_3 ), .A2(
        \SB4_6/i0[10] ), .A3(\SB4_6/i0[6] ), .ZN(
        \SB4_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_6/Component_Function_3/N4  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0[8] ), .A3(\SB4_6/i3[0] ), .ZN(
        \SB4_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_3/N3  ( .A1(\SB4_6/i1[9] ), .A2(
        \SB4_6/i1_7 ), .A3(\SB4_6/i0[10] ), .ZN(
        \SB4_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_6/Component_Function_4/N3  ( .A1(\SB4_6/i0[9] ), .A2(
        \SB4_6/i0[10] ), .A3(\SB4_6/i0_3 ), .ZN(
        \SB4_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_7/Component_Function_2/N3  ( .A1(n877), .A2(\SB4_7/i0[8] ), 
        .A3(\SB4_7/i0[9] ), .ZN(\SB4_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_7/Component_Function_2/N2  ( .A1(\SB4_7/i0_3 ), .A2(
        \SB4_7/i0[10] ), .A3(\SB4_7/i0[6] ), .ZN(
        \SB4_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_7/Component_Function_3/N4  ( .A1(\SB4_7/i1_5 ), .A2(
        \SB4_7/i0[8] ), .A3(\SB4_7/i3[0] ), .ZN(
        \SB4_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_3/N3  ( .A1(\SB4_7/i1[9] ), .A2(
        \SB4_7/i1_7 ), .A3(\SB4_7/i0[10] ), .ZN(
        \SB4_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_7/Component_Function_4/N3  ( .A1(\SB4_7/i0[9] ), .A2(
        \SB4_7/i0[10] ), .A3(n877), .ZN(
        \SB4_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_7/Component_Function_4/N1  ( .A1(\SB4_7/i0[9] ), .A2(
        \SB4_7/i0_0 ), .A3(\SB4_7/i0[8] ), .ZN(
        \SB4_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_2/N3  ( .A1(\SB4_8/i0_3 ), .A2(
        \SB4_8/i0[8] ), .A3(\SB4_8/i0[9] ), .ZN(
        \SB4_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_8/Component_Function_2/N2  ( .A1(n863), .A2(\SB4_8/i0[10] ), 
        .A3(\SB4_8/i0[6] ), .ZN(\SB4_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_8/Component_Function_2/N1  ( .A1(\SB4_8/i1_5 ), .A2(
        \SB4_8/i0[10] ), .A3(\SB4_8/i1[9] ), .ZN(
        \SB4_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_3/N4  ( .A1(\SB4_8/i1_5 ), .A2(
        \SB4_8/i0[8] ), .A3(\SB4_8/i3[0] ), .ZN(
        \SB4_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_8/Component_Function_4/N4  ( .A1(\SB4_8/i1[9] ), .A2(
        \SB4_8/i1_5 ), .A3(n1638), .ZN(
        \SB4_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_8/Component_Function_4/N3  ( .A1(\SB4_8/i0[9] ), .A2(
        \SB4_8/i0[10] ), .A3(\SB4_8/i0_3 ), .ZN(
        \SB4_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_8/Component_Function_4/N1  ( .A1(\SB4_8/i0[9] ), .A2(
        \SB4_8/i0_0 ), .A3(\SB4_8/i0[8] ), .ZN(
        \SB4_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_9/Component_Function_2/N3  ( .A1(n1663), .A2(\SB4_9/i0[8] ), 
        .A3(\SB4_9/i0[9] ), .ZN(\SB4_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_9/Component_Function_2/N2  ( .A1(\SB4_9/i0_3 ), .A2(
        \SB4_9/i0[10] ), .A3(\SB4_9/i0[6] ), .ZN(
        \SB4_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_9/Component_Function_2/N1  ( .A1(\SB4_9/i1_5 ), .A2(
        \SB4_9/i0[10] ), .A3(\SB4_9/i1[9] ), .ZN(
        \SB4_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_9/Component_Function_3/N4  ( .A1(\SB4_9/i1_5 ), .A2(
        \SB4_9/i0[8] ), .A3(\SB4_9/i3[0] ), .ZN(
        \SB4_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_3/N3  ( .A1(\SB4_9/i1[9] ), .A2(
        \SB4_9/i1_7 ), .A3(\SB4_9/i0[10] ), .ZN(
        \SB4_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_9/Component_Function_4/N4  ( .A1(\SB4_9/i1[9] ), .A2(
        \SB4_9/i1_5 ), .A3(\RI3[4][136] ), .ZN(
        \SB4_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_4/N1  ( .A1(\SB4_9/i0[9] ), .A2(
        \SB4_9/i0_0 ), .A3(\SB4_9/i0[8] ), .ZN(
        \SB4_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_10/Component_Function_2/N3  ( .A1(\SB4_10/i0_3 ), .A2(
        \SB4_10/i0[8] ), .A3(\SB4_10/i0[9] ), .ZN(
        \SB4_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_10/Component_Function_2/N2  ( .A1(\SB4_10/i0_3 ), .A2(
        \SB4_10/i0[10] ), .A3(\SB4_10/i0[6] ), .ZN(
        \SB4_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_10/Component_Function_3/N4  ( .A1(\SB4_10/i1_5 ), .A2(
        \SB4_10/i0[8] ), .A3(\SB4_10/i3[0] ), .ZN(
        \SB4_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_10/Component_Function_4/N1  ( .A1(\SB4_10/i0[9] ), .A2(
        \SB4_10/i0_0 ), .A3(\SB4_10/i0[8] ), .ZN(
        \SB4_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_11/Component_Function_2/N3  ( .A1(n841), .A2(\SB4_11/i0[8] ), 
        .A3(\SB4_11/i0[9] ), .ZN(\SB4_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_11/Component_Function_2/N2  ( .A1(\SB4_11/i0_3 ), .A2(
        \SB4_11/i0[10] ), .A3(\SB4_11/i0[6] ), .ZN(
        \SB4_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_11/Component_Function_2/N1  ( .A1(\SB4_11/i1_5 ), .A2(
        \SB4_11/i0[10] ), .A3(\SB4_11/i1[9] ), .ZN(
        \SB4_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_11/Component_Function_3/N4  ( .A1(\SB4_11/i1_5 ), .A2(
        \SB4_11/i0[8] ), .A3(\SB4_11/i3[0] ), .ZN(
        \SB4_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_11/Component_Function_4/N3  ( .A1(\SB4_11/i0[9] ), .A2(
        \SB4_11/i0[10] ), .A3(n841), .ZN(
        \SB4_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_11/Component_Function_4/N1  ( .A1(\SB4_11/i0[9] ), .A2(
        \SB4_11/i0_0 ), .A3(\SB4_11/i0[8] ), .ZN(
        \SB4_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_12/Component_Function_2/N3  ( .A1(\SB4_12/i0_3 ), .A2(
        \SB4_12/i0[8] ), .A3(\SB4_12/i0[9] ), .ZN(
        \SB4_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_12/Component_Function_2/N2  ( .A1(n828), .A2(\SB4_12/i0[10] ), 
        .A3(\SB4_12/i0[6] ), .ZN(\SB4_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_12/Component_Function_2/N1  ( .A1(\SB4_12/i1_5 ), .A2(
        \SB4_12/i0[10] ), .A3(\SB4_12/i1[9] ), .ZN(
        \SB4_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_12/Component_Function_3/N4  ( .A1(\SB4_12/i1_5 ), .A2(
        \SB4_12/i0[8] ), .A3(\SB4_12/i3[0] ), .ZN(
        \SB4_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_12/Component_Function_3/N3  ( .A1(\SB4_12/i1[9] ), .A2(
        \SB4_12/i1_7 ), .A3(\SB4_12/i0[10] ), .ZN(
        \SB4_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_12/Component_Function_4/N3  ( .A1(\SB4_12/i0[9] ), .A2(
        \SB4_12/i0[10] ), .A3(n828), .ZN(
        \SB4_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_13/Component_Function_2/N4  ( .A1(\SB4_13/i1_5 ), .A2(
        \SB4_13/i0_0 ), .A3(\SB4_13/i0_4 ), .ZN(
        \SB4_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_13/Component_Function_2/N3  ( .A1(\SB4_13/i0_3 ), .A2(
        \SB4_13/i0[8] ), .A3(\SB4_13/i0[9] ), .ZN(
        \SB4_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_13/Component_Function_2/N2  ( .A1(n2148), .A2(\SB4_13/i0[10] ), 
        .A3(\SB4_13/i0[6] ), .ZN(\SB4_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_13/Component_Function_3/N4  ( .A1(\SB4_13/i1_5 ), .A2(
        \SB4_13/i0[8] ), .A3(\SB4_13/i3[0] ), .ZN(
        \SB4_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_13/Component_Function_3/N2  ( .A1(\SB4_13/i0_0 ), .A2(n2148), 
        .A3(\SB4_13/i0_4 ), .ZN(\SB4_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_13/Component_Function_4/N3  ( .A1(\SB4_13/i0[9] ), .A2(
        \SB4_13/i0[10] ), .A3(\SB4_13/i0_3 ), .ZN(
        \SB4_13/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_13/Component_Function_4/N1  ( .A1(\SB4_13/i0[9] ), .A2(
        \SB4_13/i0_0 ), .A3(\SB4_13/i0[8] ), .ZN(
        \SB4_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_2/N3  ( .A1(\SB4_14/i0[9] ), .A2(
        \SB4_14/i0[8] ), .A3(\SB4_14/i0_3 ), .ZN(
        \SB4_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_14/Component_Function_2/N2  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i0[10] ), .A3(n806), .ZN(
        \SB4_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_14/Component_Function_2/N1  ( .A1(\SB4_14/i1_5 ), .A2(
        \SB4_14/i0[10] ), .A3(\SB4_14/i1[9] ), .ZN(
        \SB4_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_3/N4  ( .A1(\SB4_14/i1_5 ), .A2(
        \SB4_14/i0[8] ), .A3(\SB4_14/i3[0] ), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_14/Component_Function_3/N3  ( .A1(\SB4_14/i1[9] ), .A2(
        \SB4_14/i1_7 ), .A3(\SB4_14/i0[10] ), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_14/Component_Function_4/N1  ( .A1(\SB4_14/i0[9] ), .A2(
        \SB4_14/i0_0 ), .A3(\SB4_14/i0[8] ), .ZN(
        \SB4_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_15/Component_Function_2/N3  ( .A1(\SB4_15/i0_3 ), .A2(
        \SB4_15/i0[8] ), .A3(\SB4_15/i0[9] ), .ZN(
        \SB4_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_15/Component_Function_2/N2  ( .A1(n871), .A2(\SB4_15/i0[10] ), 
        .A3(\SB4_15/i0[6] ), .ZN(\SB4_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_15/Component_Function_2/N1  ( .A1(\SB4_15/i1_5 ), .A2(
        \SB4_15/i0[10] ), .A3(\SB4_15/i1[9] ), .ZN(
        \SB4_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_15/Component_Function_3/N4  ( .A1(\SB4_15/i1_5 ), .A2(
        \SB4_15/i0[8] ), .A3(\SB4_15/i3[0] ), .ZN(
        \SB4_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_15/Component_Function_4/N3  ( .A1(\SB4_15/i0[9] ), .A2(
        \SB4_15/i0[10] ), .A3(\SB4_15/i0_3 ), .ZN(
        \SB4_15/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_15/Component_Function_4/N2  ( .A1(\SB4_15/i3[0] ), .A2(
        \SB4_15/i0_0 ), .A3(\SB4_15/i1_7 ), .ZN(
        \SB4_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_15/Component_Function_4/N1  ( .A1(\SB4_15/i0[9] ), .A2(
        \SB4_15/i0_0 ), .A3(\SB4_15/i0[8] ), .ZN(
        \SB4_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_16/Component_Function_2/N3  ( .A1(\SB4_16/i0_3 ), .A2(
        \SB4_16/i0[8] ), .A3(\SB4_16/i0[9] ), .ZN(
        \SB4_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_16/Component_Function_2/N2  ( .A1(\SB4_16/i0_3 ), .A2(
        \SB4_16/i0[10] ), .A3(\SB4_16/i0[6] ), .ZN(
        \SB4_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_16/Component_Function_3/N4  ( .A1(\SB4_16/i1_5 ), .A2(
        \SB4_16/i0[8] ), .A3(\SB4_16/i3[0] ), .ZN(
        \SB4_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_16/Component_Function_3/N3  ( .A1(\SB4_16/i1[9] ), .A2(
        \SB4_16/i1_7 ), .A3(\SB4_16/i0[10] ), .ZN(
        \SB4_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_16/Component_Function_4/N4  ( .A1(\SB4_16/i1[9] ), .A2(
        \SB4_16/i1_5 ), .A3(\SB4_16/i0_4 ), .ZN(
        \SB4_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_16/Component_Function_4/N3  ( .A1(\SB4_16/i0_3 ), .A2(
        \SB4_16/i0[10] ), .A3(\SB4_16/i0[9] ), .ZN(
        \SB4_16/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_17/Component_Function_2/N3  ( .A1(n868), .A2(\SB4_17/i0[8] ), 
        .A3(\SB4_17/i0[9] ), .ZN(\SB4_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_17/Component_Function_2/N2  ( .A1(\SB4_17/i0_3 ), .A2(
        \SB4_17/i0[10] ), .A3(\SB4_17/i0[6] ), .ZN(
        \SB4_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_17/Component_Function_3/N4  ( .A1(\SB4_17/i1_5 ), .A2(
        \SB4_17/i0[8] ), .A3(\SB4_17/i3[0] ), .ZN(
        \SB4_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_3/N1  ( .A1(\SB4_17/i1[9] ), .A2(n868), 
        .A3(\SB4_17/i0[6] ), .ZN(\SB4_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_17/Component_Function_4/N4  ( .A1(\SB4_17/i1[9] ), .A2(
        \SB4_17/i1_5 ), .A3(\SB4_17/i0_4 ), .ZN(
        \SB4_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_4/N3  ( .A1(\SB4_17/i0[9] ), .A2(
        \SB4_17/i0[10] ), .A3(n868), .ZN(
        \SB4_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_2/N3  ( .A1(n870), .A2(\SB4_18/i0[8] ), 
        .A3(\SB4_18/i0[9] ), .ZN(\SB4_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_2/N2  ( .A1(\SB4_18/i0_3 ), .A2(
        \SB4_18/i0[10] ), .A3(\SB4_18/i0[6] ), .ZN(
        \SB4_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_18/Component_Function_2/N1  ( .A1(\SB4_18/i1_5 ), .A2(
        \SB4_18/i0[10] ), .A3(n2113), .ZN(
        \SB4_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_3/N4  ( .A1(\SB4_18/i1_5 ), .A2(
        \SB4_18/i0[8] ), .A3(\SB4_18/i3[0] ), .ZN(
        \SB4_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_18/Component_Function_3/N3  ( .A1(n2113), .A2(\SB4_18/i1_7 ), 
        .A3(\SB4_18/i0[10] ), .ZN(\SB4_18/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 \SB4_18/Component_Function_3/N1  ( .A1(n2113), .A2(n870), .A3(
        \SB4_18/i0[6] ), .ZN(\SB4_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_4/N3  ( .A1(\SB4_18/i0[9] ), .A2(
        \SB4_18/i0[10] ), .A3(n870), .ZN(
        \SB4_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_4/N2  ( .A1(\SB4_18/i3[0] ), .A2(
        \SB4_18/i0_0 ), .A3(\SB4_18/i1_7 ), .ZN(
        \SB4_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_18/Component_Function_4/N1  ( .A1(\SB4_18/i0[9] ), .A2(
        \SB4_18/i0_0 ), .A3(\SB4_18/i0[8] ), .ZN(
        \SB4_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_2/N3  ( .A1(\SB4_19/i0_3 ), .A2(
        \SB4_19/i0[8] ), .A3(\SB4_19/i0[9] ), .ZN(
        \SB4_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_2/N2  ( .A1(\SB4_19/i0_3 ), .A2(
        \SB4_19/i0[10] ), .A3(\SB4_19/i0[6] ), .ZN(
        \SB4_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_19/Component_Function_2/N1  ( .A1(\SB4_19/i1_5 ), .A2(
        \SB4_19/i0[10] ), .A3(\SB4_19/i1[9] ), .ZN(
        \SB4_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_3/N4  ( .A1(\SB4_19/i1_5 ), .A2(
        \SB4_19/i0[8] ), .A3(\SB4_19/i3[0] ), .ZN(
        \SB4_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_3/N3  ( .A1(\SB4_19/i1[9] ), .A2(
        \SB4_19/i1_7 ), .A3(\SB4_19/i0[10] ), .ZN(
        \SB4_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_3/N1  ( .A1(\SB4_19/i1[9] ), .A2(
        \SB4_19/i0_3 ), .A3(\SB4_19/i0[6] ), .ZN(
        \SB4_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_4/N3  ( .A1(\SB4_19/i0[9] ), .A2(
        \SB4_19/i0[10] ), .A3(\SB4_19/i0_3 ), .ZN(
        \SB4_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_20/Component_Function_2/N4  ( .A1(\SB4_20/i1_5 ), .A2(
        \SB4_20/i0_0 ), .A3(n844), .ZN(
        \SB4_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_2/N3  ( .A1(\SB4_20/i0_3 ), .A2(
        \SB4_20/i0[8] ), .A3(\SB4_20/i0[9] ), .ZN(
        \SB4_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_20/Component_Function_2/N2  ( .A1(\SB4_20/i0_3 ), .A2(
        \SB4_20/i0[10] ), .A3(\SB4_20/i0[6] ), .ZN(
        \SB4_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_20/Component_Function_3/N4  ( .A1(\SB4_20/i1_5 ), .A2(
        \SB4_20/i0[8] ), .A3(\SB4_20/i3[0] ), .ZN(
        \SB4_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_4/N4  ( .A1(\SB4_20/i1[9] ), .A2(
        \SB4_20/i1_5 ), .A3(n844), .ZN(
        \SB4_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_4/N3  ( .A1(\SB4_20/i0[9] ), .A2(
        \SB4_20/i0[10] ), .A3(\SB4_20/i0_3 ), .ZN(
        \SB4_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_20/Component_Function_4/N2  ( .A1(\SB4_20/i3[0] ), .A2(
        \SB4_20/i0_0 ), .A3(\SB4_20/i1_7 ), .ZN(
        \SB4_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_20/Component_Function_4/N1  ( .A1(\SB4_20/i0[9] ), .A2(
        \SB4_20/i0_0 ), .A3(\SB4_20/i0[8] ), .ZN(
        \SB4_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_2/N3  ( .A1(n854), .A2(\SB4_21/i0[8] ), 
        .A3(\SB4_21/i0[9] ), .ZN(\SB4_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_21/Component_Function_2/N2  ( .A1(\SB4_21/i0_3 ), .A2(
        \SB4_21/i0[10] ), .A3(\SB4_21/i0[6] ), .ZN(
        \SB4_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_21/Component_Function_2/N1  ( .A1(\SB4_21/i1_5 ), .A2(
        \SB4_21/i0[10] ), .A3(\SB4_21/i1[9] ), .ZN(
        \SB4_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_3/N4  ( .A1(\SB4_21/i1_5 ), .A2(
        \SB4_21/i0[8] ), .A3(\SB4_21/i3[0] ), .ZN(
        \SB4_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_21/Component_Function_4/N3  ( .A1(\SB4_21/i0[9] ), .A2(
        \SB4_21/i0[10] ), .A3(\SB4_21/i0_3 ), .ZN(
        \SB4_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_21/Component_Function_4/N1  ( .A1(\SB4_21/i0[9] ), .A2(
        \SB4_21/i0_0 ), .A3(\SB4_21/i0[8] ), .ZN(
        \SB4_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_22/Component_Function_2/N2  ( .A1(\SB4_22/i0_3 ), .A2(
        \SB4_22/i0[10] ), .A3(\SB4_22/i0[6] ), .ZN(
        \SB4_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_22/Component_Function_3/N4  ( .A1(\SB4_22/i1_5 ), .A2(
        \SB4_22/i0[8] ), .A3(n550), .ZN(
        \SB4_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_22/Component_Function_3/N3  ( .A1(\SB4_22/i1[9] ), .A2(
        \SB4_22/i1_7 ), .A3(\SB4_22/i0[10] ), .ZN(
        \SB4_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_23/Component_Function_2/N3  ( .A1(n848), .A2(\SB4_23/i0[8] ), 
        .A3(\SB4_23/i0[9] ), .ZN(\SB4_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_23/Component_Function_2/N2  ( .A1(n2100), .A2(\SB4_23/i0[10] ), 
        .A3(\SB4_23/i0[6] ), .ZN(\SB4_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_23/Component_Function_2/N1  ( .A1(\SB4_23/i1_5 ), .A2(
        \SB4_23/i0[10] ), .A3(\SB4_23/i1[9] ), .ZN(
        \SB4_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_23/Component_Function_3/N4  ( .A1(\SB4_23/i1_5 ), .A2(
        \SB4_23/i0[8] ), .A3(\SB4_23/i3[0] ), .ZN(
        \SB4_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_3/N3  ( .A1(\SB4_23/i1[9] ), .A2(
        \SB4_23/i1_7 ), .A3(\SB4_23/i0[10] ), .ZN(
        \SB4_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_23/Component_Function_4/N4  ( .A1(\SB4_23/i1[9] ), .A2(
        \SB4_23/i1_5 ), .A3(\SB4_23/i0_4 ), .ZN(
        \SB4_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_4/N3  ( .A1(\SB4_23/i0[9] ), .A2(
        \SB4_23/i0[10] ), .A3(n2100), .ZN(
        \SB4_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_23/Component_Function_4/N1  ( .A1(\SB4_23/i0[9] ), .A2(
        \SB4_23/i0_0 ), .A3(\SB4_23/i0[8] ), .ZN(
        \SB4_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_2/N4  ( .A1(\SB4_24/i1_5 ), .A2(
        \SB4_24/i0_0 ), .A3(\SB4_24/i0_4 ), .ZN(
        \SB4_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_2/N3  ( .A1(\SB4_24/i0_3 ), .A2(
        \SB4_24/i0[8] ), .A3(\SB4_24/i0[9] ), .ZN(
        \SB4_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_24/Component_Function_2/N2  ( .A1(n2135), .A2(\SB4_24/i0[10] ), 
        .A3(\SB4_24/i0[6] ), .ZN(\SB4_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_24/Component_Function_3/N4  ( .A1(\SB4_24/i1_5 ), .A2(
        \SB4_24/i0[8] ), .A3(\SB4_24/i3[0] ), .ZN(
        \SB4_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_4/N4  ( .A1(\SB4_24/i1[9] ), .A2(
        \SB4_24/i1_5 ), .A3(\SB4_24/i0_4 ), .ZN(
        \SB4_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_4/N1  ( .A1(\SB4_24/i0[9] ), .A2(
        \SB4_24/i0_0 ), .A3(\SB4_24/i0[8] ), .ZN(
        \SB4_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_2/N4  ( .A1(\SB4_25/i0_4 ), .A2(
        \SB4_25/i0_0 ), .A3(\SB4_25/i1_5 ), .ZN(
        \SB4_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_2/N3  ( .A1(\SB4_25/i0[9] ), .A2(
        \SB4_25/i0[8] ), .A3(\SB4_25/i0_3 ), .ZN(
        \SB4_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_25/Component_Function_2/N2  ( .A1(\SB4_25/i0_3 ), .A2(
        \SB4_25/i0[10] ), .A3(\SB4_25/i0[6] ), .ZN(
        \SB4_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_2/N1  ( .A1(\SB4_25/i1_5 ), .A2(
        \SB4_25/i0[10] ), .A3(\SB4_25/i1[9] ), .ZN(
        \SB4_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_3/N4  ( .A1(\SB4_25/i1_5 ), .A2(
        \SB4_25/i0[8] ), .A3(\SB4_25/i3[0] ), .ZN(
        \SB4_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_4/N2  ( .A1(\SB4_25/i3[0] ), .A2(
        \SB4_25/i0_0 ), .A3(\SB4_25/i1_7 ), .ZN(
        \SB4_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_4/N1  ( .A1(\SB4_25/i0[9] ), .A2(
        \SB4_25/i0_0 ), .A3(\SB4_25/i0[8] ), .ZN(
        \SB4_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_2/N3  ( .A1(\SB4_26/i0_3 ), .A2(
        \SB4_26/i0[8] ), .A3(\SB4_26/i0[9] ), .ZN(
        \SB4_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_26/Component_Function_2/N2  ( .A1(n1671), .A2(\SB4_26/i0[10] ), 
        .A3(\SB4_26/i0[6] ), .ZN(\SB4_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_26/Component_Function_3/N4  ( .A1(\SB4_26/i1_5 ), .A2(
        \SB4_26/i0[8] ), .A3(\SB4_26/i3[0] ), .ZN(
        \SB4_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_26/Component_Function_4/N4  ( .A1(\SB4_26/i1[9] ), .A2(
        \SB4_26/i1_5 ), .A3(\SB4_26/i0_4 ), .ZN(
        \SB4_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_26/Component_Function_4/N3  ( .A1(\SB4_26/i0[9] ), .A2(
        \SB4_26/i0[10] ), .A3(\SB4_26/i0_3 ), .ZN(
        \SB4_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_27/Component_Function_2/N3  ( .A1(n1949), .A2(\SB4_27/i0[8] ), 
        .A3(\SB4_27/i0[9] ), .ZN(\SB4_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_27/Component_Function_2/N2  ( .A1(n1949), .A2(\SB4_27/i0[10] ), 
        .A3(\SB4_27/i0[6] ), .ZN(\SB4_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_27/Component_Function_3/N1  ( .A1(\SB4_27/i1[9] ), .A2(n1949), 
        .A3(\SB4_27/i0[6] ), .ZN(\SB4_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_4/N3  ( .A1(\SB4_27/i0[9] ), .A2(
        \SB4_27/i0[10] ), .A3(n1949), .ZN(
        \SB4_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_27/Component_Function_4/N1  ( .A1(\SB4_27/i0[9] ), .A2(
        \SB4_27/i0_0 ), .A3(\SB4_27/i0[8] ), .ZN(
        \SB4_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_28/Component_Function_2/N3  ( .A1(n866), .A2(\SB4_28/i0[8] ), 
        .A3(\SB4_28/i0[9] ), .ZN(\SB4_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_28/Component_Function_2/N2  ( .A1(\SB4_28/i0_3 ), .A2(
        \SB4_28/i0[10] ), .A3(\SB4_28/i0[6] ), .ZN(
        \SB4_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_28/Component_Function_3/N4  ( .A1(\SB4_28/i1_5 ), .A2(
        \SB4_28/i0[8] ), .A3(\SB4_28/i3[0] ), .ZN(
        \SB4_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_28/Component_Function_3/N2  ( .A1(\SB4_28/i0_0 ), .A2(n866), 
        .A3(\SB4_28/i0_4 ), .ZN(\SB4_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_28/Component_Function_4/N3  ( .A1(\SB4_28/i0[9] ), .A2(
        \SB4_28/i0[10] ), .A3(\SB4_28/i0_3 ), .ZN(
        \SB4_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_28/Component_Function_4/N1  ( .A1(\SB4_28/i0[9] ), .A2(
        \SB4_28/i0_0 ), .A3(\SB4_28/i0[8] ), .ZN(
        \SB4_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_29/Component_Function_2/N3  ( .A1(\SB4_29/i0_3 ), .A2(
        \SB4_29/i0[8] ), .A3(n790), .ZN(
        \SB4_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_29/Component_Function_2/N2  ( .A1(\SB4_29/i0_3 ), .A2(
        \SB4_29/i0[10] ), .A3(n791), .ZN(
        \SB4_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_29/Component_Function_3/N4  ( .A1(\SB4_29/i1_5 ), .A2(
        \SB4_29/i0[8] ), .A3(n555), .ZN(
        \SB4_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_29/Component_Function_4/N2  ( .A1(n555), .A2(\SB4_29/i0_0 ), 
        .A3(n554), .ZN(\SB4_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_30/Component_Function_2/N3  ( .A1(n1668), .A2(\SB4_30/i0[8] ), 
        .A3(\SB4_30/i0[9] ), .ZN(\SB4_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_30/Component_Function_2/N2  ( .A1(\SB4_30/i0_3 ), .A2(
        \SB4_30/i0[10] ), .A3(\SB4_30/i0[6] ), .ZN(
        \SB4_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_30/Component_Function_3/N4  ( .A1(\SB4_30/i1_5 ), .A2(
        \SB4_30/i0[8] ), .A3(\SB4_30/i3[0] ), .ZN(
        \SB4_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_30/Component_Function_4/N3  ( .A1(\SB4_30/i0[9] ), .A2(
        \SB4_30/i0[10] ), .A3(\SB4_30/i0_3 ), .ZN(
        \SB4_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_30/Component_Function_4/N2  ( .A1(\SB4_30/i3[0] ), .A2(
        \SB4_30/i0_0 ), .A3(\SB4_30/i1_7 ), .ZN(
        \SB4_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_30/Component_Function_4/N1  ( .A1(\SB4_30/i0[9] ), .A2(
        \SB4_30/i0_0 ), .A3(\SB4_30/i0[8] ), .ZN(
        \SB4_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_31/Component_Function_2/N3  ( .A1(n2106), .A2(\SB4_31/i0[8] ), 
        .A3(\SB4_31/i0[9] ), .ZN(\SB4_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_31/Component_Function_2/N2  ( .A1(n1670), .A2(\SB4_31/i0[10] ), 
        .A3(\SB4_31/i0[6] ), .ZN(\SB4_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_31/Component_Function_3/N4  ( .A1(n1964), .A2(\SB4_31/i0[8] ), 
        .A3(\SB4_31/i3[0] ), .ZN(\SB4_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_31/Component_Function_3/N3  ( .A1(\SB4_31/i1[9] ), .A2(
        \SB4_31/i1_7 ), .A3(\SB4_31/i0[10] ), .ZN(
        \SB4_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB4_31/Component_Function_4/N3  ( .A1(\SB4_31/i0[9] ), .A2(
        \SB4_31/i0[10] ), .A3(n1670), .ZN(
        \SB4_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_31/Component_Function_4/N1  ( .A1(\SB4_31/i0[9] ), .A2(
        \SB4_31/i0_0 ), .A3(\SB4_31/i0[8] ), .ZN(
        \SB4_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_0/Component_Function_0/N2  ( .A1(\SB1_0_0/i0[8] ), .A2(
        \SB1_0_0/i0[7] ), .A3(\SB1_0_0/i0[6] ), .ZN(
        \SB1_0_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_0/Component_Function_0/N1  ( .A1(\SB1_0_0/i0[10] ), .A2(
        \SB1_0_0/i0[9] ), .ZN(\SB1_0_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_0/Component_Function_1/N4  ( .A1(\SB1_0_0/i1_7 ), .A2(
        \SB1_0_0/i0[8] ), .A3(\SB1_0_0/i0_4 ), .ZN(
        \SB1_0_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_1/N3  ( .A1(n380), .A2(\SB1_0_0/i0[6] ), 
        .A3(\SB1_0_0/i0[9] ), .ZN(\SB1_0_0/Component_Function_1/NAND4_in[2] )
         );
  NAND3_X1 \SB1_0_0/Component_Function_1/N2  ( .A1(\SB1_0_0/i0_3 ), .A2(
        \SB1_0_0/i1_7 ), .A3(\SB1_0_0/i0[8] ), .ZN(
        \SB1_0_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_0/Component_Function_1/N1  ( .A1(\SB1_0_0/i0_3 ), .A2(
        \SB1_0_0/i1[9] ), .ZN(\SB1_0_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_0/Component_Function_5/N4  ( .A1(\SB1_0_0/i0[9] ), .A2(
        \SB1_0_0/i0[6] ), .A3(\SB1_0_0/i0_4 ), .ZN(
        \SB1_0_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_5/N2  ( .A1(\SB1_0_0/i0_0 ), .A2(
        \SB1_0_0/i0[6] ), .A3(\SB1_0_0/i0[10] ), .ZN(
        \SB1_0_0/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_0/Component_Function_5/N1  ( .A1(\SB1_0_0/i0_0 ), .A2(
        \SB1_0_0/i3[0] ), .ZN(\SB1_0_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_0/N4  ( .A1(\SB1_0_1/i0[7] ), .A2(
        \SB1_0_1/i0_3 ), .A3(\SB1_0_1/i0_0 ), .ZN(
        \SB1_0_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_1/Component_Function_0/N3  ( .A1(\SB1_0_1/i0[10] ), .A2(
        \SB1_0_1/i0_4 ), .A3(\SB1_0_1/i0_3 ), .ZN(
        \SB1_0_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_1/Component_Function_0/N2  ( .A1(\SB1_0_1/i0[8] ), .A2(
        \SB1_0_1/i0[7] ), .A3(\SB1_0_1/i0[6] ), .ZN(
        \SB1_0_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_1/Component_Function_0/N1  ( .A1(\SB1_0_1/i0[10] ), .A2(
        \SB1_0_1/i0[9] ), .ZN(\SB1_0_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_1/N4  ( .A1(\SB1_0_1/i1_7 ), .A2(
        \SB1_0_1/i0[8] ), .A3(\SB1_0_1/i0_4 ), .ZN(
        \SB1_0_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_1/Component_Function_1/N2  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i1_7 ), .A3(\SB1_0_1/i0[8] ), .ZN(
        \SB1_0_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_1/Component_Function_1/N1  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i1[9] ), .ZN(\SB1_0_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_5/N4  ( .A1(\SB1_0_1/i0[9] ), .A2(
        \SB1_0_1/i0[6] ), .A3(\SB1_0_1/i0_4 ), .ZN(
        \SB1_0_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_1/Component_Function_5/N2  ( .A1(\SB1_0_1/i0_0 ), .A2(
        \SB1_0_1/i0[6] ), .A3(\SB1_0_1/i0[10] ), .ZN(
        \SB1_0_1/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_1/Component_Function_5/N1  ( .A1(\SB1_0_1/i0_0 ), .A2(
        \SB1_0_1/i3[0] ), .ZN(\SB1_0_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_0/N4  ( .A1(\SB1_0_2/i0[7] ), .A2(
        \SB1_0_2/i0_3 ), .A3(\SB1_0_2/i0_0 ), .ZN(
        \SB1_0_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_0/N3  ( .A1(\SB1_0_2/i0[10] ), .A2(
        \SB1_0_2/i0_4 ), .A3(\SB1_0_2/i0_3 ), .ZN(
        \SB1_0_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_2/Component_Function_0/N2  ( .A1(\SB1_0_2/i0[8] ), .A2(
        \SB1_0_2/i0[7] ), .A3(\SB1_0_2/i0[6] ), .ZN(
        \SB1_0_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_2/Component_Function_0/N1  ( .A1(\SB1_0_2/i0[10] ), .A2(
        \SB1_0_2/i0[9] ), .ZN(\SB1_0_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_1/N4  ( .A1(\SB1_0_2/i1_7 ), .A2(
        \SB1_0_2/i0[8] ), .A3(\SB1_0_2/i0_4 ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_1/N3  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[6] ), .A3(\SB1_0_2/i0[9] ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_2/Component_Function_1/N2  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i1_7 ), .A3(\SB1_0_2/i0[8] ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_2/Component_Function_1/N1  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i1[9] ), .ZN(\SB1_0_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_5/N4  ( .A1(\SB1_0_2/i0[9] ), .A2(
        \SB1_0_2/i0[6] ), .A3(\SB1_0_2/i0_4 ), .ZN(
        \SB1_0_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_5/N2  ( .A1(\SB1_0_2/i0_0 ), .A2(
        \SB1_0_2/i0[6] ), .A3(\SB1_0_2/i0[10] ), .ZN(
        \SB1_0_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_2/Component_Function_5/N1  ( .A1(\SB1_0_2/i0_0 ), .A2(
        \SB1_0_2/i3[0] ), .ZN(\SB1_0_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_0/N4  ( .A1(\SB1_0_3/i0[7] ), .A2(
        \SB1_0_3/i0_3 ), .A3(\SB1_0_3/i0_0 ), .ZN(
        \SB1_0_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_0/N3  ( .A1(\SB1_0_3/i0[10] ), .A2(
        \SB1_0_3/i0_4 ), .A3(\SB1_0_3/i0_3 ), .ZN(
        \SB1_0_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_0/N2  ( .A1(\SB1_0_3/i0[8] ), .A2(
        \SB1_0_3/i0[7] ), .A3(\SB1_0_3/i0[6] ), .ZN(
        \SB1_0_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_3/Component_Function_0/N1  ( .A1(\SB1_0_3/i0[10] ), .A2(
        \SB1_0_3/i0[9] ), .ZN(\SB1_0_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N4  ( .A1(\SB1_0_3/i1_7 ), .A2(
        \SB1_0_3/i0[8] ), .A3(\SB1_0_3/i0_4 ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N3  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[6] ), .A3(\SB1_0_3/i0[9] ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N2  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i1_7 ), .A3(\SB1_0_3/i0[8] ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_3/Component_Function_1/N1  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i1[9] ), .ZN(\SB1_0_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_5/N4  ( .A1(\SB1_0_3/i0[9] ), .A2(
        \SB1_0_3/i0[6] ), .A3(\SB1_0_3/i0_4 ), .ZN(
        \SB1_0_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_5/N2  ( .A1(\SB1_0_3/i0_0 ), .A2(
        \SB1_0_3/i0[6] ), .A3(\SB1_0_3/i0[10] ), .ZN(
        \SB1_0_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_3/Component_Function_5/N1  ( .A1(\SB1_0_3/i0_0 ), .A2(
        \SB1_0_3/i3[0] ), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_0/N3  ( .A1(\SB1_0_4/i0[10] ), .A2(
        \SB1_0_4/i0_4 ), .A3(\SB1_0_4/i0_3 ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_0/N2  ( .A1(\SB1_0_4/i0[8] ), .A2(
        \SB1_0_4/i0[7] ), .A3(\SB1_0_4/i0[6] ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_4/Component_Function_0/N1  ( .A1(\SB1_0_4/i0[10] ), .A2(
        \SB1_0_4/i0[9] ), .ZN(\SB1_0_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_1/N4  ( .A1(\SB1_0_4/i1_7 ), .A2(
        \SB1_0_4/i0[8] ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_1/N2  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i1_7 ), .A3(\SB1_0_4/i0[8] ), .ZN(
        \SB1_0_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_4/Component_Function_1/N1  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i1[9] ), .ZN(\SB1_0_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_5/N2  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i0[6] ), .A3(\SB1_0_4/i0[10] ), .ZN(
        \SB1_0_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_4/Component_Function_5/N1  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i3[0] ), .ZN(\SB1_0_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_0/N4  ( .A1(\SB1_0_5/i0[7] ), .A2(
        \SB1_0_5/i0_3 ), .A3(\SB1_0_5/i0_0 ), .ZN(
        \SB1_0_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_5/Component_Function_0/N2  ( .A1(\SB1_0_5/i0[8] ), .A2(
        \SB1_0_5/i0[7] ), .A3(\SB1_0_5/i0[6] ), .ZN(
        \SB1_0_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_5/Component_Function_0/N1  ( .A1(\SB1_0_5/i0[10] ), .A2(
        \SB1_0_5/i0[9] ), .ZN(\SB1_0_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_1/N4  ( .A1(\SB1_0_5/i1_7 ), .A2(
        \SB1_0_5/i0[8] ), .A3(\SB1_0_5/i0_4 ), .ZN(
        \SB1_0_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_5/Component_Function_1/N3  ( .A1(\SB1_0_5/i1_5 ), .A2(
        \SB1_0_5/i0[6] ), .A3(\SB1_0_5/i0[9] ), .ZN(
        \SB1_0_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_5/Component_Function_1/N2  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i1_7 ), .A3(\SB1_0_5/i0[8] ), .ZN(
        \SB1_0_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_5/Component_Function_1/N1  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i1[9] ), .ZN(\SB1_0_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_5/N4  ( .A1(\SB1_0_5/i0[9] ), .A2(
        \SB1_0_5/i0[6] ), .A3(\SB1_0_5/i0_4 ), .ZN(
        \SB1_0_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_5/Component_Function_5/N2  ( .A1(\SB1_0_5/i0_0 ), .A2(
        \SB1_0_5/i0[6] ), .A3(\SB1_0_5/i0[10] ), .ZN(
        \SB1_0_5/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_5/Component_Function_5/N1  ( .A1(\SB1_0_5/i0_0 ), .A2(
        \SB1_0_5/i3[0] ), .ZN(\SB1_0_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_0/N2  ( .A1(\SB1_0_6/i0[8] ), .A2(
        \SB1_0_6/i0[7] ), .A3(\SB1_0_6/i0[6] ), .ZN(
        \SB1_0_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_6/Component_Function_0/N1  ( .A1(\SB1_0_6/i0[10] ), .A2(
        \SB1_0_6/i0[9] ), .ZN(\SB1_0_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_1/N4  ( .A1(\SB1_0_6/i1_7 ), .A2(
        \SB1_0_6/i0[8] ), .A3(\SB1_0_6/i0_4 ), .ZN(
        \SB1_0_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_1/N3  ( .A1(\SB1_0_6/i1_5 ), .A2(
        \SB1_0_6/i0[6] ), .A3(\SB1_0_6/i0[9] ), .ZN(
        \SB1_0_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_6/Component_Function_1/N2  ( .A1(n2136), .A2(\SB1_0_6/i1_7 ), 
        .A3(\SB1_0_6/i0[8] ), .ZN(\SB1_0_6/Component_Function_1/NAND4_in[1] )
         );
  NAND2_X1 \SB1_0_6/Component_Function_1/N1  ( .A1(n2136), .A2(\SB1_0_6/i1[9] ), .ZN(\SB1_0_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_5/N4  ( .A1(\SB1_0_6/i0[9] ), .A2(
        \SB1_0_6/i0[6] ), .A3(\SB1_0_6/i0_4 ), .ZN(
        \SB1_0_6/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_6/Component_Function_5/N1  ( .A1(\SB1_0_6/i0_0 ), .A2(
        \SB1_0_6/i3[0] ), .ZN(\SB1_0_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_0/N4  ( .A1(\SB1_0_7/i0[7] ), .A2(
        \SB1_0_7/i0_3 ), .A3(\SB1_0_7/i0_0 ), .ZN(
        \SB1_0_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_0/N3  ( .A1(\SB1_0_7/i0[10] ), .A2(
        \SB1_0_7/i0_4 ), .A3(\SB1_0_7/i0_3 ), .ZN(
        \SB1_0_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_0/N2  ( .A1(\SB1_0_7/i0[8] ), .A2(
        \SB1_0_7/i0[7] ), .A3(\SB1_0_7/i0[6] ), .ZN(
        \SB1_0_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_7/Component_Function_0/N1  ( .A1(\SB1_0_7/i0[10] ), .A2(
        \SB1_0_7/i0[9] ), .ZN(\SB1_0_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N4  ( .A1(\SB1_0_7/i1_7 ), .A2(
        \SB1_0_7/i0[8] ), .A3(\SB1_0_7/i0_4 ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N3  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0[6] ), .A3(\SB1_0_7/i0[9] ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N2  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i1_7 ), .A3(\SB1_0_7/i0[8] ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_7/Component_Function_1/N1  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i1[9] ), .ZN(\SB1_0_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_5/N4  ( .A1(\SB1_0_7/i0[9] ), .A2(
        \SB1_0_7/i0[6] ), .A3(\SB1_0_7/i0_4 ), .ZN(
        \SB1_0_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_5/N2  ( .A1(\SB1_0_7/i0_0 ), .A2(
        \SB1_0_7/i0[6] ), .A3(\SB1_0_7/i0[10] ), .ZN(
        \SB1_0_7/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_7/Component_Function_5/N1  ( .A1(\SB1_0_7/i0_0 ), .A2(
        \SB1_0_7/i3[0] ), .ZN(\SB1_0_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_0/N4  ( .A1(\SB1_0_8/i0[7] ), .A2(
        \SB1_0_8/i0_3 ), .A3(\SB1_0_8/i0_0 ), .ZN(
        \SB1_0_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_0/N3  ( .A1(\SB1_0_8/i0[10] ), .A2(
        \SB1_0_8/i0_4 ), .A3(\SB1_0_8/i0_3 ), .ZN(
        \SB1_0_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_8/Component_Function_0/N2  ( .A1(\SB1_0_8/i0[8] ), .A2(
        \SB1_0_8/i0[7] ), .A3(\SB1_0_8/i0[6] ), .ZN(
        \SB1_0_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_8/Component_Function_0/N1  ( .A1(\SB1_0_8/i0[10] ), .A2(
        \SB1_0_8/i0[9] ), .ZN(\SB1_0_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N4  ( .A1(\SB1_0_8/i1_7 ), .A2(
        \SB1_0_8/i0[8] ), .A3(\SB1_0_8/i0_4 ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N3  ( .A1(\SB1_0_8/i1_5 ), .A2(
        \SB1_0_8/i0[6] ), .A3(\SB1_0_8/i0[9] ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N2  ( .A1(n1664), .A2(\SB1_0_8/i1_7 ), 
        .A3(\SB1_0_8/i0[8] ), .ZN(\SB1_0_8/Component_Function_1/NAND4_in[1] )
         );
  NAND2_X1 \SB1_0_8/Component_Function_1/N1  ( .A1(n1664), .A2(\SB1_0_8/i1[9] ), .ZN(\SB1_0_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_5/N4  ( .A1(\SB1_0_8/i0[9] ), .A2(
        \SB1_0_8/i0[6] ), .A3(\SB1_0_8/i0_4 ), .ZN(
        \SB1_0_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_5/N2  ( .A1(\SB1_0_8/i0_0 ), .A2(
        \SB1_0_8/i0[6] ), .A3(\SB1_0_8/i0[10] ), .ZN(
        \SB1_0_8/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_8/Component_Function_5/N1  ( .A1(\SB1_0_8/i0_0 ), .A2(
        \SB1_0_8/i3[0] ), .ZN(\SB1_0_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_0/N4  ( .A1(\SB1_0_9/i0[7] ), .A2(
        \SB1_0_9/i0_3 ), .A3(\SB1_0_9/i0_0 ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_0/N2  ( .A1(\SB1_0_9/i0[8] ), .A2(
        \SB1_0_9/i0[7] ), .A3(\SB1_0_9/i0[6] ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_9/Component_Function_0/N1  ( .A1(\SB1_0_9/i0[10] ), .A2(
        \SB1_0_9/i0[9] ), .ZN(\SB1_0_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_1/N4  ( .A1(\SB1_0_9/i1_7 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_1/N2  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i1_7 ), .A3(\SB1_0_9/i0[8] ), .ZN(
        \SB1_0_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_9/Component_Function_1/N1  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i1[9] ), .ZN(\SB1_0_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_5/N2  ( .A1(\SB1_0_9/i0_0 ), .A2(
        \SB1_0_9/i0[6] ), .A3(\SB1_0_9/i0[10] ), .ZN(
        \SB1_0_9/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_9/Component_Function_5/N1  ( .A1(\SB1_0_9/i0_0 ), .A2(
        \SB1_0_9/i3[0] ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_0/N4  ( .A1(\SB1_0_10/i0[7] ), .A2(
        \SB1_0_10/i0_3 ), .A3(\SB1_0_10/i0_0 ), .ZN(
        \SB1_0_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_0/N2  ( .A1(\SB1_0_10/i0[8] ), .A2(
        \SB1_0_10/i0[7] ), .A3(\SB1_0_10/i0[6] ), .ZN(
        \SB1_0_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_10/Component_Function_0/N1  ( .A1(\SB1_0_10/i0[10] ), .A2(
        \SB1_0_10/i0[9] ), .ZN(\SB1_0_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N4  ( .A1(\SB1_0_10/i1_7 ), .A2(
        \SB1_0_10/i0[8] ), .A3(\SB1_0_10/i0_4 ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N3  ( .A1(\SB1_0_10/i1_5 ), .A2(
        \SB1_0_10/i0[6] ), .A3(\SB1_0_10/i0[9] ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N2  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i1_7 ), .A3(\SB1_0_10/i0[8] ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_10/Component_Function_1/N1  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i1[9] ), .ZN(\SB1_0_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_5/N4  ( .A1(\SB1_0_10/i0[9] ), .A2(
        \SB1_0_10/i0[6] ), .A3(\SB1_0_10/i0_4 ), .ZN(
        \SB1_0_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_5/N2  ( .A1(\SB1_0_10/i0_0 ), .A2(
        \SB1_0_10/i0[6] ), .A3(\SB1_0_10/i0[10] ), .ZN(
        \SB1_0_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_10/Component_Function_5/N1  ( .A1(\SB1_0_10/i0_0 ), .A2(
        \SB1_0_10/i3[0] ), .ZN(\SB1_0_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_0/N3  ( .A1(\SB1_0_11/i0[10] ), .A2(
        \SB1_0_11/i0_4 ), .A3(\SB1_0_11/i0_3 ), .ZN(
        \SB1_0_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_0/N2  ( .A1(\SB1_0_11/i0[8] ), .A2(
        \SB1_0_11/i0[7] ), .A3(\SB1_0_11/i0[6] ), .ZN(
        \SB1_0_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_11/Component_Function_0/N1  ( .A1(\SB1_0_11/i0[10] ), .A2(
        \SB1_0_11/i0[9] ), .ZN(\SB1_0_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_1/N3  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0[6] ), .A3(\SB1_0_11/i0[9] ), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_1/N2  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i1_7 ), .A3(\SB1_0_11/i0[8] ), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_11/Component_Function_1/N1  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i1[9] ), .ZN(\SB1_0_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_5/N4  ( .A1(\SB1_0_11/i0[9] ), .A2(
        \SB1_0_11/i0[6] ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_5/N2  ( .A1(\SB1_0_11/i0_0 ), .A2(
        \SB1_0_11/i0[6] ), .A3(\SB1_0_11/i0[10] ), .ZN(
        \SB1_0_11/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_11/Component_Function_5/N1  ( .A1(\SB1_0_11/i0_0 ), .A2(
        \SB1_0_11/i3[0] ), .ZN(\SB1_0_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_0/N2  ( .A1(\SB1_0_12/i0[8] ), .A2(
        \SB1_0_12/i0[7] ), .A3(\SB1_0_12/i0[6] ), .ZN(
        \SB1_0_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_12/Component_Function_0/N1  ( .A1(\SB1_0_12/i0[10] ), .A2(
        \SB1_0_12/i0[9] ), .ZN(\SB1_0_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N4  ( .A1(\SB1_0_12/i1_7 ), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N3  ( .A1(n381), .A2(
        \SB1_0_12/i0[6] ), .A3(\SB1_0_12/i0[9] ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N2  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i1_7 ), .A3(\SB1_0_12/i0[8] ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_12/Component_Function_1/N1  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i1[9] ), .ZN(\SB1_0_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_5/N4  ( .A1(\SB1_0_12/i0[9] ), .A2(
        \SB1_0_12/i0[6] ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_5/N2  ( .A1(\SB1_0_12/i0_0 ), .A2(
        \SB1_0_12/i0[6] ), .A3(\SB1_0_12/i0[10] ), .ZN(
        \SB1_0_12/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_12/Component_Function_5/N1  ( .A1(\SB1_0_12/i0_0 ), .A2(
        \SB1_0_12/i3[0] ), .ZN(\SB1_0_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_0/N4  ( .A1(\SB1_0_13/i0[7] ), .A2(
        \SB1_0_13/i0_3 ), .A3(\SB1_0_13/i0_0 ), .ZN(
        \SB1_0_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_0/N3  ( .A1(\SB1_0_13/i0[10] ), .A2(
        \SB1_0_13/i0_4 ), .A3(\SB1_0_13/i0_3 ), .ZN(
        \SB1_0_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_13/Component_Function_0/N2  ( .A1(\SB1_0_13/i0[8] ), .A2(
        \SB1_0_13/i0[7] ), .A3(\SB1_0_13/i0[6] ), .ZN(
        \SB1_0_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_13/Component_Function_0/N1  ( .A1(\SB1_0_13/i0[10] ), .A2(
        \SB1_0_13/i0[9] ), .ZN(\SB1_0_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_1/N4  ( .A1(\SB1_0_13/i1_7 ), .A2(
        \SB1_0_13/i0[8] ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_1/N3  ( .A1(\SB1_0_13/i1_5 ), .A2(
        \SB1_0_13/i0[6] ), .A3(\SB1_0_13/i0[9] ), .ZN(
        \SB1_0_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_13/Component_Function_1/N2  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i1_7 ), .A3(\SB1_0_13/i0[8] ), .ZN(
        \SB1_0_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_13/Component_Function_1/N1  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i1[9] ), .ZN(\SB1_0_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_5/N4  ( .A1(\SB1_0_13/i0[9] ), .A2(
        \SB1_0_13/i0[6] ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_5/N2  ( .A1(\SB1_0_13/i0_0 ), .A2(
        \SB1_0_13/i0[6] ), .A3(\SB1_0_13/i0[10] ), .ZN(
        \SB1_0_13/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_13/Component_Function_5/N1  ( .A1(\SB1_0_13/i0_0 ), .A2(
        \SB1_0_13/i3[0] ), .ZN(\SB1_0_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_0/N3  ( .A1(\SB1_0_14/i0[10] ), .A2(
        \SB1_0_14/i0_4 ), .A3(n862), .ZN(
        \SB1_0_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_0/N2  ( .A1(\SB1_0_14/i0[8] ), .A2(
        \SB1_0_14/i0[7] ), .A3(\SB1_0_14/i0[6] ), .ZN(
        \SB1_0_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_14/Component_Function_0/N1  ( .A1(\SB1_0_14/i0[10] ), .A2(
        \SB1_0_14/i0[9] ), .ZN(\SB1_0_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N4  ( .A1(\SB1_0_14/i1_7 ), .A2(
        \SB1_0_14/i0[8] ), .A3(\SB1_0_14/i0_4 ), .ZN(
        \SB1_0_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N3  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[6] ), .A3(\SB1_0_14/i0[9] ), .ZN(
        \SB1_0_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N2  ( .A1(n862), .A2(\SB1_0_14/i1_7 ), .A3(\SB1_0_14/i0[8] ), .ZN(\SB1_0_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_14/Component_Function_1/N1  ( .A1(n862), .A2(
        \SB1_0_14/i1[9] ), .ZN(\SB1_0_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_5/N4  ( .A1(\SB1_0_14/i0[9] ), .A2(
        \SB1_0_14/i0[6] ), .A3(\SB1_0_14/i0_4 ), .ZN(
        \SB1_0_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_5/N2  ( .A1(\SB1_0_14/i0_0 ), .A2(
        \SB1_0_14/i0[6] ), .A3(\SB1_0_14/i0[10] ), .ZN(
        \SB1_0_14/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_14/Component_Function_5/N1  ( .A1(\SB1_0_14/i0_0 ), .A2(
        \SB1_0_14/i3[0] ), .ZN(\SB1_0_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_0/N4  ( .A1(\SB1_0_15/i0[7] ), .A2(
        \SB1_0_15/i0_3 ), .A3(\SB1_0_15/i0_0 ), .ZN(
        \SB1_0_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_0/N2  ( .A1(\SB1_0_15/i0[8] ), .A2(
        \SB1_0_15/i0[7] ), .A3(\SB1_0_15/i0[6] ), .ZN(
        \SB1_0_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_15/Component_Function_0/N1  ( .A1(\SB1_0_15/i0[10] ), .A2(
        \SB1_0_15/i0[9] ), .ZN(\SB1_0_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_1/N4  ( .A1(\SB1_0_15/i1_7 ), .A2(
        \SB1_0_15/i0[8] ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_1/N3  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0[6] ), .A3(\SB1_0_15/i0[9] ), .ZN(
        \SB1_0_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_15/Component_Function_1/N2  ( .A1(\SB1_0_15/i0_3 ), .A2(
        \SB1_0_15/i1_7 ), .A3(\SB1_0_15/i0[8] ), .ZN(
        \SB1_0_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_15/Component_Function_1/N1  ( .A1(\SB1_0_15/i0_3 ), .A2(
        \SB1_0_15/i1[9] ), .ZN(\SB1_0_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_5/N4  ( .A1(\SB1_0_15/i0[9] ), .A2(
        \SB1_0_15/i0[6] ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_5/N2  ( .A1(\SB1_0_15/i0_0 ), .A2(
        \SB1_0_15/i0[6] ), .A3(\SB1_0_15/i0[10] ), .ZN(
        \SB1_0_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_15/Component_Function_5/N1  ( .A1(\SB1_0_15/i0_0 ), .A2(
        \SB1_0_15/i3[0] ), .ZN(\SB1_0_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_0/N4  ( .A1(\SB1_0_16/i0[7] ), .A2(
        \SB1_0_16/i0_3 ), .A3(\SB1_0_16/i0_0 ), .ZN(
        \SB1_0_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_0/N3  ( .A1(\SB1_0_16/i0[10] ), .A2(
        \SB1_0_16/i0_4 ), .A3(\SB1_0_16/i0_3 ), .ZN(
        \SB1_0_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_16/Component_Function_0/N2  ( .A1(\SB1_0_16/i0[8] ), .A2(
        \SB1_0_16/i0[7] ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_16/Component_Function_0/N1  ( .A1(\SB1_0_16/i0[10] ), .A2(
        \SB1_0_16/i0[9] ), .ZN(\SB1_0_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_1/N4  ( .A1(\SB1_0_16/i1_7 ), .A2(
        \SB1_0_16/i0[8] ), .A3(\SB1_0_16/i0_4 ), .ZN(
        \SB1_0_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_1/N3  ( .A1(\SB1_0_16/i1_5 ), .A2(
        \SB1_0_16/i0[6] ), .A3(\SB1_0_16/i0[9] ), .ZN(
        \SB1_0_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_16/Component_Function_1/N2  ( .A1(\SB1_0_16/i0_3 ), .A2(
        \SB1_0_16/i1_7 ), .A3(\SB1_0_16/i0[8] ), .ZN(
        \SB1_0_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_16/Component_Function_1/N1  ( .A1(\SB1_0_16/i0_3 ), .A2(
        \SB1_0_16/i1[9] ), .ZN(\SB1_0_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_5/N4  ( .A1(\SB1_0_16/i0[9] ), .A2(
        \SB1_0_16/i0[6] ), .A3(\SB1_0_16/i0_4 ), .ZN(
        \SB1_0_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_5/N2  ( .A1(\SB1_0_16/i0_0 ), .A2(
        \SB1_0_16/i0[6] ), .A3(\SB1_0_16/i0[10] ), .ZN(
        \SB1_0_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_16/Component_Function_5/N1  ( .A1(\SB1_0_16/i0_0 ), .A2(
        \SB1_0_16/i3[0] ), .ZN(\SB1_0_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_0/N4  ( .A1(\SB1_0_17/i0[7] ), .A2(
        \SB1_0_17/i0_3 ), .A3(\SB1_0_17/i0_0 ), .ZN(
        \SB1_0_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_0/N3  ( .A1(\SB1_0_17/i0[10] ), .A2(
        \SB1_0_17/i0_4 ), .A3(\SB1_0_17/i0_3 ), .ZN(
        \SB1_0_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_17/Component_Function_0/N2  ( .A1(\SB1_0_17/i0[8] ), .A2(
        \SB1_0_17/i0[7] ), .A3(\SB1_0_17/i0[6] ), .ZN(
        \SB1_0_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_17/Component_Function_0/N1  ( .A1(\SB1_0_17/i0[10] ), .A2(
        \SB1_0_17/i0[9] ), .ZN(\SB1_0_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_1/N4  ( .A1(\SB1_0_17/i1_7 ), .A2(
        \SB1_0_17/i0[8] ), .A3(\SB1_0_17/i0_4 ), .ZN(
        \SB1_0_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_1/N3  ( .A1(\SB1_0_17/i1_5 ), .A2(
        \SB1_0_17/i0[6] ), .A3(\SB1_0_17/i0[9] ), .ZN(
        \SB1_0_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_17/Component_Function_1/N2  ( .A1(\SB1_0_17/i0_3 ), .A2(
        \SB1_0_17/i1_7 ), .A3(\SB1_0_17/i0[8] ), .ZN(
        \SB1_0_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_17/Component_Function_1/N1  ( .A1(\SB1_0_17/i0_3 ), .A2(
        \SB1_0_17/i1[9] ), .ZN(\SB1_0_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_5/N4  ( .A1(\SB1_0_17/i0[9] ), .A2(
        \SB1_0_17/i0[6] ), .A3(\SB1_0_17/i0_4 ), .ZN(
        \SB1_0_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_5/N2  ( .A1(\SB1_0_17/i0_0 ), .A2(
        \SB1_0_17/i0[6] ), .A3(\SB1_0_17/i0[10] ), .ZN(
        \SB1_0_17/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_17/Component_Function_5/N1  ( .A1(\SB1_0_17/i0_0 ), .A2(
        \SB1_0_17/i3[0] ), .ZN(\SB1_0_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_0/N4  ( .A1(\SB1_0_18/i0[7] ), .A2(
        \SB1_0_18/i0_3 ), .A3(\SB1_0_18/i0_0 ), .ZN(
        \SB1_0_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_0/N2  ( .A1(\SB1_0_18/i0[8] ), .A2(
        \SB1_0_18/i0[7] ), .A3(\SB1_0_18/i0[6] ), .ZN(
        \SB1_0_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_18/Component_Function_0/N1  ( .A1(\SB1_0_18/i0[10] ), .A2(
        \SB1_0_18/i0[9] ), .ZN(\SB1_0_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_1/N4  ( .A1(\SB1_0_18/i1_7 ), .A2(n111), .A3(\SB1_0_18/i0_4 ), .ZN(\SB1_0_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_1/N3  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0[6] ), .A3(\SB1_0_18/i0[9] ), .ZN(
        \SB1_0_18/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_18/Component_Function_1/N1  ( .A1(\SB1_0_18/i0_3 ), .A2(
        \SB1_0_18/i1[9] ), .ZN(\SB1_0_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_5/N4  ( .A1(\SB1_0_18/i0[9] ), .A2(
        \SB1_0_18/i0[6] ), .A3(\SB1_0_18/i0_4 ), .ZN(
        \SB1_0_18/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_18/Component_Function_5/N1  ( .A1(\SB1_0_18/i0_0 ), .A2(
        \SB1_0_18/i3[0] ), .ZN(\SB1_0_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_0/N4  ( .A1(\SB1_0_19/i0[7] ), .A2(
        n873), .A3(\SB1_0_19/i0_0 ), .ZN(
        \SB1_0_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_0/N3  ( .A1(\SB1_0_19/i0[10] ), .A2(
        \SB1_0_19/i0_4 ), .A3(n873), .ZN(
        \SB1_0_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_0/N2  ( .A1(\SB1_0_19/i0[8] ), .A2(
        \SB1_0_19/i0[7] ), .A3(\SB1_0_19/i0[6] ), .ZN(
        \SB1_0_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_19/Component_Function_0/N1  ( .A1(\SB1_0_19/i0[10] ), .A2(
        \SB1_0_19/i0[9] ), .ZN(\SB1_0_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_1/N4  ( .A1(\SB1_0_19/i1_7 ), .A2(
        \SB1_0_19/i0[8] ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_1/N2  ( .A1(n873), .A2(\SB1_0_19/i1_7 ), .A3(\SB1_0_19/i0[8] ), .ZN(\SB1_0_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_19/Component_Function_1/N1  ( .A1(n873), .A2(
        \SB1_0_19/i1[9] ), .ZN(\SB1_0_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_5/N2  ( .A1(\SB1_0_19/i0_0 ), .A2(
        \SB1_0_19/i0[6] ), .A3(\SB1_0_19/i0[10] ), .ZN(
        \SB1_0_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_19/Component_Function_5/N1  ( .A1(\SB1_0_19/i0_0 ), .A2(
        \SB1_0_19/i3[0] ), .ZN(\SB1_0_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_0/N3  ( .A1(\SB1_0_20/i0[10] ), .A2(
        \SB1_0_20/i0_4 ), .A3(\SB1_0_20/i0_3 ), .ZN(
        \SB1_0_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_20/Component_Function_0/N2  ( .A1(\SB1_0_20/i0[8] ), .A2(
        \SB1_0_20/i0[7] ), .A3(\SB1_0_20/i0[6] ), .ZN(
        \SB1_0_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_20/Component_Function_0/N1  ( .A1(\SB1_0_20/i0[10] ), .A2(
        \SB1_0_20/i0[9] ), .ZN(\SB1_0_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_1/N4  ( .A1(\SB1_0_20/i1_7 ), .A2(
        \SB1_0_20/i0[8] ), .A3(\SB1_0_20/i0_4 ), .ZN(
        \SB1_0_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_1/N3  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0[6] ), .A3(\SB1_0_20/i0[9] ), .ZN(
        \SB1_0_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_20/Component_Function_1/N2  ( .A1(\SB1_0_20/i0_3 ), .A2(
        \SB1_0_20/i1_7 ), .A3(\SB1_0_20/i0[8] ), .ZN(
        \SB1_0_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_20/Component_Function_1/N1  ( .A1(\SB1_0_20/i0_3 ), .A2(
        \SB1_0_20/i1[9] ), .ZN(\SB1_0_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_5/N4  ( .A1(\SB1_0_20/i0[9] ), .A2(
        \SB1_0_20/i0[6] ), .A3(\SB1_0_20/i0_4 ), .ZN(
        \SB1_0_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_5/N2  ( .A1(\SB1_0_20/i0_0 ), .A2(
        \SB1_0_20/i0[6] ), .A3(\SB1_0_20/i0[10] ), .ZN(
        \SB1_0_20/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_20/Component_Function_5/N1  ( .A1(\SB1_0_20/i0_0 ), .A2(
        \SB1_0_20/i3[0] ), .ZN(\SB1_0_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_0/N3  ( .A1(\SB1_0_21/i0[10] ), .A2(
        \SB1_0_21/i0_4 ), .A3(\SB1_0_21/i0_3 ), .ZN(
        \SB1_0_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_21/Component_Function_0/N2  ( .A1(\SB1_0_21/i0[8] ), .A2(
        \SB1_0_21/i0[7] ), .A3(\SB1_0_21/i0[6] ), .ZN(
        \SB1_0_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_21/Component_Function_0/N1  ( .A1(\SB1_0_21/i0[10] ), .A2(
        \SB1_0_21/i0[9] ), .ZN(\SB1_0_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_1/N4  ( .A1(\SB1_0_21/i1_7 ), .A2(
        \SB1_0_21/i0[8] ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_21/Component_Function_1/N3  ( .A1(\SB1_0_21/i1_5 ), .A2(
        \SB1_0_21/i0[6] ), .A3(\SB1_0_21/i0[9] ), .ZN(
        \SB1_0_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_21/Component_Function_1/N2  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i1_7 ), .A3(\SB1_0_21/i0[8] ), .ZN(
        \SB1_0_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_21/Component_Function_1/N1  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i1[9] ), .ZN(\SB1_0_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_5/N4  ( .A1(\SB1_0_21/i0[9] ), .A2(
        \SB1_0_21/i0[6] ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_21/Component_Function_5/N2  ( .A1(\SB1_0_21/i0_0 ), .A2(
        \SB1_0_21/i0[6] ), .A3(\SB1_0_21/i0[10] ), .ZN(
        \SB1_0_21/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_21/Component_Function_5/N1  ( .A1(\SB1_0_21/i0_0 ), .A2(
        \SB1_0_21/i3[0] ), .ZN(\SB1_0_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_0/N2  ( .A1(\SB1_0_22/i0[8] ), .A2(
        \SB1_0_22/i0[7] ), .A3(\SB1_0_22/i0[6] ), .ZN(
        \SB1_0_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_22/Component_Function_0/N1  ( .A1(\SB1_0_22/i0[10] ), .A2(
        \SB1_0_22/i0[9] ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_1/N3  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[6] ), .A3(\SB1_0_22/i0[9] ), .ZN(
        \SB1_0_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_22/Component_Function_1/N2  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i1_7 ), .A3(\SB1_0_22/i0[8] ), .ZN(
        \SB1_0_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_22/Component_Function_1/N1  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i1[9] ), .ZN(\SB1_0_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_5/N4  ( .A1(\SB1_0_22/i0[9] ), .A2(
        \SB1_0_22/i0[6] ), .A3(\SB1_0_22/i0_4 ), .ZN(
        \SB1_0_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_5/N2  ( .A1(\SB1_0_22/i0_0 ), .A2(
        \SB1_0_22/i0[6] ), .A3(\SB1_0_22/i0[10] ), .ZN(
        \SB1_0_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_22/Component_Function_5/N1  ( .A1(\SB1_0_22/i0_0 ), .A2(
        \SB1_0_22/i3[0] ), .ZN(\SB1_0_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_0/N2  ( .A1(\SB1_0_23/i0[8] ), .A2(
        \SB1_0_23/i0[7] ), .A3(\SB1_0_23/i0[6] ), .ZN(
        \SB1_0_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_23/Component_Function_0/N1  ( .A1(\SB1_0_23/i0[10] ), .A2(
        \SB1_0_23/i0[9] ), .ZN(\SB1_0_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_1/N4  ( .A1(\SB1_0_23/i1_7 ), .A2(
        \SB1_0_23/i0[8] ), .A3(\SB1_0_23/i0_4 ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_1/N3  ( .A1(\SB1_0_23/i1_5 ), .A2(
        \SB1_0_23/i0[6] ), .A3(\SB1_0_23/i0[9] ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_23/Component_Function_1/N2  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i1_7 ), .A3(\SB1_0_23/i0[8] ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_23/Component_Function_1/N1  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i1[9] ), .ZN(\SB1_0_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_5/N4  ( .A1(\SB1_0_23/i0[9] ), .A2(
        \SB1_0_23/i0[6] ), .A3(\SB1_0_23/i0_4 ), .ZN(
        \SB1_0_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_5/N2  ( .A1(\SB1_0_23/i0_0 ), .A2(
        \SB1_0_23/i0[6] ), .A3(\SB1_0_23/i0[10] ), .ZN(
        \SB1_0_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_24/Component_Function_0/N4  ( .A1(\SB1_0_24/i0[7] ), .A2(
        \SB1_0_24/i0_3 ), .A3(\SB1_0_24/i0_0 ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_0/N3  ( .A1(\SB1_0_24/i0[10] ), .A2(
        \SB1_0_24/i0_4 ), .A3(\SB1_0_24/i0_3 ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_24/Component_Function_0/N2  ( .A1(\SB1_0_24/i0[8] ), .A2(
        \SB1_0_24/i0[7] ), .A3(\SB1_0_24/i0[6] ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_24/Component_Function_0/N1  ( .A1(\SB1_0_24/i0[10] ), .A2(
        \SB1_0_24/i0[9] ), .ZN(\SB1_0_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_1/N4  ( .A1(\SB1_0_24/i1_7 ), .A2(
        \SB1_0_24/i0[8] ), .A3(\SB1_0_24/i0_4 ), .ZN(
        \SB1_0_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_1/N3  ( .A1(\SB1_0_24/i1_5 ), .A2(
        \SB1_0_24/i0[6] ), .A3(\SB1_0_24/i0[9] ), .ZN(
        \SB1_0_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_24/Component_Function_1/N2  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i1_7 ), .A3(\SB1_0_24/i0[8] ), .ZN(
        \SB1_0_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_24/Component_Function_1/N1  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i1[9] ), .ZN(\SB1_0_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_5/N4  ( .A1(\SB1_0_24/i0[9] ), .A2(
        \SB1_0_24/i0[6] ), .A3(\SB1_0_24/i0_4 ), .ZN(
        \SB1_0_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_5/N2  ( .A1(\SB1_0_24/i0_0 ), .A2(
        \SB1_0_24/i0[6] ), .A3(\SB1_0_24/i0[10] ), .ZN(
        \SB1_0_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_24/Component_Function_5/N1  ( .A1(\SB1_0_24/i0_0 ), .A2(
        \SB1_0_24/i3[0] ), .ZN(\SB1_0_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_0/N3  ( .A1(\SB1_0_25/i0[10] ), .A2(
        \SB1_0_25/i0_4 ), .A3(\SB1_0_25/i0_3 ), .ZN(
        \SB1_0_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_25/Component_Function_0/N2  ( .A1(\SB1_0_25/i0[8] ), .A2(
        \SB1_0_25/i0[7] ), .A3(\SB1_0_25/i0[6] ), .ZN(
        \SB1_0_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_25/Component_Function_0/N1  ( .A1(\SB1_0_25/i0[10] ), .A2(
        \SB1_0_25/i0[9] ), .ZN(\SB1_0_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_1/N4  ( .A1(\SB1_0_25/i1_7 ), .A2(
        \SB1_0_25/i0[8] ), .A3(\SB1_0_25/i0_4 ), .ZN(
        \SB1_0_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_25/Component_Function_1/N3  ( .A1(\SB1_0_25/i1_5 ), .A2(
        \SB1_0_25/i0[6] ), .A3(\SB1_0_25/i0[9] ), .ZN(
        \SB1_0_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_25/Component_Function_1/N2  ( .A1(\SB1_0_25/i0_3 ), .A2(
        \SB1_0_25/i1_7 ), .A3(\SB1_0_25/i0[8] ), .ZN(
        \SB1_0_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_25/Component_Function_1/N1  ( .A1(\SB1_0_25/i0_3 ), .A2(
        \SB1_0_25/i1[9] ), .ZN(\SB1_0_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_5/N4  ( .A1(\SB1_0_25/i0[9] ), .A2(
        \SB1_0_25/i0[6] ), .A3(\SB1_0_25/i0_4 ), .ZN(
        \SB1_0_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_25/Component_Function_5/N2  ( .A1(\SB1_0_25/i0_0 ), .A2(
        \SB1_0_25/i0[6] ), .A3(\SB1_0_25/i0[10] ), .ZN(
        \SB1_0_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_25/Component_Function_5/N1  ( .A1(\SB1_0_25/i0_0 ), .A2(
        \SB1_0_25/i3[0] ), .ZN(\SB1_0_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_0/N3  ( .A1(\SB1_0_26/i0[10] ), .A2(
        \SB1_0_26/i0_4 ), .A3(\SB1_0_26/i0_3 ), .ZN(
        \SB1_0_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_26/Component_Function_0/N2  ( .A1(\SB1_0_26/i0[8] ), .A2(
        \SB1_0_26/i0[7] ), .A3(\SB1_0_26/i0[6] ), .ZN(
        \SB1_0_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_26/Component_Function_0/N1  ( .A1(\SB1_0_26/i0[10] ), .A2(
        \SB1_0_26/i0[9] ), .ZN(\SB1_0_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_1/N4  ( .A1(\SB1_0_26/i1_7 ), .A2(
        \SB1_0_26/i0[8] ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_1/N3  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0[6] ), .A3(\SB1_0_26/i0[9] ), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_26/Component_Function_1/N2  ( .A1(\SB1_0_26/i0_3 ), .A2(
        \SB1_0_26/i1_7 ), .A3(\SB1_0_26/i0[8] ), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_26/Component_Function_1/N1  ( .A1(\SB1_0_26/i0_3 ), .A2(
        \SB1_0_26/i1[9] ), .ZN(\SB1_0_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_5/N4  ( .A1(\SB1_0_26/i0[9] ), .A2(
        \SB1_0_26/i0[6] ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_5/N2  ( .A1(\SB1_0_26/i0_0 ), .A2(
        \SB1_0_26/i0[6] ), .A3(\SB1_0_26/i0[10] ), .ZN(
        \SB1_0_26/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_26/Component_Function_5/N1  ( .A1(\SB1_0_26/i0_0 ), .A2(
        \SB1_0_26/i3[0] ), .ZN(\SB1_0_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N4  ( .A1(\SB1_0_27/i0[7] ), .A2(
        \SB1_0_27/i0_3 ), .A3(\SB1_0_27/i0_0 ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N3  ( .A1(\SB1_0_27/i0[10] ), .A2(
        \SB1_0_27/i0_4 ), .A3(\SB1_0_27/i0_3 ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N2  ( .A1(\SB1_0_27/i0[8] ), .A2(
        \SB1_0_27/i0[7] ), .A3(\SB1_0_27/i0[6] ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_27/Component_Function_0/N1  ( .A1(\SB1_0_27/i0[10] ), .A2(
        \SB1_0_27/i0[9] ), .ZN(\SB1_0_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N4  ( .A1(\SB1_0_27/i1_7 ), .A2(
        \SB1_0_27/i0[8] ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N3  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0[6] ), .A3(\SB1_0_27/i0[9] ), .ZN(
        \SB1_0_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N2  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i1_7 ), .A3(\SB1_0_27/i0[8] ), .ZN(
        \SB1_0_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_27/Component_Function_1/N1  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i1[9] ), .ZN(\SB1_0_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_5/N4  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0[6] ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_5/N2  ( .A1(\SB1_0_27/i0[10] ), .A2(
        \SB1_0_27/i0[6] ), .A3(\SB1_0_27/i0_0 ), .ZN(
        \SB1_0_27/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_27/Component_Function_5/N1  ( .A1(\SB1_0_27/i0_0 ), .A2(
        \SB1_0_27/i3[0] ), .ZN(\SB1_0_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_0/N2  ( .A1(\SB1_0_28/i0[8] ), .A2(
        \SB1_0_28/i0[7] ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_28/Component_Function_0/N1  ( .A1(\SB1_0_28/i0[10] ), .A2(
        \SB1_0_28/i0[9] ), .ZN(\SB1_0_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_1/N4  ( .A1(\SB1_0_28/i1_7 ), .A2(
        \SB1_0_28/i0[8] ), .A3(\SB1_0_28/i0_4 ), .ZN(
        \SB1_0_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_1/N3  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0[6] ), .A3(\SB1_0_28/i0[9] ), .ZN(
        \SB1_0_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_28/Component_Function_1/N2  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i1_7 ), .A3(\SB1_0_28/i0[8] ), .ZN(
        \SB1_0_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_28/Component_Function_1/N1  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i1[9] ), .ZN(\SB1_0_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_5/N4  ( .A1(\SB1_0_28/i0[9] ), .A2(
        \SB1_0_28/i0[6] ), .A3(\SB1_0_28/i0_4 ), .ZN(
        \SB1_0_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_5/N2  ( .A1(\SB1_0_28/i0_0 ), .A2(
        \SB1_0_28/i0[6] ), .A3(\SB1_0_28/i0[10] ), .ZN(
        \SB1_0_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_28/Component_Function_5/N1  ( .A1(\SB1_0_28/i0_0 ), .A2(
        \SB1_0_28/i3[0] ), .ZN(\SB1_0_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_0/N4  ( .A1(\SB1_0_29/i0[7] ), .A2(
        \SB1_0_29/i0_3 ), .A3(\SB1_0_29/i0_0 ), .ZN(
        \SB1_0_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_0/N2  ( .A1(\SB1_0_29/i0[8] ), .A2(
        \SB1_0_29/i0[7] ), .A3(\SB1_0_29/i0[6] ), .ZN(
        \SB1_0_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_29/Component_Function_0/N1  ( .A1(\SB1_0_29/i0[10] ), .A2(
        \SB1_0_29/i0[9] ), .ZN(\SB1_0_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_1/N3  ( .A1(\SB1_0_29/i1_5 ), .A2(
        \SB1_0_29/i0[6] ), .A3(\SB1_0_29/i0[9] ), .ZN(
        \SB1_0_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_29/Component_Function_1/N2  ( .A1(\SB1_0_29/i0_3 ), .A2(
        \SB1_0_29/i1_7 ), .A3(\SB1_0_29/i0[8] ), .ZN(
        \SB1_0_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_29/Component_Function_1/N1  ( .A1(\SB1_0_29/i0_3 ), .A2(
        \SB1_0_29/i1[9] ), .ZN(\SB1_0_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_5/N4  ( .A1(\SB1_0_29/i0[9] ), .A2(
        \SB1_0_29/i0[6] ), .A3(\SB1_0_29/i0_4 ), .ZN(
        \SB1_0_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_5/N2  ( .A1(\SB1_0_29/i0_0 ), .A2(
        \SB1_0_29/i0[6] ), .A3(\SB1_0_29/i0[10] ), .ZN(
        \SB1_0_29/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_29/Component_Function_5/N1  ( .A1(\SB1_0_29/i0_0 ), .A2(
        \SB1_0_29/i3[0] ), .ZN(\SB1_0_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_0/N4  ( .A1(\SB1_0_30/i0[7] ), .A2(
        \SB1_0_30/i0_3 ), .A3(\SB1_0_30/i0_0 ), .ZN(
        \SB1_0_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_0/N3  ( .A1(\SB1_0_30/i0[10] ), .A2(
        \SB1_0_30/i0_4 ), .A3(\SB1_0_30/i0_3 ), .ZN(
        \SB1_0_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_30/Component_Function_0/N2  ( .A1(\SB1_0_30/i0[8] ), .A2(
        \SB1_0_30/i0[7] ), .A3(\SB1_0_30/i0[6] ), .ZN(
        \SB1_0_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_30/Component_Function_0/N1  ( .A1(\SB1_0_30/i0[10] ), .A2(
        \SB1_0_30/i0[9] ), .ZN(\SB1_0_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_1/N4  ( .A1(\SB1_0_30/i1_7 ), .A2(
        \SB1_0_30/i0[8] ), .A3(\SB1_0_30/i0_4 ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_1/N3  ( .A1(\SB1_0_30/i1_5 ), .A2(
        \SB1_0_30/i0[6] ), .A3(\SB1_0_30/i0[9] ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_30/Component_Function_1/N1  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i1[9] ), .ZN(\SB1_0_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_5/N4  ( .A1(\SB1_0_30/i0[9] ), .A2(
        \SB1_0_30/i0[6] ), .A3(\SB1_0_30/i0_4 ), .ZN(
        \SB1_0_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_5/N2  ( .A1(\SB1_0_30/i0_0 ), .A2(
        \SB1_0_30/i0[6] ), .A3(\SB1_0_30/i0[10] ), .ZN(
        \SB1_0_30/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_30/Component_Function_5/N1  ( .A1(\SB1_0_30/i0_0 ), .A2(
        \SB1_0_30/i3[0] ), .ZN(\SB1_0_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_0/N4  ( .A1(\SB1_0_31/i0[7] ), .A2(
        \SB1_0_31/i0_3 ), .A3(\SB1_0_31/i0_0 ), .ZN(
        \SB1_0_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_0/N2  ( .A1(\SB1_0_31/i0[8] ), .A2(
        \SB1_0_31/i0[7] ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_31/Component_Function_0/N1  ( .A1(\SB1_0_31/i0[10] ), .A2(
        \SB1_0_31/i0[9] ), .ZN(\SB1_0_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N4  ( .A1(\SB1_0_31/i1_7 ), .A2(
        \SB1_0_31/i0[8] ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N3  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[6] ), .A3(\SB1_0_31/i0[9] ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N2  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i1_7 ), .A3(\SB1_0_31/i0[8] ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_31/Component_Function_1/N1  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i1[9] ), .ZN(\SB1_0_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_5/N4  ( .A1(\SB1_0_31/i0[9] ), .A2(
        \SB1_0_31/i0[6] ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_5/N2  ( .A1(\SB1_0_31/i0_0 ), .A2(
        \SB1_0_31/i0[6] ), .A3(\SB1_0_31/i0[10] ), .ZN(
        \SB1_0_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_31/Component_Function_5/N1  ( .A1(\SB1_0_31/i0_0 ), .A2(
        \SB1_0_31/i3[0] ), .ZN(\SB1_0_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_0/N4  ( .A1(\SB2_0_0/i0[7] ), .A2(
        \SB2_0_0/i0_3 ), .A3(\SB2_0_0/i0_0 ), .ZN(
        \SB2_0_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_0/Component_Function_0/N3  ( .A1(\SB2_0_0/i0[10] ), .A2(
        \SB2_0_0/i0_4 ), .A3(\SB2_0_0/i0_3 ), .ZN(
        \SB2_0_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_0/Component_Function_0/N2  ( .A1(\SB2_0_0/i0[8] ), .A2(
        \SB2_0_0/i0[7] ), .A3(\SB2_0_0/i0[6] ), .ZN(
        \SB2_0_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_0/Component_Function_0/N1  ( .A1(\SB2_0_0/i0[10] ), .A2(
        \SB2_0_0/i0[9] ), .ZN(\SB2_0_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_1/N4  ( .A1(\SB2_0_0/i1_7 ), .A2(
        \SB2_0_0/i0[8] ), .A3(\SB2_0_0/i0_4 ), .ZN(
        \SB2_0_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_0/Component_Function_1/N3  ( .A1(\SB2_0_0/i1_5 ), .A2(
        \SB2_0_0/i0[6] ), .A3(\SB2_0_0/i0[9] ), .ZN(
        \SB2_0_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_0/Component_Function_1/N2  ( .A1(\SB2_0_0/i0_3 ), .A2(
        \SB2_0_0/i1_7 ), .A3(\SB2_0_0/i0[8] ), .ZN(
        \SB2_0_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_0/Component_Function_1/N1  ( .A1(\SB2_0_0/i0_3 ), .A2(
        \SB2_0_0/i1[9] ), .ZN(\SB2_0_0/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_0/Component_Function_5/N1  ( .A1(\SB2_0_0/i0_0 ), .A2(
        \SB2_0_0/i3[0] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_0/N4  ( .A1(\SB2_0_1/i0[7] ), .A2(
        \SB2_0_1/i0_3 ), .A3(\SB2_0_1/i0_0 ), .ZN(
        \SB2_0_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_1/Component_Function_0/N3  ( .A1(\SB2_0_1/i0[10] ), .A2(
        \SB2_0_1/i0_4 ), .A3(\SB2_0_1/i0_3 ), .ZN(
        \SB2_0_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_1/Component_Function_0/N2  ( .A1(\SB2_0_1/i0[8] ), .A2(
        \SB2_0_1/i0[7] ), .A3(\SB2_0_1/i0[6] ), .ZN(
        \SB2_0_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_1/Component_Function_0/N1  ( .A1(\SB2_0_1/i0[10] ), .A2(
        \SB2_0_1/i0[9] ), .ZN(\SB2_0_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_1/N4  ( .A1(\SB2_0_1/i1_7 ), .A2(
        \SB2_0_1/i0[8] ), .A3(\SB2_0_1/i0_4 ), .ZN(
        \SB2_0_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_1/Component_Function_1/N3  ( .A1(\SB2_0_1/i1_5 ), .A2(
        \SB2_0_1/i0[6] ), .A3(\SB2_0_1/i0[9] ), .ZN(
        \SB2_0_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_1/Component_Function_1/N2  ( .A1(\SB2_0_1/i0_3 ), .A2(
        \SB2_0_1/i1_7 ), .A3(\SB2_0_1/i0[8] ), .ZN(
        \SB2_0_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_1/Component_Function_1/N1  ( .A1(\SB2_0_1/i0_3 ), .A2(
        \SB2_0_1/i1[9] ), .ZN(\SB2_0_1/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_1/Component_Function_5/N1  ( .A1(\SB2_0_1/i0_0 ), .A2(
        \SB2_0_1/i3[0] ), .ZN(\SB2_0_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_0/N3  ( .A1(\SB2_0_2/i0[10] ), .A2(
        \SB2_0_2/i0_4 ), .A3(\SB2_0_2/i0_3 ), .ZN(
        \SB2_0_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_0/N2  ( .A1(\SB2_0_2/i0[8] ), .A2(
        \SB2_0_2/i0[7] ), .A3(\SB2_0_2/i0[6] ), .ZN(
        \SB2_0_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_2/Component_Function_0/N1  ( .A1(\SB2_0_2/i0[10] ), .A2(
        \SB2_0_2/i0[9] ), .ZN(\SB2_0_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_1/N4  ( .A1(\SB2_0_2/i1_7 ), .A2(
        \SB2_0_2/i0[8] ), .A3(\SB2_0_2/i0_4 ), .ZN(
        \SB2_0_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_2/Component_Function_1/N3  ( .A1(\SB2_0_2/i1_5 ), .A2(
        \SB2_0_2/i0[6] ), .A3(\SB2_0_2/i0[9] ), .ZN(
        \SB2_0_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_1/N2  ( .A1(\SB2_0_2/i0_3 ), .A2(
        \SB2_0_2/i1_7 ), .A3(\SB2_0_2/i0[8] ), .ZN(
        \SB2_0_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_2/Component_Function_1/N1  ( .A1(\SB2_0_2/i0_3 ), .A2(
        \SB2_0_2/i1[9] ), .ZN(\SB2_0_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_5/N4  ( .A1(\SB2_0_2/i0[9] ), .A2(
        \SB2_0_2/i0[6] ), .A3(\SB2_0_2/i0_4 ), .ZN(
        \SB2_0_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_2/Component_Function_5/N3  ( .A1(\SB2_0_2/i1[9] ), .A2(
        \SB2_0_2/i0_4 ), .A3(\SB2_0_2/i0_3 ), .ZN(
        \SB2_0_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_5/N2  ( .A1(\SB2_0_2/i0_0 ), .A2(
        \SB2_0_2/i0[6] ), .A3(\SB2_0_2/i0[10] ), .ZN(
        \SB2_0_2/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_3/Component_Function_0/N3  ( .A1(\SB2_0_3/i0[10] ), .A2(
        \SB2_0_3/i0_4 ), .A3(\SB2_0_3/i0_3 ), .ZN(
        \SB2_0_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_3/Component_Function_0/N2  ( .A1(\SB2_0_3/i0[8] ), .A2(
        \SB2_0_3/i0[7] ), .A3(\SB2_0_3/i0[6] ), .ZN(
        \SB2_0_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_3/Component_Function_0/N1  ( .A1(\SB2_0_3/i0[10] ), .A2(
        \SB2_0_3/i0[9] ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_1/N4  ( .A1(\SB2_0_3/i1_7 ), .A2(
        \SB2_0_3/i0[8] ), .A3(\SB2_0_3/i0_4 ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_3/Component_Function_1/N3  ( .A1(\SB2_0_3/i1_5 ), .A2(
        \SB2_0_3/i0[6] ), .A3(\SB2_0_3/i0[9] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_3/Component_Function_1/N2  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i1_7 ), .A3(\SB2_0_3/i0[8] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_3/Component_Function_1/N1  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i1[9] ), .ZN(\SB2_0_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_5/N3  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \SB2_0_3/i0_4 ), .A3(\SB2_0_3/i0_3 ), .ZN(
        \SB2_0_3/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_3/Component_Function_5/N1  ( .A1(\SB2_0_3/i0_0 ), .A2(
        \SB2_0_3/i3[0] ), .ZN(\SB2_0_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_0/N3  ( .A1(\SB2_0_4/i0[10] ), .A2(
        \SB2_0_4/i0_4 ), .A3(\SB2_0_4/i0_3 ), .ZN(
        \SB2_0_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_4/Component_Function_0/N2  ( .A1(\SB2_0_4/i0[8] ), .A2(
        \SB2_0_4/i0[7] ), .A3(\SB2_0_4/i0[6] ), .ZN(
        \SB2_0_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_4/Component_Function_0/N1  ( .A1(\SB2_0_4/i0[10] ), .A2(
        \SB2_0_4/i0[9] ), .ZN(\SB2_0_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_1/N3  ( .A1(\SB2_0_4/i1_5 ), .A2(
        \SB2_0_4/i0[6] ), .A3(\SB2_0_4/i0[9] ), .ZN(
        \SB2_0_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_4/Component_Function_1/N2  ( .A1(\SB2_0_4/i0_3 ), .A2(
        \SB2_0_4/i1_7 ), .A3(\SB2_0_4/i0[8] ), .ZN(
        \SB2_0_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_4/Component_Function_1/N1  ( .A1(\SB2_0_4/i0_3 ), .A2(
        \SB2_0_4/i1[9] ), .ZN(\SB2_0_4/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_4/Component_Function_5/N1  ( .A1(\SB2_0_4/i0_0 ), .A2(
        \SB2_0_4/i3[0] ), .ZN(\SB2_0_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_0/N4  ( .A1(\SB2_0_5/i0[7] ), .A2(
        \SB2_0_5/i0_3 ), .A3(\SB2_0_5/i0_0 ), .ZN(
        \SB2_0_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_5/Component_Function_0/N3  ( .A1(\SB2_0_5/i0[10] ), .A2(
        \SB2_0_5/i0_4 ), .A3(\SB2_0_5/i0_3 ), .ZN(
        \SB2_0_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_5/Component_Function_0/N2  ( .A1(\SB2_0_5/i0[8] ), .A2(
        \SB2_0_5/i0[7] ), .A3(\SB2_0_5/i0[6] ), .ZN(
        \SB2_0_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_5/Component_Function_0/N1  ( .A1(\SB2_0_5/i0[10] ), .A2(
        \SB2_0_5/i0[9] ), .ZN(\SB2_0_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_1/N4  ( .A1(\SB2_0_5/i1_7 ), .A2(
        \SB2_0_5/i0[8] ), .A3(\SB2_0_5/i0_4 ), .ZN(
        \SB2_0_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_5/Component_Function_1/N3  ( .A1(\SB2_0_5/i1_5 ), .A2(
        \SB2_0_5/i0[6] ), .A3(\SB2_0_5/i0[9] ), .ZN(
        \SB2_0_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_5/Component_Function_1/N2  ( .A1(\SB2_0_5/i0_3 ), .A2(
        \SB2_0_5/i1_7 ), .A3(\SB2_0_5/i0[8] ), .ZN(
        \SB2_0_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_5/Component_Function_1/N1  ( .A1(\SB2_0_5/i0_3 ), .A2(
        \SB2_0_5/i1[9] ), .ZN(\SB2_0_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_5/N2  ( .A1(\SB2_0_5/i0_0 ), .A2(
        \RI3[0][157] ), .A3(\SB2_0_5/i0[10] ), .ZN(
        \SB2_0_5/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_5/Component_Function_5/N1  ( .A1(\SB2_0_5/i0_0 ), .A2(
        \SB2_0_5/i3[0] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_0/N4  ( .A1(\SB2_0_6/i0[7] ), .A2(
        \SB2_0_6/i0_3 ), .A3(\SB2_0_6/i0_0 ), .ZN(
        \SB2_0_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_6/Component_Function_0/N3  ( .A1(\SB2_0_6/i0[10] ), .A2(
        \SB2_0_6/i0_4 ), .A3(\SB2_0_6/i0_3 ), .ZN(
        \SB2_0_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_6/Component_Function_0/N2  ( .A1(\SB2_0_6/i0[8] ), .A2(
        \SB2_0_6/i0[7] ), .A3(\SB2_0_6/i0[6] ), .ZN(
        \SB2_0_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_6/Component_Function_0/N1  ( .A1(\SB2_0_6/i0[10] ), .A2(
        \SB2_0_6/i0[9] ), .ZN(\SB2_0_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_1/N4  ( .A1(\SB2_0_6/i1_7 ), .A2(
        \SB2_0_6/i0[8] ), .A3(\SB2_0_6/i0_4 ), .ZN(
        \SB2_0_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_6/Component_Function_1/N3  ( .A1(\SB2_0_6/i1_5 ), .A2(
        \SB2_0_6/i0[6] ), .A3(\SB2_0_6/i0[9] ), .ZN(
        \SB2_0_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_6/Component_Function_1/N2  ( .A1(\SB2_0_6/i0_3 ), .A2(
        \SB2_0_6/i1_7 ), .A3(\SB2_0_6/i0[8] ), .ZN(
        \SB2_0_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_6/Component_Function_1/N1  ( .A1(\SB2_0_6/i0_3 ), .A2(
        \SB2_0_6/i1[9] ), .ZN(\SB2_0_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_5/N2  ( .A1(\SB2_0_6/i0_0 ), .A2(
        \SB2_0_6/i0[6] ), .A3(\SB2_0_6/i0[10] ), .ZN(
        \SB2_0_6/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_6/Component_Function_5/N1  ( .A1(\SB2_0_6/i0_0 ), .A2(
        \SB2_0_6/i3[0] ), .ZN(\SB2_0_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_0/N4  ( .A1(\SB2_0_7/i0[7] ), .A2(
        \SB2_0_7/i0_3 ), .A3(\SB2_0_7/i0_0 ), .ZN(
        \SB2_0_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_7/Component_Function_0/N3  ( .A1(\SB2_0_7/i0[10] ), .A2(
        \SB2_0_7/i0_4 ), .A3(\SB2_0_7/i0_3 ), .ZN(
        \SB2_0_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_0/N2  ( .A1(\SB2_0_7/i0[8] ), .A2(
        \SB2_0_7/i0[7] ), .A3(\SB2_0_7/i0[6] ), .ZN(
        \SB2_0_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_7/Component_Function_0/N1  ( .A1(\SB2_0_7/i0[10] ), .A2(
        \SB2_0_7/i0[9] ), .ZN(\SB2_0_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_1/N4  ( .A1(\SB2_0_7/i1_7 ), .A2(
        \SB2_0_7/i0[8] ), .A3(\SB2_0_7/i0_4 ), .ZN(
        \SB2_0_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_7/Component_Function_1/N3  ( .A1(\SB2_0_7/i1_5 ), .A2(
        \SB2_0_7/i0[6] ), .A3(\SB2_0_7/i0[9] ), .ZN(
        \SB2_0_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_1/N2  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i1_7 ), .A3(\SB2_0_7/i0[8] ), .ZN(
        \SB2_0_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_7/Component_Function_1/N1  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i1[9] ), .ZN(\SB2_0_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_5/N4  ( .A1(\SB2_0_7/i0[9] ), .A2(
        \SB2_0_7/i0[6] ), .A3(\RI3[0][148] ), .ZN(
        \SB2_0_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_7/Component_Function_5/N3  ( .A1(\SB2_0_7/i1[9] ), .A2(
        \SB2_0_7/i0_4 ), .A3(\SB2_0_7/i0_3 ), .ZN(
        \SB2_0_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_5/N2  ( .A1(\SB2_0_7/i0_0 ), .A2(
        \SB2_0_7/i0[6] ), .A3(\SB2_0_7/i0[10] ), .ZN(
        \SB2_0_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_8/Component_Function_0/N3  ( .A1(\SB2_0_8/i0[10] ), .A2(
        \SB2_0_8/i0_4 ), .A3(\SB2_0_8/i0_3 ), .ZN(
        \SB2_0_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_8/Component_Function_0/N2  ( .A1(\SB2_0_8/i0[8] ), .A2(
        \SB2_0_8/i0[7] ), .A3(\SB2_0_8/i0[6] ), .ZN(
        \SB2_0_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_8/Component_Function_0/N1  ( .A1(\SB2_0_8/i0[10] ), .A2(
        \SB2_0_8/i0[9] ), .ZN(\SB2_0_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_1/N4  ( .A1(\SB2_0_8/i1_7 ), .A2(
        \SB2_0_8/i0[8] ), .A3(\SB2_0_8/i0_4 ), .ZN(
        \SB2_0_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_8/Component_Function_1/N3  ( .A1(\SB2_0_8/i1_5 ), .A2(
        \SB2_0_8/i0[6] ), .A3(\SB2_0_8/i0[9] ), .ZN(
        \SB2_0_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_8/Component_Function_1/N2  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i1_7 ), .A3(\SB2_0_8/i0[8] ), .ZN(
        \SB2_0_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_8/Component_Function_1/N1  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i1[9] ), .ZN(\SB2_0_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_5/N4  ( .A1(\SB2_0_8/i0[9] ), .A2(
        \SB2_0_8/i0[6] ), .A3(\SB2_0_8/i0_4 ), .ZN(
        \SB2_0_8/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_8/Component_Function_5/N1  ( .A1(\SB2_0_8/i0_0 ), .A2(
        \SB2_0_8/i3[0] ), .ZN(\SB2_0_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_0/N4  ( .A1(\SB2_0_9/i0[7] ), .A2(
        \SB2_0_9/i0_3 ), .A3(\SB2_0_9/i0_0 ), .ZN(
        \SB2_0_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_9/Component_Function_0/N3  ( .A1(\SB2_0_9/i0[10] ), .A2(
        \SB2_0_9/i0_4 ), .A3(\SB2_0_9/i0_3 ), .ZN(
        \SB2_0_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_0/N2  ( .A1(\SB2_0_9/i0[8] ), .A2(
        \SB2_0_9/i0[7] ), .A3(\SB2_0_9/i0[6] ), .ZN(
        \SB2_0_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_9/Component_Function_0/N1  ( .A1(\SB2_0_9/i0[10] ), .A2(
        \SB2_0_9/i0[9] ), .ZN(\SB2_0_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N4  ( .A1(\SB2_0_9/i1_7 ), .A2(
        \SB2_0_9/i0[8] ), .A3(\SB2_0_9/i0_4 ), .ZN(
        \SB2_0_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N3  ( .A1(\SB2_0_9/i1_5 ), .A2(
        \SB2_0_9/i0[6] ), .A3(\SB2_0_9/i0[9] ), .ZN(
        \SB2_0_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N2  ( .A1(\SB2_0_9/i0_3 ), .A2(
        \SB2_0_9/i1_7 ), .A3(\SB2_0_9/i0[8] ), .ZN(
        \SB2_0_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_9/Component_Function_1/N1  ( .A1(\SB2_0_9/i0_3 ), .A2(
        \SB2_0_9/i1[9] ), .ZN(\SB2_0_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_5/N2  ( .A1(\SB2_0_9/i0_0 ), .A2(
        \SB2_0_9/i0[6] ), .A3(\SB2_0_9/i0[10] ), .ZN(
        \SB2_0_9/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_9/Component_Function_5/N1  ( .A1(\SB2_0_9/i0_0 ), .A2(
        \SB2_0_9/i3[0] ), .ZN(\SB2_0_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_0/N4  ( .A1(\SB2_0_10/i0[7] ), .A2(
        \SB2_0_10/i0_3 ), .A3(\SB2_0_10/i0_0 ), .ZN(
        \SB2_0_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_0/N3  ( .A1(\SB2_0_10/i0[10] ), .A2(
        \SB2_0_10/i0_4 ), .A3(\SB2_0_10/i0_3 ), .ZN(
        \SB2_0_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_10/Component_Function_0/N2  ( .A1(\SB2_0_10/i0[8] ), .A2(
        \SB2_0_10/i0[7] ), .A3(\SB2_0_10/i0[6] ), .ZN(
        \SB2_0_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_10/Component_Function_0/N1  ( .A1(\SB2_0_10/i0[10] ), .A2(
        \SB2_0_10/i0[9] ), .ZN(\SB2_0_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_1/N4  ( .A1(\SB2_0_10/i1_7 ), .A2(
        \SB2_0_10/i0[8] ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_1/N3  ( .A1(\SB2_0_10/i1_5 ), .A2(
        \SB2_0_10/i0[6] ), .A3(\SB2_0_10/i0[9] ), .ZN(
        \SB2_0_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_10/Component_Function_1/N2  ( .A1(\SB2_0_10/i0_3 ), .A2(
        \SB2_0_10/i1_7 ), .A3(\SB2_0_10/i0[8] ), .ZN(
        \SB2_0_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_10/Component_Function_1/N1  ( .A1(\SB2_0_10/i0_3 ), .A2(
        \SB2_0_10/i1[9] ), .ZN(\SB2_0_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_5/N4  ( .A1(\SB2_0_10/i0[9] ), .A2(
        \SB2_0_10/i0[6] ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_5/N3  ( .A1(\SB2_0_10/i1[9] ), .A2(
        \SB2_0_10/i0_4 ), .A3(\SB2_0_10/i0_3 ), .ZN(
        \SB2_0_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_0/N3  ( .A1(\SB2_0_11/i0[10] ), .A2(
        \SB2_0_11/i0_4 ), .A3(\SB2_0_11/i0_3 ), .ZN(
        \SB2_0_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_0/N2  ( .A1(\SB2_0_11/i0[8] ), .A2(
        \SB2_0_11/i0[7] ), .A3(\SB2_0_11/i0[6] ), .ZN(
        \SB2_0_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_11/Component_Function_0/N1  ( .A1(\SB2_0_11/i0[10] ), .A2(
        \SB2_0_11/i0[9] ), .ZN(\SB2_0_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_1/N4  ( .A1(\SB2_0_11/i1_7 ), .A2(
        \SB2_0_11/i0[8] ), .A3(\SB2_0_11/i0_4 ), .ZN(
        \SB2_0_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_1/N3  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \SB2_0_11/i0[6] ), .A3(\SB2_0_11/i0[9] ), .ZN(
        \SB2_0_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_1/N2  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i1_7 ), .A3(\SB2_0_11/i0[8] ), .ZN(
        \SB2_0_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_11/Component_Function_1/N1  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i1[9] ), .ZN(\SB2_0_11/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_11/Component_Function_5/N1  ( .A1(\SB2_0_11/i0_0 ), .A2(
        \SB2_0_11/i3[0] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N4  ( .A1(\SB2_0_12/i0[7] ), .A2(
        \SB2_0_12/i0_3 ), .A3(\SB2_0_12/i0_0 ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N3  ( .A1(\SB2_0_12/i0[10] ), .A2(
        \SB2_0_12/i0_4 ), .A3(\SB2_0_12/i0_3 ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N2  ( .A1(\SB2_0_12/i0[8] ), .A2(
        \SB2_0_12/i0[7] ), .A3(\SB2_0_12/i0[6] ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_12/Component_Function_0/N1  ( .A1(\SB2_0_12/i0[10] ), .A2(
        \SB2_0_12/i0[9] ), .ZN(\SB2_0_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N4  ( .A1(\SB2_0_12/i1_7 ), .A2(
        \SB2_0_12/i0[8] ), .A3(\SB2_0_12/i0_4 ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N3  ( .A1(\SB2_0_12/i1_5 ), .A2(
        \SB2_0_12/i0[6] ), .A3(\SB2_0_12/i0[9] ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N2  ( .A1(\SB2_0_12/i0_3 ), .A2(
        \SB2_0_12/i1_7 ), .A3(\SB2_0_12/i0[8] ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_12/Component_Function_1/N1  ( .A1(\SB2_0_12/i0_3 ), .A2(
        \SB2_0_12/i1[9] ), .ZN(\SB2_0_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_5/N4  ( .A1(\SB2_0_12/i0[9] ), .A2(
        \SB2_0_12/i0[6] ), .A3(\SB2_0_12/i0_4 ), .ZN(
        \SB2_0_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_5/N3  ( .A1(\SB2_0_12/i1[9] ), .A2(
        \SB2_0_12/i0_4 ), .A3(\SB2_0_12/i0_3 ), .ZN(
        \SB2_0_12/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_5/N2  ( .A1(\SB2_0_12/i0_0 ), .A2(
        \SB2_0_12/i0[6] ), .A3(\SB2_0_12/i0[10] ), .ZN(
        \SB2_0_12/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_12/Component_Function_5/N1  ( .A1(\SB2_0_12/i0_0 ), .A2(
        \SB2_0_12/i3[0] ), .ZN(\SB2_0_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_0/N4  ( .A1(\SB2_0_13/i0[7] ), .A2(
        \SB2_0_13/i0_3 ), .A3(\SB2_0_13/i0_0 ), .ZN(
        \SB2_0_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_13/Component_Function_0/N3  ( .A1(\SB2_0_13/i0[10] ), .A2(
        \SB2_0_13/i0_4 ), .A3(\SB2_0_13/i0_3 ), .ZN(
        \SB2_0_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_13/Component_Function_0/N2  ( .A1(\SB2_0_13/i0[8] ), .A2(
        \SB2_0_13/i0[7] ), .A3(\SB2_0_13/i0[6] ), .ZN(
        \SB2_0_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_13/Component_Function_0/N1  ( .A1(\SB2_0_13/i0[10] ), .A2(
        \SB2_0_13/i0[9] ), .ZN(\SB2_0_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_1/N4  ( .A1(\SB2_0_13/i1_7 ), .A2(
        \SB2_0_13/i0[8] ), .A3(\SB2_0_13/i0_4 ), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_13/Component_Function_1/N3  ( .A1(\SB2_0_13/i1_5 ), .A2(
        \SB2_0_13/i0[6] ), .A3(\SB2_0_13/i0[9] ), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_13/Component_Function_1/N2  ( .A1(\SB2_0_13/i0_3 ), .A2(
        \SB2_0_13/i1_7 ), .A3(\SB2_0_13/i0[8] ), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_13/Component_Function_1/N1  ( .A1(\SB2_0_13/i0_3 ), .A2(
        \SB2_0_13/i1[9] ), .ZN(\SB2_0_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_5/N4  ( .A1(\SB2_0_13/i0[9] ), .A2(
        \SB2_0_13/i0[6] ), .A3(\SB2_0_13/i0_4 ), .ZN(
        \SB2_0_13/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_13/Component_Function_5/N1  ( .A1(\SB2_0_13/i0_0 ), .A2(
        \SB2_0_13/i3[0] ), .ZN(\SB2_0_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_0/N4  ( .A1(\SB2_0_14/i0[7] ), .A2(
        \SB2_0_14/i0_3 ), .A3(\SB2_0_14/i0_0 ), .ZN(
        \SB2_0_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_0/N3  ( .A1(\SB2_0_14/i0[10] ), .A2(
        \SB2_0_14/i0_4 ), .A3(\SB2_0_14/i0_3 ), .ZN(
        \SB2_0_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_14/Component_Function_0/N2  ( .A1(\SB2_0_14/i0[8] ), .A2(
        \SB2_0_14/i0[7] ), .A3(\SB2_0_14/i0[6] ), .ZN(
        \SB2_0_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_14/Component_Function_0/N1  ( .A1(\SB2_0_14/i0[10] ), .A2(
        \SB2_0_14/i0[9] ), .ZN(\SB2_0_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_1/N4  ( .A1(\SB2_0_14/i1_7 ), .A2(
        \SB2_0_14/i0[8] ), .A3(\SB2_0_14/i0_4 ), .ZN(
        \SB2_0_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_1/N3  ( .A1(\SB2_0_14/i1_5 ), .A2(
        \SB2_0_14/i0[6] ), .A3(\SB2_0_14/i0[9] ), .ZN(
        \SB2_0_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_14/Component_Function_1/N2  ( .A1(\SB2_0_14/i0_3 ), .A2(
        \SB2_0_14/i1_7 ), .A3(\SB2_0_14/i0[8] ), .ZN(
        \SB2_0_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_14/Component_Function_1/N1  ( .A1(\SB2_0_14/i0_3 ), .A2(
        \SB2_0_14/i1[9] ), .ZN(\SB2_0_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_5/N4  ( .A1(\SB2_0_14/i0[9] ), .A2(
        \RI3[0][103] ), .A3(\SB2_0_14/i0_4 ), .ZN(
        \SB2_0_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_5/N2  ( .A1(\SB2_0_14/i0_0 ), .A2(
        \SB2_0_14/i0[6] ), .A3(\SB2_0_14/i0[10] ), .ZN(
        \SB2_0_14/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_14/Component_Function_5/N1  ( .A1(\SB2_0_14/i0_0 ), .A2(
        \SB2_0_14/i3[0] ), .ZN(\SB2_0_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_0/N3  ( .A1(\SB2_0_15/i0[10] ), .A2(
        \SB2_0_15/i0_4 ), .A3(\SB2_0_15/i0_3 ), .ZN(
        \SB2_0_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_15/Component_Function_0/N2  ( .A1(\SB2_0_15/i0[8] ), .A2(
        \SB2_0_15/i0[7] ), .A3(\SB2_0_15/i0[6] ), .ZN(
        \SB2_0_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_15/Component_Function_0/N1  ( .A1(\SB2_0_15/i0[10] ), .A2(
        \SB2_0_15/i0[9] ), .ZN(\SB2_0_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_1/N4  ( .A1(\SB2_0_15/i1_7 ), .A2(
        \SB2_0_15/i0[8] ), .A3(\SB2_0_15/i0_4 ), .ZN(
        \SB2_0_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_15/Component_Function_1/N3  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB2_0_15/i0[6] ), .A3(\SB2_0_15/i0[9] ), .ZN(
        \SB2_0_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_15/Component_Function_1/N2  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i1_7 ), .A3(\SB2_0_15/i0[8] ), .ZN(
        \SB2_0_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_15/Component_Function_1/N1  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i1[9] ), .ZN(\SB2_0_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_5/N4  ( .A1(\SB2_0_15/i0[9] ), .A2(
        \SB2_0_15/i0[6] ), .A3(\SB2_0_15/i0_4 ), .ZN(
        \SB2_0_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_15/Component_Function_5/N3  ( .A1(\SB2_0_15/i1[9] ), .A2(
        \SB2_0_15/i0_4 ), .A3(\SB2_0_15/i0_3 ), .ZN(
        \SB2_0_15/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_15/Component_Function_5/N2  ( .A1(\SB2_0_15/i0_0 ), .A2(
        \SB2_0_15/i0[6] ), .A3(\SB2_0_15/i0[10] ), .ZN(
        \SB2_0_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_15/Component_Function_5/N1  ( .A1(\SB2_0_15/i0_0 ), .A2(
        \SB2_0_15/i3[0] ), .ZN(\SB2_0_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_0/N3  ( .A1(\SB2_0_16/i0[10] ), .A2(
        \SB2_0_16/i0_4 ), .A3(\SB2_0_16/i0_3 ), .ZN(
        \SB2_0_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_16/Component_Function_0/N2  ( .A1(\SB2_0_16/i0[8] ), .A2(
        \SB2_0_16/i0[7] ), .A3(\SB2_0_16/i0[6] ), .ZN(
        \SB2_0_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_16/Component_Function_0/N1  ( .A1(\SB2_0_16/i0[10] ), .A2(
        \SB2_0_16/i0[9] ), .ZN(\SB2_0_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_1/N4  ( .A1(\SB2_0_16/i1_7 ), .A2(
        \SB2_0_16/i0[8] ), .A3(\SB2_0_16/i0_4 ), .ZN(
        \SB2_0_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_1/N3  ( .A1(\SB2_0_16/i1_5 ), .A2(
        \SB2_0_16/i0[6] ), .A3(\SB2_0_16/i0[9] ), .ZN(
        \SB2_0_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_16/Component_Function_1/N2  ( .A1(\SB2_0_16/i0_3 ), .A2(
        \SB2_0_16/i1_7 ), .A3(\SB2_0_16/i0[8] ), .ZN(
        \SB2_0_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_16/Component_Function_1/N1  ( .A1(\SB2_0_16/i0_3 ), .A2(
        \SB2_0_16/i1[9] ), .ZN(\SB2_0_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_5/N4  ( .A1(\SB2_0_16/i0[9] ), .A2(
        \SB2_0_16/i0[6] ), .A3(\SB2_0_16/i0_4 ), .ZN(
        \SB2_0_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_5/N2  ( .A1(\SB2_0_16/i0_0 ), .A2(
        \SB2_0_16/i0[6] ), .A3(\SB2_0_16/i0[10] ), .ZN(
        \SB2_0_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_16/Component_Function_5/N1  ( .A1(\SB2_0_16/i0_0 ), .A2(
        \SB2_0_16/i3[0] ), .ZN(\SB2_0_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_0/N4  ( .A1(\SB2_0_17/i0[7] ), .A2(
        \SB2_0_17/i0_3 ), .A3(\SB2_0_17/i0_0 ), .ZN(
        \SB2_0_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_0/N3  ( .A1(\SB2_0_17/i0[10] ), .A2(
        \SB2_0_17/i0_4 ), .A3(\SB2_0_17/i0_3 ), .ZN(
        \SB2_0_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_17/Component_Function_0/N2  ( .A1(\SB2_0_17/i0[8] ), .A2(
        \SB2_0_17/i0[7] ), .A3(\SB2_0_17/i0[6] ), .ZN(
        \SB2_0_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_17/Component_Function_0/N1  ( .A1(\SB2_0_17/i0[10] ), .A2(
        \SB2_0_17/i0[9] ), .ZN(\SB2_0_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_1/N4  ( .A1(\SB2_0_17/i1_7 ), .A2(
        \SB2_0_17/i0[8] ), .A3(\SB2_0_17/i0_4 ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_1/N3  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0[6] ), .A3(\SB2_0_17/i0[9] ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_17/Component_Function_1/N2  ( .A1(\SB2_0_17/i0_3 ), .A2(
        \SB2_0_17/i1_7 ), .A3(\SB2_0_17/i0[8] ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_17/Component_Function_1/N1  ( .A1(\SB2_0_17/i0_3 ), .A2(
        \SB2_0_17/i1[9] ), .ZN(\SB2_0_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_5/N3  ( .A1(\SB2_0_17/i1[9] ), .A2(
        \SB2_0_17/i0_4 ), .A3(\SB2_0_17/i0_3 ), .ZN(
        \SB2_0_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_17/Component_Function_5/N2  ( .A1(\SB2_0_17/i0_0 ), .A2(
        \SB2_0_17/i0[6] ), .A3(\SB2_0_17/i0[10] ), .ZN(
        \SB2_0_17/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_17/Component_Function_5/N1  ( .A1(\SB2_0_17/i0_0 ), .A2(
        \SB2_0_17/i3[0] ), .ZN(\SB2_0_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_18/Component_Function_0/N4  ( .A1(\SB2_0_18/i0[7] ), .A2(
        \SB2_0_18/i0_3 ), .A3(\SB2_0_18/i0_0 ), .ZN(
        \SB2_0_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_18/Component_Function_0/N3  ( .A1(\SB2_0_18/i0[10] ), .A2(
        \SB2_0_18/i0_4 ), .A3(\SB2_0_18/i0_3 ), .ZN(
        \SB2_0_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_18/Component_Function_0/N2  ( .A1(\SB2_0_18/i0[8] ), .A2(
        \SB2_0_18/i0[7] ), .A3(\SB2_0_18/i0[6] ), .ZN(
        \SB2_0_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_18/Component_Function_0/N1  ( .A1(\SB2_0_18/i0[10] ), .A2(
        \SB2_0_18/i0[9] ), .ZN(\SB2_0_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_18/Component_Function_1/N4  ( .A1(\SB2_0_18/i1_7 ), .A2(
        \SB2_0_18/i0[8] ), .A3(\SB2_0_18/i0_4 ), .ZN(
        \SB2_0_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_18/Component_Function_1/N3  ( .A1(\SB2_0_18/i1_5 ), .A2(
        \SB2_0_18/i0[6] ), .A3(\SB2_0_18/i0[9] ), .ZN(
        \SB2_0_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_18/Component_Function_1/N2  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i1_7 ), .A3(\SB2_0_18/i0[8] ), .ZN(
        \SB2_0_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_18/Component_Function_1/N1  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i1[9] ), .ZN(\SB2_0_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_18/Component_Function_5/N2  ( .A1(\SB2_0_18/i0_0 ), .A2(
        \RI3[0][79] ), .A3(\SB2_0_18/i0[10] ), .ZN(
        \SB2_0_18/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_18/Component_Function_5/N1  ( .A1(\SB2_0_18/i0_0 ), .A2(
        \SB2_0_18/i3[0] ), .ZN(\SB2_0_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_0/N4  ( .A1(\SB2_0_19/i0[7] ), .A2(
        \SB2_0_19/i0_3 ), .A3(\SB2_0_19/i0_0 ), .ZN(
        \SB2_0_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_19/Component_Function_0/N3  ( .A1(\SB2_0_19/i0[10] ), .A2(
        \SB2_0_19/i0_4 ), .A3(\SB2_0_19/i0_3 ), .ZN(
        \SB2_0_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_19/Component_Function_0/N2  ( .A1(\SB2_0_19/i0[8] ), .A2(
        \SB2_0_19/i0[7] ), .A3(\SB2_0_19/i0[6] ), .ZN(
        \SB2_0_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_19/Component_Function_0/N1  ( .A1(\SB2_0_19/i0[10] ), .A2(
        \SB2_0_19/i0[9] ), .ZN(\SB2_0_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_1/N4  ( .A1(\SB2_0_19/i1_7 ), .A2(
        \SB2_0_19/i0[8] ), .A3(\SB2_0_19/i0_4 ), .ZN(
        \SB2_0_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_19/Component_Function_1/N3  ( .A1(\SB2_0_19/i1_5 ), .A2(
        \SB2_0_19/i0[6] ), .A3(\SB2_0_19/i0[9] ), .ZN(
        \SB2_0_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_19/Component_Function_1/N2  ( .A1(\SB2_0_19/i0_3 ), .A2(
        \SB2_0_19/i1_7 ), .A3(\SB2_0_19/i0[8] ), .ZN(
        \SB2_0_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_19/Component_Function_1/N1  ( .A1(\SB2_0_19/i0_3 ), .A2(
        \SB2_0_19/i1[9] ), .ZN(\SB2_0_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_5/N4  ( .A1(\SB2_0_19/i0[9] ), .A2(
        \SB2_0_19/i0[6] ), .A3(\SB2_0_19/i0_4 ), .ZN(
        \SB2_0_19/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_19/Component_Function_5/N1  ( .A1(\SB2_0_19/i0_0 ), .A2(
        \SB2_0_19/i3[0] ), .ZN(\SB2_0_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_20/Component_Function_0/N3  ( .A1(\SB2_0_20/i0[10] ), .A2(
        \SB2_0_20/i0_4 ), .A3(\SB2_0_20/i0_3 ), .ZN(
        \SB2_0_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_20/Component_Function_0/N2  ( .A1(\SB2_0_20/i0[8] ), .A2(
        \SB2_0_20/i0[7] ), .A3(\SB2_0_20/i0[6] ), .ZN(
        \SB2_0_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_20/Component_Function_0/N1  ( .A1(\SB2_0_20/i0[10] ), .A2(
        \SB2_0_20/i0[9] ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_20/Component_Function_1/N4  ( .A1(\SB2_0_20/i1_7 ), .A2(
        \SB2_0_20/i0[8] ), .A3(\SB2_0_20/i0_4 ), .ZN(
        \SB2_0_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_20/Component_Function_1/N3  ( .A1(\SB2_0_20/i1_5 ), .A2(
        \SB2_0_20/i0[6] ), .A3(\SB2_0_20/i0[9] ), .ZN(
        \SB2_0_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_20/Component_Function_1/N2  ( .A1(\SB2_0_20/i0_3 ), .A2(
        \SB2_0_20/i1_7 ), .A3(\SB2_0_20/i0[8] ), .ZN(
        \SB2_0_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_20/Component_Function_1/N1  ( .A1(\SB2_0_20/i0_3 ), .A2(
        \SB2_0_20/i1[9] ), .ZN(\SB2_0_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_20/Component_Function_5/N2  ( .A1(\SB2_0_20/i0_0 ), .A2(
        \SB2_0_20/i0[6] ), .A3(\SB2_0_20/i0[10] ), .ZN(
        \SB2_0_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_21/Component_Function_0/N3  ( .A1(\SB2_0_21/i0[10] ), .A2(
        \SB2_0_21/i0_4 ), .A3(\SB2_0_21/i0_3 ), .ZN(
        \SB2_0_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_21/Component_Function_0/N2  ( .A1(\SB2_0_21/i0[8] ), .A2(
        \SB2_0_21/i0[7] ), .A3(\SB2_0_21/i0[6] ), .ZN(
        \SB2_0_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_21/Component_Function_0/N1  ( .A1(\SB2_0_21/i0[10] ), .A2(
        \SB2_0_21/i0[9] ), .ZN(\SB2_0_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_21/Component_Function_1/N4  ( .A1(\SB2_0_21/i1_7 ), .A2(
        \SB2_0_21/i0[8] ), .A3(\SB2_0_21/i0_4 ), .ZN(
        \SB2_0_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_21/Component_Function_1/N3  ( .A1(\SB2_0_21/i1_5 ), .A2(
        \SB2_0_21/i0[6] ), .A3(\SB2_0_21/i0[9] ), .ZN(
        \SB2_0_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_21/Component_Function_1/N2  ( .A1(\SB2_0_21/i0_3 ), .A2(
        \SB2_0_21/i1_7 ), .A3(\SB2_0_21/i0[8] ), .ZN(
        \SB2_0_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_21/Component_Function_1/N1  ( .A1(\SB2_0_21/i0_3 ), .A2(
        \SB2_0_21/i1[9] ), .ZN(\SB2_0_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_21/Component_Function_5/N4  ( .A1(\SB2_0_21/i0[9] ), .A2(
        \SB2_0_21/i0[6] ), .A3(\SB2_0_21/i0_4 ), .ZN(
        \SB2_0_21/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_21/Component_Function_5/N1  ( .A1(\SB2_0_21/i0_0 ), .A2(
        \SB2_0_21/i3[0] ), .ZN(\SB2_0_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_22/Component_Function_0/N4  ( .A1(\SB2_0_22/i0[7] ), .A2(
        \SB2_0_22/i0_3 ), .A3(\SB2_0_22/i0_0 ), .ZN(
        \SB2_0_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_22/Component_Function_0/N3  ( .A1(\SB2_0_22/i0[10] ), .A2(
        \SB2_0_22/i0_4 ), .A3(\SB2_0_22/i0_3 ), .ZN(
        \SB2_0_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_22/Component_Function_0/N2  ( .A1(\SB2_0_22/i0[8] ), .A2(
        \SB2_0_22/i0[7] ), .A3(\SB2_0_22/i0[6] ), .ZN(
        \SB2_0_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_22/Component_Function_0/N1  ( .A1(\SB2_0_22/i0[10] ), .A2(
        \SB2_0_22/i0[9] ), .ZN(\SB2_0_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_22/Component_Function_1/N4  ( .A1(\SB2_0_22/i1_7 ), .A2(
        \SB2_0_22/i0[8] ), .A3(\SB2_0_22/i0_4 ), .ZN(
        \SB2_0_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_22/Component_Function_1/N3  ( .A1(\SB2_0_22/i1_5 ), .A2(
        \SB2_0_22/i0[6] ), .A3(\SB2_0_22/i0[9] ), .ZN(
        \SB2_0_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_22/Component_Function_1/N2  ( .A1(\SB2_0_22/i0_3 ), .A2(
        \SB2_0_22/i1_7 ), .A3(\SB2_0_22/i0[8] ), .ZN(
        \SB2_0_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_22/Component_Function_1/N1  ( .A1(\SB2_0_22/i0_3 ), .A2(
        \SB2_0_22/i1[9] ), .ZN(\SB2_0_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_22/Component_Function_5/N3  ( .A1(\SB2_0_22/i1[9] ), .A2(
        \SB2_0_22/i0_4 ), .A3(\SB2_0_22/i0_3 ), .ZN(
        \SB2_0_22/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_22/Component_Function_5/N2  ( .A1(\SB2_0_22/i0_0 ), .A2(
        \SB2_0_22/i0[6] ), .A3(\SB2_0_22/i0[10] ), .ZN(
        \SB2_0_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_22/Component_Function_5/N1  ( .A1(\SB2_0_22/i0_0 ), .A2(
        \SB2_0_22/i3[0] ), .ZN(\SB2_0_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_0/N4  ( .A1(\SB2_0_23/i0[7] ), .A2(
        \SB2_0_23/i0_3 ), .A3(\SB2_0_23/i0_0 ), .ZN(
        \SB2_0_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_23/Component_Function_0/N2  ( .A1(\SB2_0_23/i0[8] ), .A2(
        \SB2_0_23/i0[7] ), .A3(\SB2_0_23/i0[6] ), .ZN(
        \SB2_0_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_23/Component_Function_1/N4  ( .A1(\SB2_0_23/i1_7 ), .A2(
        \SB2_0_23/i0[8] ), .A3(\SB2_0_23/i0_4 ), .ZN(
        \SB2_0_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_23/Component_Function_1/N3  ( .A1(\SB2_0_23/i1_5 ), .A2(
        \SB2_0_23/i0[6] ), .A3(\SB2_0_23/i0[9] ), .ZN(
        \SB2_0_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_23/Component_Function_1/N2  ( .A1(\SB2_0_23/i0_3 ), .A2(
        \SB2_0_23/i1_7 ), .A3(\SB2_0_23/i0[8] ), .ZN(
        \SB2_0_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_23/Component_Function_1/N1  ( .A1(\SB2_0_23/i0_3 ), .A2(
        \SB2_0_23/i1[9] ), .ZN(\SB2_0_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_5/N4  ( .A1(\RI3[0][48] ), .A2(
        \RI3[0][49] ), .A3(\SB2_0_23/i0_4 ), .ZN(
        \SB2_0_23/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_23/Component_Function_5/N1  ( .A1(\SB2_0_23/i0_0 ), .A2(
        \SB2_0_23/i3[0] ), .ZN(\SB2_0_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_0/N4  ( .A1(\SB2_0_24/i0[7] ), .A2(
        \SB2_0_24/i0_3 ), .A3(\SB2_0_24/i0_0 ), .ZN(
        \SB2_0_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_24/Component_Function_0/N3  ( .A1(\SB2_0_24/i0[10] ), .A2(
        \SB2_0_24/i0_4 ), .A3(\SB2_0_24/i0_3 ), .ZN(
        \SB2_0_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_0/N2  ( .A1(\SB2_0_24/i0[8] ), .A2(
        \SB2_0_24/i0[7] ), .A3(\SB2_0_24/i0[6] ), .ZN(
        \SB2_0_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_24/Component_Function_0/N1  ( .A1(\SB2_0_24/i0[10] ), .A2(
        \SB2_0_24/i0[9] ), .ZN(\SB2_0_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N4  ( .A1(\SB2_0_24/i1_7 ), .A2(
        \SB2_0_24/i0[8] ), .A3(\SB2_0_24/i0_4 ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N3  ( .A1(\SB2_0_24/i1_5 ), .A2(
        \SB2_0_24/i0[6] ), .A3(\SB2_0_24/i0[9] ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N2  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i1_7 ), .A3(\SB2_0_24/i0[8] ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_24/Component_Function_1/N1  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i1[9] ), .ZN(\SB2_0_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_5/N2  ( .A1(\SB2_0_24/i0_0 ), .A2(
        \SB2_0_24/i0[6] ), .A3(\SB2_0_24/i0[10] ), .ZN(
        \SB2_0_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_24/Component_Function_5/N1  ( .A1(\SB2_0_24/i0_0 ), .A2(
        \SB2_0_24/i3[0] ), .ZN(\SB2_0_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_0/N3  ( .A1(\SB2_0_25/i0[10] ), .A2(
        \SB2_0_25/i0_4 ), .A3(\SB2_0_25/i0_3 ), .ZN(
        \SB2_0_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_25/Component_Function_0/N2  ( .A1(\SB2_0_25/i0[8] ), .A2(
        \SB2_0_25/i0[7] ), .A3(\SB2_0_25/i0[6] ), .ZN(
        \SB2_0_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_25/Component_Function_0/N1  ( .A1(\SB2_0_25/i0[10] ), .A2(
        \SB2_0_25/i0[9] ), .ZN(\SB2_0_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_1/N4  ( .A1(\SB2_0_25/i1_7 ), .A2(
        \SB2_0_25/i0[8] ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_25/Component_Function_1/N3  ( .A1(\SB2_0_25/i1_5 ), .A2(
        \SB2_0_25/i0[6] ), .A3(\SB2_0_25/i0[9] ), .ZN(
        \SB2_0_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_25/Component_Function_1/N2  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i1_7 ), .A3(\SB2_0_25/i0[8] ), .ZN(
        \SB2_0_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_25/Component_Function_1/N1  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i1[9] ), .ZN(\SB2_0_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_5/N4  ( .A1(\SB2_0_25/i0[9] ), .A2(
        \SB2_0_25/i0[6] ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_25/Component_Function_5/N1  ( .A1(\SB2_0_25/i0_0 ), .A2(
        \SB2_0_25/i3[0] ), .ZN(\SB2_0_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_0/N3  ( .A1(\SB2_0_26/i0[10] ), .A2(
        \SB2_0_26/i0_4 ), .A3(\SB2_0_26/i0_3 ), .ZN(
        \SB2_0_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_26/Component_Function_0/N2  ( .A1(\SB2_0_26/i0[8] ), .A2(
        \SB2_0_26/i0[7] ), .A3(\SB2_0_26/i0[6] ), .ZN(
        \SB2_0_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_26/Component_Function_0/N1  ( .A1(\SB2_0_26/i0[10] ), .A2(
        n2132), .ZN(\SB2_0_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_1/N4  ( .A1(\SB2_0_26/i1_7 ), .A2(
        \SB2_0_26/i0[8] ), .A3(\SB2_0_26/i0_4 ), .ZN(
        \SB2_0_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_26/Component_Function_1/N3  ( .A1(\SB2_0_26/i1_5 ), .A2(
        \SB2_0_26/i0[6] ), .A3(n2132), .ZN(
        \SB2_0_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_26/Component_Function_1/N2  ( .A1(\SB2_0_26/i0_3 ), .A2(
        \SB2_0_26/i1_7 ), .A3(\SB2_0_26/i0[8] ), .ZN(
        \SB2_0_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_26/Component_Function_1/N1  ( .A1(\SB2_0_26/i0_3 ), .A2(
        \SB2_0_26/i1[9] ), .ZN(\SB2_0_26/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_26/Component_Function_5/N1  ( .A1(\SB2_0_26/i0_0 ), .A2(
        \SB2_0_26/i3[0] ), .ZN(\SB2_0_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_0/N3  ( .A1(\SB2_0_27/i0[10] ), .A2(
        \SB2_0_27/i0_4 ), .A3(\SB2_0_27/i0_3 ), .ZN(
        \SB2_0_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_27/Component_Function_0/N2  ( .A1(\SB2_0_27/i0[8] ), .A2(
        \SB2_0_27/i0[7] ), .A3(\SB2_0_27/i0[6] ), .ZN(
        \SB2_0_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_27/Component_Function_0/N1  ( .A1(\SB2_0_27/i0[10] ), .A2(
        \SB2_0_27/i0[9] ), .ZN(\SB2_0_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_1/N4  ( .A1(\SB2_0_27/i1_7 ), .A2(
        \SB2_0_27/i0[8] ), .A3(\SB2_0_27/i0_4 ), .ZN(
        \SB2_0_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_27/Component_Function_1/N3  ( .A1(\SB2_0_27/i1_5 ), .A2(
        \SB2_0_27/i0[6] ), .A3(\SB2_0_27/i0[9] ), .ZN(
        \SB2_0_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_27/Component_Function_1/N2  ( .A1(\SB2_0_27/i0_3 ), .A2(
        \SB2_0_27/i1_7 ), .A3(\SB2_0_27/i0[8] ), .ZN(
        \SB2_0_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_27/Component_Function_1/N1  ( .A1(\SB2_0_27/i0_3 ), .A2(
        \SB2_0_27/i1[9] ), .ZN(\SB2_0_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_5/N4  ( .A1(\SB2_0_27/i0[9] ), .A2(
        \SB2_0_27/i0[6] ), .A3(\SB2_0_27/i0_4 ), .ZN(
        \SB2_0_27/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_27/Component_Function_5/N1  ( .A1(\SB2_0_27/i0_0 ), .A2(
        \SB2_0_27/i3[0] ), .ZN(\SB2_0_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_0/N4  ( .A1(\SB2_0_28/i0[7] ), .A2(
        \SB2_0_28/i0_3 ), .A3(\SB2_0_28/i0_0 ), .ZN(
        \SB2_0_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_28/Component_Function_0/N3  ( .A1(\SB2_0_28/i0[10] ), .A2(
        \SB2_0_28/i0_4 ), .A3(\SB2_0_28/i0_3 ), .ZN(
        \SB2_0_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_28/Component_Function_0/N2  ( .A1(\SB2_0_28/i0[8] ), .A2(
        \SB2_0_28/i0[7] ), .A3(\SB2_0_28/i0[6] ), .ZN(
        \SB2_0_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_28/Component_Function_0/N1  ( .A1(\SB2_0_28/i0[10] ), .A2(
        \SB2_0_28/i0[9] ), .ZN(\SB2_0_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_1/N4  ( .A1(\SB2_0_28/i1_7 ), .A2(
        \SB2_0_28/i0[8] ), .A3(\SB2_0_28/i0_4 ), .ZN(
        \SB2_0_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_28/Component_Function_1/N3  ( .A1(\SB2_0_28/i1_5 ), .A2(
        \SB2_0_28/i0[6] ), .A3(\SB2_0_28/i0[9] ), .ZN(
        \SB2_0_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_28/Component_Function_1/N2  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i1_7 ), .A3(\SB2_0_28/i0[8] ), .ZN(
        \SB2_0_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_28/Component_Function_1/N1  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i1[9] ), .ZN(\SB2_0_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_5/N2  ( .A1(\SB2_0_28/i0_0 ), .A2(
        \SB2_0_28/i0[6] ), .A3(\SB2_0_28/i0[10] ), .ZN(
        \SB2_0_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_28/Component_Function_5/N1  ( .A1(\SB2_0_28/i0_0 ), .A2(
        \SB2_0_28/i3[0] ), .ZN(\SB2_0_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_0/N4  ( .A1(\SB2_0_29/i0[7] ), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0_0 ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_0/N3  ( .A1(\SB2_0_29/i0[10] ), .A2(
        \SB2_0_29/i0_4 ), .A3(\SB2_0_29/i0_3 ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_0/N2  ( .A1(\SB2_0_29/i0[8] ), .A2(
        \SB2_0_29/i0[7] ), .A3(\SB2_0_29/i0[6] ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_29/Component_Function_0/N1  ( .A1(\SB2_0_29/i0[10] ), .A2(
        \SB2_0_29/i0[9] ), .ZN(\SB2_0_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_1/N4  ( .A1(\SB2_0_29/i1_7 ), .A2(
        \SB2_0_29/i0[8] ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_1/N3  ( .A1(\SB2_0_29/i1_5 ), .A2(
        \SB2_0_29/i0[6] ), .A3(\SB2_0_29/i0[9] ), .ZN(
        \SB2_0_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_1/N2  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i1_7 ), .A3(\SB2_0_29/i0[8] ), .ZN(
        \SB2_0_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_29/Component_Function_1/N1  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i1[9] ), .ZN(\SB2_0_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_5/N4  ( .A1(\SB2_0_29/i0[9] ), .A2(
        \SB2_0_29/i0[6] ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_5/N3  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i0_4 ), .A3(\SB2_0_29/i0_3 ), .ZN(
        \SB2_0_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_5/N2  ( .A1(\SB2_0_29/i0_0 ), .A2(
        \SB2_0_29/i0[6] ), .A3(\SB2_0_29/i0[10] ), .ZN(
        \SB2_0_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_30/Component_Function_0/N3  ( .A1(\SB2_0_30/i0[10] ), .A2(
        \SB2_0_30/i0_4 ), .A3(\SB2_0_30/i0_3 ), .ZN(
        \SB2_0_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_30/Component_Function_0/N2  ( .A1(\SB2_0_30/i0[8] ), .A2(
        \SB2_0_30/i0[7] ), .A3(\SB2_0_30/i0[6] ), .ZN(
        \SB2_0_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_30/Component_Function_0/N1  ( .A1(\SB2_0_30/i0[10] ), .A2(
        \SB2_0_30/i0[9] ), .ZN(\SB2_0_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_1/N4  ( .A1(\SB2_0_30/i1_7 ), .A2(
        \SB2_0_30/i0[8] ), .A3(\SB2_0_30/i0_4 ), .ZN(
        \SB2_0_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_30/Component_Function_1/N3  ( .A1(\SB2_0_30/i1_5 ), .A2(
        \SB2_0_30/i0[6] ), .A3(\SB2_0_30/i0[9] ), .ZN(
        \SB2_0_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_30/Component_Function_1/N2  ( .A1(\SB2_0_30/i0_3 ), .A2(
        \SB2_0_30/i1_7 ), .A3(\SB2_0_30/i0[8] ), .ZN(
        \SB2_0_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_30/Component_Function_1/N1  ( .A1(\SB2_0_30/i0_3 ), .A2(
        \SB2_0_30/i1[9] ), .ZN(\SB2_0_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_0/N3  ( .A1(\SB2_0_31/i0[10] ), .A2(
        \SB2_0_31/i0_4 ), .A3(\SB2_0_31/i0_3 ), .ZN(
        \SB2_0_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_0/N2  ( .A1(\SB2_0_31/i0[8] ), .A2(
        \SB2_0_31/i0[7] ), .A3(\SB2_0_31/i0[6] ), .ZN(
        \SB2_0_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_31/Component_Function_0/N1  ( .A1(\SB2_0_31/i0[10] ), .A2(
        \SB2_0_31/i0[9] ), .ZN(\SB2_0_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N4  ( .A1(\SB2_0_31/i1_7 ), .A2(
        \SB2_0_31/i0[8] ), .A3(\SB2_0_31/i0_4 ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N3  ( .A1(\SB2_0_31/i1_5 ), .A2(
        \SB2_0_31/i0[6] ), .A3(\SB2_0_31/i0[9] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N2  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i1_7 ), .A3(\SB2_0_31/i0[8] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_31/Component_Function_1/N1  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i1[9] ), .ZN(\SB2_0_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_5/N4  ( .A1(\SB2_0_31/i0[9] ), .A2(
        \SB2_0_31/i0[6] ), .A3(\SB2_0_31/i0_4 ), .ZN(
        \SB2_0_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_5/N3  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i0_4 ), .A3(\SB2_0_31/i1[9] ), .ZN(
        \SB2_0_31/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_31/Component_Function_5/N1  ( .A1(\SB2_0_31/i0_0 ), .A2(
        \SB2_0_31/i3[0] ), .ZN(\SB2_0_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_0/N4  ( .A1(\SB1_1_0/i0[7] ), .A2(
        \SB1_1_0/i0_3 ), .A3(\SB1_1_0/i0_0 ), .ZN(
        \SB1_1_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_0/Component_Function_0/N3  ( .A1(\SB1_1_0/i0[10] ), .A2(
        \SB1_1_0/i0_4 ), .A3(\SB1_1_0/i0_3 ), .ZN(
        \SB1_1_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_0/Component_Function_0/N2  ( .A1(\SB1_1_0/i0[8] ), .A2(
        \SB1_1_0/i0[7] ), .A3(\SB1_1_0/i0[6] ), .ZN(
        \SB1_1_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_0/Component_Function_0/N1  ( .A1(\SB1_1_0/i0[10] ), .A2(
        \SB1_1_0/i0[9] ), .ZN(\SB1_1_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_1/N4  ( .A1(\SB1_1_0/i1_7 ), .A2(
        \SB1_1_0/i0[8] ), .A3(\SB1_1_0/i0_4 ), .ZN(
        \SB1_1_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_0/Component_Function_1/N3  ( .A1(\SB1_1_0/i1_5 ), .A2(
        \SB1_1_0/i0[6] ), .A3(\SB1_1_0/i0[9] ), .ZN(
        \SB1_1_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_0/Component_Function_1/N2  ( .A1(\SB1_1_0/i0_3 ), .A2(
        \SB1_1_0/i1_7 ), .A3(\SB1_1_0/i0[8] ), .ZN(
        \SB1_1_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_0/Component_Function_1/N1  ( .A1(\SB1_1_0/i0_3 ), .A2(
        \SB1_1_0/i1[9] ), .ZN(\SB1_1_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_5/N4  ( .A1(\SB1_1_0/i0[9] ), .A2(
        \SB1_1_0/i0[6] ), .A3(\SB1_1_0/i0_4 ), .ZN(
        \SB1_1_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_0/Component_Function_5/N2  ( .A1(\SB1_1_0/i0_0 ), .A2(
        \SB1_1_0/i0[6] ), .A3(\SB1_1_0/i0[10] ), .ZN(
        \SB1_1_0/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_0/Component_Function_5/N1  ( .A1(\SB1_1_0/i0_0 ), .A2(
        \SB1_1_0/i3[0] ), .ZN(\SB1_1_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_0/N3  ( .A1(\SB1_1_1/i0[10] ), .A2(
        \SB1_1_1/i0_4 ), .A3(\SB1_1_1/i0_3 ), .ZN(
        \SB1_1_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_1/Component_Function_0/N2  ( .A1(\SB1_1_1/i0[8] ), .A2(
        \SB1_1_1/i0[7] ), .A3(\SB1_1_1/i0[6] ), .ZN(
        \SB1_1_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_1/Component_Function_0/N1  ( .A1(\SB1_1_1/i0[10] ), .A2(
        \SB1_1_1/i0[9] ), .ZN(\SB1_1_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_1/N4  ( .A1(\SB1_1_1/i1_7 ), .A2(
        \SB1_1_1/i0[8] ), .A3(\SB1_1_1/i0_4 ), .ZN(
        \SB1_1_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_1/Component_Function_1/N3  ( .A1(\SB1_1_1/i1_5 ), .A2(
        \SB1_1_1/i0[6] ), .A3(\SB1_1_1/i0[9] ), .ZN(
        \SB1_1_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_1/Component_Function_1/N2  ( .A1(\SB1_1_1/i0_3 ), .A2(
        \SB1_1_1/i1_7 ), .A3(\SB1_1_1/i0[8] ), .ZN(
        \SB1_1_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_1/Component_Function_1/N1  ( .A1(\SB1_1_1/i0_3 ), .A2(
        \SB1_1_1/i1[9] ), .ZN(\SB1_1_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_5/N4  ( .A1(\SB1_1_1/i0[9] ), .A2(
        \SB1_1_1/i0[6] ), .A3(\SB1_1_1/i0_4 ), .ZN(
        \SB1_1_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_1/Component_Function_5/N2  ( .A1(\SB1_1_1/i0_0 ), .A2(
        \SB1_1_1/i0[6] ), .A3(\SB1_1_1/i0[10] ), .ZN(
        \SB1_1_1/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_1/Component_Function_5/N1  ( .A1(\SB1_1_1/i0_0 ), .A2(
        \SB1_1_1/i3[0] ), .ZN(\SB1_1_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_0/N4  ( .A1(\SB1_1_2/i0[7] ), .A2(
        \SB1_1_2/i0_3 ), .A3(\SB1_1_2/i0_0 ), .ZN(
        \SB1_1_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_2/Component_Function_0/N3  ( .A1(\SB1_1_2/i0[10] ), .A2(
        \SB1_1_2/i0_4 ), .A3(\SB1_1_2/i0_3 ), .ZN(
        \SB1_1_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_2/Component_Function_0/N2  ( .A1(\SB1_1_2/i0[8] ), .A2(
        \SB1_1_2/i0[7] ), .A3(\SB1_1_2/i0[6] ), .ZN(
        \SB1_1_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_2/Component_Function_0/N1  ( .A1(\SB1_1_2/i0[10] ), .A2(
        \SB1_1_2/i0[9] ), .ZN(\SB1_1_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_1/N3  ( .A1(\SB1_1_2/i1_5 ), .A2(
        \SB1_1_2/i0[6] ), .A3(\SB1_1_2/i0[9] ), .ZN(
        \SB1_1_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_2/Component_Function_1/N2  ( .A1(\SB1_1_2/i0_3 ), .A2(
        \SB1_1_2/i1_7 ), .A3(\SB1_1_2/i0[8] ), .ZN(
        \SB1_1_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_2/Component_Function_1/N1  ( .A1(\SB1_1_2/i0_3 ), .A2(
        \SB1_1_2/i1[9] ), .ZN(\SB1_1_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_5/N2  ( .A1(\SB1_1_2/i0_0 ), .A2(
        \SB1_1_2/i0[6] ), .A3(\SB1_1_2/i0[10] ), .ZN(
        \SB1_1_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_2/Component_Function_5/N1  ( .A1(\SB1_1_2/i0_0 ), .A2(
        \SB1_1_2/i3[0] ), .ZN(\SB1_1_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_0/N4  ( .A1(\SB1_1_3/i0[7] ), .A2(
        \SB1_1_3/i0_3 ), .A3(\SB1_1_3/i0_0 ), .ZN(
        \SB1_1_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_3/Component_Function_0/N2  ( .A1(\SB1_1_3/i0[8] ), .A2(
        \SB1_1_3/i0[7] ), .A3(\SB1_1_3/i0[6] ), .ZN(
        \SB1_1_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_3/Component_Function_0/N1  ( .A1(\SB1_1_3/i0[10] ), .A2(
        \SB1_1_3/i0[9] ), .ZN(\SB1_1_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_1/N4  ( .A1(\SB1_1_3/i1_7 ), .A2(
        \SB1_1_3/i0[8] ), .A3(\SB1_1_3/i0_4 ), .ZN(
        \SB1_1_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_3/Component_Function_1/N3  ( .A1(\SB1_1_3/i1_5 ), .A2(
        \SB1_1_3/i0[6] ), .A3(\SB1_1_3/i0[9] ), .ZN(
        \SB1_1_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_3/Component_Function_1/N2  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i1_7 ), .A3(\SB1_1_3/i0[8] ), .ZN(
        \SB1_1_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_3/Component_Function_1/N1  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i1[9] ), .ZN(\SB1_1_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_5/N2  ( .A1(\SB1_1_3/i0_0 ), .A2(
        \SB1_1_3/i0[6] ), .A3(\SB1_1_3/i0[10] ), .ZN(
        \SB1_1_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_3/Component_Function_5/N1  ( .A1(\SB1_1_3/i0_0 ), .A2(
        \SB1_1_3/i3[0] ), .ZN(\SB1_1_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_0/N3  ( .A1(\SB1_1_4/i0[10] ), .A2(
        \SB1_1_4/i0_4 ), .A3(\SB1_1_4/i0_3 ), .ZN(
        \SB1_1_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_4/Component_Function_0/N2  ( .A1(\SB1_1_4/i0[8] ), .A2(
        \SB1_1_4/i0[7] ), .A3(\SB1_1_4/i0[6] ), .ZN(
        \SB1_1_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_4/Component_Function_0/N1  ( .A1(\SB1_1_4/i0[10] ), .A2(
        \SB1_1_4/i0[9] ), .ZN(\SB1_1_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_1/N3  ( .A1(\SB1_1_4/i1_5 ), .A2(
        \SB1_1_4/i0[6] ), .A3(\SB1_1_4/i0[9] ), .ZN(
        \SB1_1_4/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_4/Component_Function_1/N1  ( .A1(n2149), .A2(\SB1_1_4/i1[9] ), .ZN(\SB1_1_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_5/N4  ( .A1(\SB1_1_4/i0[9] ), .A2(
        \SB1_1_4/i0[6] ), .A3(\SB1_1_4/i0_4 ), .ZN(
        \SB1_1_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_4/Component_Function_5/N2  ( .A1(\SB1_1_4/i0_0 ), .A2(
        \SB1_1_4/i0[6] ), .A3(\SB1_1_4/i0[10] ), .ZN(
        \SB1_1_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_4/Component_Function_5/N1  ( .A1(\SB1_1_4/i0_0 ), .A2(
        \SB1_1_4/i3[0] ), .ZN(\SB1_1_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N4  ( .A1(\SB1_1_5/i0[7] ), .A2(
        \SB1_1_5/i0_3 ), .A3(\SB1_1_5/i0_0 ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N3  ( .A1(\SB1_1_5/i0[10] ), .A2(
        \SB1_1_5/i0_4 ), .A3(\SB1_1_5/i0_3 ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N2  ( .A1(\SB1_1_5/i0[8] ), .A2(
        \SB1_1_5/i0[7] ), .A3(\SB1_1_5/i0[6] ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_5/Component_Function_0/N1  ( .A1(\SB1_1_5/i0[10] ), .A2(
        \SB1_1_5/i0[9] ), .ZN(\SB1_1_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_1/N4  ( .A1(\SB1_1_5/i1_7 ), .A2(
        \SB1_1_5/i0[8] ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_1/N3  ( .A1(\SB1_1_5/i1_5 ), .A2(
        \SB1_1_5/i0[6] ), .A3(\SB1_1_5/i0[9] ), .ZN(
        \SB1_1_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_5/Component_Function_1/N2  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i1_7 ), .A3(\SB1_1_5/i0[8] ), .ZN(
        \SB1_1_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_5/Component_Function_1/N1  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i1[9] ), .ZN(\SB1_1_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_5/N4  ( .A1(\SB1_1_5/i0[9] ), .A2(
        \SB1_1_5/i0[6] ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_5/N2  ( .A1(\SB1_1_5/i0_0 ), .A2(
        \SB1_1_5/i0[6] ), .A3(\SB1_1_5/i0[10] ), .ZN(
        \SB1_1_5/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_5/Component_Function_5/N1  ( .A1(\SB1_1_5/i0_0 ), .A2(
        \SB1_1_5/i3[0] ), .ZN(\SB1_1_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_0/N2  ( .A1(\SB1_1_6/i0[8] ), .A2(
        \SB1_1_6/i0[7] ), .A3(\SB1_1_6/i0[6] ), .ZN(
        \SB1_1_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_6/Component_Function_0/N1  ( .A1(\SB1_1_6/i0[10] ), .A2(
        \SB1_1_6/i0[9] ), .ZN(\SB1_1_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_1/N4  ( .A1(\SB1_1_6/i1_7 ), .A2(
        \SB1_1_6/i0[8] ), .A3(\SB1_1_6/i0_4 ), .ZN(
        \SB1_1_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_6/Component_Function_1/N3  ( .A1(\SB1_1_6/i1_5 ), .A2(
        \SB1_1_6/i0[6] ), .A3(\SB1_1_6/i0[9] ), .ZN(
        \SB1_1_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_6/Component_Function_1/N2  ( .A1(\SB1_1_6/i0_3 ), .A2(
        \SB1_1_6/i1_7 ), .A3(\SB1_1_6/i0[8] ), .ZN(
        \SB1_1_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_6/Component_Function_1/N1  ( .A1(\SB1_1_6/i0_3 ), .A2(
        \SB1_1_6/i1[9] ), .ZN(\SB1_1_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_5/N4  ( .A1(\SB1_1_6/i0[9] ), .A2(
        \SB1_1_6/i0[6] ), .A3(\SB1_1_6/i0_4 ), .ZN(
        \SB1_1_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_6/Component_Function_5/N2  ( .A1(\SB1_1_6/i0_0 ), .A2(
        \SB1_1_6/i0[6] ), .A3(\SB1_1_6/i0[10] ), .ZN(
        \SB1_1_6/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_6/Component_Function_5/N1  ( .A1(\SB1_1_6/i0_0 ), .A2(
        \SB1_1_6/i3[0] ), .ZN(\SB1_1_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_0/N4  ( .A1(\SB1_1_7/i0[7] ), .A2(
        \SB1_1_7/i0_3 ), .A3(\SB1_1_7/i0_0 ), .ZN(
        \SB1_1_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_7/Component_Function_0/N2  ( .A1(\SB1_1_7/i0[8] ), .A2(
        \SB1_1_7/i0[7] ), .A3(\SB1_1_7/i0[6] ), .ZN(
        \SB1_1_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_7/Component_Function_0/N1  ( .A1(\SB1_1_7/i0[10] ), .A2(
        \SB1_1_7/i0[9] ), .ZN(\SB1_1_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_1/N4  ( .A1(\SB1_1_7/i1_7 ), .A2(
        \SB1_1_7/i0[8] ), .A3(\SB1_1_7/i0_4 ), .ZN(
        \SB1_1_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_7/Component_Function_1/N3  ( .A1(\SB1_1_7/i1_5 ), .A2(
        \SB1_1_7/i0[6] ), .A3(\SB1_1_7/i0[9] ), .ZN(
        \SB1_1_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_7/Component_Function_1/N2  ( .A1(\SB1_1_7/i0_3 ), .A2(
        \SB1_1_7/i1_7 ), .A3(\SB1_1_7/i0[8] ), .ZN(
        \SB1_1_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_7/Component_Function_1/N1  ( .A1(\SB1_1_7/i0_3 ), .A2(
        \SB1_1_7/i1[9] ), .ZN(\SB1_1_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_5/N4  ( .A1(\SB1_1_7/i0[9] ), .A2(
        \SB1_1_7/i0[6] ), .A3(\SB1_1_7/i0_4 ), .ZN(
        \SB1_1_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_7/Component_Function_5/N2  ( .A1(\SB1_1_7/i0_0 ), .A2(
        \SB1_1_7/i0[6] ), .A3(\SB1_1_7/i0[10] ), .ZN(
        \SB1_1_7/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_7/Component_Function_5/N1  ( .A1(\SB1_1_7/i0_0 ), .A2(
        \SB1_1_7/i3[0] ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_8/Component_Function_0/N4  ( .A1(\SB1_1_8/i0[7] ), .A2(
        \SB1_1_8/i0_3 ), .A3(\SB1_1_8/i0_0 ), .ZN(
        \SB1_1_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_8/Component_Function_0/N3  ( .A1(\SB1_1_8/i0[10] ), .A2(
        \SB1_1_8/i0_4 ), .A3(\SB1_1_8/i0_3 ), .ZN(
        \SB1_1_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_8/Component_Function_0/N2  ( .A1(\SB1_1_8/i0[8] ), .A2(
        \SB1_1_8/i0[7] ), .A3(\SB1_1_8/i0[6] ), .ZN(
        \SB1_1_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_8/Component_Function_0/N1  ( .A1(\SB1_1_8/i0[10] ), .A2(
        \SB1_1_8/i0[9] ), .ZN(\SB1_1_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_8/Component_Function_1/N3  ( .A1(\SB1_1_8/i1_5 ), .A2(
        \SB1_1_8/i0[6] ), .A3(\SB1_1_8/i0[9] ), .ZN(
        \SB1_1_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_8/Component_Function_1/N2  ( .A1(\SB1_1_8/i0_3 ), .A2(
        \SB1_1_8/i1_7 ), .A3(\SB1_1_8/i0[8] ), .ZN(
        \SB1_1_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_8/Component_Function_1/N1  ( .A1(\SB1_1_8/i0_3 ), .A2(
        \SB1_1_8/i1[9] ), .ZN(\SB1_1_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_8/Component_Function_5/N4  ( .A1(\SB1_1_8/i0[9] ), .A2(
        \SB1_1_8/i0[6] ), .A3(\SB1_1_8/i0_4 ), .ZN(
        \SB1_1_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_8/Component_Function_5/N2  ( .A1(\SB1_1_8/i0_0 ), .A2(
        \SB1_1_8/i0[6] ), .A3(\SB1_1_8/i0[10] ), .ZN(
        \SB1_1_8/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_8/Component_Function_5/N1  ( .A1(\SB1_1_8/i0_0 ), .A2(
        \SB1_1_8/i3[0] ), .ZN(\SB1_1_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_0/N2  ( .A1(\SB1_1_9/i0[8] ), .A2(
        \SB1_1_9/i0[7] ), .A3(\SB1_1_9/i0[6] ), .ZN(
        \SB1_1_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_9/Component_Function_0/N1  ( .A1(\SB1_1_9/i0[10] ), .A2(
        \SB1_1_9/i0[9] ), .ZN(\SB1_1_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_1/N4  ( .A1(\SB1_1_9/i1_7 ), .A2(
        \SB1_1_9/i0[8] ), .A3(\SB1_1_9/i0_4 ), .ZN(
        \SB1_1_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_9/Component_Function_1/N2  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i1_7 ), .A3(\SB1_1_9/i0[8] ), .ZN(
        \SB1_1_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_9/Component_Function_1/N1  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i1[9] ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_5/N3  ( .A1(\SB1_1_9/i1[9] ), .A2(
        \SB1_1_9/i0_4 ), .A3(\SB1_1_9/i0_3 ), .ZN(
        \SB1_1_9/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_9/Component_Function_5/N1  ( .A1(\SB1_1_9/i0_0 ), .A2(
        \SB1_1_9/i3[0] ), .ZN(\SB1_1_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_0/N4  ( .A1(\SB1_1_10/i0[7] ), .A2(
        n826), .A3(\SB1_1_10/i0_0 ), .ZN(
        \SB1_1_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_0/N2  ( .A1(\SB1_1_10/i0[8] ), .A2(
        \SB1_1_10/i0[7] ), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_10/Component_Function_0/N1  ( .A1(\SB1_1_10/i0[10] ), .A2(
        \SB1_1_10/i0[9] ), .ZN(\SB1_1_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N4  ( .A1(\SB1_1_10/i1_7 ), .A2(
        \SB1_1_10/i0[8] ), .A3(\SB1_1_10/i0_4 ), .ZN(
        \SB1_1_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N3  ( .A1(\SB1_1_10/i1_5 ), .A2(
        \SB1_1_10/i0[6] ), .A3(\SB1_1_10/i0[9] ), .ZN(
        \SB1_1_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N2  ( .A1(n826), .A2(\SB1_1_10/i1_7 ), .A3(\SB1_1_10/i0[8] ), .ZN(\SB1_1_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_10/Component_Function_1/N1  ( .A1(n826), .A2(
        \SB1_1_10/i1[9] ), .ZN(\SB1_1_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_5/N4  ( .A1(\SB1_1_10/i0[9] ), .A2(
        \SB1_1_10/i0[6] ), .A3(\SB1_1_10/i0_4 ), .ZN(
        \SB1_1_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_5/N2  ( .A1(\SB1_1_10/i0_0 ), .A2(
        \SB1_1_10/i0[6] ), .A3(\SB1_1_10/i0[10] ), .ZN(
        \SB1_1_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_10/Component_Function_5/N1  ( .A1(\SB1_1_10/i0_0 ), .A2(
        \SB1_1_10/i3[0] ), .ZN(\SB1_1_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_0/N2  ( .A1(\SB1_1_11/i0[8] ), .A2(
        \SB1_1_11/i0[7] ), .A3(\SB1_1_11/i0[6] ), .ZN(
        \SB1_1_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_11/Component_Function_0/N1  ( .A1(\SB1_1_11/i0[10] ), .A2(
        \SB1_1_11/i0[9] ), .ZN(\SB1_1_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_1/N2  ( .A1(\SB1_1_11/i0_3 ), .A2(
        \SB1_1_11/i1_7 ), .A3(\SB1_1_11/i0[8] ), .ZN(
        \SB1_1_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_11/Component_Function_1/N1  ( .A1(n2141), .A2(
        \SB1_1_11/i1[9] ), .ZN(\SB1_1_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_5/N4  ( .A1(\SB1_1_11/i0[9] ), .A2(
        \SB1_1_11/i0[6] ), .A3(\SB1_1_11/i0_4 ), .ZN(
        \SB1_1_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_11/Component_Function_5/N2  ( .A1(\SB1_1_11/i0_0 ), .A2(
        \SB1_1_11/i0[6] ), .A3(\SB1_1_11/i0[10] ), .ZN(
        \SB1_1_11/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_11/Component_Function_5/N1  ( .A1(\SB1_1_11/i0_0 ), .A2(
        \SB1_1_11/i3[0] ), .ZN(\SB1_1_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_0/N4  ( .A1(\SB1_1_12/i0[7] ), .A2(
        \SB1_1_12/i0_3 ), .A3(\SB1_1_12/i0_0 ), .ZN(
        \SB1_1_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_12/Component_Function_0/N2  ( .A1(\SB1_1_12/i0[8] ), .A2(
        \SB1_1_12/i0[7] ), .A3(\SB1_1_12/i0[6] ), .ZN(
        \SB1_1_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_12/Component_Function_0/N1  ( .A1(\SB1_1_12/i0[10] ), .A2(
        \SB1_1_12/i0[9] ), .ZN(\SB1_1_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_1/N3  ( .A1(\SB1_1_12/i1_5 ), .A2(
        \SB1_1_12/i0[6] ), .A3(\SB1_1_12/i0[9] ), .ZN(
        \SB1_1_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_12/Component_Function_1/N2  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i1_7 ), .A3(\SB1_1_12/i0[8] ), .ZN(
        \SB1_1_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_12/Component_Function_1/N1  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i1[9] ), .ZN(\SB1_1_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_5/N4  ( .A1(\SB1_1_12/i0[9] ), .A2(
        \SB1_1_12/i0[6] ), .A3(\SB1_1_12/i0_4 ), .ZN(
        \SB1_1_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_12/Component_Function_5/N2  ( .A1(\SB1_1_12/i0_0 ), .A2(
        \SB1_1_12/i0[6] ), .A3(\SB1_1_12/i0[10] ), .ZN(
        \SB1_1_12/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_12/Component_Function_5/N1  ( .A1(\SB1_1_12/i0_0 ), .A2(
        \SB1_1_12/i3[0] ), .ZN(\SB1_1_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N4  ( .A1(\SB1_1_13/i0[7] ), .A2(
        \SB1_1_13/i0_3 ), .A3(\SB1_1_13/i0_0 ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N2  ( .A1(\SB1_1_13/i0[8] ), .A2(
        \SB1_1_13/i0[7] ), .A3(\SB1_1_13/i0[6] ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_13/Component_Function_0/N1  ( .A1(\SB1_1_13/i0[10] ), .A2(
        \SB1_1_13/i0[9] ), .ZN(\SB1_1_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_1/N4  ( .A1(\SB1_1_13/i1_7 ), .A2(
        \SB1_1_13/i0[8] ), .A3(\SB1_1_13/i0_4 ), .ZN(
        \SB1_1_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_13/Component_Function_1/N3  ( .A1(\SB1_1_13/i1_5 ), .A2(
        \SB1_1_13/i0[6] ), .A3(\SB1_1_13/i0[9] ), .ZN(
        \SB1_1_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_13/Component_Function_1/N2  ( .A1(\SB1_1_13/i0_3 ), .A2(
        \SB1_1_13/i1_7 ), .A3(\SB1_1_13/i0[8] ), .ZN(
        \SB1_1_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_13/Component_Function_1/N1  ( .A1(\SB1_1_13/i0_3 ), .A2(
        \SB1_1_13/i1[9] ), .ZN(\SB1_1_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_5/N4  ( .A1(\SB1_1_13/i0[9] ), .A2(
        \SB1_1_13/i0[6] ), .A3(\SB1_1_13/i0_4 ), .ZN(
        \SB1_1_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_13/Component_Function_5/N2  ( .A1(\SB1_1_13/i0_0 ), .A2(
        \SB1_1_13/i0[6] ), .A3(\SB1_1_13/i0[10] ), .ZN(
        \SB1_1_13/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_13/Component_Function_5/N1  ( .A1(\SB1_1_13/i0_0 ), .A2(
        \SB1_1_13/i3[0] ), .ZN(\SB1_1_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_0/N2  ( .A1(\SB1_1_14/i0[8] ), .A2(
        \SB1_1_14/i0[7] ), .A3(\SB1_1_14/i0[6] ), .ZN(
        \SB1_1_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_14/Component_Function_0/N1  ( .A1(\SB1_1_14/i0[10] ), .A2(
        \SB1_1_14/i0[9] ), .ZN(\SB1_1_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_1/N4  ( .A1(\SB1_1_14/i1_7 ), .A2(
        \SB1_1_14/i0[8] ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_14/Component_Function_1/N3  ( .A1(\SB1_1_14/i1_5 ), .A2(
        \SB1_1_14/i0[6] ), .A3(\SB1_1_14/i0[9] ), .ZN(
        \SB1_1_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_14/Component_Function_1/N2  ( .A1(\SB1_1_14/i0_3 ), .A2(
        \SB1_1_14/i1_7 ), .A3(\SB1_1_14/i0[8] ), .ZN(
        \SB1_1_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_14/Component_Function_1/N1  ( .A1(\SB1_1_14/i0_3 ), .A2(
        \SB1_1_14/i1[9] ), .ZN(\SB1_1_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_5/N4  ( .A1(\SB1_1_14/i0[9] ), .A2(
        \SB1_1_14/i0[6] ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_14/Component_Function_5/N2  ( .A1(\SB1_1_14/i0_0 ), .A2(
        \SB1_1_14/i0[6] ), .A3(\SB1_1_14/i0[10] ), .ZN(
        \SB1_1_14/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_14/Component_Function_5/N1  ( .A1(\SB1_1_14/i0_0 ), .A2(
        \SB1_1_14/i3[0] ), .ZN(\SB1_1_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_0/N4  ( .A1(\SB1_1_15/i0[7] ), .A2(
        \SB1_1_15/i0_3 ), .A3(\SB1_1_15/i0_0 ), .ZN(
        \SB1_1_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_15/Component_Function_0/N2  ( .A1(\SB1_1_15/i0[8] ), .A2(
        \SB1_1_15/i0[7] ), .A3(\SB1_1_15/i0[6] ), .ZN(
        \SB1_1_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_15/Component_Function_0/N1  ( .A1(\SB1_1_15/i0[10] ), .A2(
        \SB1_1_15/i0[9] ), .ZN(\SB1_1_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_1/N4  ( .A1(\SB1_1_15/i1_7 ), .A2(
        \SB1_1_15/i0[8] ), .A3(\SB1_1_15/i0_4 ), .ZN(
        \SB1_1_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_15/Component_Function_1/N3  ( .A1(\SB1_1_15/i1_5 ), .A2(
        \SB1_1_15/i0[6] ), .A3(\SB1_1_15/i0[9] ), .ZN(
        \SB1_1_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_15/Component_Function_1/N2  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i1_7 ), .A3(\SB1_1_15/i0[8] ), .ZN(
        \SB1_1_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_15/Component_Function_1/N1  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i1[9] ), .ZN(\SB1_1_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_5/N4  ( .A1(\SB1_1_15/i0[9] ), .A2(
        \SB1_1_15/i0[6] ), .A3(\SB1_1_15/i0_4 ), .ZN(
        \SB1_1_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_15/Component_Function_5/N2  ( .A1(\SB1_1_15/i0_0 ), .A2(
        \SB1_1_15/i0[6] ), .A3(\SB1_1_15/i0[10] ), .ZN(
        \SB1_1_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_15/Component_Function_5/N1  ( .A1(\SB1_1_15/i0_0 ), .A2(
        \SB1_1_15/i3[0] ), .ZN(\SB1_1_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_0/N4  ( .A1(\SB1_1_16/i0[7] ), .A2(
        \SB1_1_16/i0_3 ), .A3(\SB1_1_16/i0_0 ), .ZN(
        \SB1_1_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_16/Component_Function_0/N3  ( .A1(\SB1_1_16/i0[10] ), .A2(
        \SB1_1_16/i0_4 ), .A3(\SB1_1_16/i0_3 ), .ZN(
        \SB1_1_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_16/Component_Function_0/N2  ( .A1(\SB1_1_16/i0[8] ), .A2(
        \SB1_1_16/i0[7] ), .A3(\SB1_1_16/i0[6] ), .ZN(
        \SB1_1_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_16/Component_Function_0/N1  ( .A1(\SB1_1_16/i0[10] ), .A2(
        \SB1_1_16/i0[9] ), .ZN(\SB1_1_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_1/N4  ( .A1(\SB1_1_16/i1_7 ), .A2(
        \SB1_1_16/i0[8] ), .A3(\SB1_1_16/i0_4 ), .ZN(
        \SB1_1_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_16/Component_Function_1/N3  ( .A1(\SB1_1_16/i1_5 ), .A2(
        \SB1_1_16/i0[6] ), .A3(\SB1_1_16/i0[9] ), .ZN(
        \SB1_1_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_16/Component_Function_1/N2  ( .A1(\SB1_1_16/i0_3 ), .A2(
        \SB1_1_16/i1_7 ), .A3(\SB1_1_16/i0[8] ), .ZN(
        \SB1_1_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_16/Component_Function_1/N1  ( .A1(\SB1_1_16/i0_3 ), .A2(
        \SB1_1_16/i1[9] ), .ZN(\SB1_1_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_5/N3  ( .A1(\SB1_1_16/i1[9] ), .A2(
        \SB1_1_16/i0_4 ), .A3(\SB1_1_16/i0_3 ), .ZN(
        \SB1_1_16/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_16/Component_Function_5/N1  ( .A1(\SB1_1_16/i0_0 ), .A2(
        \SB1_1_16/i3[0] ), .ZN(\SB1_1_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_0/N4  ( .A1(\SB1_1_17/i0[7] ), .A2(
        n789), .A3(\SB1_1_17/i0_0 ), .ZN(
        \SB1_1_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_17/Component_Function_0/N3  ( .A1(\SB1_1_17/i0[10] ), .A2(
        \SB1_1_17/i0_4 ), .A3(n789), .ZN(
        \SB1_1_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_17/Component_Function_0/N2  ( .A1(\SB1_1_17/i0[8] ), .A2(
        \SB1_1_17/i0[7] ), .A3(\SB1_1_17/i0[6] ), .ZN(
        \SB1_1_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_17/Component_Function_0/N1  ( .A1(\SB1_1_17/i0[10] ), .A2(
        \SB1_1_17/i0[9] ), .ZN(\SB1_1_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_1/N4  ( .A1(\SB1_1_17/i1_7 ), .A2(
        \SB1_1_17/i0[8] ), .A3(\SB1_1_17/i0_4 ), .ZN(
        \SB1_1_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_17/Component_Function_1/N3  ( .A1(\SB1_1_17/i1_5 ), .A2(
        \SB1_1_17/i0[6] ), .A3(\SB1_1_17/i0[9] ), .ZN(
        \SB1_1_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_17/Component_Function_1/N2  ( .A1(n789), .A2(\SB1_1_17/i1_7 ), .A3(\SB1_1_17/i0[8] ), .ZN(\SB1_1_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_17/Component_Function_1/N1  ( .A1(n789), .A2(
        \SB1_1_17/i1[9] ), .ZN(\SB1_1_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_5/N4  ( .A1(\SB1_1_17/i0[9] ), .A2(
        \SB1_1_17/i0[6] ), .A3(\SB1_1_17/i0_4 ), .ZN(
        \SB1_1_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_17/Component_Function_5/N2  ( .A1(\SB1_1_17/i0_0 ), .A2(
        \SB1_1_17/i0[6] ), .A3(\SB1_1_17/i0[10] ), .ZN(
        \SB1_1_17/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_17/Component_Function_5/N1  ( .A1(\SB1_1_17/i0_0 ), .A2(
        \SB1_1_17/i3[0] ), .ZN(\SB1_1_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_0/N4  ( .A1(\SB1_1_18/i0[7] ), .A2(
        \SB1_1_18/i0_3 ), .A3(\SB1_1_18/i0_0 ), .ZN(
        \SB1_1_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_18/Component_Function_0/N2  ( .A1(\SB1_1_18/i0[8] ), .A2(
        \SB1_1_18/i0[7] ), .A3(\SB1_1_18/i0[6] ), .ZN(
        \SB1_1_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_18/Component_Function_0/N1  ( .A1(\SB1_1_18/i0[10] ), .A2(
        \SB1_1_18/i0[9] ), .ZN(\SB1_1_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_1/N4  ( .A1(\SB1_1_18/i1_7 ), .A2(
        \SB1_1_18/i0[8] ), .A3(\SB1_1_18/i0_4 ), .ZN(
        \SB1_1_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_18/Component_Function_1/N3  ( .A1(\SB1_1_18/i1_5 ), .A2(
        \SB1_1_18/i0[6] ), .A3(\SB1_1_18/i0[9] ), .ZN(
        \SB1_1_18/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_18/Component_Function_1/N1  ( .A1(\SB1_1_18/i0_3 ), .A2(
        \SB1_1_18/i1[9] ), .ZN(\SB1_1_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_5/N4  ( .A1(\SB1_1_18/i0[9] ), .A2(
        \SB1_1_18/i0[6] ), .A3(\SB1_1_18/i0_4 ), .ZN(
        \SB1_1_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_18/Component_Function_5/N2  ( .A1(\SB1_1_18/i0_0 ), .A2(
        \SB1_1_18/i0[6] ), .A3(\SB1_1_18/i0[10] ), .ZN(
        \SB1_1_18/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_18/Component_Function_5/N1  ( .A1(\SB1_1_18/i0_0 ), .A2(
        \SB1_1_18/i3[0] ), .ZN(\SB1_1_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_0/N4  ( .A1(\SB1_1_19/i0[7] ), .A2(
        \SB1_1_19/i0_3 ), .A3(\SB1_1_19/i0_0 ), .ZN(
        \SB1_1_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_0/N3  ( .A1(\SB1_1_19/i0[10] ), .A2(
        \SB1_1_19/i0_4 ), .A3(\SB1_1_19/i0_3 ), .ZN(
        \SB1_1_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_19/Component_Function_0/N2  ( .A1(\SB1_1_19/i0[8] ), .A2(
        \SB1_1_19/i0[7] ), .A3(\SB1_1_19/i0[6] ), .ZN(
        \SB1_1_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_19/Component_Function_0/N1  ( .A1(\SB1_1_19/i0[10] ), .A2(
        \SB1_1_19/i0[9] ), .ZN(\SB1_1_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_1/N4  ( .A1(\SB1_1_19/i1_7 ), .A2(
        \SB1_1_19/i0[8] ), .A3(\SB1_1_19/i0_4 ), .ZN(
        \SB1_1_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_1/N3  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0[6] ), .A3(\SB1_1_19/i0[9] ), .ZN(
        \SB1_1_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_19/Component_Function_1/N2  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i1_7 ), .A3(\SB1_1_19/i0[8] ), .ZN(
        \SB1_1_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_19/Component_Function_1/N1  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i1[9] ), .ZN(\SB1_1_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_5/N4  ( .A1(\SB1_1_19/i0[9] ), .A2(
        \SB1_1_19/i0[6] ), .A3(\SB1_1_19/i0_4 ), .ZN(
        \SB1_1_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_5/N2  ( .A1(\SB1_1_19/i0_0 ), .A2(
        \SB1_1_19/i0[6] ), .A3(\SB1_1_19/i0[10] ), .ZN(
        \SB1_1_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_19/Component_Function_5/N1  ( .A1(\SB1_1_19/i0_0 ), .A2(
        \SB1_1_19/i3[0] ), .ZN(\SB1_1_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_0/N4  ( .A1(\SB1_1_20/i0[7] ), .A2(
        \SB1_1_20/i0_3 ), .A3(\SB1_1_20/i0_0 ), .ZN(
        \SB1_1_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_20/Component_Function_0/N2  ( .A1(\SB1_1_20/i0[8] ), .A2(
        \SB1_1_20/i0[7] ), .A3(\SB1_1_20/i0[6] ), .ZN(
        \SB1_1_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_20/Component_Function_0/N1  ( .A1(\SB1_1_20/i0[10] ), .A2(
        \SB1_1_20/i0[9] ), .ZN(\SB1_1_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_1/N4  ( .A1(\SB1_1_20/i1_7 ), .A2(
        \SB1_1_20/i0[8] ), .A3(\SB1_1_20/i0_4 ), .ZN(
        \SB1_1_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_20/Component_Function_1/N2  ( .A1(\SB1_1_20/i0_3 ), .A2(
        \SB1_1_20/i1_7 ), .A3(\SB1_1_20/i0[8] ), .ZN(
        \SB1_1_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_20/Component_Function_1/N1  ( .A1(\SB1_1_20/i0_3 ), .A2(
        \SB1_1_20/i1[9] ), .ZN(\SB1_1_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_5/N2  ( .A1(\SB1_1_20/i0_0 ), .A2(
        \SB1_1_20/i0[6] ), .A3(\SB1_1_20/i0[10] ), .ZN(
        \SB1_1_20/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_20/Component_Function_5/N1  ( .A1(\SB1_1_20/i0_0 ), .A2(
        \SB1_1_20/i3[0] ), .ZN(\SB1_1_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_0/N4  ( .A1(\SB1_1_21/i0[7] ), .A2(
        \SB1_1_21/i0_3 ), .A3(\SB1_1_21/i0_0 ), .ZN(
        \SB1_1_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_0/N2  ( .A1(\SB1_1_21/i0[8] ), .A2(
        \SB1_1_21/i0[7] ), .A3(\SB1_1_21/i0[6] ), .ZN(
        \SB1_1_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_21/Component_Function_0/N1  ( .A1(\SB1_1_21/i0[10] ), .A2(
        \SB1_1_21/i0[9] ), .ZN(\SB1_1_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_1/N4  ( .A1(\SB1_1_21/i1_7 ), .A2(
        \SB1_1_21/i0[8] ), .A3(\SB1_1_21/i0_4 ), .ZN(
        \SB1_1_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_1/N2  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i1_7 ), .A3(\SB1_1_21/i0[8] ), .ZN(
        \SB1_1_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_21/Component_Function_1/N1  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i1[9] ), .ZN(\SB1_1_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_5/N2  ( .A1(\SB1_1_21/i0_0 ), .A2(
        \SB1_1_21/i0[6] ), .A3(\SB1_1_21/i0[10] ), .ZN(
        \SB1_1_21/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_21/Component_Function_5/N1  ( .A1(\SB1_1_21/i0_0 ), .A2(
        \SB1_1_21/i3[0] ), .ZN(\SB1_1_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_0/N4  ( .A1(\SB1_1_22/i0[7] ), .A2(
        \SB1_1_22/i0_3 ), .A3(\SB1_1_22/i0_0 ), .ZN(
        \SB1_1_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_22/Component_Function_0/N2  ( .A1(\SB1_1_22/i0[8] ), .A2(
        \SB1_1_22/i0[7] ), .A3(\SB1_1_22/i0[6] ), .ZN(
        \SB1_1_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_22/Component_Function_0/N1  ( .A1(\SB1_1_22/i0[10] ), .A2(
        \SB1_1_22/i0[9] ), .ZN(\SB1_1_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_1/N4  ( .A1(\SB1_1_22/i1_7 ), .A2(
        \SB1_1_22/i0[8] ), .A3(\SB1_1_22/i0_4 ), .ZN(
        \SB1_1_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_22/Component_Function_1/N3  ( .A1(\SB1_1_22/i1_5 ), .A2(
        \SB1_1_22/i0[6] ), .A3(\SB1_1_22/i0[9] ), .ZN(
        \SB1_1_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_22/Component_Function_1/N2  ( .A1(\SB1_1_22/i0_3 ), .A2(
        \SB1_1_22/i1_7 ), .A3(\SB1_1_22/i0[8] ), .ZN(
        \SB1_1_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_22/Component_Function_1/N1  ( .A1(\SB1_1_22/i0_3 ), .A2(
        \SB1_1_22/i1[9] ), .ZN(\SB1_1_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_5/N4  ( .A1(\SB1_1_22/i0[9] ), .A2(
        \SB1_1_22/i0[6] ), .A3(\SB1_1_22/i0_4 ), .ZN(
        \SB1_1_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_22/Component_Function_5/N2  ( .A1(\SB1_1_22/i0_0 ), .A2(
        \SB1_1_22/i0[6] ), .A3(\SB1_1_22/i0[10] ), .ZN(
        \SB1_1_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_22/Component_Function_5/N1  ( .A1(\SB1_1_22/i0_0 ), .A2(
        \SB1_1_22/i3[0] ), .ZN(\SB1_1_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_0/N4  ( .A1(\SB1_1_23/i0[7] ), .A2(
        \SB1_1_23/i0_3 ), .A3(\SB1_1_23/i0_0 ), .ZN(
        \SB1_1_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_23/Component_Function_0/N3  ( .A1(\SB1_1_23/i0[10] ), .A2(
        \SB1_1_23/i0_4 ), .A3(\SB1_1_23/i0_3 ), .ZN(
        \SB1_1_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_23/Component_Function_0/N2  ( .A1(\SB1_1_23/i0[8] ), .A2(
        \SB1_1_23/i0[7] ), .A3(\SB1_1_23/i0[6] ), .ZN(
        \SB1_1_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_23/Component_Function_0/N1  ( .A1(\SB1_1_23/i0[10] ), .A2(
        \SB1_1_23/i0[9] ), .ZN(\SB1_1_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_1/N4  ( .A1(\SB1_1_23/i1_7 ), .A2(
        \SB1_1_23/i0[8] ), .A3(\SB1_1_23/i0_4 ), .ZN(
        \SB1_1_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_23/Component_Function_1/N3  ( .A1(\SB1_1_23/i1_5 ), .A2(
        \SB1_1_23/i0[6] ), .A3(\SB1_1_23/i0[9] ), .ZN(
        \SB1_1_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_23/Component_Function_1/N2  ( .A1(\SB1_1_23/i0_3 ), .A2(
        \SB1_1_23/i1_7 ), .A3(\SB1_1_23/i0[8] ), .ZN(
        \SB1_1_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_23/Component_Function_1/N1  ( .A1(\SB1_1_23/i0_3 ), .A2(
        \SB1_1_23/i1[9] ), .ZN(\SB1_1_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_5/N4  ( .A1(\SB1_1_23/i0[9] ), .A2(
        \SB1_1_23/i0[6] ), .A3(\SB1_1_23/i0_4 ), .ZN(
        \SB1_1_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_23/Component_Function_5/N2  ( .A1(\SB1_1_23/i0_0 ), .A2(
        \SB1_1_23/i0[6] ), .A3(\SB1_1_23/i0[10] ), .ZN(
        \SB1_1_23/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_23/Component_Function_5/N1  ( .A1(\SB1_1_23/i0_0 ), .A2(
        \SB1_1_23/i3[0] ), .ZN(\SB1_1_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_0/N4  ( .A1(\SB1_1_24/i0[7] ), .A2(
        \SB1_1_24/i0_3 ), .A3(\SB1_1_24/i0_0 ), .ZN(
        \SB1_1_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_24/Component_Function_0/N3  ( .A1(\SB1_1_24/i0[10] ), .A2(
        \SB1_1_24/i0_4 ), .A3(\SB1_1_24/i0_3 ), .ZN(
        \SB1_1_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_24/Component_Function_0/N2  ( .A1(\SB1_1_24/i0[8] ), .A2(
        \SB1_1_24/i0[7] ), .A3(\SB1_1_24/i0[6] ), .ZN(
        \SB1_1_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_24/Component_Function_0/N1  ( .A1(\SB1_1_24/i0[10] ), .A2(
        \SB1_1_24/i0[9] ), .ZN(\SB1_1_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_1/N3  ( .A1(\SB1_1_24/i1_5 ), .A2(
        \SB1_1_24/i0[6] ), .A3(\SB1_1_24/i0[9] ), .ZN(
        \SB1_1_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_24/Component_Function_1/N2  ( .A1(\SB1_1_24/i0_3 ), .A2(
        \SB1_1_24/i1_7 ), .A3(\SB1_1_24/i0[8] ), .ZN(
        \SB1_1_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_24/Component_Function_1/N1  ( .A1(\SB1_1_24/i0_3 ), .A2(
        \SB1_1_24/i1[9] ), .ZN(\SB1_1_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_5/N4  ( .A1(\SB1_1_24/i0[9] ), .A2(
        \SB1_1_24/i0[6] ), .A3(\SB1_1_24/i0_4 ), .ZN(
        \SB1_1_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_24/Component_Function_5/N2  ( .A1(\SB1_1_24/i0_0 ), .A2(
        \SB1_1_24/i0[6] ), .A3(\SB1_1_24/i0[10] ), .ZN(
        \SB1_1_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_24/Component_Function_5/N1  ( .A1(\SB1_1_24/i0_0 ), .A2(
        \SB1_1_24/i3[0] ), .ZN(\SB1_1_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_0/N4  ( .A1(\SB1_1_25/i0[7] ), .A2(
        \SB1_1_25/i0_3 ), .A3(\SB1_1_25/i0_0 ), .ZN(
        \SB1_1_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_0/N3  ( .A1(\SB1_1_25/i0[10] ), .A2(
        \SB1_1_25/i0_4 ), .A3(\SB1_1_25/i0_3 ), .ZN(
        \SB1_1_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_25/Component_Function_0/N2  ( .A1(\SB1_1_25/i0[8] ), .A2(
        \SB1_1_25/i0[7] ), .A3(\SB1_1_25/i0[6] ), .ZN(
        \SB1_1_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_25/Component_Function_0/N1  ( .A1(\SB1_1_25/i0[10] ), .A2(
        \SB1_1_25/i0[9] ), .ZN(\SB1_1_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_1/N4  ( .A1(\SB1_1_25/i1_7 ), .A2(
        \SB1_1_25/i0[8] ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_1/N3  ( .A1(\SB1_1_25/i1_5 ), .A2(
        \SB1_1_25/i0[6] ), .A3(\SB1_1_25/i0[9] ), .ZN(
        \SB1_1_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_25/Component_Function_1/N2  ( .A1(\SB1_1_25/i0_3 ), .A2(
        \SB1_1_25/i1_7 ), .A3(\SB1_1_25/i0[8] ), .ZN(
        \SB1_1_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_25/Component_Function_1/N1  ( .A1(\SB1_1_25/i0_3 ), .A2(
        \SB1_1_25/i1[9] ), .ZN(\SB1_1_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_5/N4  ( .A1(\SB1_1_25/i0[9] ), .A2(
        \SB1_1_25/i0[6] ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_5/N2  ( .A1(\SB1_1_25/i0_0 ), .A2(
        \SB1_1_25/i0[6] ), .A3(\SB1_1_25/i0[10] ), .ZN(
        \SB1_1_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_25/Component_Function_5/N1  ( .A1(\SB1_1_25/i0_0 ), .A2(
        \SB1_1_25/i3[0] ), .ZN(\SB1_1_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_0/N2  ( .A1(\SB1_1_26/i0[8] ), .A2(
        \SB1_1_26/i0[7] ), .A3(\SB1_1_26/i0[6] ), .ZN(
        \SB1_1_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_26/Component_Function_0/N1  ( .A1(\SB1_1_26/i0[10] ), .A2(
        \SB1_1_26/i0[9] ), .ZN(\SB1_1_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_1/N4  ( .A1(\SB1_1_26/i1_7 ), .A2(
        \SB1_1_26/i0[8] ), .A3(\SB1_1_26/i0_4 ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_26/Component_Function_1/N3  ( .A1(\SB1_1_26/i1_5 ), .A2(
        \SB1_1_26/i0[6] ), .A3(\SB1_1_26/i0[9] ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_26/Component_Function_1/N2  ( .A1(\SB1_1_26/i0_3 ), .A2(
        \SB1_1_26/i1_7 ), .A3(\SB1_1_26/i0[8] ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_26/Component_Function_1/N1  ( .A1(\SB1_1_26/i0_3 ), .A2(
        \SB1_1_26/i1[9] ), .ZN(\SB1_1_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_5/N4  ( .A1(\SB1_1_26/i0[9] ), .A2(
        \SB1_1_26/i0[6] ), .A3(\SB1_1_26/i0_4 ), .ZN(
        \SB1_1_26/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_26/Component_Function_5/N1  ( .A1(\SB1_1_26/i0_0 ), .A2(
        \SB1_1_26/i3[0] ), .ZN(\SB1_1_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_0/N4  ( .A1(\SB1_1_27/i0[7] ), .A2(
        \SB1_1_27/i0_3 ), .A3(\SB1_1_27/i0_0 ), .ZN(
        \SB1_1_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_0/N3  ( .A1(\SB1_1_27/i0[10] ), .A2(
        \SB1_1_27/i0_4 ), .A3(\SB1_1_27/i0_3 ), .ZN(
        \SB1_1_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_27/Component_Function_0/N2  ( .A1(\SB1_1_27/i0[8] ), .A2(
        \SB1_1_27/i0[7] ), .A3(\SB1_1_27/i0[6] ), .ZN(
        \SB1_1_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_27/Component_Function_0/N1  ( .A1(\SB1_1_27/i0[10] ), .A2(
        \SB1_1_27/i0[9] ), .ZN(\SB1_1_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_1/N4  ( .A1(\SB1_1_27/i1_7 ), .A2(
        \SB1_1_27/i0[8] ), .A3(\SB1_1_27/i0_4 ), .ZN(
        \SB1_1_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_1/N3  ( .A1(\SB1_1_27/i1_5 ), .A2(
        \SB1_1_27/i0[6] ), .A3(\SB1_1_27/i0[9] ), .ZN(
        \SB1_1_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_27/Component_Function_1/N2  ( .A1(\SB1_1_27/i0_3 ), .A2(
        \SB1_1_27/i1_7 ), .A3(\SB1_1_27/i0[8] ), .ZN(
        \SB1_1_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_27/Component_Function_1/N1  ( .A1(\SB1_1_27/i0_3 ), .A2(
        \SB1_1_27/i1[9] ), .ZN(\SB1_1_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_5/N4  ( .A1(\SB1_1_27/i0[9] ), .A2(
        \SB1_1_27/i0[6] ), .A3(\SB1_1_27/i0_4 ), .ZN(
        \SB1_1_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_5/N2  ( .A1(\SB1_1_27/i0_0 ), .A2(
        \SB1_1_27/i0[6] ), .A3(\SB1_1_27/i0[10] ), .ZN(
        \SB1_1_27/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_27/Component_Function_5/N1  ( .A1(\SB1_1_27/i0_0 ), .A2(
        \SB1_1_27/i3[0] ), .ZN(\SB1_1_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_0/N4  ( .A1(\SB1_1_28/i0[7] ), .A2(
        \SB1_1_28/i0_3 ), .A3(\SB1_1_28/i0_0 ), .ZN(
        \SB1_1_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_0/N2  ( .A1(\SB1_1_28/i0[8] ), .A2(
        \SB1_1_28/i0[7] ), .A3(\SB1_1_28/i0[6] ), .ZN(
        \SB1_1_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_28/Component_Function_0/N1  ( .A1(\SB1_1_28/i0[10] ), .A2(
        \SB1_1_28/i0[9] ), .ZN(\SB1_1_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_1/N4  ( .A1(\SB1_1_28/i1_7 ), .A2(
        \SB1_1_28/i0[8] ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_1/N3  ( .A1(\SB1_1_28/i1_5 ), .A2(
        \SB1_1_28/i0[6] ), .A3(\SB1_1_28/i0[9] ), .ZN(
        \SB1_1_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_28/Component_Function_1/N2  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i1_7 ), .A3(\SB1_1_28/i0[8] ), .ZN(
        \SB1_1_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_28/Component_Function_1/N1  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i1[9] ), .ZN(\SB1_1_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_5/N4  ( .A1(\SB1_1_28/i0[9] ), .A2(
        \SB1_1_28/i0[6] ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_5/N2  ( .A1(\SB1_1_28/i0_0 ), .A2(
        \SB1_1_28/i0[6] ), .A3(\SB1_1_28/i0[10] ), .ZN(
        \SB1_1_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_28/Component_Function_5/N1  ( .A1(\SB1_1_28/i0_0 ), .A2(
        \SB1_1_28/i3[0] ), .ZN(\SB1_1_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N4  ( .A1(\SB1_1_29/i0[7] ), .A2(
        \SB1_1_29/i0_3 ), .A3(\SB1_1_29/i0_0 ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N3  ( .A1(\SB1_1_29/i0[10] ), .A2(
        \SB1_1_29/i0_4 ), .A3(\SB1_1_29/i0_3 ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N2  ( .A1(\SB1_1_29/i0[8] ), .A2(
        \SB1_1_29/i0[7] ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_29/Component_Function_0/N1  ( .A1(\SB1_1_29/i0[10] ), .A2(
        \SB1_1_29/i0[9] ), .ZN(\SB1_1_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_1/N4  ( .A1(\SB1_1_29/i1_7 ), .A2(
        \SB1_1_29/i0[8] ), .A3(\SB1_1_29/i0_4 ), .ZN(
        \SB1_1_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_29/Component_Function_1/N2  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i1_7 ), .A3(\SB1_1_29/i0[8] ), .ZN(
        \SB1_1_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_29/Component_Function_1/N1  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i1[9] ), .ZN(\SB1_1_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_5/N4  ( .A1(\SB1_1_29/i0[9] ), .A2(
        \SB1_1_29/i0[6] ), .A3(\SB1_1_29/i0_4 ), .ZN(
        \SB1_1_29/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_29/Component_Function_5/N1  ( .A1(\SB1_1_29/i0_0 ), .A2(
        \SB1_1_29/i3[0] ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_0/N4  ( .A1(\SB1_1_30/i0[7] ), .A2(
        \SB1_1_30/i0_3 ), .A3(\SB1_1_30/i0_0 ), .ZN(
        \SB1_1_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_30/Component_Function_0/N3  ( .A1(\SB1_1_30/i0[10] ), .A2(
        \SB1_1_30/i0_4 ), .A3(\SB1_1_30/i0_3 ), .ZN(
        \SB1_1_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_30/Component_Function_0/N2  ( .A1(\SB1_1_30/i0[8] ), .A2(
        \SB1_1_30/i0[7] ), .A3(\SB1_1_30/i0[6] ), .ZN(
        \SB1_1_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_30/Component_Function_0/N1  ( .A1(\SB1_1_30/i0[10] ), .A2(
        \SB1_1_30/i0[9] ), .ZN(\SB1_1_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_1/N3  ( .A1(\SB1_1_30/i1_5 ), .A2(
        \SB1_1_30/i0[6] ), .A3(\SB1_1_30/i0[9] ), .ZN(
        \SB1_1_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_30/Component_Function_1/N2  ( .A1(\SB1_1_30/i0_3 ), .A2(
        \SB1_1_30/i1_7 ), .A3(\SB1_1_30/i0[8] ), .ZN(
        \SB1_1_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_30/Component_Function_1/N1  ( .A1(\SB1_1_30/i0_3 ), .A2(
        \SB1_1_30/i1[9] ), .ZN(\SB1_1_30/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_30/Component_Function_5/N1  ( .A1(\SB1_1_30/i0_0 ), .A2(
        \SB1_1_30/i3[0] ), .ZN(\SB1_1_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_0/N4  ( .A1(\SB1_1_31/i0[7] ), .A2(
        \SB1_1_31/i0_3 ), .A3(\SB1_1_31/i0_0 ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_31/Component_Function_0/N2  ( .A1(\SB1_1_31/i0[8] ), .A2(
        \SB1_1_31/i0[7] ), .A3(\SB1_1_31/i0[6] ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_31/Component_Function_0/N1  ( .A1(\SB1_1_31/i0[10] ), .A2(
        \SB1_1_31/i0[9] ), .ZN(\SB1_1_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_1/N4  ( .A1(\SB1_1_31/i1_7 ), .A2(
        \SB1_1_31/i0[8] ), .A3(\SB1_1_31/i0_4 ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_31/Component_Function_1/N3  ( .A1(\SB1_1_31/i1_5 ), .A2(
        \SB1_1_31/i0[6] ), .A3(\SB1_1_31/i0[9] ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_31/Component_Function_1/N2  ( .A1(\SB1_1_31/i0_3 ), .A2(
        \SB1_1_31/i1_7 ), .A3(\SB1_1_31/i0[8] ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_31/Component_Function_1/N1  ( .A1(\SB1_1_31/i0_3 ), .A2(
        \SB1_1_31/i1[9] ), .ZN(\SB1_1_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_5/N4  ( .A1(\SB1_1_31/i0[9] ), .A2(
        \SB1_1_31/i0[6] ), .A3(\SB1_1_31/i0_4 ), .ZN(
        \SB1_1_31/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_31/Component_Function_5/N1  ( .A1(\SB1_1_31/i0_0 ), .A2(
        \SB1_1_31/i3[0] ), .ZN(\SB1_1_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_0/Component_Function_0/N4  ( .A1(\SB2_1_0/i0[7] ), .A2(
        \SB2_1_0/i0_3 ), .A3(\SB2_1_0/i0_0 ), .ZN(
        \SB2_1_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_0/Component_Function_0/N3  ( .A1(\SB2_1_0/i0[10] ), .A2(
        \SB2_1_0/i0_4 ), .A3(\SB2_1_0/i0_3 ), .ZN(
        \SB2_1_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_0/Component_Function_0/N2  ( .A1(\SB2_1_0/i0[8] ), .A2(
        \SB2_1_0/i0[7] ), .A3(\SB2_1_0/i0[6] ), .ZN(
        \SB2_1_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_0/Component_Function_0/N1  ( .A1(\SB2_1_0/i0[10] ), .A2(
        \SB2_1_0/i0[9] ), .ZN(\SB2_1_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_0/Component_Function_1/N4  ( .A1(\SB2_1_0/i1_7 ), .A2(
        \SB2_1_0/i0[8] ), .A3(\SB2_1_0/i0_4 ), .ZN(
        \SB2_1_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_0/Component_Function_1/N3  ( .A1(\SB2_1_0/i1_5 ), .A2(
        \SB2_1_0/i0[6] ), .A3(\SB2_1_0/i0[9] ), .ZN(
        \SB2_1_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_0/Component_Function_1/N2  ( .A1(\SB2_1_0/i0_3 ), .A2(
        \SB2_1_0/i1_7 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        \SB2_1_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_0/Component_Function_1/N1  ( .A1(\SB2_1_0/i0_3 ), .A2(
        \SB2_1_0/i1[9] ), .ZN(\SB2_1_0/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_0/Component_Function_5/N1  ( .A1(\SB2_1_0/i0_0 ), .A2(
        \SB2_1_0/i3[0] ), .ZN(\SB2_1_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_0/N4  ( .A1(\SB2_1_1/i0[7] ), .A2(
        \SB2_1_1/i0_3 ), .A3(\SB2_1_1/i0_0 ), .ZN(
        \SB2_1_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_1/Component_Function_0/N3  ( .A1(\SB2_1_1/i0[10] ), .A2(
        \SB2_1_1/i0_4 ), .A3(\SB2_1_1/i0_3 ), .ZN(
        \SB2_1_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_1/Component_Function_0/N2  ( .A1(\SB2_1_1/i0[8] ), .A2(
        \SB2_1_1/i0[7] ), .A3(\SB2_1_1/i0[6] ), .ZN(
        \SB2_1_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_1/Component_Function_0/N1  ( .A1(\SB2_1_1/i0[10] ), .A2(
        \SB2_1_1/i0[9] ), .ZN(\SB2_1_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_1/N4  ( .A1(\SB2_1_1/i1_7 ), .A2(
        \SB2_1_1/i0[8] ), .A3(\SB2_1_1/i0_4 ), .ZN(
        \SB2_1_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_1/Component_Function_1/N3  ( .A1(\SB2_1_1/i1_5 ), .A2(
        \SB2_1_1/i0[6] ), .A3(\SB2_1_1/i0[9] ), .ZN(
        \SB2_1_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_1/Component_Function_1/N2  ( .A1(\SB2_1_1/i0_3 ), .A2(
        \SB2_1_1/i1_7 ), .A3(\SB2_1_1/i0[8] ), .ZN(
        \SB2_1_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_1/Component_Function_1/N1  ( .A1(\SB2_1_1/i0_3 ), .A2(
        \SB2_1_1/i1[9] ), .ZN(\SB2_1_1/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_1/Component_Function_5/N1  ( .A1(\SB2_1_1/i0_0 ), .A2(
        \SB2_1_1/i3[0] ), .ZN(\SB2_1_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_0/N4  ( .A1(\SB2_1_2/i0[7] ), .A2(
        \SB2_1_2/i0_3 ), .A3(\SB2_1_2/i0_0 ), .ZN(
        \SB2_1_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_2/Component_Function_0/N3  ( .A1(\SB2_1_2/i0[10] ), .A2(
        \SB2_1_2/i0_4 ), .A3(\SB2_1_2/i0_3 ), .ZN(
        \SB2_1_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_2/Component_Function_0/N2  ( .A1(\SB2_1_2/i0[8] ), .A2(
        \SB2_1_2/i0[7] ), .A3(\SB2_1_2/i0[6] ), .ZN(
        \SB2_1_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_2/Component_Function_0/N1  ( .A1(\SB2_1_2/i0[10] ), .A2(
        \SB2_1_2/i0[9] ), .ZN(\SB2_1_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_1/N3  ( .A1(\SB2_1_2/i1_5 ), .A2(
        \SB2_1_2/i0[6] ), .A3(\SB2_1_2/i0[9] ), .ZN(
        \SB2_1_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_2/Component_Function_1/N2  ( .A1(\SB2_1_2/i0_3 ), .A2(
        \SB2_1_2/i1_7 ), .A3(\SB2_1_2/i0[8] ), .ZN(
        \SB2_1_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_2/Component_Function_1/N1  ( .A1(\SB2_1_2/i0_3 ), .A2(
        \SB2_1_2/i1[9] ), .ZN(\SB2_1_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_5/N2  ( .A1(\SB2_1_2/i0_0 ), .A2(
        \SB2_1_2/i0[6] ), .A3(\SB2_1_2/i0[10] ), .ZN(
        \SB2_1_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_2/Component_Function_5/N1  ( .A1(\SB2_1_2/i0_0 ), .A2(
        \SB2_1_2/i3[0] ), .ZN(\SB2_1_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_0/N4  ( .A1(\SB2_1_3/i0[7] ), .A2(
        \SB2_1_3/i0_3 ), .A3(\SB2_1_3/i0_0 ), .ZN(
        \SB2_1_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_3/Component_Function_0/N3  ( .A1(\SB2_1_3/i0[10] ), .A2(
        \SB2_1_3/i0_4 ), .A3(\SB2_1_3/i0_3 ), .ZN(
        \SB2_1_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_3/Component_Function_0/N2  ( .A1(\SB2_1_3/i0[8] ), .A2(
        \SB2_1_3/i0[7] ), .A3(\SB2_1_3/i0[6] ), .ZN(
        \SB2_1_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_3/Component_Function_0/N1  ( .A1(\SB2_1_3/i0[10] ), .A2(
        \SB2_1_3/i0[9] ), .ZN(\SB2_1_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_1/N3  ( .A1(\SB2_1_3/i1_5 ), .A2(
        \SB2_1_3/i0[6] ), .A3(\SB2_1_3/i0[9] ), .ZN(
        \SB2_1_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_3/Component_Function_1/N2  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i1_7 ), .A3(\SB2_1_3/i0[8] ), .ZN(
        \SB2_1_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_3/Component_Function_1/N1  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i1[9] ), .ZN(\SB2_1_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_5/N3  ( .A1(\SB2_1_3/i1[9] ), .A2(
        \SB2_1_3/i0_4 ), .A3(\SB2_1_3/i0_3 ), .ZN(
        \SB2_1_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_0/N4  ( .A1(\SB2_1_4/i0[7] ), .A2(
        \SB2_1_4/i0_3 ), .A3(\SB2_1_4/i0_0 ), .ZN(
        \SB2_1_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_0/N3  ( .A1(\SB2_1_4/i0[10] ), .A2(
        \SB2_1_4/i0_4 ), .A3(\SB2_1_4/i0_3 ), .ZN(
        \SB2_1_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_0/N2  ( .A1(\SB2_1_4/i0[8] ), .A2(
        \SB2_1_4/i0[7] ), .A3(\SB2_1_4/i0[6] ), .ZN(
        \SB2_1_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_4/Component_Function_0/N1  ( .A1(\SB2_1_4/i0[10] ), .A2(
        \SB2_1_4/i0[9] ), .ZN(\SB2_1_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_1/N4  ( .A1(\SB2_1_4/i1_7 ), .A2(
        \SB2_1_4/i0[8] ), .A3(\SB2_1_4/i0_4 ), .ZN(
        \SB2_1_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_1/N3  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB2_1_4/i0[6] ), .A3(\SB2_1_4/i0[9] ), .ZN(
        \SB2_1_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_1/N2  ( .A1(\SB2_1_4/i0_3 ), .A2(
        \SB2_1_4/i1_7 ), .A3(\SB2_1_4/i0[8] ), .ZN(
        \SB2_1_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_4/Component_Function_1/N1  ( .A1(\SB2_1_4/i0_3 ), .A2(
        \SB2_1_4/i1[9] ), .ZN(\SB2_1_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_5/N3  ( .A1(\SB2_1_4/i1[9] ), .A2(
        \SB2_1_4/i0_4 ), .A3(\SB2_1_4/i0_3 ), .ZN(
        \SB2_1_4/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_4/Component_Function_5/N1  ( .A1(\SB2_1_4/i0_0 ), .A2(
        \SB2_1_4/i3[0] ), .ZN(\SB2_1_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_0/N4  ( .A1(\SB2_1_5/i0[7] ), .A2(
        \SB2_1_5/i0_3 ), .A3(\SB2_1_5/i0_0 ), .ZN(
        \SB2_1_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_5/Component_Function_0/N3  ( .A1(\SB2_1_5/i0[10] ), .A2(
        \SB2_1_5/i0_4 ), .A3(\SB2_1_5/i0_3 ), .ZN(
        \SB2_1_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_5/Component_Function_0/N2  ( .A1(\SB2_1_5/i0[8] ), .A2(
        \SB2_1_5/i0[7] ), .A3(\SB2_1_5/i0[6] ), .ZN(
        \SB2_1_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_5/Component_Function_0/N1  ( .A1(\SB2_1_5/i0[10] ), .A2(
        \SB2_1_5/i0[9] ), .ZN(\SB2_1_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_1/N3  ( .A1(\SB2_1_5/i1_5 ), .A2(
        \SB2_1_5/i0[6] ), .A3(\SB2_1_5/i0[9] ), .ZN(
        \SB2_1_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_5/Component_Function_1/N2  ( .A1(\SB2_1_5/i0_3 ), .A2(
        \SB2_1_5/i1_7 ), .A3(\SB2_1_5/i0[8] ), .ZN(
        \SB2_1_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_5/Component_Function_1/N1  ( .A1(\SB2_1_5/i0_3 ), .A2(
        \SB2_1_5/i1[9] ), .ZN(\SB2_1_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_5/N3  ( .A1(\SB2_1_5/i1[9] ), .A2(
        \SB2_1_5/i0_4 ), .A3(\SB2_1_5/i0_3 ), .ZN(
        \SB2_1_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_5/Component_Function_5/N2  ( .A1(\SB2_1_5/i0_0 ), .A2(
        \SB2_1_5/i0[6] ), .A3(\SB2_1_5/i0[10] ), .ZN(
        \SB2_1_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_6/Component_Function_0/N4  ( .A1(\SB2_1_6/i0[7] ), .A2(
        \SB2_1_6/i0_3 ), .A3(\SB2_1_6/i0_0 ), .ZN(
        \SB2_1_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_6/Component_Function_0/N3  ( .A1(\SB2_1_6/i0[10] ), .A2(
        \SB2_1_6/i0_4 ), .A3(\SB2_1_6/i0_3 ), .ZN(
        \SB2_1_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_6/Component_Function_0/N2  ( .A1(\SB2_1_6/i0[8] ), .A2(
        \SB2_1_6/i0[7] ), .A3(\SB2_1_6/i0[6] ), .ZN(
        \SB2_1_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_6/Component_Function_0/N1  ( .A1(\SB2_1_6/i0[10] ), .A2(
        \SB2_1_6/i0[9] ), .ZN(\SB2_1_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_1/N4  ( .A1(\SB2_1_6/i1_7 ), .A2(
        \SB2_1_6/i0[8] ), .A3(\SB2_1_6/i0_4 ), .ZN(
        \SB2_1_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_6/Component_Function_1/N3  ( .A1(\SB2_1_6/i1_5 ), .A2(
        \SB2_1_6/i0[6] ), .A3(\SB2_1_6/i0[9] ), .ZN(
        \SB2_1_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_6/Component_Function_1/N2  ( .A1(\SB2_1_6/i0_3 ), .A2(
        \SB2_1_6/i1_7 ), .A3(\SB2_1_6/i0[8] ), .ZN(
        \SB2_1_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_6/Component_Function_1/N1  ( .A1(\SB2_1_6/i0_3 ), .A2(
        \SB2_1_6/i1[9] ), .ZN(\SB2_1_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_5/N2  ( .A1(\SB2_1_6/i0_0 ), .A2(
        \SB2_1_6/i0[6] ), .A3(\SB2_1_6/i0[10] ), .ZN(
        \SB2_1_6/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_6/Component_Function_5/N1  ( .A1(\SB2_1_6/i0_0 ), .A2(
        \SB2_1_6/i3[0] ), .ZN(\SB2_1_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_0/N4  ( .A1(\SB2_1_7/i0[7] ), .A2(
        \SB2_1_7/i0_3 ), .A3(\SB2_1_7/i0_0 ), .ZN(
        \SB2_1_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_7/Component_Function_0/N3  ( .A1(\SB2_1_7/i0[10] ), .A2(
        \SB2_1_7/i0_4 ), .A3(\SB2_1_7/i0_3 ), .ZN(
        \SB2_1_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_7/Component_Function_0/N2  ( .A1(\SB2_1_7/i0[8] ), .A2(
        \SB2_1_7/i0[7] ), .A3(\SB2_1_7/i0[6] ), .ZN(
        \SB2_1_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_7/Component_Function_0/N1  ( .A1(\SB2_1_7/i0[10] ), .A2(
        \SB2_1_7/i0[9] ), .ZN(\SB2_1_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_1/N3  ( .A1(\SB2_1_7/i1_5 ), .A2(
        \SB2_1_7/i0[6] ), .A3(\SB2_1_7/i0[9] ), .ZN(
        \SB2_1_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_7/Component_Function_1/N2  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i1_7 ), .A3(\SB2_1_7/i0[8] ), .ZN(
        \SB2_1_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_7/Component_Function_1/N1  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i1[9] ), .ZN(\SB2_1_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_7/Component_Function_5/N1  ( .A1(\SB2_1_7/i0_0 ), .A2(
        \SB2_1_7/i3[0] ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_0/N4  ( .A1(\SB2_1_8/i0[7] ), .A2(
        \SB2_1_8/i0_3 ), .A3(\SB2_1_8/i0_0 ), .ZN(
        \SB2_1_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_8/Component_Function_0/N3  ( .A1(\SB2_1_8/i0[10] ), .A2(
        \SB2_1_8/i0_4 ), .A3(\SB2_1_8/i0_3 ), .ZN(
        \SB2_1_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_8/Component_Function_0/N2  ( .A1(\SB2_1_8/i0[8] ), .A2(
        \SB2_1_8/i0[7] ), .A3(\SB2_1_8/i0[6] ), .ZN(
        \SB2_1_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_8/Component_Function_0/N1  ( .A1(\SB2_1_8/i0[10] ), .A2(
        \SB2_1_8/i0[9] ), .ZN(\SB2_1_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_1/N4  ( .A1(\SB2_1_8/i1_7 ), .A2(
        \SB2_1_8/i0[8] ), .A3(\SB2_1_8/i0_4 ), .ZN(
        \SB2_1_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_8/Component_Function_1/N3  ( .A1(\SB2_1_8/i1_5 ), .A2(
        \SB2_1_8/i0[6] ), .A3(\SB2_1_8/i0[9] ), .ZN(
        \SB2_1_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_8/Component_Function_1/N2  ( .A1(\SB2_1_8/i0_3 ), .A2(
        \SB2_1_8/i1_7 ), .A3(\SB2_1_8/i0[8] ), .ZN(
        \SB2_1_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_8/Component_Function_1/N1  ( .A1(\SB2_1_8/i0_3 ), .A2(
        \SB2_1_8/i1[9] ), .ZN(\SB2_1_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_8/Component_Function_5/N1  ( .A1(\SB2_1_8/i0_0 ), .A2(
        \SB2_1_8/i3[0] ), .ZN(\SB2_1_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_9/Component_Function_0/N4  ( .A1(\SB2_1_9/i0[7] ), .A2(
        \SB2_1_9/i0_3 ), .A3(\SB2_1_9/i0_0 ), .ZN(
        \SB2_1_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_9/Component_Function_0/N3  ( .A1(\SB2_1_9/i0[10] ), .A2(
        \SB2_1_9/i0_4 ), .A3(\SB2_1_9/i0_3 ), .ZN(
        \SB2_1_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_9/Component_Function_0/N2  ( .A1(\SB2_1_9/i0[8] ), .A2(
        \SB2_1_9/i0[7] ), .A3(\SB2_1_9/i0[6] ), .ZN(
        \SB2_1_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_9/Component_Function_0/N1  ( .A1(\SB2_1_9/i0[10] ), .A2(
        \SB2_1_9/i0[9] ), .ZN(\SB2_1_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_9/Component_Function_1/N4  ( .A1(\SB2_1_9/i1_7 ), .A2(
        \SB2_1_9/i0[8] ), .A3(\SB2_1_9/i0_4 ), .ZN(
        \SB2_1_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_9/Component_Function_1/N3  ( .A1(\SB2_1_9/i1_5 ), .A2(
        \SB2_1_9/i0[6] ), .A3(\SB2_1_9/i0[9] ), .ZN(
        \SB2_1_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_9/Component_Function_1/N2  ( .A1(\SB2_1_9/i0_3 ), .A2(
        \SB2_1_9/i1_7 ), .A3(\SB2_1_9/i0[8] ), .ZN(
        \SB2_1_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_9/Component_Function_1/N1  ( .A1(\SB2_1_9/i0_3 ), .A2(
        \SB2_1_9/i1[9] ), .ZN(\SB2_1_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_9/Component_Function_5/N3  ( .A1(\SB2_1_9/i1[9] ), .A2(
        \SB2_1_9/i0_4 ), .A3(\SB2_1_9/i0_3 ), .ZN(
        \SB2_1_9/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_9/Component_Function_5/N1  ( .A1(\SB2_1_9/i0_0 ), .A2(
        \SB2_1_9/i3[0] ), .ZN(\SB2_1_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_10/Component_Function_0/N4  ( .A1(\SB2_1_10/i0[7] ), .A2(
        \SB2_1_10/i0_3 ), .A3(\SB2_1_10/i0_0 ), .ZN(
        \SB2_1_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_10/Component_Function_0/N3  ( .A1(\SB2_1_10/i0[10] ), .A2(
        \SB2_1_10/i0_4 ), .A3(\SB2_1_10/i0_3 ), .ZN(
        \SB2_1_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_10/Component_Function_0/N2  ( .A1(\SB2_1_10/i0[8] ), .A2(
        \SB2_1_10/i0[7] ), .A3(\SB2_1_10/i0[6] ), .ZN(
        \SB2_1_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_10/Component_Function_0/N1  ( .A1(\SB2_1_10/i0[10] ), .A2(
        \SB2_1_10/i0[9] ), .ZN(\SB2_1_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N4  ( .A1(\SB2_1_10/i1_7 ), .A2(
        \SB2_1_10/i0[8] ), .A3(\SB2_1_10/i0_4 ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N3  ( .A1(\SB2_1_10/i1_5 ), .A2(
        \SB2_1_10/i0[6] ), .A3(\SB2_1_10/i0[9] ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N2  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i1_7 ), .A3(\SB2_1_10/i0[8] ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_10/Component_Function_1/N1  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i1[9] ), .ZN(\SB2_1_10/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_10/Component_Function_5/N1  ( .A1(\SB2_1_10/i0_0 ), .A2(
        \SB2_1_10/i3[0] ), .ZN(\SB2_1_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_0/N4  ( .A1(\SB2_1_11/i0[7] ), .A2(
        \SB2_1_11/i0_3 ), .A3(\SB2_1_11/i0_0 ), .ZN(
        \SB2_1_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_11/Component_Function_0/N3  ( .A1(\SB2_1_11/i0[10] ), .A2(
        \SB2_1_11/i0_4 ), .A3(\SB2_1_11/i0_3 ), .ZN(
        \SB2_1_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_11/Component_Function_0/N2  ( .A1(\SB2_1_11/i0[8] ), .A2(
        \SB2_1_11/i0[7] ), .A3(\SB2_1_11/i0[6] ), .ZN(
        \SB2_1_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_11/Component_Function_0/N1  ( .A1(\SB2_1_11/i0[10] ), .A2(
        \SB2_1_11/i0[9] ), .ZN(\SB2_1_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_1/N4  ( .A1(\SB2_1_11/i1_7 ), .A2(
        \SB2_1_11/i0[8] ), .A3(\SB2_1_11/i0_4 ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_11/Component_Function_1/N3  ( .A1(\SB2_1_11/i1_5 ), .A2(
        \SB2_1_11/i0[6] ), .A3(\SB2_1_11/i0[9] ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_11/Component_Function_1/N2  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i1_7 ), .A3(\SB2_1_11/i0[8] ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_11/Component_Function_1/N1  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i1[9] ), .ZN(\SB2_1_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_0/N4  ( .A1(\SB2_1_12/i0[7] ), .A2(
        \SB2_1_12/i0_3 ), .A3(\SB2_1_12/i0_0 ), .ZN(
        \SB2_1_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_12/Component_Function_0/N3  ( .A1(\SB2_1_12/i0[10] ), .A2(
        \SB2_1_12/i0_4 ), .A3(\SB2_1_12/i0_3 ), .ZN(
        \SB2_1_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_12/Component_Function_0/N2  ( .A1(\SB2_1_12/i0[8] ), .A2(
        \SB2_1_12/i0[7] ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_12/Component_Function_0/N1  ( .A1(\SB2_1_12/i0[10] ), .A2(
        \SB2_1_12/i0[9] ), .ZN(\SB2_1_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_1/N3  ( .A1(\SB2_1_12/i1_5 ), .A2(
        \SB2_1_12/i0[6] ), .A3(\SB2_1_12/i0[9] ), .ZN(
        \SB2_1_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_12/Component_Function_1/N2  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i1_7 ), .A3(\SB2_1_12/i0[8] ), .ZN(
        \SB2_1_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_12/Component_Function_1/N1  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i1[9] ), .ZN(\SB2_1_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_0/N4  ( .A1(\SB2_1_13/i0[7] ), .A2(
        \SB2_1_13/i0_3 ), .A3(\SB2_1_13/i0_0 ), .ZN(
        \SB2_1_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_13/Component_Function_0/N3  ( .A1(\SB2_1_13/i0[10] ), .A2(
        \SB2_1_13/i0_4 ), .A3(\SB2_1_13/i0_3 ), .ZN(
        \SB2_1_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_13/Component_Function_0/N2  ( .A1(\SB2_1_13/i0[8] ), .A2(
        \SB2_1_13/i0[7] ), .A3(\SB2_1_13/i0[6] ), .ZN(
        \SB2_1_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_13/Component_Function_0/N1  ( .A1(\SB2_1_13/i0[10] ), .A2(
        \SB2_1_13/i0[9] ), .ZN(\SB2_1_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_1/N3  ( .A1(\SB2_1_13/i1_5 ), .A2(
        \SB2_1_13/i0[6] ), .A3(\SB2_1_13/i0[9] ), .ZN(
        \SB2_1_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_13/Component_Function_1/N2  ( .A1(\SB2_1_13/i0_3 ), .A2(
        \SB2_1_13/i1_7 ), .A3(\SB2_1_13/i0[8] ), .ZN(
        \SB2_1_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_13/Component_Function_1/N1  ( .A1(\SB2_1_13/i1[9] ), .A2(
        \SB2_1_13/i0_3 ), .ZN(\SB2_1_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_5/N4  ( .A1(\SB2_1_13/i0[9] ), .A2(
        \SB2_1_13/i0[6] ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_13/Component_Function_5/N1  ( .A1(\SB2_1_13/i0_0 ), .A2(
        \SB2_1_13/i3[0] ), .ZN(\SB2_1_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_0/N4  ( .A1(\SB2_1_14/i0[7] ), .A2(
        \SB2_1_14/i0_3 ), .A3(\SB2_1_14/i0_0 ), .ZN(
        \SB2_1_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_14/Component_Function_0/N3  ( .A1(\SB2_1_14/i0[10] ), .A2(
        \SB2_1_14/i0_4 ), .A3(\SB2_1_14/i0_3 ), .ZN(
        \SB2_1_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_14/Component_Function_0/N2  ( .A1(\SB2_1_14/i0[8] ), .A2(
        \SB2_1_14/i0[7] ), .A3(\SB2_1_14/i0[6] ), .ZN(
        \SB2_1_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_14/Component_Function_0/N1  ( .A1(\SB2_1_14/i0[10] ), .A2(
        \SB2_1_14/i0[9] ), .ZN(\SB2_1_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_1/N3  ( .A1(\SB2_1_14/i1_5 ), .A2(
        \SB2_1_14/i0[6] ), .A3(\SB2_1_14/i0[9] ), .ZN(
        \SB2_1_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_14/Component_Function_1/N2  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i1_7 ), .A3(\SB2_1_14/i0[8] ), .ZN(
        \SB2_1_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_14/Component_Function_1/N1  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_5/N3  ( .A1(\SB2_1_14/i1[9] ), .A2(
        \SB2_1_14/i0_4 ), .A3(\SB2_1_14/i0_3 ), .ZN(
        \SB2_1_14/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_14/Component_Function_5/N1  ( .A1(\SB2_1_14/i0_0 ), .A2(
        \SB2_1_14/i3[0] ), .ZN(\SB2_1_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_15/Component_Function_0/N4  ( .A1(\SB2_1_15/i0[7] ), .A2(
        \SB2_1_15/i0_3 ), .A3(\SB2_1_15/i0_0 ), .ZN(
        \SB2_1_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_15/Component_Function_0/N3  ( .A1(\SB2_1_15/i0[10] ), .A2(
        \SB2_1_15/i0_4 ), .A3(\SB2_1_15/i0_3 ), .ZN(
        \SB2_1_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_15/Component_Function_0/N2  ( .A1(\SB2_1_15/i0[8] ), .A2(
        \SB2_1_15/i0[7] ), .A3(\SB2_1_15/i0[6] ), .ZN(
        \SB2_1_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_15/Component_Function_0/N1  ( .A1(\SB2_1_15/i0[10] ), .A2(
        \SB2_1_15/i0[9] ), .ZN(\SB2_1_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_15/Component_Function_1/N3  ( .A1(\SB2_1_15/i1_5 ), .A2(
        \SB2_1_15/i0[6] ), .A3(\SB2_1_15/i0[9] ), .ZN(
        \SB2_1_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_15/Component_Function_1/N2  ( .A1(\SB2_1_15/i0_3 ), .A2(
        \SB2_1_15/i1_7 ), .A3(\SB2_1_15/i0[8] ), .ZN(
        \SB2_1_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_15/Component_Function_1/N1  ( .A1(\SB2_1_15/i0_3 ), .A2(
        \SB2_1_15/i1[9] ), .ZN(\SB2_1_15/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_15/Component_Function_5/N1  ( .A1(\SB2_1_15/i0_0 ), .A2(
        \SB2_1_15/i3[0] ), .ZN(\SB2_1_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_16/Component_Function_0/N4  ( .A1(\SB2_1_16/i0[7] ), .A2(
        \SB2_1_16/i0_3 ), .A3(\SB2_1_16/i0_0 ), .ZN(
        \SB2_1_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_16/Component_Function_0/N3  ( .A1(\SB2_1_16/i0[10] ), .A2(
        \SB2_1_16/i0_4 ), .A3(\SB2_1_16/i0_3 ), .ZN(
        \SB2_1_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_16/Component_Function_0/N2  ( .A1(\SB2_1_16/i0[8] ), .A2(
        \SB2_1_16/i0[7] ), .A3(\SB2_1_16/i0[6] ), .ZN(
        \SB2_1_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_16/Component_Function_0/N1  ( .A1(\SB2_1_16/i0[10] ), .A2(
        \SB2_1_16/i0[9] ), .ZN(\SB2_1_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_16/Component_Function_1/N3  ( .A1(\SB2_1_16/i1_5 ), .A2(
        \SB2_1_16/i0[6] ), .A3(\SB2_1_16/i0[9] ), .ZN(
        \SB2_1_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_16/Component_Function_1/N2  ( .A1(\SB2_1_16/i0_3 ), .A2(
        \SB2_1_16/i1_7 ), .A3(\SB2_1_16/i0[8] ), .ZN(
        \SB2_1_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_16/Component_Function_1/N1  ( .A1(\SB2_1_16/i0_3 ), .A2(
        \SB2_1_16/i1[9] ), .ZN(\SB2_1_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_16/Component_Function_5/N3  ( .A1(\SB2_1_16/i1[9] ), .A2(
        \SB2_1_16/i0_4 ), .A3(\SB2_1_16/i0_3 ), .ZN(
        \SB2_1_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_16/Component_Function_5/N2  ( .A1(\SB2_1_16/i0_0 ), .A2(
        \SB2_1_16/i0[6] ), .A3(\SB2_1_16/i0[10] ), .ZN(
        \SB2_1_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_16/Component_Function_5/N1  ( .A1(\SB2_1_16/i0_0 ), .A2(
        \SB2_1_16/i3[0] ), .ZN(\SB2_1_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_0/N4  ( .A1(\SB2_1_17/i0[7] ), .A2(
        \SB2_1_17/i0_3 ), .A3(\SB2_1_17/i0_0 ), .ZN(
        \SB2_1_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_17/Component_Function_0/N3  ( .A1(\SB2_1_17/i0[10] ), .A2(
        \SB2_1_17/i0_4 ), .A3(\SB2_1_17/i0_3 ), .ZN(
        \SB2_1_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_17/Component_Function_0/N2  ( .A1(\SB2_1_17/i0[8] ), .A2(
        \SB2_1_17/i0[7] ), .A3(\SB2_1_17/i0[6] ), .ZN(
        \SB2_1_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_17/Component_Function_0/N1  ( .A1(\SB2_1_17/i0[10] ), .A2(
        \SB2_1_17/i0[9] ), .ZN(\SB2_1_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_1/N4  ( .A1(\SB2_1_17/i1_7 ), .A2(
        \SB2_1_17/i0[8] ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_17/Component_Function_1/N3  ( .A1(\SB2_1_17/i1_5 ), .A2(
        \SB2_1_17/i0[6] ), .A3(\SB2_1_17/i0[9] ), .ZN(
        \SB2_1_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_17/Component_Function_1/N2  ( .A1(\SB2_1_17/i0_3 ), .A2(
        \SB2_1_17/i1_7 ), .A3(\SB2_1_17/i0[8] ), .ZN(
        \SB2_1_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_17/Component_Function_1/N1  ( .A1(\SB2_1_17/i1[9] ), .A2(
        \SB2_1_17/i0_3 ), .ZN(\SB2_1_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_17/Component_Function_5/N1  ( .A1(\SB2_1_17/i0_0 ), .A2(
        \SB2_1_17/i3[0] ), .ZN(\SB2_1_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_0/N4  ( .A1(\SB2_1_18/i0[7] ), .A2(
        \SB2_1_18/i0_3 ), .A3(\SB2_1_18/i0_0 ), .ZN(
        \SB2_1_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_18/Component_Function_0/N3  ( .A1(\SB2_1_18/i0[10] ), .A2(
        \SB2_1_18/i0_4 ), .A3(\SB2_1_18/i0_3 ), .ZN(
        \SB2_1_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_18/Component_Function_0/N2  ( .A1(\SB2_1_18/i0[8] ), .A2(
        \SB2_1_18/i0[7] ), .A3(\SB2_1_18/i0[6] ), .ZN(
        \SB2_1_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_18/Component_Function_0/N1  ( .A1(\SB2_1_18/i0[10] ), .A2(
        \SB2_1_18/i0[9] ), .ZN(\SB2_1_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_1/N3  ( .A1(\SB2_1_18/i1_5 ), .A2(
        \SB2_1_18/i0[6] ), .A3(\SB2_1_18/i0[9] ), .ZN(
        \SB2_1_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_18/Component_Function_1/N2  ( .A1(\SB2_1_18/i0_3 ), .A2(
        \SB2_1_18/i1_7 ), .A3(\SB2_1_18/i0[8] ), .ZN(
        \SB2_1_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_18/Component_Function_1/N1  ( .A1(\SB2_1_18/i0_3 ), .A2(
        \SB2_1_18/i1[9] ), .ZN(\SB2_1_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_5/N3  ( .A1(\SB2_1_18/i1[9] ), .A2(
        \SB2_1_18/i0_4 ), .A3(\SB2_1_18/i0_3 ), .ZN(
        \SB2_1_18/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_18/Component_Function_5/N1  ( .A1(\SB2_1_18/i0_0 ), .A2(
        \SB2_1_18/i3[0] ), .ZN(\SB2_1_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_19/Component_Function_0/N4  ( .A1(\SB2_1_19/i0[7] ), .A2(
        \SB2_1_19/i0_3 ), .A3(\SB2_1_19/i0_0 ), .ZN(
        \SB2_1_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_19/Component_Function_0/N3  ( .A1(\SB2_1_19/i0[10] ), .A2(
        \SB2_1_19/i0_4 ), .A3(\SB2_1_19/i0_3 ), .ZN(
        \SB2_1_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_19/Component_Function_0/N2  ( .A1(\SB2_1_19/i0[8] ), .A2(
        \SB2_1_19/i0[7] ), .A3(\SB2_1_19/i0[6] ), .ZN(
        \SB2_1_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_19/Component_Function_0/N1  ( .A1(\SB2_1_19/i0[10] ), .A2(
        \SB2_1_19/i0[9] ), .ZN(\SB2_1_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_19/Component_Function_1/N3  ( .A1(\SB2_1_19/i1_5 ), .A2(
        \SB2_1_19/i0[6] ), .A3(\SB2_1_19/i0[9] ), .ZN(
        \SB2_1_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_19/Component_Function_1/N2  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i1_7 ), .A3(\SB2_1_19/i0[8] ), .ZN(
        \SB2_1_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_19/Component_Function_1/N1  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i1[9] ), .ZN(\SB2_1_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_19/Component_Function_5/N1  ( .A1(\SB2_1_19/i0_0 ), .A2(
        \SB2_1_19/i3[0] ), .ZN(\SB2_1_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_20/Component_Function_0/N3  ( .A1(\SB2_1_20/i0[10] ), .A2(
        \SB2_1_20/i0_4 ), .A3(\SB2_1_20/i0_3 ), .ZN(
        \SB2_1_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_20/Component_Function_0/N2  ( .A1(\SB2_1_20/i0[8] ), .A2(
        \SB2_1_20/i0[7] ), .A3(\SB2_1_20/i0[6] ), .ZN(
        \SB2_1_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_20/Component_Function_0/N1  ( .A1(\SB2_1_20/i0[10] ), .A2(
        \SB2_1_20/i0[9] ), .ZN(\SB2_1_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_20/Component_Function_1/N4  ( .A1(\SB2_1_20/i1_7 ), .A2(
        \SB2_1_20/i0[8] ), .A3(\SB2_1_20/i0_4 ), .ZN(
        \SB2_1_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_20/Component_Function_1/N3  ( .A1(\SB2_1_20/i1_5 ), .A2(
        \SB2_1_20/i0[6] ), .A3(\SB2_1_20/i0[9] ), .ZN(
        \SB2_1_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_20/Component_Function_1/N2  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i1_7 ), .A3(\SB2_1_20/i0[8] ), .ZN(
        \SB2_1_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_20/Component_Function_1/N1  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i1[9] ), .ZN(\SB2_1_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_20/Component_Function_5/N4  ( .A1(\RI3[1][66] ), .A2(
        \SB2_1_20/i0[6] ), .A3(\RI3[1][70] ), .ZN(
        \SB2_1_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_21/Component_Function_0/N4  ( .A1(\SB2_1_21/i0[7] ), .A2(
        \SB2_1_21/i0_3 ), .A3(\SB2_1_21/i0_0 ), .ZN(
        \SB2_1_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_21/Component_Function_0/N3  ( .A1(\SB2_1_21/i0[10] ), .A2(
        \SB2_1_21/i0_4 ), .A3(\SB2_1_21/i0_3 ), .ZN(
        \SB2_1_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_21/Component_Function_0/N2  ( .A1(\SB2_1_21/i0[8] ), .A2(
        \SB2_1_21/i0[7] ), .A3(\SB2_1_21/i0[6] ), .ZN(
        \SB2_1_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_21/Component_Function_0/N1  ( .A1(\SB2_1_21/i0[10] ), .A2(
        \SB2_1_21/i0[9] ), .ZN(\SB2_1_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_21/Component_Function_1/N4  ( .A1(\SB2_1_21/i1_7 ), .A2(
        \SB2_1_21/i0[8] ), .A3(\SB2_1_21/i0_4 ), .ZN(
        \SB2_1_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_21/Component_Function_1/N3  ( .A1(\SB2_1_21/i1_5 ), .A2(
        \SB2_1_21/i0[6] ), .A3(\SB2_1_21/i0[9] ), .ZN(
        \SB2_1_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_21/Component_Function_1/N2  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i1_7 ), .A3(\SB2_1_21/i0[8] ), .ZN(
        \SB2_1_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_21/Component_Function_1/N1  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i1[9] ), .ZN(\SB2_1_21/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_21/Component_Function_5/N1  ( .A1(\SB2_1_21/i0_0 ), .A2(
        \SB2_1_21/i3[0] ), .ZN(\SB2_1_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_0/N4  ( .A1(\SB2_1_22/i0[7] ), .A2(
        \SB2_1_22/i0_3 ), .A3(\SB2_1_22/i0_0 ), .ZN(
        \SB2_1_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_22/Component_Function_0/N3  ( .A1(\SB2_1_22/i0[10] ), .A2(
        \SB2_1_22/i0_4 ), .A3(\SB2_1_22/i0_3 ), .ZN(
        \SB2_1_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_22/Component_Function_0/N2  ( .A1(\SB2_1_22/i0[8] ), .A2(
        \SB2_1_22/i0[7] ), .A3(\SB2_1_22/i0[6] ), .ZN(
        \SB2_1_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_22/Component_Function_0/N1  ( .A1(\SB2_1_22/i0[10] ), .A2(
        \SB2_1_22/i0[9] ), .ZN(\SB2_1_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_1/N4  ( .A1(\SB2_1_22/i1_7 ), .A2(
        \SB2_1_22/i0[8] ), .A3(\SB2_1_22/i0_4 ), .ZN(
        \SB2_1_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_22/Component_Function_1/N3  ( .A1(\SB2_1_22/i1_5 ), .A2(
        \SB2_1_22/i0[6] ), .A3(\SB2_1_22/i0[9] ), .ZN(
        \SB2_1_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_22/Component_Function_1/N2  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i1_7 ), .A3(\SB2_1_22/i0[8] ), .ZN(
        \SB2_1_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_22/Component_Function_1/N1  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i1[9] ), .ZN(\SB2_1_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_5/N4  ( .A1(\SB2_1_22/i0[9] ), .A2(
        \SB2_1_22/i0[6] ), .A3(\SB2_1_22/i0_4 ), .ZN(
        \SB2_1_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_22/Component_Function_5/N2  ( .A1(\SB2_1_22/i0_0 ), .A2(
        \SB2_1_22/i0[6] ), .A3(\SB2_1_22/i0[10] ), .ZN(
        \SB2_1_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_22/Component_Function_5/N1  ( .A1(\SB2_1_22/i0_0 ), .A2(
        \SB2_1_22/i3[0] ), .ZN(\SB2_1_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_0/N4  ( .A1(\SB2_1_23/i0[7] ), .A2(
        \SB2_1_23/i0_3 ), .A3(\SB2_1_23/i0_0 ), .ZN(
        \SB2_1_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_23/Component_Function_0/N3  ( .A1(\SB2_1_23/i0[10] ), .A2(
        \SB2_1_23/i0_4 ), .A3(\SB2_1_23/i0_3 ), .ZN(
        \SB2_1_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_23/Component_Function_0/N2  ( .A1(\SB2_1_23/i0[8] ), .A2(
        \SB2_1_23/i0[7] ), .A3(\SB2_1_23/i0[6] ), .ZN(
        \SB2_1_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_23/Component_Function_0/N1  ( .A1(\SB2_1_23/i0[10] ), .A2(
        \SB2_1_23/i0[9] ), .ZN(\SB2_1_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_1/N4  ( .A1(\SB2_1_23/i1_7 ), .A2(
        \SB2_1_23/i0[8] ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_23/Component_Function_1/N3  ( .A1(\SB2_1_23/i1_5 ), .A2(
        \SB2_1_23/i0[6] ), .A3(\SB2_1_23/i0[9] ), .ZN(
        \SB2_1_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_23/Component_Function_1/N2  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i1_7 ), .A3(\SB2_1_23/i0[8] ), .ZN(
        \SB2_1_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_23/Component_Function_1/N1  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i1[9] ), .ZN(\SB2_1_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_5/N4  ( .A1(\SB2_1_23/i0[9] ), .A2(
        \SB2_1_23/i0[6] ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_23/Component_Function_5/N1  ( .A1(\SB2_1_23/i0_0 ), .A2(
        \SB2_1_23/i3[0] ), .ZN(\SB2_1_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_0/N4  ( .A1(\SB2_1_24/i0[7] ), .A2(
        \SB2_1_24/i0_3 ), .A3(\SB2_1_24/i0_0 ), .ZN(
        \SB2_1_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_24/Component_Function_0/N3  ( .A1(\SB2_1_24/i0[10] ), .A2(
        \SB2_1_24/i0_4 ), .A3(\SB2_1_24/i0_3 ), .ZN(
        \SB2_1_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_24/Component_Function_0/N2  ( .A1(\SB2_1_24/i0[8] ), .A2(
        \SB2_1_24/i0[7] ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_24/Component_Function_0/N1  ( .A1(\SB2_1_24/i0[10] ), .A2(
        \SB2_1_24/i0[9] ), .ZN(\SB2_1_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_1/N4  ( .A1(\SB2_1_24/i1_7 ), .A2(
        \SB2_1_24/i0[8] ), .A3(\SB2_1_24/i0_4 ), .ZN(
        \SB2_1_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_24/Component_Function_1/N3  ( .A1(\SB2_1_24/i1_5 ), .A2(
        \SB2_1_24/i0[6] ), .A3(\SB2_1_24/i0[9] ), .ZN(
        \SB2_1_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_24/Component_Function_1/N2  ( .A1(\SB2_1_24/i0_3 ), .A2(
        \SB2_1_24/i1_7 ), .A3(\SB2_1_24/i0[8] ), .ZN(
        \SB2_1_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_24/Component_Function_1/N1  ( .A1(\SB2_1_24/i0_3 ), .A2(
        \SB2_1_24/i1[9] ), .ZN(\SB2_1_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_0/N3  ( .A1(\SB2_1_25/i0[10] ), .A2(
        \SB2_1_25/i0_4 ), .A3(\SB2_1_25/i0_3 ), .ZN(
        \SB2_1_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_25/Component_Function_0/N2  ( .A1(\SB2_1_25/i0[8] ), .A2(
        \SB2_1_25/i0[7] ), .A3(\SB2_1_25/i0[6] ), .ZN(
        \SB2_1_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_25/Component_Function_0/N1  ( .A1(\SB2_1_25/i0[10] ), .A2(
        \SB2_1_25/i0[9] ), .ZN(\SB2_1_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_1/N3  ( .A1(\SB2_1_25/i1_5 ), .A2(
        \SB2_1_25/i0[6] ), .A3(\SB2_1_25/i0[9] ), .ZN(
        \SB2_1_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_25/Component_Function_1/N2  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i1_7 ), .A3(\SB2_1_25/i0[8] ), .ZN(
        \SB2_1_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_25/Component_Function_1/N1  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i1[9] ), .ZN(\SB2_1_25/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_25/Component_Function_5/N1  ( .A1(\SB2_1_25/i0_0 ), .A2(
        \SB2_1_25/i3[0] ), .ZN(\SB2_1_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_0/N4  ( .A1(\SB2_1_26/i0[7] ), .A2(
        \SB2_1_26/i0_3 ), .A3(\SB2_1_26/i0_0 ), .ZN(
        \SB2_1_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_26/Component_Function_0/N3  ( .A1(\SB2_1_26/i0[10] ), .A2(
        \SB2_1_26/i0_4 ), .A3(\SB2_1_26/i0_3 ), .ZN(
        \SB2_1_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_26/Component_Function_0/N2  ( .A1(\SB2_1_26/i0[8] ), .A2(
        \SB2_1_26/i0[7] ), .A3(\SB2_1_26/i0[6] ), .ZN(
        \SB2_1_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_26/Component_Function_0/N1  ( .A1(\SB2_1_26/i0[10] ), .A2(
        \SB2_1_26/i0[9] ), .ZN(\SB2_1_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_1/N3  ( .A1(\SB2_1_26/i1_5 ), .A2(
        \SB2_1_26/i0[6] ), .A3(\SB2_1_26/i0[9] ), .ZN(
        \SB2_1_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_26/Component_Function_1/N2  ( .A1(\SB2_1_26/i0_3 ), .A2(
        \SB2_1_26/i1_7 ), .A3(\SB2_1_26/i0[8] ), .ZN(
        \SB2_1_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_26/Component_Function_1/N1  ( .A1(\SB2_1_26/i0_3 ), .A2(
        \SB2_1_26/i1[9] ), .ZN(\SB2_1_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_5/N3  ( .A1(\SB2_1_26/i1[9] ), .A2(
        \SB2_1_26/i0_4 ), .A3(\SB2_1_26/i0_3 ), .ZN(
        \SB2_1_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_26/Component_Function_5/N2  ( .A1(\SB2_1_26/i0_0 ), .A2(
        \SB2_1_26/i0[6] ), .A3(\SB2_1_26/i0[10] ), .ZN(
        \SB2_1_26/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_26/Component_Function_5/N1  ( .A1(\SB2_1_26/i0_0 ), .A2(
        \SB2_1_26/i3[0] ), .ZN(\SB2_1_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_0/N4  ( .A1(\SB2_1_27/i0[7] ), .A2(
        \SB2_1_27/i0_3 ), .A3(\SB2_1_27/i0_0 ), .ZN(
        \SB2_1_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_27/Component_Function_0/N3  ( .A1(\SB2_1_27/i0[10] ), .A2(
        \SB2_1_27/i0_4 ), .A3(\SB2_1_27/i0_3 ), .ZN(
        \SB2_1_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_27/Component_Function_0/N2  ( .A1(\SB2_1_27/i0[8] ), .A2(
        \SB2_1_27/i0[7] ), .A3(\SB2_1_27/i0[6] ), .ZN(
        \SB2_1_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_27/Component_Function_0/N1  ( .A1(\SB2_1_27/i0[10] ), .A2(
        \SB2_1_27/i0[9] ), .ZN(\SB2_1_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_1/N4  ( .A1(\SB2_1_27/i0[8] ), .A2(
        \SB2_1_27/i1_7 ), .A3(\SB2_1_27/i0_4 ), .ZN(
        \SB2_1_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_27/Component_Function_1/N3  ( .A1(\SB2_1_27/i1_5 ), .A2(
        \SB2_1_27/i0[6] ), .A3(\SB2_1_27/i0[9] ), .ZN(
        \SB2_1_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_27/Component_Function_1/N2  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i1_7 ), .A3(\SB2_1_27/i0[8] ), .ZN(
        \SB2_1_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_27/Component_Function_1/N1  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i1[9] ), .ZN(\SB2_1_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_5/N4  ( .A1(\SB2_1_27/i0[9] ), .A2(
        \SB2_1_27/i0[6] ), .A3(\SB2_1_27/i0_4 ), .ZN(
        \SB2_1_27/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_27/Component_Function_5/N1  ( .A1(\SB2_1_27/i0_0 ), .A2(
        \SB2_1_27/i3[0] ), .ZN(\SB2_1_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_0/N4  ( .A1(\SB2_1_28/i0[7] ), .A2(
        \SB2_1_28/i0_3 ), .A3(\SB2_1_28/i0_0 ), .ZN(
        \SB2_1_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_28/Component_Function_0/N3  ( .A1(\SB2_1_28/i0[10] ), .A2(
        \SB2_1_28/i0_4 ), .A3(\SB2_1_28/i0_3 ), .ZN(
        \SB2_1_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_28/Component_Function_0/N2  ( .A1(\SB2_1_28/i0[8] ), .A2(
        \SB2_1_28/i0[7] ), .A3(\SB2_1_28/i0[6] ), .ZN(
        \SB2_1_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_28/Component_Function_0/N1  ( .A1(\SB2_1_28/i0[10] ), .A2(
        \SB2_1_28/i0[9] ), .ZN(\SB2_1_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_1/N3  ( .A1(\SB2_1_28/i1_5 ), .A2(
        \SB2_1_28/i0[6] ), .A3(\SB2_1_28/i0[9] ), .ZN(
        \SB2_1_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_28/Component_Function_1/N2  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i1_7 ), .A3(\SB2_1_28/i0[8] ), .ZN(
        \SB2_1_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_28/Component_Function_1/N1  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i1[9] ), .ZN(\SB2_1_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_5/N2  ( .A1(\SB2_1_28/i0_0 ), .A2(
        \SB2_1_28/i0[6] ), .A3(\SB2_1_28/i0[10] ), .ZN(
        \SB2_1_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_29/Component_Function_0/N3  ( .A1(\SB2_1_29/i0[10] ), .A2(
        \SB2_1_29/i0_4 ), .A3(\SB2_1_29/i0_3 ), .ZN(
        \SB2_1_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_29/Component_Function_0/N2  ( .A1(\SB2_1_29/i0[8] ), .A2(
        \SB2_1_29/i0[7] ), .A3(\SB2_1_29/i0[6] ), .ZN(
        \SB2_1_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_29/Component_Function_0/N1  ( .A1(\SB2_1_29/i0[10] ), .A2(
        \SB2_1_29/i0[9] ), .ZN(\SB2_1_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_1/N3  ( .A1(\SB2_1_29/i1_5 ), .A2(
        \SB2_1_29/i0[6] ), .A3(\SB2_1_29/i0[9] ), .ZN(
        \SB2_1_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_29/Component_Function_1/N2  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i1_7 ), .A3(\SB2_1_29/i0[8] ), .ZN(
        \SB2_1_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_29/Component_Function_1/N1  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i1[9] ), .ZN(\SB2_1_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_5/N4  ( .A1(\SB2_1_29/i0[9] ), .A2(
        \SB2_1_29/i0[6] ), .A3(\RI3[1][16] ), .ZN(
        \SB2_1_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_29/Component_Function_5/N3  ( .A1(\SB2_1_29/i1[9] ), .A2(
        \SB2_1_29/i0_4 ), .A3(\SB2_1_29/i0_3 ), .ZN(
        \SB2_1_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_29/Component_Function_5/N2  ( .A1(\SB2_1_29/i0_0 ), .A2(
        \SB2_1_29/i0[6] ), .A3(\SB2_1_29/i0[10] ), .ZN(
        \SB2_1_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_30/Component_Function_0/N4  ( .A1(\SB2_1_30/i0[7] ), .A2(
        \SB2_1_30/i0_3 ), .A3(\SB2_1_30/i0_0 ), .ZN(
        \SB2_1_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_30/Component_Function_0/N3  ( .A1(\SB2_1_30/i0[10] ), .A2(
        \SB2_1_30/i0_4 ), .A3(\SB2_1_30/i0_3 ), .ZN(
        \SB2_1_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_30/Component_Function_0/N2  ( .A1(\SB2_1_30/i0[8] ), .A2(
        \SB2_1_30/i0[7] ), .A3(\SB2_1_30/i0[6] ), .ZN(
        \SB2_1_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_30/Component_Function_0/N1  ( .A1(\SB2_1_30/i0[10] ), .A2(
        \SB2_1_30/i0[9] ), .ZN(\SB2_1_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_1/N3  ( .A1(\SB2_1_30/i1_5 ), .A2(
        \SB2_1_30/i0[6] ), .A3(\SB2_1_30/i0[9] ), .ZN(
        \SB2_1_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_30/Component_Function_1/N2  ( .A1(\SB2_1_30/i0_3 ), .A2(
        \SB2_1_30/i1_7 ), .A3(\SB2_1_30/i0[8] ), .ZN(
        \SB2_1_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_30/Component_Function_1/N1  ( .A1(\SB2_1_30/i0_3 ), .A2(
        \SB2_1_30/i1[9] ), .ZN(\SB2_1_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_5/N3  ( .A1(\SB2_1_30/i1[9] ), .A2(
        \SB2_1_30/i0_4 ), .A3(\SB2_1_30/i0_3 ), .ZN(
        \SB2_1_30/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_30/Component_Function_5/N1  ( .A1(\SB2_1_30/i0_0 ), .A2(
        \SB2_1_30/i3[0] ), .ZN(\SB2_1_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_0/N3  ( .A1(\SB2_1_31/i0[10] ), .A2(
        \SB2_1_31/i0_4 ), .A3(\SB2_1_31/i0_3 ), .ZN(
        \SB2_1_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_31/Component_Function_0/N2  ( .A1(\SB2_1_31/i0[8] ), .A2(
        \SB2_1_31/i0[7] ), .A3(\SB2_1_31/i0[6] ), .ZN(
        \SB2_1_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_31/Component_Function_0/N1  ( .A1(\SB2_1_31/i0[10] ), .A2(
        \SB2_1_31/i0[9] ), .ZN(\SB2_1_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_1/N3  ( .A1(\SB2_1_31/i1_5 ), .A2(
        \SB2_1_31/i0[6] ), .A3(\SB2_1_31/i0[9] ), .ZN(
        \SB2_1_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_31/Component_Function_1/N2  ( .A1(\SB2_1_31/i0_3 ), .A2(
        \SB2_1_31/i1_7 ), .A3(\SB2_1_31/i0[8] ), .ZN(
        \SB2_1_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_31/Component_Function_1/N1  ( .A1(\SB2_1_31/i0_3 ), .A2(
        \SB2_1_31/i1[9] ), .ZN(\SB2_1_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_5/N4  ( .A1(\SB2_1_31/i0[9] ), .A2(
        \SB2_1_31/i0[6] ), .A3(\SB2_1_31/i0_4 ), .ZN(
        \SB2_1_31/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_31/Component_Function_5/N1  ( .A1(\SB2_1_31/i0_0 ), .A2(
        \SB2_1_31/i3[0] ), .ZN(\SB2_1_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_0/N4  ( .A1(\SB1_2_0/i0[7] ), .A2(
        \SB1_2_0/i0_3 ), .A3(\SB1_2_0/i0_0 ), .ZN(
        \SB1_2_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_0/Component_Function_0/N2  ( .A1(\SB1_2_0/i0[8] ), .A2(
        \SB1_2_0/i0[7] ), .A3(\SB1_2_0/i0[6] ), .ZN(
        \SB1_2_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_0/Component_Function_0/N1  ( .A1(\SB1_2_0/i0[10] ), .A2(
        \SB1_2_0/i0[9] ), .ZN(\SB1_2_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_1/N4  ( .A1(\SB1_2_0/i1_7 ), .A2(
        \SB1_2_0/i0[8] ), .A3(\SB1_2_0/i0_4 ), .ZN(
        \SB1_2_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_0/Component_Function_1/N3  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[6] ), .A3(\SB1_2_0/i0[9] ), .ZN(
        \SB1_2_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_0/Component_Function_1/N2  ( .A1(\SB1_2_0/i0_3 ), .A2(
        \SB1_2_0/i1_7 ), .A3(\SB1_2_0/i0[8] ), .ZN(
        \SB1_2_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_0/Component_Function_1/N1  ( .A1(\SB1_2_0/i0_3 ), .A2(
        \SB1_2_0/i1[9] ), .ZN(\SB1_2_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_5/N4  ( .A1(\SB1_2_0/i0[9] ), .A2(
        \SB1_2_0/i0[6] ), .A3(\SB1_2_0/i0_4 ), .ZN(
        \SB1_2_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_0/Component_Function_5/N2  ( .A1(\SB1_2_0/i0_0 ), .A2(
        \SB1_2_0/i0[6] ), .A3(\SB1_2_0/i0[10] ), .ZN(
        \SB1_2_0/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_0/Component_Function_5/N1  ( .A1(\SB1_2_0/i0_0 ), .A2(
        \SB1_2_0/i3[0] ), .ZN(\SB1_2_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_0/N4  ( .A1(\SB1_2_1/i0[7] ), .A2(
        \SB1_2_1/i0_3 ), .A3(\SB1_2_1/i0_0 ), .ZN(
        \SB1_2_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_1/Component_Function_0/N3  ( .A1(\SB1_2_1/i0[10] ), .A2(
        \SB1_2_1/i0_4 ), .A3(\SB1_2_1/i0_3 ), .ZN(
        \SB1_2_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_1/Component_Function_0/N2  ( .A1(\SB1_2_1/i0[8] ), .A2(
        \SB1_2_1/i0[7] ), .A3(\SB1_2_1/i0[6] ), .ZN(
        \SB1_2_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_1/Component_Function_0/N1  ( .A1(\SB1_2_1/i0[10] ), .A2(
        \SB1_2_1/i0[9] ), .ZN(\SB1_2_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_1/N4  ( .A1(\SB1_2_1/i1_7 ), .A2(
        \SB1_2_1/i0[8] ), .A3(\SB1_2_1/i0_4 ), .ZN(
        \SB1_2_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_1/Component_Function_1/N3  ( .A1(\SB1_2_1/i1_5 ), .A2(
        \SB1_2_1/i0[6] ), .A3(\SB1_2_1/i0[9] ), .ZN(
        \SB1_2_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_1/Component_Function_1/N2  ( .A1(\SB1_2_1/i0_3 ), .A2(
        \SB1_2_1/i1_7 ), .A3(\SB1_2_1/i0[8] ), .ZN(
        \SB1_2_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_1/Component_Function_1/N1  ( .A1(\SB1_2_1/i0_3 ), .A2(
        \SB1_2_1/i1[9] ), .ZN(\SB1_2_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_5/N4  ( .A1(\SB1_2_1/i0[9] ), .A2(
        \SB1_2_1/i0[6] ), .A3(\SB1_2_1/i0_4 ), .ZN(
        \SB1_2_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_1/Component_Function_5/N2  ( .A1(\SB1_2_1/i0_0 ), .A2(
        \SB1_2_1/i0[6] ), .A3(\SB1_2_1/i0[10] ), .ZN(
        \SB1_2_1/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_1/Component_Function_5/N1  ( .A1(\SB1_2_1/i0_0 ), .A2(
        \SB1_2_1/i3[0] ), .ZN(\SB1_2_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_0/N4  ( .A1(\SB1_2_2/i0[7] ), .A2(n1648), .A3(\SB1_2_2/i0_0 ), .ZN(\SB1_2_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_0/N2  ( .A1(\SB1_2_2/i0[8] ), .A2(
        \SB1_2_2/i0[7] ), .A3(\SB1_2_2/i0[6] ), .ZN(
        \SB1_2_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_2/Component_Function_0/N1  ( .A1(\SB1_2_2/i0[10] ), .A2(
        \SB1_2_2/i0[9] ), .ZN(\SB1_2_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_1/N4  ( .A1(\SB1_2_2/i1_7 ), .A2(
        \SB1_2_2/i0[8] ), .A3(\SB1_2_2/i0_4 ), .ZN(
        \SB1_2_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_1/N2  ( .A1(n1648), .A2(\SB1_2_2/i1_7 ), 
        .A3(\SB1_2_2/i0[8] ), .ZN(\SB1_2_2/Component_Function_1/NAND4_in[1] )
         );
  NAND2_X1 \SB1_2_2/Component_Function_1/N1  ( .A1(n1648), .A2(\SB1_2_2/i1[9] ), .ZN(\SB1_2_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_5/N4  ( .A1(\SB1_2_2/i0[9] ), .A2(
        \SB1_2_2/i0[6] ), .A3(\SB1_2_2/i0_4 ), .ZN(
        \SB1_2_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_5/N2  ( .A1(\SB1_2_2/i0_0 ), .A2(
        \SB1_2_2/i0[6] ), .A3(\SB1_2_2/i0[10] ), .ZN(
        \SB1_2_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_2/Component_Function_5/N1  ( .A1(\SB1_2_2/i0_0 ), .A2(
        \SB1_2_2/i3[0] ), .ZN(\SB1_2_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_0/N4  ( .A1(\SB1_2_3/i0[7] ), .A2(
        \SB1_2_3/i0_3 ), .A3(\SB1_2_3/i0_0 ), .ZN(
        \SB1_2_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_3/Component_Function_0/N2  ( .A1(\SB1_2_3/i0[8] ), .A2(
        \SB1_2_3/i0[7] ), .A3(\SB1_2_3/i0[6] ), .ZN(
        \SB1_2_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_3/Component_Function_0/N1  ( .A1(\SB1_2_3/i0[10] ), .A2(
        \SB1_2_3/i0[9] ), .ZN(\SB1_2_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_1/N4  ( .A1(\SB1_2_3/i1_7 ), .A2(
        \SB1_2_3/i0[8] ), .A3(\SB1_2_3/i0_4 ), .ZN(
        \SB1_2_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_3/Component_Function_1/N3  ( .A1(\SB1_2_3/i1_5 ), .A2(
        \SB1_2_3/i0[6] ), .A3(\SB1_2_3/i0[9] ), .ZN(
        \SB1_2_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_3/Component_Function_1/N2  ( .A1(\SB1_2_3/i0_3 ), .A2(
        \SB1_2_3/i1_7 ), .A3(\SB1_2_3/i0[8] ), .ZN(
        \SB1_2_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_3/Component_Function_1/N1  ( .A1(\SB1_2_3/i0_3 ), .A2(
        \SB1_2_3/i1[9] ), .ZN(\SB1_2_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_5/N4  ( .A1(\SB1_2_3/i0[9] ), .A2(
        \SB1_2_3/i0[6] ), .A3(\SB1_2_3/i0_4 ), .ZN(
        \SB1_2_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_3/Component_Function_5/N2  ( .A1(\SB1_2_3/i0_0 ), .A2(
        \SB1_2_3/i0[6] ), .A3(\SB1_2_3/i0[10] ), .ZN(
        \SB1_2_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_3/Component_Function_5/N1  ( .A1(\SB1_2_3/i0_0 ), .A2(
        \SB1_2_3/i3[0] ), .ZN(\SB1_2_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_0/N4  ( .A1(\SB1_2_4/i0[7] ), .A2(
        \SB1_2_4/i0_3 ), .A3(\SB1_2_4/i0_0 ), .ZN(
        \SB1_2_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_4/Component_Function_0/N2  ( .A1(\SB1_2_4/i0[8] ), .A2(
        \SB1_2_4/i0[7] ), .A3(\SB1_2_4/i0[6] ), .ZN(
        \SB1_2_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_4/Component_Function_0/N1  ( .A1(\SB1_2_4/i0[10] ), .A2(
        \SB1_2_4/i0[9] ), .ZN(\SB1_2_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_1/N4  ( .A1(\SB1_2_4/i1_7 ), .A2(
        \SB1_2_4/i0[8] ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_4/Component_Function_1/N3  ( .A1(\SB1_2_4/i1_5 ), .A2(
        \SB1_2_4/i0[6] ), .A3(\SB1_2_4/i0[9] ), .ZN(
        \SB1_2_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_4/Component_Function_1/N2  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i1_7 ), .A3(\SB1_2_4/i0[8] ), .ZN(
        \SB1_2_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_4/Component_Function_1/N1  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i1[9] ), .ZN(\SB1_2_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_5/N4  ( .A1(\SB1_2_4/i0[9] ), .A2(
        \SB1_2_4/i0[6] ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_4/Component_Function_5/N2  ( .A1(\SB1_2_4/i0_0 ), .A2(
        \SB1_2_4/i0[6] ), .A3(\SB1_2_4/i0[10] ), .ZN(
        \SB1_2_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_4/Component_Function_5/N1  ( .A1(\SB1_2_4/i0_0 ), .A2(
        \SB1_2_4/i3[0] ), .ZN(\SB1_2_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_0/N4  ( .A1(\SB1_2_5/i0[7] ), .A2(
        \SB1_2_5/i0_3 ), .A3(\SB1_2_5/i0_0 ), .ZN(
        \SB1_2_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_5/Component_Function_0/N3  ( .A1(\SB1_2_5/i0[10] ), .A2(
        \SB1_2_5/i0_4 ), .A3(\SB1_2_5/i0_3 ), .ZN(
        \SB1_2_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_5/Component_Function_0/N2  ( .A1(\SB1_2_5/i0[8] ), .A2(
        \SB1_2_5/i0[7] ), .A3(\SB1_2_5/i0[6] ), .ZN(
        \SB1_2_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_5/Component_Function_0/N1  ( .A1(\SB1_2_5/i0[10] ), .A2(
        \SB1_2_5/i0[9] ), .ZN(\SB1_2_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_1/N4  ( .A1(\SB1_2_5/i1_7 ), .A2(
        \SB1_2_5/i0[8] ), .A3(\SB1_2_5/i0_4 ), .ZN(
        \SB1_2_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_5/Component_Function_1/N3  ( .A1(\SB1_2_5/i1_5 ), .A2(
        \SB1_2_5/i0[6] ), .A3(\SB1_2_5/i0[9] ), .ZN(
        \SB1_2_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_5/Component_Function_1/N2  ( .A1(\SB1_2_5/i0_3 ), .A2(
        \SB1_2_5/i1_7 ), .A3(\SB1_2_5/i0[8] ), .ZN(
        \SB1_2_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_5/Component_Function_1/N1  ( .A1(\SB1_2_5/i0_3 ), .A2(
        \SB1_2_5/i1[9] ), .ZN(\SB1_2_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_5/N2  ( .A1(\SB1_2_5/i0_0 ), .A2(
        \SB1_2_5/i0[6] ), .A3(\SB1_2_5/i0[10] ), .ZN(
        \SB1_2_5/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_5/Component_Function_5/N1  ( .A1(\SB1_2_5/i0_0 ), .A2(
        \SB1_2_5/i3[0] ), .ZN(\SB1_2_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_0/N4  ( .A1(\SB1_2_6/i0[7] ), .A2(
        \SB1_2_6/i0_3 ), .A3(\SB1_2_6/i0_0 ), .ZN(
        \SB1_2_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_6/Component_Function_0/N3  ( .A1(\SB1_2_6/i0[10] ), .A2(
        \SB1_2_6/i0_4 ), .A3(\SB1_2_6/i0_3 ), .ZN(
        \SB1_2_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_6/Component_Function_0/N2  ( .A1(\SB1_2_6/i0[8] ), .A2(
        \SB1_2_6/i0[7] ), .A3(\SB1_2_6/i0[6] ), .ZN(
        \SB1_2_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_6/Component_Function_0/N1  ( .A1(\SB1_2_6/i0[10] ), .A2(
        \SB1_2_6/i0[9] ), .ZN(\SB1_2_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_1/N4  ( .A1(\SB1_2_6/i1_7 ), .A2(
        \SB1_2_6/i0[8] ), .A3(\SB1_2_6/i0_4 ), .ZN(
        \SB1_2_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_6/Component_Function_1/N3  ( .A1(\SB1_2_6/i1_5 ), .A2(
        \SB1_2_6/i0[6] ), .A3(\SB1_2_6/i0[9] ), .ZN(
        \SB1_2_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_6/Component_Function_1/N2  ( .A1(\SB1_2_6/i0_3 ), .A2(
        \SB1_2_6/i1_7 ), .A3(\SB1_2_6/i0[8] ), .ZN(
        \SB1_2_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_6/Component_Function_1/N1  ( .A1(\SB1_2_6/i0_3 ), .A2(
        \SB1_2_6/i1[9] ), .ZN(\SB1_2_6/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_6/Component_Function_5/N1  ( .A1(\SB1_2_6/i0_0 ), .A2(
        \SB1_2_6/i3[0] ), .ZN(\SB1_2_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_0/N4  ( .A1(\SB1_2_7/i0[7] ), .A2(
        \SB1_2_7/i0_3 ), .A3(\SB1_2_7/i0_0 ), .ZN(
        \SB1_2_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_7/Component_Function_0/N3  ( .A1(\SB1_2_7/i0[10] ), .A2(
        \SB1_2_7/i0_4 ), .A3(\SB1_2_7/i0_3 ), .ZN(
        \SB1_2_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_7/Component_Function_0/N2  ( .A1(\SB1_2_7/i0[8] ), .A2(
        \SB1_2_7/i0[7] ), .A3(\SB1_2_7/i0[6] ), .ZN(
        \SB1_2_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_7/Component_Function_0/N1  ( .A1(\SB1_2_7/i0[10] ), .A2(
        \SB1_2_7/i0[9] ), .ZN(\SB1_2_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_1/N4  ( .A1(\SB1_2_7/i1_7 ), .A2(
        \SB1_2_7/i0[8] ), .A3(\SB1_2_7/i0_4 ), .ZN(
        \SB1_2_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_7/Component_Function_1/N3  ( .A1(\SB1_2_7/i1_5 ), .A2(
        \SB1_2_7/i0[6] ), .A3(\SB1_2_7/i0[9] ), .ZN(
        \SB1_2_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_7/Component_Function_1/N2  ( .A1(\SB1_2_7/i0_3 ), .A2(
        \SB1_2_7/i1_7 ), .A3(\SB1_2_7/i0[8] ), .ZN(
        \SB1_2_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_7/Component_Function_1/N1  ( .A1(\SB1_2_7/i0_3 ), .A2(
        \SB1_2_7/i1[9] ), .ZN(\SB1_2_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_5/N4  ( .A1(\SB1_2_7/i0[9] ), .A2(
        \SB1_2_7/i0[6] ), .A3(\SB1_2_7/i0_4 ), .ZN(
        \SB1_2_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_7/Component_Function_5/N2  ( .A1(\SB1_2_7/i0_0 ), .A2(
        \SB1_2_7/i0[6] ), .A3(\SB1_2_7/i0[10] ), .ZN(
        \SB1_2_7/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_7/Component_Function_5/N1  ( .A1(\SB1_2_7/i0_0 ), .A2(
        \SB1_2_7/i3[0] ), .ZN(\SB1_2_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_0/N3  ( .A1(\SB1_2_8/i0[10] ), .A2(
        \SB1_2_8/i0_4 ), .A3(\SB1_2_8/i0_3 ), .ZN(
        \SB1_2_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_8/Component_Function_0/N2  ( .A1(\SB1_2_8/i0[8] ), .A2(
        \SB1_2_8/i0[7] ), .A3(\SB1_2_8/i0[6] ), .ZN(
        \SB1_2_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_8/Component_Function_0/N1  ( .A1(\SB1_2_8/i0[10] ), .A2(
        \SB1_2_8/i0[9] ), .ZN(\SB1_2_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_1/N4  ( .A1(\SB1_2_8/i1_7 ), .A2(
        \SB1_2_8/i0[8] ), .A3(\SB1_2_8/i0_4 ), .ZN(
        \SB1_2_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_8/Component_Function_1/N3  ( .A1(\SB1_2_8/i1_5 ), .A2(
        \SB1_2_8/i0[6] ), .A3(\SB1_2_8/i0[9] ), .ZN(
        \SB1_2_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_8/Component_Function_1/N2  ( .A1(\SB1_2_8/i0_3 ), .A2(
        \SB1_2_8/i1_7 ), .A3(\SB1_2_8/i0[8] ), .ZN(
        \SB1_2_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_8/Component_Function_1/N1  ( .A1(\SB1_2_8/i0_3 ), .A2(
        \SB1_2_8/i1[9] ), .ZN(\SB1_2_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_5/N2  ( .A1(\SB1_2_8/i0_0 ), .A2(
        \SB1_2_8/i0[6] ), .A3(\SB1_2_8/i0[10] ), .ZN(
        \SB1_2_8/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_8/Component_Function_5/N1  ( .A1(\SB1_2_8/i0_0 ), .A2(
        \SB1_2_8/i3[0] ), .ZN(\SB1_2_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_0/N4  ( .A1(\SB1_2_9/i0[7] ), .A2(
        \SB1_2_9/i0_0 ), .A3(n1657), .ZN(
        \SB1_2_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_9/Component_Function_0/N3  ( .A1(\SB1_2_9/i0[10] ), .A2(
        \SB1_2_9/i0_4 ), .A3(n1657), .ZN(
        \SB1_2_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_9/Component_Function_0/N2  ( .A1(\SB1_2_9/i0[8] ), .A2(
        \SB1_2_9/i0[7] ), .A3(\SB1_2_9/i0[6] ), .ZN(
        \SB1_2_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_9/Component_Function_0/N1  ( .A1(\SB1_2_9/i0[10] ), .A2(
        \SB1_2_9/i0[9] ), .ZN(\SB1_2_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_1/N4  ( .A1(\SB1_2_9/i1_7 ), .A2(
        \SB1_2_9/i0[8] ), .A3(\SB1_2_9/i0_4 ), .ZN(
        \SB1_2_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_9/Component_Function_1/N3  ( .A1(\SB1_2_9/i1_5 ), .A2(
        \SB1_2_9/i0[6] ), .A3(\SB1_2_9/i0[9] ), .ZN(
        \SB1_2_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_9/Component_Function_1/N2  ( .A1(n1657), .A2(\SB1_2_9/i1_7 ), 
        .A3(\SB1_2_9/i0[8] ), .ZN(\SB1_2_9/Component_Function_1/NAND4_in[1] )
         );
  NAND2_X1 \SB1_2_9/Component_Function_1/N1  ( .A1(n1657), .A2(\SB1_2_9/i1[9] ), .ZN(\SB1_2_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_5/N4  ( .A1(\SB1_2_9/i0[9] ), .A2(
        \SB1_2_9/i0[6] ), .A3(\SB1_2_9/i0_4 ), .ZN(
        \SB1_2_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_9/Component_Function_5/N2  ( .A1(\SB1_2_9/i0_0 ), .A2(
        \SB1_2_9/i0[6] ), .A3(\SB1_2_9/i0[10] ), .ZN(
        \SB1_2_9/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_9/Component_Function_5/N1  ( .A1(\SB1_2_9/i0_0 ), .A2(
        \SB1_2_9/i3[0] ), .ZN(\SB1_2_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_0/N4  ( .A1(\SB1_2_10/i0[7] ), .A2(
        \SB1_2_10/i0_3 ), .A3(\SB1_2_10/i0_0 ), .ZN(
        \SB1_2_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_10/Component_Function_0/N2  ( .A1(\SB1_2_10/i0[8] ), .A2(
        \SB1_2_10/i0[7] ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_10/Component_Function_0/N1  ( .A1(\SB1_2_10/i0[10] ), .A2(
        \SB1_2_10/i0[9] ), .ZN(\SB1_2_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_1/N4  ( .A1(\SB1_2_10/i1_7 ), .A2(
        \SB1_2_10/i0[8] ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_10/Component_Function_1/N3  ( .A1(\SB1_2_10/i1_5 ), .A2(
        \SB1_2_10/i0[6] ), .A3(\SB1_2_10/i0[9] ), .ZN(
        \SB1_2_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_10/Component_Function_1/N2  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i1_7 ), .A3(\SB1_2_10/i0[8] ), .ZN(
        \SB1_2_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_10/Component_Function_1/N1  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i1[9] ), .ZN(\SB1_2_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_5/N4  ( .A1(\SB1_2_10/i0[9] ), .A2(
        \SB1_2_10/i0[6] ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_10/Component_Function_5/N2  ( .A1(\SB1_2_10/i0_0 ), .A2(
        \SB1_2_10/i0[6] ), .A3(\SB1_2_10/i0[10] ), .ZN(
        \SB1_2_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_10/Component_Function_5/N1  ( .A1(\SB1_2_10/i0_0 ), .A2(
        \SB1_2_10/i3[0] ), .ZN(\SB1_2_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_0/N4  ( .A1(\SB1_2_11/i0[7] ), .A2(
        \SB1_2_11/i0_3 ), .A3(\SB1_2_11/i0_0 ), .ZN(
        \SB1_2_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_11/Component_Function_0/N3  ( .A1(\SB1_2_11/i0[10] ), .A2(
        \SB1_2_11/i0_4 ), .A3(\SB1_2_11/i0_3 ), .ZN(
        \SB1_2_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_11/Component_Function_0/N2  ( .A1(\SB1_2_11/i0[8] ), .A2(
        \SB1_2_11/i0[7] ), .A3(\SB1_2_11/i0[6] ), .ZN(
        \SB1_2_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_11/Component_Function_0/N1  ( .A1(\SB1_2_11/i0[10] ), .A2(
        \SB1_2_11/i0[9] ), .ZN(\SB1_2_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_1/N4  ( .A1(\SB1_2_11/i1_7 ), .A2(
        \SB1_2_11/i0[8] ), .A3(\SB1_2_11/i0_4 ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_11/Component_Function_1/N3  ( .A1(\SB1_2_11/i1_5 ), .A2(
        \SB1_2_11/i0[6] ), .A3(\SB1_2_11/i0[9] ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_11/Component_Function_1/N2  ( .A1(\SB1_2_11/i0_3 ), .A2(
        \SB1_2_11/i1_7 ), .A3(\SB1_2_11/i0[8] ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_11/Component_Function_1/N1  ( .A1(\SB1_2_11/i0_3 ), .A2(
        \SB1_2_11/i1[9] ), .ZN(\SB1_2_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_5/N4  ( .A1(\SB1_2_11/i0[9] ), .A2(
        \SB1_2_11/i0[6] ), .A3(\SB1_2_11/i0_4 ), .ZN(
        \SB1_2_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_11/Component_Function_5/N2  ( .A1(\SB1_2_11/i0_0 ), .A2(
        \SB1_2_11/i0[6] ), .A3(\SB1_2_11/i0[10] ), .ZN(
        \SB1_2_11/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_11/Component_Function_5/N1  ( .A1(\SB1_2_11/i0_0 ), .A2(
        \SB1_2_11/i3[0] ), .ZN(\SB1_2_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_0/N2  ( .A1(\SB1_2_12/i0[8] ), .A2(
        \SB1_2_12/i0[7] ), .A3(\SB1_2_12/i0[6] ), .ZN(
        \SB1_2_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_12/Component_Function_0/N1  ( .A1(\SB1_2_12/i0[10] ), .A2(
        \SB1_2_12/i0[9] ), .ZN(\SB1_2_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_1/N4  ( .A1(\SB1_2_12/i1_7 ), .A2(
        \SB1_2_12/i0[8] ), .A3(\SB1_2_12/i0_4 ), .ZN(
        \SB1_2_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_12/Component_Function_1/N3  ( .A1(\SB1_2_12/i1_5 ), .A2(
        \SB1_2_12/i0[6] ), .A3(\SB1_2_12/i0[9] ), .ZN(
        \SB1_2_12/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_12/Component_Function_1/N1  ( .A1(\SB1_2_12/i0_3 ), .A2(
        \SB1_2_12/i1[9] ), .ZN(\SB1_2_12/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_12/Component_Function_5/N1  ( .A1(\SB1_2_12/i0_0 ), .A2(
        \SB1_2_12/i3[0] ), .ZN(\SB1_2_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_0/N4  ( .A1(\SB1_2_13/i0[7] ), .A2(
        \SB1_2_13/i0_3 ), .A3(\SB1_2_13/i0_0 ), .ZN(
        \SB1_2_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_13/Component_Function_0/N3  ( .A1(\SB1_2_13/i0[10] ), .A2(
        \SB1_2_13/i0_4 ), .A3(\SB1_2_13/i0_3 ), .ZN(
        \SB1_2_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_13/Component_Function_0/N2  ( .A1(\SB1_2_13/i0[8] ), .A2(
        \SB1_2_13/i0[7] ), .A3(\SB1_2_13/i0[6] ), .ZN(
        \SB1_2_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_13/Component_Function_0/N1  ( .A1(\SB1_2_13/i0[10] ), .A2(
        \SB1_2_13/i0[9] ), .ZN(\SB1_2_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_1/N3  ( .A1(\SB1_2_13/i1_5 ), .A2(
        \SB1_2_13/i0[6] ), .A3(\SB1_2_13/i0[9] ), .ZN(
        \SB1_2_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_13/Component_Function_1/N2  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i1_7 ), .A3(\SB1_2_13/i0[8] ), .ZN(
        \SB1_2_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_13/Component_Function_1/N1  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i1[9] ), .ZN(\SB1_2_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_5/N4  ( .A1(\SB1_2_13/i0[9] ), .A2(
        \SB1_2_13/i0[6] ), .A3(\SB1_2_13/i0_4 ), .ZN(
        \SB1_2_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_13/Component_Function_5/N2  ( .A1(\SB1_2_13/i0_0 ), .A2(
        \SB1_2_13/i0[6] ), .A3(\SB1_2_13/i0[10] ), .ZN(
        \SB1_2_13/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_13/Component_Function_5/N1  ( .A1(\SB1_2_13/i0_0 ), .A2(
        \SB1_2_13/i3[0] ), .ZN(\SB1_2_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_0/N4  ( .A1(\SB1_2_14/i0[7] ), .A2(
        \SB1_2_14/i0_3 ), .A3(\SB1_2_14/i0_0 ), .ZN(
        \SB1_2_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_14/Component_Function_0/N2  ( .A1(\SB1_2_14/i0[8] ), .A2(
        \SB1_2_14/i0[7] ), .A3(\SB1_2_14/i0[6] ), .ZN(
        \SB1_2_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_14/Component_Function_0/N1  ( .A1(\SB1_2_14/i0[10] ), .A2(
        \SB1_2_14/i0[9] ), .ZN(\SB1_2_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_1/N4  ( .A1(\SB1_2_14/i1_7 ), .A2(
        \SB1_2_14/i0[8] ), .A3(\SB1_2_14/i0_4 ), .ZN(
        \SB1_2_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_14/Component_Function_1/N3  ( .A1(\SB1_2_14/i1_5 ), .A2(
        \SB1_2_14/i0[6] ), .A3(\SB1_2_14/i0[9] ), .ZN(
        \SB1_2_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_14/Component_Function_1/N2  ( .A1(\SB1_2_14/i0_3 ), .A2(
        \SB1_2_14/i1_7 ), .A3(\SB1_2_14/i0[8] ), .ZN(
        \SB1_2_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_14/Component_Function_1/N1  ( .A1(\SB1_2_14/i0_3 ), .A2(
        \SB1_2_14/i1[9] ), .ZN(\SB1_2_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_5/N4  ( .A1(\SB1_2_14/i0[9] ), .A2(
        \SB1_2_14/i0[6] ), .A3(\SB1_2_14/i0_4 ), .ZN(
        \SB1_2_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_14/Component_Function_5/N2  ( .A1(\SB1_2_14/i0_0 ), .A2(
        \SB1_2_14/i0[6] ), .A3(\SB1_2_14/i0[10] ), .ZN(
        \SB1_2_14/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_14/Component_Function_5/N1  ( .A1(\SB1_2_14/i0_0 ), .A2(
        \SB1_2_14/i3[0] ), .ZN(\SB1_2_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_0/N3  ( .A1(\SB1_2_15/i0[10] ), .A2(
        \SB1_2_15/i0_4 ), .A3(\SB1_2_15/i0_3 ), .ZN(
        \SB1_2_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_15/Component_Function_0/N2  ( .A1(\SB1_2_15/i0[8] ), .A2(
        \SB1_2_15/i0[7] ), .A3(\SB1_2_15/i0[6] ), .ZN(
        \SB1_2_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_15/Component_Function_0/N1  ( .A1(\SB1_2_15/i0[10] ), .A2(
        \SB1_2_15/i0[9] ), .ZN(\SB1_2_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_1/N4  ( .A1(\SB1_2_15/i1_7 ), .A2(
        \SB1_2_15/i0[8] ), .A3(\SB1_2_15/i0_4 ), .ZN(
        \SB1_2_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_15/Component_Function_1/N3  ( .A1(\SB1_2_15/i1_5 ), .A2(
        \SB1_2_15/i0[6] ), .A3(\SB1_2_15/i0[9] ), .ZN(
        \SB1_2_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_15/Component_Function_1/N2  ( .A1(\SB1_2_15/i0_3 ), .A2(
        \SB1_2_15/i1_7 ), .A3(\SB1_2_15/i0[8] ), .ZN(
        \SB1_2_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_15/Component_Function_1/N1  ( .A1(\SB1_2_15/i0_3 ), .A2(
        \SB1_2_15/i1[9] ), .ZN(\SB1_2_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_5/N4  ( .A1(\SB1_2_15/i0[9] ), .A2(
        \SB1_2_15/i0[6] ), .A3(\SB1_2_15/i0_4 ), .ZN(
        \SB1_2_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_15/Component_Function_5/N2  ( .A1(\SB1_2_15/i0_0 ), .A2(
        \SB1_2_15/i0[6] ), .A3(\SB1_2_15/i0[10] ), .ZN(
        \SB1_2_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_15/Component_Function_5/N1  ( .A1(\SB1_2_15/i0_0 ), .A2(
        \SB1_2_15/i3[0] ), .ZN(\SB1_2_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_0/N4  ( .A1(\SB1_2_16/i0[7] ), .A2(
        \SB1_2_16/i0_3 ), .A3(\SB1_2_16/i0_0 ), .ZN(
        \SB1_2_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_16/Component_Function_0/N3  ( .A1(\SB1_2_16/i0[10] ), .A2(
        \SB1_2_16/i0_4 ), .A3(\SB1_2_16/i0_3 ), .ZN(
        \SB1_2_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_16/Component_Function_0/N2  ( .A1(\SB1_2_16/i0[8] ), .A2(
        \SB1_2_16/i0[7] ), .A3(\SB1_2_16/i0[6] ), .ZN(
        \SB1_2_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_16/Component_Function_0/N1  ( .A1(\SB1_2_16/i0[10] ), .A2(
        \SB1_2_16/i0[9] ), .ZN(\SB1_2_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_1/N4  ( .A1(\SB1_2_16/i1_7 ), .A2(
        \SB1_2_16/i0[8] ), .A3(\SB1_2_16/i0_4 ), .ZN(
        \SB1_2_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_16/Component_Function_1/N3  ( .A1(\SB1_2_16/i1_5 ), .A2(
        \SB1_2_16/i0[6] ), .A3(\SB1_2_16/i0[9] ), .ZN(
        \SB1_2_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_16/Component_Function_1/N2  ( .A1(\SB1_2_16/i0_3 ), .A2(
        \SB1_2_16/i1_7 ), .A3(\SB1_2_16/i0[8] ), .ZN(
        \SB1_2_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_16/Component_Function_1/N1  ( .A1(\SB1_2_16/i0_3 ), .A2(
        \SB1_2_16/i1[9] ), .ZN(\SB1_2_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_5/N4  ( .A1(\SB1_2_16/i0[9] ), .A2(
        \SB1_2_16/i0[6] ), .A3(\SB1_2_16/i0_4 ), .ZN(
        \SB1_2_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_16/Component_Function_5/N2  ( .A1(\SB1_2_16/i0_0 ), .A2(
        \SB1_2_16/i0[6] ), .A3(\SB1_2_16/i0[10] ), .ZN(
        \SB1_2_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_16/Component_Function_5/N1  ( .A1(\SB1_2_16/i0_0 ), .A2(
        \SB1_2_16/i3[0] ), .ZN(\SB1_2_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_0/N4  ( .A1(\SB1_2_17/i0[7] ), .A2(
        \SB1_2_17/i0_3 ), .A3(\SB1_2_17/i0_0 ), .ZN(
        \SB1_2_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_17/Component_Function_0/N3  ( .A1(\SB1_2_17/i0[10] ), .A2(
        \SB1_2_17/i0_4 ), .A3(\SB1_2_17/i0_3 ), .ZN(
        \SB1_2_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_17/Component_Function_0/N2  ( .A1(\SB1_2_17/i0[8] ), .A2(
        \SB1_2_17/i0[7] ), .A3(\SB1_2_17/i0[6] ), .ZN(
        \SB1_2_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_17/Component_Function_0/N1  ( .A1(\SB1_2_17/i0[10] ), .A2(
        \SB1_2_17/i0[9] ), .ZN(\SB1_2_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_1/N4  ( .A1(\SB1_2_17/i1_7 ), .A2(
        \SB1_2_17/i0[8] ), .A3(\SB1_2_17/i0_4 ), .ZN(
        \SB1_2_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_17/Component_Function_1/N3  ( .A1(\SB1_2_17/i1_5 ), .A2(
        \SB1_2_17/i0[6] ), .A3(\SB1_2_17/i0[9] ), .ZN(
        \SB1_2_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_17/Component_Function_1/N2  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i1_7 ), .A3(\SB1_2_17/i0[8] ), .ZN(
        \SB1_2_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_17/Component_Function_1/N1  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i1[9] ), .ZN(\SB1_2_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_17/Component_Function_5/N1  ( .A1(\SB1_2_17/i0_0 ), .A2(
        \SB1_2_17/i3[0] ), .ZN(\SB1_2_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_0/N4  ( .A1(\SB1_2_18/i0[7] ), .A2(
        \SB1_2_18/i0_3 ), .A3(\SB1_2_18/i0_0 ), .ZN(
        \SB1_2_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_18/Component_Function_0/N3  ( .A1(\SB1_2_18/i0[10] ), .A2(
        \SB1_2_18/i0_4 ), .A3(\SB1_2_18/i0_3 ), .ZN(
        \SB1_2_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_18/Component_Function_0/N2  ( .A1(\SB1_2_18/i0[8] ), .A2(
        \SB1_2_18/i0[7] ), .A3(\SB1_2_18/i0[6] ), .ZN(
        \SB1_2_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_18/Component_Function_0/N1  ( .A1(\SB1_2_18/i0[10] ), .A2(
        \SB1_2_18/i0[9] ), .ZN(\SB1_2_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_1/N4  ( .A1(\SB1_2_18/i1_7 ), .A2(
        \SB1_2_18/i0[8] ), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_18/Component_Function_1/N3  ( .A1(\SB1_2_18/i1_5 ), .A2(
        \SB1_2_18/i0[6] ), .A3(\SB1_2_18/i0[9] ), .ZN(
        \SB1_2_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_18/Component_Function_1/N2  ( .A1(\SB1_2_18/i0_3 ), .A2(
        \SB1_2_18/i1_7 ), .A3(\SB1_2_18/i0[8] ), .ZN(
        \SB1_2_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_18/Component_Function_1/N1  ( .A1(\SB1_2_18/i0_3 ), .A2(
        \SB1_2_18/i1[9] ), .ZN(\SB1_2_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_5/N4  ( .A1(\SB1_2_18/i0[9] ), .A2(
        \SB1_2_18/i0[6] ), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_18/Component_Function_5/N2  ( .A1(\SB1_2_18/i0_0 ), .A2(
        \SB1_2_18/i0[6] ), .A3(\SB1_2_18/i0[10] ), .ZN(
        \SB1_2_18/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_18/Component_Function_5/N1  ( .A1(\SB1_2_18/i0_0 ), .A2(
        \SB1_2_18/i3[0] ), .ZN(\SB1_2_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N4  ( .A1(\SB1_2_19/i0[7] ), .A2(
        n1649), .A3(\SB1_2_19/i0_0 ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N3  ( .A1(\SB1_2_19/i0[10] ), .A2(
        \SB1_2_19/i0_4 ), .A3(\SB1_2_19/i0_3 ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N2  ( .A1(\SB1_2_19/i0[8] ), .A2(
        \SB1_2_19/i0[7] ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_19/Component_Function_0/N1  ( .A1(\SB1_2_19/i0[10] ), .A2(
        \SB1_2_19/i0[9] ), .ZN(\SB1_2_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_1/N4  ( .A1(\SB1_2_19/i1_7 ), .A2(
        \SB1_2_19/i0[8] ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_1/N3  ( .A1(\SB1_2_19/i1_5 ), .A2(
        \SB1_2_19/i0[6] ), .A3(\SB1_2_19/i0[9] ), .ZN(
        \SB1_2_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_19/Component_Function_1/N2  ( .A1(\SB1_2_19/i0_3 ), .A2(
        \SB1_2_19/i1_7 ), .A3(\SB1_2_19/i0[8] ), .ZN(
        \SB1_2_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_19/Component_Function_1/N1  ( .A1(n1649), .A2(
        \SB1_2_19/i1[9] ), .ZN(\SB1_2_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_5/N4  ( .A1(\SB1_2_19/i0[9] ), .A2(
        \SB1_2_19/i0[6] ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_5/N2  ( .A1(\SB1_2_19/i0_0 ), .A2(
        \SB1_2_19/i0[6] ), .A3(\SB1_2_19/i0[10] ), .ZN(
        \SB1_2_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_19/Component_Function_5/N1  ( .A1(\SB1_2_19/i0_0 ), .A2(
        \SB1_2_19/i3[0] ), .ZN(\SB1_2_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_0/N4  ( .A1(\SB1_2_20/i0[7] ), .A2(
        n1644), .A3(\SB1_2_20/i0_0 ), .ZN(
        \SB1_2_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_0/N3  ( .A1(\SB1_2_20/i0[10] ), .A2(
        \SB1_2_20/i0_4 ), .A3(n1644), .ZN(
        \SB1_2_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_20/Component_Function_0/N2  ( .A1(\SB1_2_20/i0[8] ), .A2(
        \SB1_2_20/i0[7] ), .A3(\SB1_2_20/i0[6] ), .ZN(
        \SB1_2_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_20/Component_Function_0/N1  ( .A1(\SB1_2_20/i0[10] ), .A2(
        \SB1_2_20/i0[9] ), .ZN(\SB1_2_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_1/N3  ( .A1(\SB1_2_20/i1_5 ), .A2(
        \SB1_2_20/i0[6] ), .A3(\SB1_2_20/i0[9] ), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_20/Component_Function_1/N2  ( .A1(\SB1_2_20/i0_3 ), .A2(
        \SB1_2_20/i1_7 ), .A3(\SB1_2_20/i0[8] ), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_20/Component_Function_1/N1  ( .A1(n1644), .A2(
        \SB1_2_20/i1[9] ), .ZN(\SB1_2_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_5/N4  ( .A1(\SB1_2_20/i0[9] ), .A2(
        \SB1_2_20/i0[6] ), .A3(\SB1_2_20/i0_4 ), .ZN(
        \SB1_2_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_5/N2  ( .A1(\SB1_2_20/i0_0 ), .A2(
        \SB1_2_20/i0[6] ), .A3(\SB1_2_20/i0[10] ), .ZN(
        \SB1_2_20/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_20/Component_Function_5/N1  ( .A1(\SB1_2_20/i0_0 ), .A2(
        \SB1_2_20/i3[0] ), .ZN(\SB1_2_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_0/N4  ( .A1(\SB1_2_21/i0[7] ), .A2(
        \SB1_2_21/i0_3 ), .A3(\SB1_2_21/i0_0 ), .ZN(
        \SB1_2_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_21/Component_Function_0/N2  ( .A1(\SB1_2_21/i0[8] ), .A2(
        \SB1_2_21/i0[7] ), .A3(\SB1_2_21/i0[6] ), .ZN(
        \SB1_2_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_21/Component_Function_0/N1  ( .A1(\SB1_2_21/i0[10] ), .A2(
        \SB1_2_21/i0[9] ), .ZN(\SB1_2_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_1/N3  ( .A1(\SB1_2_21/i1_5 ), .A2(
        \SB1_2_21/i0[6] ), .A3(\SB1_2_21/i0[9] ), .ZN(
        \SB1_2_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_21/Component_Function_1/N2  ( .A1(\SB1_2_21/i0_3 ), .A2(
        \SB1_2_21/i1_7 ), .A3(\SB1_2_21/i0[8] ), .ZN(
        \SB1_2_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_21/Component_Function_1/N1  ( .A1(\SB1_2_21/i0_3 ), .A2(
        \SB1_2_21/i1[9] ), .ZN(\SB1_2_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_5/N4  ( .A1(\SB1_2_21/i0[9] ), .A2(
        \SB1_2_21/i0[6] ), .A3(\SB1_2_21/i0_4 ), .ZN(
        \SB1_2_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_21/Component_Function_5/N2  ( .A1(\SB1_2_21/i0_0 ), .A2(
        \SB1_2_21/i0[6] ), .A3(\SB1_2_21/i0[10] ), .ZN(
        \SB1_2_21/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_21/Component_Function_5/N1  ( .A1(\SB1_2_21/i0_0 ), .A2(
        \SB1_2_21/i3[0] ), .ZN(\SB1_2_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_0/N4  ( .A1(\SB1_2_22/i0[7] ), .A2(
        \SB1_2_22/i0_3 ), .A3(\SB1_2_22/i0_0 ), .ZN(
        \SB1_2_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_22/Component_Function_0/N3  ( .A1(\SB1_2_22/i0[10] ), .A2(
        \SB1_2_22/i0_4 ), .A3(\SB1_2_22/i0_3 ), .ZN(
        \SB1_2_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_22/Component_Function_0/N2  ( .A1(\SB1_2_22/i0[8] ), .A2(
        \SB1_2_22/i0[7] ), .A3(\SB1_2_22/i0[6] ), .ZN(
        \SB1_2_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_22/Component_Function_0/N1  ( .A1(\SB1_2_22/i0[10] ), .A2(
        \SB1_2_22/i0[9] ), .ZN(\SB1_2_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_1/N3  ( .A1(\SB1_2_22/i1_5 ), .A2(
        \SB1_2_22/i0[6] ), .A3(\SB1_2_22/i0[9] ), .ZN(
        \SB1_2_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_22/Component_Function_1/N2  ( .A1(\SB1_2_22/i0_3 ), .A2(
        \SB1_2_22/i1_7 ), .A3(\SB1_2_22/i0[8] ), .ZN(
        \SB1_2_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_22/Component_Function_1/N1  ( .A1(\SB1_2_22/i0_3 ), .A2(
        \SB1_2_22/i1[9] ), .ZN(\SB1_2_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_5/N4  ( .A1(\SB1_2_22/i0[9] ), .A2(
        \SB1_2_22/i0[6] ), .A3(\SB1_2_22/i0_4 ), .ZN(
        \SB1_2_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_22/Component_Function_5/N2  ( .A1(\SB1_2_22/i0[10] ), .A2(
        \SB1_2_22/i0[6] ), .A3(\SB1_2_22/i0_0 ), .ZN(
        \SB1_2_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_22/Component_Function_5/N1  ( .A1(\SB1_2_22/i0_0 ), .A2(
        \SB1_2_22/i3[0] ), .ZN(\SB1_2_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N4  ( .A1(\SB1_2_23/i0[7] ), .A2(
        \SB1_2_23/i0_3 ), .A3(\SB1_2_23/i0_0 ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N3  ( .A1(\SB1_2_23/i0[10] ), .A2(
        \SB1_2_23/i0_4 ), .A3(\SB1_2_23/i0_3 ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N2  ( .A1(\SB1_2_23/i0[8] ), .A2(
        \SB1_2_23/i0[7] ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_23/Component_Function_0/N1  ( .A1(\SB1_2_23/i0[10] ), .A2(
        \SB1_2_23/i0[9] ), .ZN(\SB1_2_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_1/N4  ( .A1(\SB1_2_23/i1_7 ), .A2(
        \SB1_2_23/i0[8] ), .A3(\SB1_2_23/i0_4 ), .ZN(
        \SB1_2_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_23/Component_Function_1/N3  ( .A1(\SB1_2_23/i1_5 ), .A2(
        \SB1_2_23/i0[6] ), .A3(\SB1_2_23/i0[9] ), .ZN(
        \SB1_2_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_23/Component_Function_1/N2  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i1_7 ), .A3(\SB1_2_23/i0[8] ), .ZN(
        \SB1_2_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_23/Component_Function_1/N1  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i1[9] ), .ZN(\SB1_2_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_5/N4  ( .A1(\SB1_2_23/i0[9] ), .A2(
        \SB1_2_23/i0[6] ), .A3(\SB1_2_23/i0_4 ), .ZN(
        \SB1_2_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_23/Component_Function_5/N2  ( .A1(\SB1_2_23/i0_0 ), .A2(
        \SB1_2_23/i0[6] ), .A3(\SB1_2_23/i0[10] ), .ZN(
        \SB1_2_23/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_23/Component_Function_5/N1  ( .A1(\SB1_2_23/i0_0 ), .A2(
        \SB1_2_23/i3[0] ), .ZN(\SB1_2_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_0/N4  ( .A1(\SB1_2_24/i0[7] ), .A2(
        \SB1_2_24/i0_3 ), .A3(\SB1_2_24/i0_0 ), .ZN(
        \SB1_2_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_24/Component_Function_0/N3  ( .A1(\SB1_2_24/i0[10] ), .A2(
        \SB1_2_24/i0_4 ), .A3(\SB1_2_24/i0_3 ), .ZN(
        \SB1_2_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_24/Component_Function_0/N2  ( .A1(\SB1_2_24/i0[8] ), .A2(
        \SB1_2_24/i0[7] ), .A3(\SB1_2_24/i0[6] ), .ZN(
        \SB1_2_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_24/Component_Function_0/N1  ( .A1(\SB1_2_24/i0[10] ), .A2(
        \SB1_2_24/i0[9] ), .ZN(\SB1_2_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_1/N4  ( .A1(\SB1_2_24/i1_7 ), .A2(
        \SB1_2_24/i0[8] ), .A3(\SB1_2_24/i0_4 ), .ZN(
        \SB1_2_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_24/Component_Function_1/N3  ( .A1(\SB1_2_24/i1_5 ), .A2(
        \SB1_2_24/i0[6] ), .A3(\SB1_2_24/i0[9] ), .ZN(
        \SB1_2_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_24/Component_Function_1/N2  ( .A1(\SB1_2_24/i0_3 ), .A2(
        \SB1_2_24/i1_7 ), .A3(\SB1_2_24/i0[8] ), .ZN(
        \SB1_2_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_24/Component_Function_1/N1  ( .A1(\SB1_2_24/i0_3 ), .A2(
        \SB1_2_24/i1[9] ), .ZN(\SB1_2_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_5/N4  ( .A1(\SB1_2_24/i0[9] ), .A2(
        \SB1_2_24/i0[6] ), .A3(\SB1_2_24/i0_4 ), .ZN(
        \SB1_2_24/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_24/Component_Function_5/N1  ( .A1(\SB1_2_24/i0_0 ), .A2(
        \SB1_2_24/i3[0] ), .ZN(\SB1_2_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N4  ( .A1(\SB1_2_25/i0[7] ), .A2(
        \SB1_2_25/i0_3 ), .A3(\SB1_2_25/i0_0 ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N3  ( .A1(\SB1_2_25/i0[10] ), .A2(
        \SB1_2_25/i0_4 ), .A3(\SB1_2_25/i0_3 ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N2  ( .A1(\SB1_2_25/i0[8] ), .A2(
        \SB1_2_25/i0[7] ), .A3(\SB1_2_25/i0[6] ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_25/Component_Function_0/N1  ( .A1(\SB1_2_25/i0[10] ), .A2(
        \SB1_2_25/i0[9] ), .ZN(\SB1_2_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_1/N4  ( .A1(\SB1_2_25/i1_7 ), .A2(
        \SB1_2_25/i0[8] ), .A3(\SB1_2_25/i0_4 ), .ZN(
        \SB1_2_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_1/N3  ( .A1(\SB1_2_25/i1_5 ), .A2(
        \SB1_2_25/i0[6] ), .A3(\SB1_2_25/i0[9] ), .ZN(
        \SB1_2_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_1/N2  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i1_7 ), .A3(\SB1_2_25/i0[8] ), .ZN(
        \SB1_2_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_25/Component_Function_1/N1  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i1[9] ), .ZN(\SB1_2_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_5/N4  ( .A1(\SB1_2_25/i0[9] ), .A2(
        \SB1_2_25/i0[6] ), .A3(\SB1_2_25/i0_4 ), .ZN(
        \SB1_2_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_5/N2  ( .A1(\SB1_2_25/i0_0 ), .A2(
        \SB1_2_25/i0[6] ), .A3(\SB1_2_25/i0[10] ), .ZN(
        \SB1_2_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_25/Component_Function_5/N1  ( .A1(\SB1_2_25/i0_0 ), .A2(
        \SB1_2_25/i3[0] ), .ZN(\SB1_2_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_0/N4  ( .A1(\SB1_2_26/i0_0 ), .A2(
        \SB1_2_26/i0_3 ), .A3(\SB1_2_26/i0[7] ), .ZN(
        \SB1_2_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_26/Component_Function_0/N2  ( .A1(\SB1_2_26/i0[8] ), .A2(
        \SB1_2_26/i0[7] ), .A3(\SB1_2_26/i0[6] ), .ZN(
        \SB1_2_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_26/Component_Function_0/N1  ( .A1(\SB1_2_26/i0[10] ), .A2(
        \SB1_2_26/i0[9] ), .ZN(\SB1_2_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_1/N4  ( .A1(\SB1_2_26/i1_7 ), .A2(
        \SB1_2_26/i0[8] ), .A3(\SB1_2_26/i0_4 ), .ZN(
        \SB1_2_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_26/Component_Function_1/N3  ( .A1(\SB1_2_26/i1_5 ), .A2(
        \SB1_2_26/i0[6] ), .A3(\SB1_2_26/i0[9] ), .ZN(
        \SB1_2_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_26/Component_Function_1/N2  ( .A1(\SB1_2_26/i0_3 ), .A2(
        \SB1_2_26/i1_7 ), .A3(\SB1_2_26/i0[8] ), .ZN(
        \SB1_2_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_26/Component_Function_1/N1  ( .A1(\SB1_2_26/i0_3 ), .A2(
        \SB1_2_26/i1[9] ), .ZN(\SB1_2_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_5/N4  ( .A1(\SB1_2_26/i0[9] ), .A2(
        \SB1_2_26/i0[6] ), .A3(\SB1_2_26/i0_4 ), .ZN(
        \SB1_2_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_26/Component_Function_5/N2  ( .A1(\SB1_2_26/i0_0 ), .A2(
        \SB1_2_26/i0[6] ), .A3(\SB1_2_26/i0[10] ), .ZN(
        \SB1_2_26/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_26/Component_Function_5/N1  ( .A1(\SB1_2_26/i0_0 ), .A2(
        \SB1_2_26/i3[0] ), .ZN(\SB1_2_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N4  ( .A1(\SB1_2_27/i0[7] ), .A2(
        \SB1_2_27/i0_3 ), .A3(\SB1_2_27/i0_0 ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N3  ( .A1(\SB1_2_27/i0[10] ), .A2(
        \SB1_2_27/i0_4 ), .A3(\SB1_2_27/i0_3 ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N2  ( .A1(\SB1_2_27/i0[8] ), .A2(
        \SB1_2_27/i0[7] ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_27/Component_Function_0/N1  ( .A1(\SB1_2_27/i0[10] ), .A2(
        \SB1_2_27/i0[9] ), .ZN(\SB1_2_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N4  ( .A1(\SB1_2_27/i1_7 ), .A2(
        \SB1_2_27/i0[8] ), .A3(\SB1_2_27/i0_4 ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N3  ( .A1(\SB1_2_27/i1_5 ), .A2(
        \SB1_2_27/i0[6] ), .A3(\SB1_2_27/i0[9] ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N2  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i1_7 ), .A3(\SB1_2_27/i0[8] ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_27/Component_Function_1/N1  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i1[9] ), .ZN(\SB1_2_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_5/N4  ( .A1(\SB1_2_27/i0[9] ), .A2(
        \SB1_2_27/i0[6] ), .A3(\SB1_2_27/i0_4 ), .ZN(
        \SB1_2_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_5/N2  ( .A1(\SB1_2_27/i0_0 ), .A2(
        \SB1_2_27/i0[6] ), .A3(\SB1_2_27/i0[10] ), .ZN(
        \SB1_2_27/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_27/Component_Function_5/N1  ( .A1(\SB1_2_27/i0_0 ), .A2(
        \SB1_2_27/i3[0] ), .ZN(\SB1_2_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N4  ( .A1(\SB1_2_28/i0[7] ), .A2(
        \SB1_2_28/i0_3 ), .A3(\SB1_2_28/i0_0 ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N3  ( .A1(\SB1_2_28/i0[10] ), .A2(
        \SB1_2_28/i0_4 ), .A3(\SB1_2_28/i0_3 ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N2  ( .A1(\SB1_2_28/i0[8] ), .A2(
        \SB1_2_28/i0[7] ), .A3(\SB1_2_28/i0[6] ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_28/Component_Function_0/N1  ( .A1(\SB1_2_28/i0[10] ), .A2(
        \SB1_2_28/i0[9] ), .ZN(\SB1_2_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_1/N4  ( .A1(\SB1_2_28/i1_7 ), .A2(
        \SB1_2_28/i0[8] ), .A3(\SB1_2_28/i0_4 ), .ZN(
        \SB1_2_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_1/N3  ( .A1(\SB1_2_28/i1_5 ), .A2(
        \SB1_2_28/i0[6] ), .A3(\SB1_2_28/i0[9] ), .ZN(
        \SB1_2_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_28/Component_Function_1/N2  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i1_7 ), .A3(\SB1_2_28/i0[8] ), .ZN(
        \SB1_2_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_28/Component_Function_1/N1  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i1[9] ), .ZN(\SB1_2_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_5/N4  ( .A1(\SB1_2_28/i0[9] ), .A2(
        \SB1_2_28/i0[6] ), .A3(\SB1_2_28/i0_4 ), .ZN(
        \SB1_2_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_5/N2  ( .A1(\SB1_2_28/i0_0 ), .A2(
        \SB1_2_28/i0[6] ), .A3(\SB1_2_28/i0[10] ), .ZN(
        \SB1_2_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_28/Component_Function_5/N1  ( .A1(\SB1_2_28/i0_0 ), .A2(
        \SB1_2_28/i3[0] ), .ZN(\SB1_2_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_0/N4  ( .A1(\SB1_2_29/i0[7] ), .A2(
        n814), .A3(\SB1_2_29/i0_0 ), .ZN(
        \SB1_2_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_29/Component_Function_0/N3  ( .A1(\SB1_2_29/i0[10] ), .A2(
        \SB1_2_29/i0_4 ), .A3(\SB1_2_29/i0_3 ), .ZN(
        \SB1_2_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_29/Component_Function_0/N2  ( .A1(\SB1_2_29/i0[8] ), .A2(
        \SB1_2_29/i0[7] ), .A3(\SB1_2_29/i0[6] ), .ZN(
        \SB1_2_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_29/Component_Function_0/N1  ( .A1(\SB1_2_29/i0[10] ), .A2(
        \SB1_2_29/i0[9] ), .ZN(\SB1_2_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_1/N3  ( .A1(\SB1_2_29/i1_5 ), .A2(
        \SB1_2_29/i0[6] ), .A3(\SB1_2_29/i0[9] ), .ZN(
        \SB1_2_29/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_29/Component_Function_1/N1  ( .A1(n814), .A2(
        \SB1_2_29/i1[9] ), .ZN(\SB1_2_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_5/N4  ( .A1(\SB1_2_29/i0[9] ), .A2(
        \SB1_2_29/i0[6] ), .A3(\SB1_2_29/i0_4 ), .ZN(
        \SB1_2_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_29/Component_Function_5/N2  ( .A1(\SB1_2_29/i0_0 ), .A2(
        \SB1_2_29/i0[6] ), .A3(\SB1_2_29/i0[10] ), .ZN(
        \SB1_2_29/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_29/Component_Function_5/N1  ( .A1(\SB1_2_29/i0_0 ), .A2(
        \SB1_2_29/i3[0] ), .ZN(\SB1_2_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_0/N4  ( .A1(\SB1_2_30/i0[7] ), .A2(
        \SB1_2_30/i0_3 ), .A3(\SB1_2_30/i0_0 ), .ZN(
        \SB1_2_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_30/Component_Function_0/N3  ( .A1(\SB1_2_30/i0[10] ), .A2(
        \SB1_2_30/i0_4 ), .A3(\SB1_2_30/i0_3 ), .ZN(
        \SB1_2_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_30/Component_Function_0/N2  ( .A1(\SB1_2_30/i0[8] ), .A2(
        \SB1_2_30/i0[7] ), .A3(\SB1_2_30/i0[6] ), .ZN(
        \SB1_2_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_30/Component_Function_0/N1  ( .A1(\SB1_2_30/i0[10] ), .A2(
        \SB1_2_30/i0[9] ), .ZN(\SB1_2_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_1/N4  ( .A1(\SB1_2_30/i1_7 ), .A2(
        \SB1_2_30/i0[8] ), .A3(\SB1_2_30/i0_4 ), .ZN(
        \SB1_2_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_30/Component_Function_1/N3  ( .A1(\SB1_2_30/i1_5 ), .A2(
        \SB1_2_30/i0[6] ), .A3(\SB1_2_30/i0[9] ), .ZN(
        \SB1_2_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_30/Component_Function_1/N2  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i1_7 ), .A3(\SB1_2_30/i0[8] ), .ZN(
        \SB1_2_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_30/Component_Function_1/N1  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i1[9] ), .ZN(\SB1_2_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_5/N4  ( .A1(\SB1_2_30/i0[9] ), .A2(
        \SB1_2_30/i0[6] ), .A3(\SB1_2_30/i0_4 ), .ZN(
        \SB1_2_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_30/Component_Function_5/N2  ( .A1(\SB1_2_30/i0_0 ), .A2(
        \SB1_2_30/i0[6] ), .A3(\SB1_2_30/i0[10] ), .ZN(
        \SB1_2_30/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_30/Component_Function_5/N1  ( .A1(\SB1_2_30/i0_0 ), .A2(
        \SB1_2_30/i3[0] ), .ZN(\SB1_2_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_0/N4  ( .A1(\SB1_2_31/i0[7] ), .A2(
        \SB1_2_31/i0_3 ), .A3(\SB1_2_31/i0_0 ), .ZN(
        \SB1_2_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_31/Component_Function_0/N3  ( .A1(\SB1_2_31/i0[10] ), .A2(
        \SB1_2_31/i0_4 ), .A3(\SB1_2_31/i0_3 ), .ZN(
        \SB1_2_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_31/Component_Function_0/N2  ( .A1(\SB1_2_31/i0[8] ), .A2(
        \SB1_2_31/i0[7] ), .A3(\SB1_2_31/i0[6] ), .ZN(
        \SB1_2_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_31/Component_Function_0/N1  ( .A1(\SB1_2_31/i0[10] ), .A2(
        \SB1_2_31/i0[9] ), .ZN(\SB1_2_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_1/N3  ( .A1(\SB1_2_31/i1_5 ), .A2(
        \SB1_2_31/i0[6] ), .A3(\SB1_2_31/i0[9] ), .ZN(
        \SB1_2_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_31/Component_Function_1/N2  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i1_7 ), .A3(\SB1_2_31/i0[8] ), .ZN(
        \SB1_2_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_31/Component_Function_1/N1  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i1[9] ), .ZN(\SB1_2_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_5/N4  ( .A1(\SB1_2_31/i0[9] ), .A2(
        \SB1_2_31/i0[6] ), .A3(\SB1_2_31/i0_4 ), .ZN(
        \SB1_2_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_31/Component_Function_5/N2  ( .A1(\SB1_2_31/i0_0 ), .A2(
        \SB1_2_31/i0[6] ), .A3(\SB1_2_31/i0[10] ), .ZN(
        \SB1_2_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_31/Component_Function_5/N1  ( .A1(\SB1_2_31/i0_0 ), .A2(
        \SB1_2_31/i3[0] ), .ZN(\SB1_2_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_0/N3  ( .A1(\SB2_2_0/i0[10] ), .A2(
        \SB2_2_0/i0_4 ), .A3(\SB2_2_0/i0_3 ), .ZN(
        \SB2_2_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_0/Component_Function_0/N2  ( .A1(\SB2_2_0/i0[8] ), .A2(
        \SB2_2_0/i0[7] ), .A3(\SB2_2_0/i0[6] ), .ZN(
        \SB2_2_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_0/Component_Function_0/N1  ( .A1(\SB2_2_0/i0[10] ), .A2(
        \SB2_2_0/i0[9] ), .ZN(\SB2_2_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_1/N4  ( .A1(\SB2_2_0/i1_7 ), .A2(
        \SB2_2_0/i0[8] ), .A3(\SB2_2_0/i0_4 ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_0/Component_Function_1/N3  ( .A1(\SB2_2_0/i1_5 ), .A2(
        \SB2_2_0/i0[6] ), .A3(\SB2_2_0/i0[9] ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_0/Component_Function_1/N2  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i1_7 ), .A3(\SB2_2_0/i0[8] ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_0/Component_Function_1/N1  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i1[9] ), .ZN(\SB2_2_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_5/N4  ( .A1(\SB2_2_0/i0[9] ), .A2(
        \SB2_2_0/i0[6] ), .A3(\SB2_2_0/i0_4 ), .ZN(
        \SB2_2_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_0/Component_Function_5/N3  ( .A1(\SB2_2_0/i1[9] ), .A2(
        \SB2_2_0/i0_4 ), .A3(\SB2_2_0/i0_3 ), .ZN(
        \SB2_2_0/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_0/Component_Function_5/N1  ( .A1(\SB2_2_0/i0_0 ), .A2(
        \SB2_2_0/i3[0] ), .ZN(\SB2_2_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_0/N4  ( .A1(\SB2_2_1/i0[7] ), .A2(
        \SB2_2_1/i0_3 ), .A3(\SB2_2_1/i0_0 ), .ZN(
        \SB2_2_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_1/Component_Function_0/N3  ( .A1(\SB2_2_1/i0_3 ), .A2(
        \SB2_2_1/i0_4 ), .A3(\SB2_2_1/i0[10] ), .ZN(
        \SB2_2_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_1/Component_Function_0/N2  ( .A1(\SB2_2_1/i0[8] ), .A2(
        \SB2_2_1/i0[7] ), .A3(\SB2_2_1/i0[6] ), .ZN(
        \SB2_2_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_1/Component_Function_0/N1  ( .A1(\SB2_2_1/i0[10] ), .A2(
        \SB2_2_1/i0[9] ), .ZN(\SB2_2_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_1/N3  ( .A1(\SB2_2_1/i1_5 ), .A2(
        \SB2_2_1/i0[6] ), .A3(\SB2_2_1/i0[9] ), .ZN(
        \SB2_2_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_1/Component_Function_1/N2  ( .A1(\SB2_2_1/i0_3 ), .A2(
        \SB2_2_1/i1_7 ), .A3(\SB2_2_1/i0[8] ), .ZN(
        \SB2_2_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_1/Component_Function_1/N1  ( .A1(\SB2_2_1/i0_3 ), .A2(
        \SB2_2_1/i1[9] ), .ZN(\SB2_2_1/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_1/Component_Function_5/N1  ( .A1(\SB2_2_1/i0_0 ), .A2(
        \SB2_2_1/i3[0] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_0/N4  ( .A1(\SB2_2_2/i0[7] ), .A2(
        \SB2_2_2/i0_3 ), .A3(\SB2_2_2/i0_0 ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_2/Component_Function_0/N3  ( .A1(\SB2_2_2/i0[10] ), .A2(
        \SB2_2_2/i0_4 ), .A3(\SB2_2_2/i0_3 ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_2/Component_Function_0/N2  ( .A1(\SB2_2_2/i0[8] ), .A2(
        \SB2_2_2/i0[7] ), .A3(\SB2_2_2/i0[6] ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_2/Component_Function_0/N1  ( .A1(\SB2_2_2/i0[10] ), .A2(
        \SB2_2_2/i0[9] ), .ZN(\SB2_2_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_1/N4  ( .A1(\SB2_2_2/i1_7 ), .A2(
        \SB2_2_2/i0[8] ), .A3(\SB2_2_2/i0_4 ), .ZN(
        \SB2_2_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_2/Component_Function_1/N3  ( .A1(\SB2_2_2/i1_5 ), .A2(
        \SB2_2_2/i0[6] ), .A3(\SB2_2_2/i0[9] ), .ZN(
        \SB2_2_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_2/Component_Function_1/N2  ( .A1(\SB2_2_2/i0_3 ), .A2(
        \SB2_2_2/i1_7 ), .A3(\SB2_2_2/i0[8] ), .ZN(
        \SB2_2_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_2/Component_Function_1/N1  ( .A1(\SB2_2_2/i0_3 ), .A2(
        \SB2_2_2/i1[9] ), .ZN(\SB2_2_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_5/N4  ( .A1(\SB2_2_2/i0[9] ), .A2(
        \SB2_2_2/i0[6] ), .A3(\SB2_2_2/i0_4 ), .ZN(
        \SB2_2_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_2/Component_Function_5/N3  ( .A1(\SB2_2_2/i1[9] ), .A2(
        \SB2_2_2/i0_4 ), .A3(\SB2_2_2/i0_3 ), .ZN(
        \SB2_2_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_2/Component_Function_5/N2  ( .A1(\SB2_2_2/i0_0 ), .A2(
        \SB2_2_2/i0[6] ), .A3(\SB2_2_2/i0[10] ), .ZN(
        \SB2_2_2/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_3/Component_Function_0/N4  ( .A1(\SB2_2_3/i0[7] ), .A2(
        \SB2_2_3/i0_3 ), .A3(\SB2_2_3/i0_0 ), .ZN(
        \SB2_2_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_3/Component_Function_0/N3  ( .A1(\SB2_2_3/i0[10] ), .A2(
        \SB2_2_3/i0_4 ), .A3(\SB2_2_3/i0_3 ), .ZN(
        \SB2_2_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_3/Component_Function_0/N2  ( .A1(\SB2_2_3/i0[8] ), .A2(
        \SB2_2_3/i0[7] ), .A3(\SB2_2_3/i0[6] ), .ZN(
        \SB2_2_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_3/Component_Function_0/N1  ( .A1(\SB2_2_3/i0[10] ), .A2(
        \SB2_2_3/i0[9] ), .ZN(\SB2_2_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_3/Component_Function_1/N4  ( .A1(\SB2_2_3/i1_7 ), .A2(
        \SB2_2_3/i0[8] ), .A3(\SB2_2_3/i0_4 ), .ZN(
        \SB2_2_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_3/Component_Function_1/N3  ( .A1(\SB2_2_3/i1_5 ), .A2(
        \SB2_2_3/i0[6] ), .A3(\SB2_2_3/i0[9] ), .ZN(
        \SB2_2_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_3/Component_Function_1/N2  ( .A1(\SB2_2_3/i0_3 ), .A2(
        \SB2_2_3/i1_7 ), .A3(\SB2_2_3/i0[8] ), .ZN(
        \SB2_2_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_3/Component_Function_1/N1  ( .A1(\SB2_2_3/i0_3 ), .A2(
        \SB2_2_3/i1[9] ), .ZN(\SB2_2_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_3/Component_Function_5/N4  ( .A1(\SB2_2_3/i0[9] ), .A2(
        \SB2_2_3/i0[6] ), .A3(\SB2_2_3/i0_4 ), .ZN(
        \SB2_2_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_3/Component_Function_5/N3  ( .A1(\SB2_2_3/i1[9] ), .A2(
        \SB2_2_3/i0_4 ), .A3(\SB2_2_3/i0_3 ), .ZN(
        \SB2_2_3/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_3/Component_Function_5/N1  ( .A1(\SB2_2_3/i0_0 ), .A2(
        \SB2_2_3/i3[0] ), .ZN(\SB2_2_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_0/N4  ( .A1(\SB2_2_4/i0[7] ), .A2(
        \SB2_2_4/i0_3 ), .A3(\SB2_2_4/i0_0 ), .ZN(
        \SB2_2_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_4/Component_Function_0/N3  ( .A1(\SB2_2_4/i0[10] ), .A2(
        \SB2_2_4/i0_4 ), .A3(\SB2_2_4/i0_3 ), .ZN(
        \SB2_2_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_4/Component_Function_0/N2  ( .A1(\SB2_2_4/i0[8] ), .A2(
        \SB2_2_4/i0[7] ), .A3(\SB2_2_4/i0[6] ), .ZN(
        \SB2_2_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_4/Component_Function_0/N1  ( .A1(\SB2_2_4/i0[10] ), .A2(
        \SB2_2_4/i0[9] ), .ZN(\SB2_2_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_1/N4  ( .A1(\SB2_2_4/i1_7 ), .A2(
        \SB2_2_4/i0[8] ), .A3(\SB2_2_4/i0_4 ), .ZN(
        \SB2_2_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_4/Component_Function_1/N3  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0[6] ), .A3(\SB2_2_4/i0[9] ), .ZN(
        \SB2_2_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_4/Component_Function_1/N2  ( .A1(\SB2_2_4/i0_3 ), .A2(
        \SB2_2_4/i1_7 ), .A3(\SB2_2_4/i0[8] ), .ZN(
        \SB2_2_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_4/Component_Function_1/N1  ( .A1(\SB2_2_4/i0_3 ), .A2(
        \SB2_2_4/i1[9] ), .ZN(\SB2_2_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_5/N2  ( .A1(\SB2_2_4/i0_0 ), .A2(
        \SB2_2_4/i0[6] ), .A3(\SB2_2_4/i0[10] ), .ZN(
        \SB2_2_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_4/Component_Function_5/N1  ( .A1(\SB2_2_4/i0_0 ), .A2(
        \SB2_2_4/i3[0] ), .ZN(\SB2_2_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_0/N4  ( .A1(\SB2_2_5/i0[7] ), .A2(
        \SB2_2_5/i0_3 ), .A3(\SB2_2_5/i0_0 ), .ZN(
        \SB2_2_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_5/Component_Function_0/N3  ( .A1(\SB2_2_5/i0[10] ), .A2(
        \SB2_2_5/i0_4 ), .A3(\SB2_2_5/i0_3 ), .ZN(
        \SB2_2_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_5/Component_Function_0/N2  ( .A1(\SB2_2_5/i0[8] ), .A2(
        \SB2_2_5/i0[7] ), .A3(\SB2_2_5/i0[6] ), .ZN(
        \SB2_2_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_5/Component_Function_0/N1  ( .A1(\SB2_2_5/i0[10] ), .A2(
        \SB2_2_5/i0[9] ), .ZN(\SB2_2_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_1/N4  ( .A1(\SB2_2_5/i1_7 ), .A2(
        \SB2_2_5/i0[8] ), .A3(\SB2_2_5/i0_4 ), .ZN(
        \SB2_2_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_5/Component_Function_1/N3  ( .A1(\SB2_2_5/i1_5 ), .A2(
        \SB2_2_5/i0[6] ), .A3(\SB2_2_5/i0[9] ), .ZN(
        \SB2_2_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_5/Component_Function_1/N2  ( .A1(\SB2_2_5/i0_3 ), .A2(
        \SB2_2_5/i1_7 ), .A3(\SB2_2_5/i0[8] ), .ZN(
        \SB2_2_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_5/Component_Function_1/N1  ( .A1(\SB2_2_5/i0_3 ), .A2(
        \SB2_2_5/i1[9] ), .ZN(\SB2_2_5/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_5/Component_Function_5/N1  ( .A1(\SB2_2_5/i0_0 ), .A2(
        \SB2_2_5/i3[0] ), .ZN(\SB2_2_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_0/N4  ( .A1(\SB2_2_6/i0[7] ), .A2(
        \SB2_2_6/i0_3 ), .A3(\SB2_2_6/i0_0 ), .ZN(
        \SB2_2_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_6/Component_Function_0/N3  ( .A1(\SB2_2_6/i0[10] ), .A2(
        \SB2_2_6/i0_4 ), .A3(\SB2_2_6/i0_3 ), .ZN(
        \SB2_2_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_6/Component_Function_0/N2  ( .A1(\SB2_2_6/i0[8] ), .A2(
        \SB2_2_6/i0[7] ), .A3(\SB2_2_6/i0[6] ), .ZN(
        \SB2_2_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_6/Component_Function_0/N1  ( .A1(\SB2_2_6/i0[10] ), .A2(
        \SB2_2_6/i0[9] ), .ZN(\SB2_2_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_1/N4  ( .A1(\SB2_2_6/i1_7 ), .A2(
        \SB2_2_6/i0[8] ), .A3(\SB2_2_6/i0_4 ), .ZN(
        \SB2_2_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_6/Component_Function_1/N3  ( .A1(\SB2_2_6/i1_5 ), .A2(
        \SB2_2_6/i0[6] ), .A3(\SB2_2_6/i0[9] ), .ZN(
        \SB2_2_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_6/Component_Function_1/N2  ( .A1(\SB2_2_6/i0_3 ), .A2(
        \SB2_2_6/i1_7 ), .A3(\SB2_2_6/i0[8] ), .ZN(
        \SB2_2_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_6/Component_Function_1/N1  ( .A1(\SB2_2_6/i0_3 ), .A2(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_5/N4  ( .A1(\SB2_2_6/i0[9] ), .A2(
        \SB2_2_6/i0[6] ), .A3(\SB2_2_6/i0_4 ), .ZN(
        \SB2_2_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_6/Component_Function_5/N2  ( .A1(\SB2_2_6/i0_0 ), .A2(
        \SB2_2_6/i0[6] ), .A3(\SB2_2_6/i0[10] ), .ZN(
        \SB2_2_6/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_6/Component_Function_5/N1  ( .A1(\SB2_2_6/i0_0 ), .A2(
        \SB2_2_6/i3[0] ), .ZN(\SB2_2_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_7/Component_Function_0/N4  ( .A1(\SB2_2_7/i0[7] ), .A2(
        \SB2_2_7/i0_3 ), .A3(\SB2_2_7/i0_0 ), .ZN(
        \SB2_2_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_7/Component_Function_0/N3  ( .A1(\SB2_2_7/i0[10] ), .A2(
        \SB2_2_7/i0_4 ), .A3(\SB2_2_7/i0_3 ), .ZN(
        \SB2_2_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_7/Component_Function_0/N2  ( .A1(\SB2_2_7/i0[8] ), .A2(
        \SB2_2_7/i0[7] ), .A3(\SB2_2_7/i0[6] ), .ZN(
        \SB2_2_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_7/Component_Function_0/N1  ( .A1(\SB2_2_7/i0[10] ), .A2(
        \SB2_2_7/i0[9] ), .ZN(\SB2_2_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_7/Component_Function_1/N4  ( .A1(\SB2_2_7/i1_7 ), .A2(
        \SB2_2_7/i0[8] ), .A3(\SB2_2_7/i0_4 ), .ZN(
        \SB2_2_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_7/Component_Function_1/N3  ( .A1(\SB2_2_7/i1_5 ), .A2(
        \SB2_2_7/i0[6] ), .A3(\SB2_2_7/i0[9] ), .ZN(
        \SB2_2_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_7/Component_Function_1/N2  ( .A1(\SB2_2_7/i0_3 ), .A2(
        \SB2_2_7/i1_7 ), .A3(\SB2_2_7/i0[8] ), .ZN(
        \SB2_2_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_7/Component_Function_1/N1  ( .A1(\SB2_2_7/i0_3 ), .A2(
        \SB2_2_7/i1[9] ), .ZN(\SB2_2_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_7/Component_Function_5/N2  ( .A1(\SB2_2_7/i0_0 ), .A2(
        \SB2_2_7/i0[6] ), .A3(\SB2_2_7/i0[10] ), .ZN(
        \SB2_2_7/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_7/Component_Function_5/N1  ( .A1(\SB2_2_7/i0_0 ), .A2(
        \SB2_2_7/i3[0] ), .ZN(\SB2_2_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_8/Component_Function_0/N3  ( .A1(\SB2_2_8/i0[10] ), .A2(
        \SB2_2_8/i0_4 ), .A3(\SB2_2_8/i0_3 ), .ZN(
        \SB2_2_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_8/Component_Function_0/N2  ( .A1(\SB2_2_8/i0[8] ), .A2(
        \SB2_2_8/i0[7] ), .A3(\SB2_2_8/i0[6] ), .ZN(
        \SB2_2_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_8/Component_Function_0/N1  ( .A1(\SB2_2_8/i0[10] ), .A2(
        \SB2_2_8/i0[9] ), .ZN(\SB2_2_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_8/Component_Function_1/N4  ( .A1(\SB2_2_8/i1_7 ), .A2(
        \SB2_2_8/i0[8] ), .A3(\SB2_2_8/i0_4 ), .ZN(
        \SB2_2_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_8/Component_Function_1/N3  ( .A1(\SB2_2_8/i1_5 ), .A2(
        \SB2_2_8/i0[6] ), .A3(\SB2_2_8/i0[9] ), .ZN(
        \SB2_2_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_8/Component_Function_1/N2  ( .A1(\SB2_2_8/i0_3 ), .A2(
        \SB2_2_8/i1_7 ), .A3(\SB2_2_8/i0[8] ), .ZN(
        \SB2_2_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_8/Component_Function_1/N1  ( .A1(\SB2_2_8/i0_3 ), .A2(
        \SB2_2_8/i1[9] ), .ZN(\SB2_2_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_8/Component_Function_5/N1  ( .A1(\SB2_2_8/i0_0 ), .A2(
        \SB2_2_8/i3[0] ), .ZN(\SB2_2_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_0/N4  ( .A1(\SB2_2_9/i0[7] ), .A2(
        \SB2_2_9/i0_3 ), .A3(\SB2_2_9/i0_0 ), .ZN(
        \SB2_2_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_9/Component_Function_0/N3  ( .A1(\SB2_2_9/i0[10] ), .A2(
        \SB2_2_9/i0_4 ), .A3(\SB2_2_9/i0_3 ), .ZN(
        \SB2_2_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_9/Component_Function_0/N2  ( .A1(\SB2_2_9/i0[8] ), .A2(
        \SB2_2_9/i0[7] ), .A3(\SB2_2_9/i0[6] ), .ZN(
        \SB2_2_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_9/Component_Function_0/N1  ( .A1(\SB2_2_9/i0[10] ), .A2(
        \SB2_2_9/i0[9] ), .ZN(\SB2_2_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_1/N4  ( .A1(\SB2_2_9/i1_7 ), .A2(
        \SB2_2_9/i0[8] ), .A3(\SB2_2_9/i0_4 ), .ZN(
        \SB2_2_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_9/Component_Function_1/N3  ( .A1(\SB2_2_9/i1_5 ), .A2(
        \SB2_2_9/i0[6] ), .A3(\SB2_2_9/i0[9] ), .ZN(
        \SB2_2_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_9/Component_Function_1/N2  ( .A1(\SB2_2_9/i0_3 ), .A2(
        \SB2_2_9/i1_7 ), .A3(\SB2_2_9/i0[8] ), .ZN(
        \SB2_2_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_9/Component_Function_1/N1  ( .A1(\SB2_2_9/i0_3 ), .A2(
        \SB2_2_9/i1[9] ), .ZN(\SB2_2_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_5/N3  ( .A1(\SB2_2_9/i1[9] ), .A2(
        \SB2_2_9/i0_4 ), .A3(\SB2_2_9/i0_3 ), .ZN(
        \SB2_2_9/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_10/Component_Function_0/N4  ( .A1(\SB2_2_10/i0[7] ), .A2(
        \SB2_2_10/i0_3 ), .A3(\SB2_2_10/i0_0 ), .ZN(
        \SB2_2_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_10/Component_Function_0/N3  ( .A1(\SB2_2_10/i0[10] ), .A2(
        \SB2_2_10/i0_4 ), .A3(\SB2_2_10/i0_3 ), .ZN(
        \SB2_2_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_10/Component_Function_0/N2  ( .A1(\SB2_2_10/i0[8] ), .A2(
        \SB2_2_10/i0[7] ), .A3(\SB2_2_10/i0[6] ), .ZN(
        \SB2_2_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_10/Component_Function_0/N1  ( .A1(\SB2_2_10/i0[10] ), .A2(
        \SB2_2_10/i0[9] ), .ZN(\SB2_2_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_10/Component_Function_1/N3  ( .A1(\SB2_2_10/i1_5 ), .A2(
        \SB2_2_10/i0[6] ), .A3(\SB2_2_10/i0[9] ), .ZN(
        \SB2_2_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_10/Component_Function_1/N2  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i1_7 ), .A3(\SB2_2_10/i0[8] ), .ZN(
        \SB2_2_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_10/Component_Function_1/N1  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i1[9] ), .ZN(\SB2_2_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_10/Component_Function_5/N4  ( .A1(\SB2_2_10/i0[9] ), .A2(
        \SB2_2_10/i0[6] ), .A3(\RI3[2][130] ), .ZN(
        \SB2_2_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_10/Component_Function_5/N2  ( .A1(\SB2_2_10/i0_0 ), .A2(
        \SB2_2_10/i0[6] ), .A3(\SB2_2_10/i0[10] ), .ZN(
        \SB2_2_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_10/Component_Function_5/N1  ( .A1(\SB2_2_10/i0_0 ), .A2(
        \SB2_2_10/i3[0] ), .ZN(\SB2_2_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_0/N4  ( .A1(\SB2_2_11/i0[7] ), .A2(
        \SB2_2_11/i0_3 ), .A3(\SB2_2_11/i0_0 ), .ZN(
        \SB2_2_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_11/Component_Function_0/N3  ( .A1(\SB2_2_11/i0[10] ), .A2(
        \SB2_2_11/i0_4 ), .A3(\SB2_2_11/i0_3 ), .ZN(
        \SB2_2_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_11/Component_Function_0/N2  ( .A1(\SB2_2_11/i0[8] ), .A2(
        \SB2_2_11/i0[7] ), .A3(\SB2_2_11/i0[6] ), .ZN(
        \SB2_2_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_11/Component_Function_0/N1  ( .A1(\SB2_2_11/i0[10] ), .A2(
        \SB2_2_11/i0[9] ), .ZN(\SB2_2_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_1/N4  ( .A1(\SB2_2_11/i1_7 ), .A2(
        \SB2_2_11/i0[8] ), .A3(\SB2_2_11/i0_4 ), .ZN(
        \SB2_2_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_11/Component_Function_1/N3  ( .A1(\SB2_2_11/i1_5 ), .A2(
        \SB2_2_11/i0[6] ), .A3(\SB2_2_11/i0[9] ), .ZN(
        \SB2_2_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_11/Component_Function_1/N2  ( .A1(\SB2_2_11/i0_3 ), .A2(
        \SB2_2_11/i1_7 ), .A3(\SB2_2_11/i0[8] ), .ZN(
        \SB2_2_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_11/Component_Function_1/N1  ( .A1(\SB2_2_11/i0_3 ), .A2(
        \SB2_2_11/i1[9] ), .ZN(\SB2_2_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_0/N3  ( .A1(\SB2_2_12/i0[10] ), .A2(
        \SB2_2_12/i0_4 ), .A3(\SB2_2_12/i0_3 ), .ZN(
        \SB2_2_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_12/Component_Function_0/N2  ( .A1(\SB2_2_12/i0[8] ), .A2(
        \SB2_2_12/i0[7] ), .A3(\SB2_2_12/i0[6] ), .ZN(
        \SB2_2_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_12/Component_Function_0/N1  ( .A1(\SB2_2_12/i0[10] ), .A2(
        \SB2_2_12/i0[9] ), .ZN(\SB2_2_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_1/N4  ( .A1(\SB2_2_12/i1_7 ), .A2(
        \SB2_2_12/i0[8] ), .A3(\SB2_2_12/i0_4 ), .ZN(
        \SB2_2_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_12/Component_Function_1/N3  ( .A1(\SB2_2_12/i1_5 ), .A2(
        \SB2_2_12/i0[6] ), .A3(\SB2_2_12/i0[9] ), .ZN(
        \SB2_2_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_12/Component_Function_1/N2  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i1_7 ), .A3(\SB2_2_12/i0[8] ), .ZN(
        \SB2_2_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_12/Component_Function_1/N1  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i1[9] ), .ZN(\SB2_2_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_5/N4  ( .A1(\SB2_2_12/i0[9] ), .A2(
        \SB2_2_12/i0[6] ), .A3(\SB2_2_12/i0_4 ), .ZN(
        \SB2_2_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_12/Component_Function_5/N3  ( .A1(\SB2_2_12/i1[9] ), .A2(
        \SB2_2_12/i0_4 ), .A3(\SB2_2_12/i0_3 ), .ZN(
        \SB2_2_12/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_12/Component_Function_5/N1  ( .A1(\SB2_2_12/i0_0 ), .A2(
        \SB2_2_12/i3[0] ), .ZN(\SB2_2_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_0/N4  ( .A1(\SB2_2_13/i0[7] ), .A2(
        \SB2_2_13/i0_3 ), .A3(\SB2_2_13/i0_0 ), .ZN(
        \SB2_2_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_13/Component_Function_0/N3  ( .A1(\SB2_2_13/i0[10] ), .A2(
        \SB2_2_13/i0_4 ), .A3(\SB2_2_13/i0_3 ), .ZN(
        \SB2_2_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_13/Component_Function_0/N2  ( .A1(\SB2_2_13/i0[8] ), .A2(
        \SB2_2_13/i0[7] ), .A3(\SB2_2_13/i0[6] ), .ZN(
        \SB2_2_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_13/Component_Function_0/N1  ( .A1(\SB2_2_13/i0[10] ), .A2(
        \SB2_2_13/i0[9] ), .ZN(\SB2_2_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_1/N4  ( .A1(\SB2_2_13/i1_7 ), .A2(
        \SB2_2_13/i0[8] ), .A3(\SB2_2_13/i0_4 ), .ZN(
        \SB2_2_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_13/Component_Function_1/N3  ( .A1(\SB2_2_13/i1_5 ), .A2(
        \SB2_2_13/i0[6] ), .A3(\SB2_2_13/i0[9] ), .ZN(
        \SB2_2_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_13/Component_Function_1/N2  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i1_7 ), .A3(\SB2_2_13/i0[8] ), .ZN(
        \SB2_2_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_13/Component_Function_1/N1  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i1[9] ), .ZN(\SB2_2_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_5/N4  ( .A1(\SB2_2_13/i0[9] ), .A2(
        \SB2_2_13/i0[6] ), .A3(\SB2_2_13/i0_4 ), .ZN(
        \SB2_2_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_13/Component_Function_5/N2  ( .A1(\SB2_2_13/i0_0 ), .A2(
        \SB2_2_13/i0[6] ), .A3(\SB2_2_13/i0[10] ), .ZN(
        \SB2_2_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_14/Component_Function_0/N3  ( .A1(\SB2_2_14/i0[10] ), .A2(
        \SB2_2_14/i0_4 ), .A3(\SB2_2_14/i0_3 ), .ZN(
        \SB2_2_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_14/Component_Function_0/N2  ( .A1(\SB2_2_14/i0[8] ), .A2(
        \SB2_2_14/i0[7] ), .A3(\SB2_2_14/i0[6] ), .ZN(
        \SB2_2_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_14/Component_Function_0/N1  ( .A1(\SB2_2_14/i0[10] ), .A2(
        \SB2_2_14/i0[9] ), .ZN(\SB2_2_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_1/N3  ( .A1(\SB2_2_14/i1_5 ), .A2(
        \SB2_2_14/i0[6] ), .A3(\SB2_2_14/i0[9] ), .ZN(
        \SB2_2_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_14/Component_Function_1/N2  ( .A1(\SB2_2_14/i0_3 ), .A2(
        \SB2_2_14/i1_7 ), .A3(\SB2_2_14/i0[8] ), .ZN(
        \SB2_2_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_14/Component_Function_1/N1  ( .A1(\SB2_2_14/i0_3 ), .A2(
        \SB2_2_14/i1[9] ), .ZN(\SB2_2_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_5/N3  ( .A1(\SB2_2_14/i1[9] ), .A2(
        \SB2_2_14/i0_4 ), .A3(\SB2_2_14/i0_3 ), .ZN(
        \SB2_2_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_14/Component_Function_5/N2  ( .A1(\SB2_2_14/i0_0 ), .A2(
        \SB2_2_14/i0[6] ), .A3(\SB2_2_14/i0[10] ), .ZN(
        \SB2_2_14/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_14/Component_Function_5/N1  ( .A1(\SB2_2_14/i0_0 ), .A2(
        \SB2_2_14/i3[0] ), .ZN(\SB2_2_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_15/Component_Function_0/N4  ( .A1(\SB2_2_15/i0[7] ), .A2(
        \SB2_2_15/i0_3 ), .A3(\SB2_2_15/i0_0 ), .ZN(
        \SB2_2_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_15/Component_Function_0/N3  ( .A1(\SB2_2_15/i0[10] ), .A2(
        \SB2_2_15/i0_4 ), .A3(\SB2_2_15/i0_3 ), .ZN(
        \SB2_2_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_15/Component_Function_0/N2  ( .A1(\SB2_2_15/i0[8] ), .A2(
        \SB2_2_15/i0[7] ), .A3(\SB2_2_15/i0[6] ), .ZN(
        \SB2_2_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_15/Component_Function_0/N1  ( .A1(\SB2_2_15/i0[10] ), .A2(
        \SB2_2_15/i0[9] ), .ZN(\SB2_2_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_15/Component_Function_1/N4  ( .A1(\SB2_2_15/i1_7 ), .A2(
        \SB2_2_15/i0[8] ), .A3(\SB2_2_15/i0_4 ), .ZN(
        \SB2_2_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_15/Component_Function_1/N3  ( .A1(\SB2_2_15/i1_5 ), .A2(
        \SB2_2_15/i0[6] ), .A3(\SB2_2_15/i0[9] ), .ZN(
        \SB2_2_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_15/Component_Function_1/N2  ( .A1(\SB2_2_15/i0_3 ), .A2(
        \SB2_2_15/i1_7 ), .A3(\SB2_2_15/i0[8] ), .ZN(
        \SB2_2_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_15/Component_Function_1/N1  ( .A1(\SB2_2_15/i0_3 ), .A2(
        \SB2_2_15/i1[9] ), .ZN(\SB2_2_15/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_15/Component_Function_5/N1  ( .A1(\SB2_2_15/i0_0 ), .A2(
        \SB2_2_15/i3[0] ), .ZN(\SB2_2_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_0/N4  ( .A1(\SB2_2_16/i0[7] ), .A2(
        \SB2_2_16/i0_3 ), .A3(\SB2_2_16/i0_0 ), .ZN(
        \SB2_2_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_16/Component_Function_0/N3  ( .A1(\SB2_2_16/i0[10] ), .A2(
        \SB2_2_16/i0_4 ), .A3(\SB2_2_16/i0_3 ), .ZN(
        \SB2_2_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_16/Component_Function_0/N2  ( .A1(\SB2_2_16/i0[8] ), .A2(
        \SB2_2_16/i0[7] ), .A3(\SB2_2_16/i0[6] ), .ZN(
        \SB2_2_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_16/Component_Function_0/N1  ( .A1(\SB2_2_16/i0[10] ), .A2(
        \SB2_2_16/i0[9] ), .ZN(\SB2_2_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_1/N3  ( .A1(\SB2_2_16/i1_5 ), .A2(
        \SB2_2_16/i0[6] ), .A3(\SB2_2_16/i0[9] ), .ZN(
        \SB2_2_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_16/Component_Function_1/N2  ( .A1(\SB2_2_16/i0_3 ), .A2(
        \SB2_2_16/i1_7 ), .A3(\SB2_2_16/i0[8] ), .ZN(
        \SB2_2_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_16/Component_Function_1/N1  ( .A1(\SB2_2_16/i0_3 ), .A2(
        \SB2_2_16/i1[9] ), .ZN(\SB2_2_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_16/Component_Function_5/N1  ( .A1(\SB2_2_16/i0_0 ), .A2(
        \SB2_2_16/i3[0] ), .ZN(\SB2_2_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_0/N3  ( .A1(\SB2_2_17/i0[10] ), .A2(
        \SB2_2_17/i0_4 ), .A3(\SB2_2_17/i0_3 ), .ZN(
        \SB2_2_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_17/Component_Function_0/N2  ( .A1(\SB2_2_17/i0[8] ), .A2(
        \SB2_2_17/i0[7] ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_17/Component_Function_0/N1  ( .A1(\SB2_2_17/i0[10] ), .A2(
        \SB2_2_17/i0[9] ), .ZN(\SB2_2_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_1/N4  ( .A1(\SB2_2_17/i1_7 ), .A2(
        \SB2_2_17/i0[8] ), .A3(\SB2_2_17/i0_4 ), .ZN(
        \SB2_2_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_17/Component_Function_1/N3  ( .A1(\SB2_2_17/i1_5 ), .A2(
        \SB2_2_17/i0[6] ), .A3(\SB2_2_17/i0[9] ), .ZN(
        \SB2_2_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_17/Component_Function_1/N2  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i1_7 ), .A3(\SB2_2_17/i0[8] ), .ZN(
        \SB2_2_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_17/Component_Function_1/N1  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i1[9] ), .ZN(\SB2_2_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_17/Component_Function_5/N1  ( .A1(\SB2_2_17/i0_0 ), .A2(
        \SB2_2_17/i3[0] ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_0/N4  ( .A1(\SB2_2_18/i0[7] ), .A2(
        \SB2_2_18/i0_3 ), .A3(\SB2_2_18/i0_0 ), .ZN(
        \SB2_2_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_18/Component_Function_0/N3  ( .A1(\SB2_2_18/i0[10] ), .A2(
        \SB2_2_18/i0_4 ), .A3(\SB2_2_18/i0_3 ), .ZN(
        \SB2_2_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_18/Component_Function_0/N2  ( .A1(\SB2_2_18/i0[8] ), .A2(
        \SB2_2_18/i0[7] ), .A3(\SB2_2_18/i0[6] ), .ZN(
        \SB2_2_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_18/Component_Function_0/N1  ( .A1(\SB2_2_18/i0[10] ), .A2(
        \SB2_2_18/i0[9] ), .ZN(\SB2_2_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_1/N4  ( .A1(\SB2_2_18/i1_7 ), .A2(
        \SB2_2_18/i0[8] ), .A3(\SB2_2_18/i0_4 ), .ZN(
        \SB2_2_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_18/Component_Function_1/N2  ( .A1(\SB2_2_18/i0_3 ), .A2(
        \SB2_2_18/i1_7 ), .A3(\SB2_2_18/i0[8] ), .ZN(
        \SB2_2_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_18/Component_Function_1/N1  ( .A1(\SB2_2_18/i0_3 ), .A2(
        \SB2_2_18/i1[9] ), .ZN(\SB2_2_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_5/N3  ( .A1(\SB2_2_18/i1[9] ), .A2(
        \SB2_2_18/i0_4 ), .A3(\SB2_2_18/i0_3 ), .ZN(
        \SB2_2_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_18/Component_Function_5/N2  ( .A1(\SB2_2_18/i0_0 ), .A2(
        \SB2_2_18/i0[6] ), .A3(\SB2_2_18/i0[10] ), .ZN(
        \SB2_2_18/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_18/Component_Function_5/N1  ( .A1(\SB2_2_18/i0_0 ), .A2(
        \SB2_2_18/i3[0] ), .ZN(\SB2_2_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_0/N4  ( .A1(\SB2_2_19/i0[7] ), .A2(
        \SB2_2_19/i0_3 ), .A3(\SB2_2_19/i0_0 ), .ZN(
        \SB2_2_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_19/Component_Function_0/N3  ( .A1(\SB2_2_19/i0[10] ), .A2(
        \SB2_2_19/i0_4 ), .A3(\SB2_2_19/i0_3 ), .ZN(
        \SB2_2_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_19/Component_Function_0/N2  ( .A1(\SB2_2_19/i0[8] ), .A2(
        \SB2_2_19/i0[7] ), .A3(\SB2_2_19/i0[6] ), .ZN(
        \SB2_2_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_19/Component_Function_0/N1  ( .A1(\SB2_2_19/i0[10] ), .A2(
        \SB2_2_19/i0[9] ), .ZN(\SB2_2_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_1/N4  ( .A1(\SB2_2_19/i1_7 ), .A2(
        \SB2_2_19/i0[8] ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_19/Component_Function_1/N3  ( .A1(\SB2_2_19/i1_5 ), .A2(
        \SB2_2_19/i0[6] ), .A3(\SB2_2_19/i0[9] ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_19/Component_Function_1/N2  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i1_7 ), .A3(\SB2_2_19/i0[8] ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_19/Component_Function_1/N1  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i1[9] ), .ZN(\SB2_2_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_5/N4  ( .A1(\SB2_2_19/i0[9] ), .A2(
        \SB2_2_19/i0[6] ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_19/Component_Function_5/N2  ( .A1(\SB2_2_19/i0_0 ), .A2(
        \SB2_2_19/i0[6] ), .A3(\SB2_2_19/i0[10] ), .ZN(
        \SB2_2_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_19/Component_Function_5/N1  ( .A1(\SB2_2_19/i0_0 ), .A2(
        \SB2_2_19/i3[0] ), .ZN(\SB2_2_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_0/N4  ( .A1(\SB2_2_20/i0[7] ), .A2(
        \SB2_2_20/i0_3 ), .A3(\SB2_2_20/i0_0 ), .ZN(
        \SB2_2_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_20/Component_Function_0/N3  ( .A1(\SB2_2_20/i0[10] ), .A2(
        \SB2_2_20/i0_4 ), .A3(\SB2_2_20/i0_3 ), .ZN(
        \SB2_2_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_20/Component_Function_0/N2  ( .A1(\SB2_2_20/i0[8] ), .A2(
        \SB2_2_20/i0[7] ), .A3(\SB2_2_20/i0[6] ), .ZN(
        \SB2_2_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_20/Component_Function_0/N1  ( .A1(\SB2_2_20/i0[10] ), .A2(
        \SB2_2_20/i0[9] ), .ZN(\SB2_2_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_1/N4  ( .A1(\SB2_2_20/i1_7 ), .A2(
        \SB2_2_20/i0[8] ), .A3(\SB2_2_20/i0_4 ), .ZN(
        \SB2_2_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_20/Component_Function_1/N3  ( .A1(\SB2_2_20/i1_5 ), .A2(
        \SB2_2_20/i0[6] ), .A3(\SB2_2_20/i0[9] ), .ZN(
        \SB2_2_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_20/Component_Function_1/N2  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i1_7 ), .A3(\SB2_2_20/i0[8] ), .ZN(
        \SB2_2_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_20/Component_Function_1/N1  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i1[9] ), .ZN(\SB2_2_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_5/N3  ( .A1(\SB2_2_20/i1[9] ), .A2(
        \SB2_2_20/i0_4 ), .A3(\SB2_2_20/i0_3 ), .ZN(
        \SB2_2_20/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_20/Component_Function_5/N1  ( .A1(\SB2_2_20/i0_0 ), .A2(
        \SB2_2_20/i3[0] ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_0/N4  ( .A1(\SB2_2_21/i0[7] ), .A2(
        \SB2_2_21/i0_3 ), .A3(\SB2_2_21/i0_0 ), .ZN(
        \SB2_2_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_21/Component_Function_0/N3  ( .A1(\SB2_2_21/i0[10] ), .A2(
        \SB2_2_21/i0_4 ), .A3(\SB2_2_21/i0_3 ), .ZN(
        \SB2_2_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_21/Component_Function_0/N2  ( .A1(\SB2_2_21/i0[8] ), .A2(
        \SB2_2_21/i0[7] ), .A3(\SB2_2_21/i0[6] ), .ZN(
        \SB2_2_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_21/Component_Function_0/N1  ( .A1(\SB2_2_21/i0[10] ), .A2(
        \SB2_2_21/i0[9] ), .ZN(\SB2_2_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_1/N4  ( .A1(\SB2_2_21/i1_7 ), .A2(
        \SB2_2_21/i0[8] ), .A3(\SB2_2_21/i0_4 ), .ZN(
        \SB2_2_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_21/Component_Function_1/N3  ( .A1(\SB2_2_21/i1_5 ), .A2(
        \SB2_2_21/i0[6] ), .A3(\SB2_2_21/i0[9] ), .ZN(
        \SB2_2_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_21/Component_Function_1/N2  ( .A1(\SB2_2_21/i0_3 ), .A2(
        \SB2_2_21/i1_7 ), .A3(\SB2_2_21/i0[8] ), .ZN(
        \SB2_2_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_21/Component_Function_1/N1  ( .A1(\SB2_2_21/i0_3 ), .A2(
        \SB2_2_21/i1[9] ), .ZN(\SB2_2_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_5/N3  ( .A1(\SB2_2_21/i1[9] ), .A2(
        \SB2_2_21/i0_4 ), .A3(\SB2_2_21/i0_3 ), .ZN(
        \SB2_2_21/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_21/Component_Function_5/N1  ( .A1(\SB2_2_21/i0_0 ), .A2(
        \SB2_2_21/i3[0] ), .ZN(\SB2_2_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_22/Component_Function_0/N4  ( .A1(\SB2_2_22/i0[7] ), .A2(
        \SB2_2_22/i0_3 ), .A3(\SB2_2_22/i0_0 ), .ZN(
        \SB2_2_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_22/Component_Function_0/N3  ( .A1(\SB2_2_22/i0[10] ), .A2(
        \SB2_2_22/i0_4 ), .A3(\SB2_2_22/i0_3 ), .ZN(
        \SB2_2_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_22/Component_Function_0/N2  ( .A1(\SB2_2_22/i0[8] ), .A2(
        \SB2_2_22/i0[7] ), .A3(\SB2_2_22/i0[6] ), .ZN(
        \SB2_2_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_22/Component_Function_0/N1  ( .A1(\SB2_2_22/i0[10] ), .A2(
        \SB2_2_22/i0[9] ), .ZN(\SB2_2_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_22/Component_Function_1/N3  ( .A1(\SB2_2_22/i1_5 ), .A2(
        \SB2_2_22/i0[6] ), .A3(\SB2_2_22/i0[9] ), .ZN(
        \SB2_2_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_22/Component_Function_1/N2  ( .A1(\SB2_2_22/i0_3 ), .A2(
        \SB2_2_22/i1_7 ), .A3(\SB2_2_22/i0[8] ), .ZN(
        \SB2_2_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_22/Component_Function_1/N1  ( .A1(\SB2_2_22/i0_3 ), .A2(
        \SB2_2_22/i1[9] ), .ZN(\SB2_2_22/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_22/Component_Function_5/N1  ( .A1(\SB2_2_22/i0_0 ), .A2(
        \SB2_2_22/i3[0] ), .ZN(\SB2_2_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_23/Component_Function_0/N4  ( .A1(\SB2_2_23/i0[7] ), .A2(
        \SB2_2_23/i0_3 ), .A3(\SB2_2_23/i0_0 ), .ZN(
        \SB2_2_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_23/Component_Function_0/N3  ( .A1(\SB2_2_23/i0[10] ), .A2(
        \SB2_2_23/i0_4 ), .A3(\SB2_2_23/i0_3 ), .ZN(
        \SB2_2_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_23/Component_Function_0/N2  ( .A1(\SB2_2_23/i0[8] ), .A2(
        \SB2_2_23/i0[7] ), .A3(\SB2_2_23/i0[6] ), .ZN(
        \SB2_2_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_23/Component_Function_0/N1  ( .A1(\SB2_2_23/i0[10] ), .A2(
        \SB2_2_23/i0[9] ), .ZN(\SB2_2_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_23/Component_Function_1/N4  ( .A1(\SB2_2_23/i1_7 ), .A2(
        \SB2_2_23/i0[8] ), .A3(\SB2_2_23/i0_4 ), .ZN(
        \SB2_2_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_23/Component_Function_1/N3  ( .A1(\SB2_2_23/i1_5 ), .A2(
        \SB2_2_23/i0[6] ), .A3(\SB2_2_23/i0[9] ), .ZN(
        \SB2_2_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_23/Component_Function_1/N2  ( .A1(\SB2_2_23/i0_3 ), .A2(
        \SB2_2_23/i1_7 ), .A3(\SB2_2_23/i0[8] ), .ZN(
        \SB2_2_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_23/Component_Function_1/N1  ( .A1(\SB2_2_23/i0_3 ), .A2(
        \SB2_2_23/i1[9] ), .ZN(\SB2_2_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_23/Component_Function_5/N4  ( .A1(\SB2_2_23/i0[9] ), .A2(
        \SB2_2_23/i0[6] ), .A3(\SB2_2_23/i0_4 ), .ZN(
        \SB2_2_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_23/Component_Function_5/N2  ( .A1(\SB2_2_23/i0_0 ), .A2(
        \SB2_2_23/i0[6] ), .A3(\SB2_2_23/i0[10] ), .ZN(
        \SB2_2_23/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_23/Component_Function_5/N1  ( .A1(\SB2_2_23/i0_0 ), .A2(
        \SB2_2_23/i3[0] ), .ZN(\SB2_2_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_0/N3  ( .A1(\SB2_2_24/i0[10] ), .A2(
        \SB2_2_24/i0_4 ), .A3(\SB2_2_24/i0_3 ), .ZN(
        \SB2_2_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_24/Component_Function_0/N2  ( .A1(\SB2_2_24/i0[8] ), .A2(
        \SB2_2_24/i0[7] ), .A3(\SB2_2_24/i0[6] ), .ZN(
        \SB2_2_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_24/Component_Function_0/N1  ( .A1(\SB2_2_24/i0[10] ), .A2(
        \SB2_2_24/i0[9] ), .ZN(\SB2_2_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_1/N4  ( .A1(\SB2_2_24/i1_7 ), .A2(
        \SB2_2_24/i0[8] ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_24/Component_Function_1/N3  ( .A1(\SB2_2_24/i1_5 ), .A2(
        \SB2_2_24/i0[6] ), .A3(\SB2_2_24/i0[9] ), .ZN(
        \SB2_2_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_24/Component_Function_1/N2  ( .A1(\SB2_2_24/i0_3 ), .A2(
        \SB2_2_24/i1_7 ), .A3(\SB2_2_24/i0[8] ), .ZN(
        \SB2_2_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_24/Component_Function_1/N1  ( .A1(\SB2_2_24/i0_3 ), .A2(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_5/N4  ( .A1(\SB2_2_24/i0[9] ), .A2(
        \SB2_2_24/i0[6] ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_24/Component_Function_5/N2  ( .A1(\SB2_2_24/i0_0 ), .A2(
        \SB2_2_24/i0[6] ), .A3(\SB2_2_24/i0[10] ), .ZN(
        \SB2_2_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_24/Component_Function_5/N1  ( .A1(\SB2_2_24/i0_0 ), .A2(
        \SB2_2_24/i3[0] ), .ZN(\SB2_2_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_0/N4  ( .A1(\SB2_2_25/i0[7] ), .A2(
        \SB2_2_25/i0_3 ), .A3(\SB2_2_25/i0_0 ), .ZN(
        \SB2_2_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_25/Component_Function_0/N3  ( .A1(\SB2_2_25/i0[10] ), .A2(
        \SB2_2_25/i0_4 ), .A3(\SB2_2_25/i0_3 ), .ZN(
        \SB2_2_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_25/Component_Function_0/N2  ( .A1(\SB2_2_25/i0[8] ), .A2(
        \SB2_2_25/i0[7] ), .A3(\SB2_2_25/i0[6] ), .ZN(
        \SB2_2_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_25/Component_Function_0/N1  ( .A1(\SB2_2_25/i0[10] ), .A2(
        \SB2_2_25/i0[9] ), .ZN(\SB2_2_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_1/N3  ( .A1(\SB2_2_25/i1_5 ), .A2(
        \SB2_2_25/i0[6] ), .A3(\SB2_2_25/i0[9] ), .ZN(
        \SB2_2_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_25/Component_Function_1/N2  ( .A1(\SB2_2_25/i0_3 ), .A2(
        \SB2_2_25/i1_7 ), .A3(\SB2_2_25/i0[8] ), .ZN(
        \SB2_2_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_25/Component_Function_1/N1  ( .A1(\SB2_2_25/i0_3 ), .A2(
        \SB2_2_25/i1[9] ), .ZN(\SB2_2_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_5/N2  ( .A1(\SB2_2_25/i0_0 ), .A2(
        \SB2_2_25/i0[6] ), .A3(\SB2_2_25/i0[10] ), .ZN(
        \SB2_2_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_25/Component_Function_5/N1  ( .A1(\SB2_2_25/i0_0 ), .A2(
        \SB2_2_25/i3[0] ), .ZN(\SB2_2_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_0/N4  ( .A1(\SB2_2_26/i0[7] ), .A2(
        \SB2_2_26/i0_3 ), .A3(\SB2_2_26/i0_0 ), .ZN(
        \SB2_2_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_26/Component_Function_0/N3  ( .A1(\SB2_2_26/i0[10] ), .A2(
        \SB2_2_26/i0_4 ), .A3(\SB2_2_26/i0_3 ), .ZN(
        \SB2_2_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_26/Component_Function_0/N2  ( .A1(\SB2_2_26/i0[8] ), .A2(
        \SB2_2_26/i0[7] ), .A3(\SB2_2_26/i0[6] ), .ZN(
        \SB2_2_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_26/Component_Function_0/N1  ( .A1(\SB2_2_26/i0[10] ), .A2(
        \SB2_2_26/i0[9] ), .ZN(\SB2_2_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_1/N4  ( .A1(\SB2_2_26/i1_7 ), .A2(
        \SB2_2_26/i0[8] ), .A3(\SB2_2_26/i0_4 ), .ZN(
        \SB2_2_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_26/Component_Function_1/N3  ( .A1(\SB2_2_26/i1_5 ), .A2(
        \SB2_2_26/i0[6] ), .A3(\SB2_2_26/i0[9] ), .ZN(
        \SB2_2_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_26/Component_Function_1/N2  ( .A1(\SB2_2_26/i0_3 ), .A2(
        \SB2_2_26/i1_7 ), .A3(\SB2_2_26/i0[8] ), .ZN(
        \SB2_2_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_26/Component_Function_1/N1  ( .A1(\SB2_2_26/i1[9] ), .A2(
        \SB2_2_26/i0_3 ), .ZN(\SB2_2_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_5/N4  ( .A1(\SB2_2_26/i0[9] ), .A2(
        \SB2_2_26/i0[6] ), .A3(\RI3[2][34] ), .ZN(
        \SB2_2_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_26/Component_Function_5/N2  ( .A1(\SB2_2_26/i0_0 ), .A2(
        \SB2_2_26/i0[6] ), .A3(\SB2_2_26/i0[10] ), .ZN(
        \SB2_2_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_27/Component_Function_0/N4  ( .A1(\SB2_2_27/i0[7] ), .A2(
        \SB2_2_27/i0_3 ), .A3(\SB2_2_27/i0_0 ), .ZN(
        \SB2_2_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_27/Component_Function_0/N3  ( .A1(\SB2_2_27/i0[10] ), .A2(
        \SB2_2_27/i0_4 ), .A3(\SB2_2_27/i0_3 ), .ZN(
        \SB2_2_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_27/Component_Function_0/N2  ( .A1(\SB2_2_27/i0[8] ), .A2(
        \SB2_2_27/i0[7] ), .A3(\SB2_2_27/i0[6] ), .ZN(
        \SB2_2_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_27/Component_Function_0/N1  ( .A1(\SB2_2_27/i0[10] ), .A2(
        \SB2_2_27/i0[9] ), .ZN(\SB2_2_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_27/Component_Function_1/N4  ( .A1(\SB2_2_27/i1_7 ), .A2(
        \SB2_2_27/i0[8] ), .A3(\SB2_2_27/i0_4 ), .ZN(
        \SB2_2_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_27/Component_Function_1/N3  ( .A1(\SB2_2_27/i1_5 ), .A2(
        \SB2_2_27/i0[6] ), .A3(\SB2_2_27/i0[9] ), .ZN(
        \SB2_2_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_27/Component_Function_1/N2  ( .A1(\SB2_2_27/i0_3 ), .A2(
        \SB2_2_27/i1_7 ), .A3(\SB2_2_27/i0[8] ), .ZN(
        \SB2_2_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_27/Component_Function_1/N1  ( .A1(\SB2_2_27/i0_3 ), .A2(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_27/Component_Function_5/N1  ( .A1(\SB2_2_27/i0_0 ), .A2(
        \SB2_2_27/i3[0] ), .ZN(\SB2_2_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_0/N3  ( .A1(\SB2_2_28/i0[10] ), .A2(
        \SB2_2_28/i0_4 ), .A3(\SB2_2_28/i0_3 ), .ZN(
        \SB2_2_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_28/Component_Function_0/N2  ( .A1(\SB2_2_28/i0[8] ), .A2(
        \SB2_2_28/i0[7] ), .A3(\SB2_2_28/i0[6] ), .ZN(
        \SB2_2_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_28/Component_Function_0/N1  ( .A1(\SB2_2_28/i0[10] ), .A2(
        \SB2_2_28/i0[9] ), .ZN(\SB2_2_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_1/N4  ( .A1(\SB2_2_28/i1_7 ), .A2(
        \SB2_2_28/i0[8] ), .A3(\SB2_2_28/i0_4 ), .ZN(
        \SB2_2_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_28/Component_Function_1/N3  ( .A1(\SB2_2_28/i1_5 ), .A2(
        \SB2_2_28/i0[6] ), .A3(\SB2_2_28/i0[9] ), .ZN(
        \SB2_2_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_28/Component_Function_1/N2  ( .A1(\SB2_2_28/i0_3 ), .A2(
        \SB2_2_28/i1_7 ), .A3(\SB2_2_28/i0[8] ), .ZN(
        \SB2_2_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_28/Component_Function_1/N1  ( .A1(\SB2_2_28/i0_3 ), .A2(
        \SB2_2_28/i1[9] ), .ZN(\SB2_2_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_5/N4  ( .A1(\SB2_2_28/i0[9] ), .A2(
        \SB2_2_28/i0[6] ), .A3(\SB2_2_28/i0_4 ), .ZN(
        \SB2_2_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_28/Component_Function_5/N3  ( .A1(\SB2_2_28/i1[9] ), .A2(
        \SB2_2_28/i0_4 ), .A3(\SB2_2_28/i0_3 ), .ZN(
        \SB2_2_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_28/Component_Function_5/N2  ( .A1(\SB2_2_28/i0_0 ), .A2(
        \SB2_2_28/i0[6] ), .A3(\SB2_2_28/i0[10] ), .ZN(
        \SB2_2_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_28/Component_Function_5/N1  ( .A1(\SB2_2_28/i0_0 ), .A2(
        \SB2_2_28/i3[0] ), .ZN(\SB2_2_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_0/N4  ( .A1(\SB2_2_29/i0[7] ), .A2(
        \SB2_2_29/i0_3 ), .A3(\SB2_2_29/i0_0 ), .ZN(
        \SB2_2_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_29/Component_Function_0/N3  ( .A1(\SB2_2_29/i0[10] ), .A2(
        \SB2_2_29/i0_4 ), .A3(\SB2_2_29/i0_3 ), .ZN(
        \SB2_2_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_29/Component_Function_0/N2  ( .A1(\SB2_2_29/i0[8] ), .A2(
        \SB2_2_29/i0[7] ), .A3(\SB2_2_29/i0[6] ), .ZN(
        \SB2_2_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_29/Component_Function_0/N1  ( .A1(\SB2_2_29/i0[10] ), .A2(
        \SB2_2_29/i0[9] ), .ZN(\SB2_2_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_1/N4  ( .A1(\SB2_2_29/i1_7 ), .A2(
        \SB2_2_29/i0[8] ), .A3(\SB2_2_29/i0_4 ), .ZN(
        \SB2_2_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_29/Component_Function_1/N3  ( .A1(\SB2_2_29/i1_5 ), .A2(
        \SB2_2_29/i0[6] ), .A3(\SB2_2_29/i0[9] ), .ZN(
        \SB2_2_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_29/Component_Function_1/N2  ( .A1(\SB2_2_29/i0_3 ), .A2(
        \SB2_2_29/i1_7 ), .A3(\SB2_2_29/i0[8] ), .ZN(
        \SB2_2_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_29/Component_Function_1/N1  ( .A1(\SB2_2_29/i0_3 ), .A2(
        \SB2_2_29/i1[9] ), .ZN(\SB2_2_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_5/N2  ( .A1(\SB2_2_29/i0_0 ), .A2(
        \SB2_2_29/i0[6] ), .A3(\SB2_2_29/i0[10] ), .ZN(
        \SB2_2_29/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_29/Component_Function_5/N1  ( .A1(\SB2_2_29/i0_0 ), .A2(
        \SB2_2_29/i3[0] ), .ZN(\SB2_2_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_0/N4  ( .A1(\SB2_2_30/i0[7] ), .A2(
        \SB2_2_30/i0_3 ), .A3(\SB2_2_30/i0_0 ), .ZN(
        \SB2_2_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_30/Component_Function_0/N3  ( .A1(\SB2_2_30/i0[10] ), .A2(
        \SB2_2_30/i0_4 ), .A3(\SB2_2_30/i0_3 ), .ZN(
        \SB2_2_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_30/Component_Function_0/N2  ( .A1(\SB2_2_30/i0[8] ), .A2(
        \SB2_2_30/i0[7] ), .A3(\SB2_2_30/i0[6] ), .ZN(
        \SB2_2_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_30/Component_Function_0/N1  ( .A1(\SB2_2_30/i0[10] ), .A2(
        \SB2_2_30/i0[9] ), .ZN(\SB2_2_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_1/N4  ( .A1(\SB2_2_30/i1_7 ), .A2(
        \SB2_2_30/i0[8] ), .A3(\SB2_2_30/i0_4 ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_30/Component_Function_1/N3  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0[6] ), .A3(\SB2_2_30/i0[9] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_30/Component_Function_1/N2  ( .A1(\SB2_2_30/i0_3 ), .A2(
        \SB2_2_30/i1_7 ), .A3(\SB2_2_30/i0[8] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_30/Component_Function_1/N1  ( .A1(\SB2_2_30/i0_3 ), .A2(
        n2118), .ZN(\SB2_2_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_5/N3  ( .A1(n2118), .A2(
        \SB2_2_30/i0_4 ), .A3(\SB2_2_30/i0_3 ), .ZN(
        \SB2_2_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_30/Component_Function_5/N2  ( .A1(\SB2_2_30/i0_0 ), .A2(
        \SB2_2_30/i0[6] ), .A3(\SB2_2_30/i0[10] ), .ZN(
        \SB2_2_30/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_31/Component_Function_0/N4  ( .A1(\SB2_2_31/i0[7] ), .A2(
        \SB2_2_31/i0_3 ), .A3(\SB2_2_31/i0_0 ), .ZN(
        \SB2_2_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_31/Component_Function_0/N3  ( .A1(\SB2_2_31/i0[10] ), .A2(
        \SB2_2_31/i0_4 ), .A3(\SB2_2_31/i0_3 ), .ZN(
        \SB2_2_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_31/Component_Function_0/N2  ( .A1(\SB2_2_31/i0[8] ), .A2(
        \SB2_2_31/i0[7] ), .A3(\SB2_2_31/i0[6] ), .ZN(
        \SB2_2_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_31/Component_Function_0/N1  ( .A1(\SB2_2_31/i0[10] ), .A2(
        \SB2_2_31/i0[9] ), .ZN(\SB2_2_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_31/Component_Function_1/N3  ( .A1(\SB2_2_31/i1_5 ), .A2(
        \SB2_2_31/i0[6] ), .A3(\SB2_2_31/i0[9] ), .ZN(
        \SB2_2_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_31/Component_Function_1/N2  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i1_7 ), .A3(\SB2_2_31/i0[8] ), .ZN(
        \SB2_2_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_31/Component_Function_1/N1  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i1[9] ), .ZN(\SB2_2_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_31/Component_Function_5/N4  ( .A1(\RI3[2][0] ), .A2(
        \SB2_2_31/i0[6] ), .A3(\SB2_2_31/i0_4 ), .ZN(
        \SB2_2_31/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_31/Component_Function_5/N1  ( .A1(\SB2_2_31/i0_0 ), .A2(
        \SB2_2_31/i3[0] ), .ZN(\SB2_2_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_0/N4  ( .A1(\SB1_3_0/i0[7] ), .A2(n809), 
        .A3(\SB1_3_0/i0_0 ), .ZN(\SB1_3_0/Component_Function_0/NAND4_in[3] )
         );
  NAND3_X1 \SB1_3_0/Component_Function_0/N2  ( .A1(\SB1_3_0/i0[8] ), .A2(
        \SB1_3_0/i0[7] ), .A3(\SB1_3_0/i0[6] ), .ZN(
        \SB1_3_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_0/Component_Function_0/N1  ( .A1(\SB1_3_0/i0[10] ), .A2(
        \SB1_3_0/i0[9] ), .ZN(\SB1_3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_1/N4  ( .A1(\SB1_3_0/i1_7 ), .A2(
        \SB1_3_0/i0[8] ), .A3(\SB1_3_0/i0_4 ), .ZN(
        \SB1_3_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_0/Component_Function_1/N3  ( .A1(\SB1_3_0/i1_5 ), .A2(
        \SB1_3_0/i0[6] ), .A3(\SB1_3_0/i0[9] ), .ZN(
        \SB1_3_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_0/Component_Function_1/N2  ( .A1(n809), .A2(\SB1_3_0/i1_7 ), 
        .A3(\SB1_3_0/i0[8] ), .ZN(\SB1_3_0/Component_Function_1/NAND4_in[1] )
         );
  NAND2_X1 \SB1_3_0/Component_Function_1/N1  ( .A1(n809), .A2(\SB1_3_0/i1[9] ), 
        .ZN(\SB1_3_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_5/N4  ( .A1(\SB1_3_0/i0[9] ), .A2(
        \SB1_3_0/i0[6] ), .A3(\SB1_3_0/i0_4 ), .ZN(
        \SB1_3_0/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_3_0/Component_Function_5/N1  ( .A1(\SB1_3_0/i0_0 ), .A2(
        \SB1_3_0/i3[0] ), .ZN(\SB1_3_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_0/N4  ( .A1(\SB1_3_1/i0[7] ), .A2(
        \SB1_3_1/i0_3 ), .A3(\SB1_3_1/i0_0 ), .ZN(
        \SB1_3_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_1/Component_Function_0/N3  ( .A1(\SB1_3_1/i0[10] ), .A2(
        \SB1_3_1/i0_4 ), .A3(\SB1_3_1/i0_3 ), .ZN(
        \SB1_3_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_1/Component_Function_0/N2  ( .A1(\SB1_3_1/i0[8] ), .A2(
        \SB1_3_1/i0[7] ), .A3(\SB1_3_1/i0[6] ), .ZN(
        \SB1_3_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_1/Component_Function_0/N1  ( .A1(\SB1_3_1/i0[10] ), .A2(
        \SB1_3_1/i0[9] ), .ZN(\SB1_3_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_1/N4  ( .A1(\SB1_3_1/i1_7 ), .A2(
        \SB1_3_1/i0[8] ), .A3(\SB1_3_1/i0_4 ), .ZN(
        \SB1_3_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_1/Component_Function_1/N3  ( .A1(\SB1_3_1/i1_5 ), .A2(
        \SB1_3_1/i0[6] ), .A3(\SB1_3_1/i0[9] ), .ZN(
        \SB1_3_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_1/Component_Function_1/N2  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i1_7 ), .A3(\SB1_3_1/i0[8] ), .ZN(
        \SB1_3_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_1/Component_Function_1/N1  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i1[9] ), .ZN(\SB1_3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_5/N4  ( .A1(\SB1_3_1/i0[9] ), .A2(
        \SB1_3_1/i0[6] ), .A3(\SB1_3_1/i0_4 ), .ZN(
        \SB1_3_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_1/Component_Function_5/N2  ( .A1(\SB1_3_1/i0_0 ), .A2(
        \SB1_3_1/i0[6] ), .A3(\SB1_3_1/i0[10] ), .ZN(
        \SB1_3_1/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_1/Component_Function_5/N1  ( .A1(\SB1_3_1/i0_0 ), .A2(
        \SB1_3_1/i3[0] ), .ZN(\SB1_3_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_0/N4  ( .A1(\SB1_3_2/i0[7] ), .A2(
        \SB1_3_2/i0_3 ), .A3(\SB1_3_2/i0_0 ), .ZN(
        \SB1_3_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_2/Component_Function_0/N3  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i0_4 ), .A3(\SB1_3_2/i0[10] ), .ZN(
        \SB1_3_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_2/Component_Function_0/N2  ( .A1(\SB1_3_2/i0[8] ), .A2(
        \SB1_3_2/i0[7] ), .A3(\SB1_3_2/i0[6] ), .ZN(
        \SB1_3_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_2/Component_Function_0/N1  ( .A1(\SB1_3_2/i0[10] ), .A2(
        \SB1_3_2/i0[9] ), .ZN(\SB1_3_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_1/N4  ( .A1(\SB1_3_2/i1_7 ), .A2(
        \SB1_3_2/i0[8] ), .A3(\SB1_3_2/i0_4 ), .ZN(
        \SB1_3_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_2/Component_Function_1/N3  ( .A1(\SB1_3_2/i1_5 ), .A2(
        \SB1_3_2/i0[6] ), .A3(\SB1_3_2/i0[9] ), .ZN(
        \SB1_3_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_2/Component_Function_1/N2  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i1_7 ), .A3(\SB1_3_2/i0[8] ), .ZN(
        \SB1_3_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_2/Component_Function_1/N1  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i1[9] ), .ZN(\SB1_3_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_5/N2  ( .A1(\SB1_3_2/i0_0 ), .A2(
        \SB1_3_2/i0[6] ), .A3(\SB1_3_2/i0[10] ), .ZN(
        \SB1_3_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_2/Component_Function_5/N1  ( .A1(\SB1_3_2/i0_0 ), .A2(
        \SB1_3_2/i3[0] ), .ZN(\SB1_3_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N4  ( .A1(\SB1_3_3/i0[7] ), .A2(
        \SB1_3_3/i0_3 ), .A3(\SB1_3_3/i0_0 ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N3  ( .A1(\SB1_3_3/i0[10] ), .A2(
        \SB1_3_3/i0_4 ), .A3(\SB1_3_3/i0_3 ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N2  ( .A1(\SB1_3_3/i0[8] ), .A2(
        \SB1_3_3/i0[7] ), .A3(\SB1_3_3/i0[6] ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_3/Component_Function_0/N1  ( .A1(\SB1_3_3/i0[10] ), .A2(
        \SB1_3_3/i0[9] ), .ZN(\SB1_3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_1/N3  ( .A1(\SB1_3_3/i1_5 ), .A2(
        \SB1_3_3/i0[6] ), .A3(\SB1_3_3/i0[9] ), .ZN(
        \SB1_3_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_3/Component_Function_1/N2  ( .A1(\SB1_3_3/i0_3 ), .A2(
        \SB1_3_3/i1_7 ), .A3(\SB1_3_3/i0[8] ), .ZN(
        \SB1_3_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_3/Component_Function_1/N1  ( .A1(\SB1_3_3/i0_3 ), .A2(
        \SB1_3_3/i1[9] ), .ZN(\SB1_3_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_5/N4  ( .A1(\SB1_3_3/i0[9] ), .A2(
        \SB1_3_3/i0[6] ), .A3(\SB1_3_3/i0_4 ), .ZN(
        \SB1_3_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_3/Component_Function_5/N2  ( .A1(\SB1_3_3/i0_0 ), .A2(
        \SB1_3_3/i0[6] ), .A3(\SB1_3_3/i0[10] ), .ZN(
        \SB1_3_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_3/Component_Function_5/N1  ( .A1(\SB1_3_3/i0_0 ), .A2(
        \SB1_3_3/i3[0] ), .ZN(\SB1_3_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_0/N4  ( .A1(\SB1_3_4/i0[7] ), .A2(
        \SB1_3_4/i0_3 ), .A3(\SB1_3_4/i0_0 ), .ZN(
        \SB1_3_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_4/Component_Function_0/N3  ( .A1(\SB1_3_4/i0[10] ), .A2(
        \SB1_3_4/i0_4 ), .A3(\SB1_3_4/i0_3 ), .ZN(
        \SB1_3_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_4/Component_Function_0/N2  ( .A1(\SB1_3_4/i0[8] ), .A2(
        \SB1_3_4/i0[7] ), .A3(\SB1_3_4/i0[6] ), .ZN(
        \SB1_3_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_4/Component_Function_0/N1  ( .A1(\SB1_3_4/i0[10] ), .A2(
        \SB1_3_4/i0[9] ), .ZN(\SB1_3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_1/N4  ( .A1(\SB1_3_4/i1_7 ), .A2(
        \SB1_3_4/i0[8] ), .A3(\SB1_3_4/i0_4 ), .ZN(
        \SB1_3_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_4/Component_Function_1/N3  ( .A1(\SB1_3_4/i1_5 ), .A2(
        \SB1_3_4/i0[6] ), .A3(\SB1_3_4/i0[9] ), .ZN(
        \SB1_3_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_4/Component_Function_1/N2  ( .A1(\SB1_3_4/i0_3 ), .A2(
        \SB1_3_4/i1_7 ), .A3(\SB1_3_4/i0[8] ), .ZN(
        \SB1_3_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_4/Component_Function_1/N1  ( .A1(\SB1_3_4/i0_3 ), .A2(
        \SB1_3_4/i1[9] ), .ZN(\SB1_3_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_5/N4  ( .A1(\SB1_3_4/i0[9] ), .A2(
        \SB1_3_4/i0[6] ), .A3(\SB1_3_4/i0_4 ), .ZN(
        \SB1_3_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_4/Component_Function_5/N2  ( .A1(\SB1_3_4/i0_0 ), .A2(
        \SB1_3_4/i0[6] ), .A3(\SB1_3_4/i0[10] ), .ZN(
        \SB1_3_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_4/Component_Function_5/N1  ( .A1(\SB1_3_4/i0_0 ), .A2(
        \SB1_3_4/i3[0] ), .ZN(\SB1_3_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N4  ( .A1(\SB1_3_5/i0[7] ), .A2(
        \SB1_3_5/i0_3 ), .A3(\SB1_3_5/i0_0 ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N3  ( .A1(\SB1_3_5/i0[10] ), .A2(
        \SB1_3_5/i0_4 ), .A3(\SB1_3_5/i0_3 ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N2  ( .A1(\SB1_3_5/i0[8] ), .A2(
        \SB1_3_5/i0[7] ), .A3(\SB1_3_5/i0[6] ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_5/Component_Function_0/N1  ( .A1(\SB1_3_5/i0[10] ), .A2(
        \SB1_3_5/i0[9] ), .ZN(\SB1_3_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_1/N4  ( .A1(\SB1_3_5/i1_7 ), .A2(
        \SB1_3_5/i0[8] ), .A3(\SB1_3_5/i0_4 ), .ZN(
        \SB1_3_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_5/Component_Function_1/N3  ( .A1(\SB1_3_5/i1_5 ), .A2(
        \SB1_3_5/i0[6] ), .A3(\SB1_3_5/i0[9] ), .ZN(
        \SB1_3_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_5/Component_Function_1/N2  ( .A1(\SB1_3_5/i0_3 ), .A2(
        \SB1_3_5/i1_7 ), .A3(\SB1_3_5/i0[8] ), .ZN(
        \SB1_3_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_5/Component_Function_1/N1  ( .A1(\SB1_3_5/i0_3 ), .A2(
        \SB1_3_5/i1[9] ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_5/Component_Function_5/N1  ( .A1(\SB1_3_5/i0_0 ), .A2(
        \SB1_3_5/i3[0] ), .ZN(\SB1_3_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_0/N4  ( .A1(\SB1_3_6/i0[7] ), .A2(
        \SB1_3_6/i0_3 ), .A3(\SB1_3_6/i0_0 ), .ZN(
        \SB1_3_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_6/Component_Function_0/N3  ( .A1(\SB1_3_6/i0[10] ), .A2(
        \SB1_3_6/i0_4 ), .A3(\SB1_3_6/i0_3 ), .ZN(
        \SB1_3_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_6/Component_Function_0/N2  ( .A1(\SB1_3_6/i0[8] ), .A2(
        \SB1_3_6/i0[7] ), .A3(\SB1_3_6/i0[6] ), .ZN(
        \SB1_3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_6/Component_Function_0/N1  ( .A1(\SB1_3_6/i0[10] ), .A2(
        \SB1_3_6/i0[9] ), .ZN(\SB1_3_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_1/N4  ( .A1(\SB1_3_6/i1_7 ), .A2(
        \SB1_3_6/i0[8] ), .A3(\SB1_3_6/i0_4 ), .ZN(
        \SB1_3_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_6/Component_Function_1/N3  ( .A1(\SB1_3_6/i1_5 ), .A2(
        \SB1_3_6/i0[6] ), .A3(\SB1_3_6/i0[9] ), .ZN(
        \SB1_3_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_6/Component_Function_1/N2  ( .A1(\SB1_3_6/i0_3 ), .A2(
        \SB1_3_6/i1_7 ), .A3(\SB1_3_6/i0[8] ), .ZN(
        \SB1_3_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_6/Component_Function_1/N1  ( .A1(\SB1_3_6/i0_3 ), .A2(
        \SB1_3_6/i1[9] ), .ZN(\SB1_3_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_5/N2  ( .A1(\SB1_3_6/i0_0 ), .A2(
        \SB1_3_6/i0[6] ), .A3(\SB1_3_6/i0[10] ), .ZN(
        \SB1_3_6/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_6/Component_Function_5/N1  ( .A1(\SB1_3_6/i0_0 ), .A2(
        \SB1_3_6/i3[0] ), .ZN(\SB1_3_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_0/N4  ( .A1(\SB1_3_7/i0[7] ), .A2(
        \SB1_3_7/i0_3 ), .A3(\SB1_3_7/i0_0 ), .ZN(
        \SB1_3_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_7/Component_Function_0/N3  ( .A1(\SB1_3_7/i0[10] ), .A2(
        \SB1_3_7/i0_4 ), .A3(\SB1_3_7/i0_3 ), .ZN(
        \SB1_3_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_7/Component_Function_0/N2  ( .A1(\SB1_3_7/i0[8] ), .A2(
        \SB1_3_7/i0[7] ), .A3(\SB1_3_7/i0[6] ), .ZN(
        \SB1_3_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_7/Component_Function_0/N1  ( .A1(\SB1_3_7/i0[10] ), .A2(
        \SB1_3_7/i0[9] ), .ZN(\SB1_3_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_1/N3  ( .A1(\SB1_3_7/i1_5 ), .A2(
        \SB1_3_7/i0[6] ), .A3(\SB1_3_7/i0[9] ), .ZN(
        \SB1_3_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_7/Component_Function_1/N2  ( .A1(\SB1_3_7/i0_3 ), .A2(
        \SB1_3_7/i1_7 ), .A3(\SB1_3_7/i0[8] ), .ZN(
        \SB1_3_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_7/Component_Function_1/N1  ( .A1(\SB1_3_7/i0_3 ), .A2(
        \SB1_3_7/i1[9] ), .ZN(\SB1_3_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_5/N4  ( .A1(\SB1_3_7/i0[9] ), .A2(
        \SB1_3_7/i0[6] ), .A3(\SB1_3_7/i0_4 ), .ZN(
        \SB1_3_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_7/Component_Function_5/N2  ( .A1(\SB1_3_7/i0_0 ), .A2(
        \SB1_3_7/i0[6] ), .A3(\SB1_3_7/i0[10] ), .ZN(
        \SB1_3_7/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_7/Component_Function_5/N1  ( .A1(\SB1_3_7/i0_0 ), .A2(
        \SB1_3_7/i3[0] ), .ZN(\SB1_3_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_0/N4  ( .A1(\SB1_3_8/i0[7] ), .A2(
        \SB1_3_8/i0_3 ), .A3(\SB1_3_8/i0_0 ), .ZN(
        \SB1_3_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_8/Component_Function_0/N3  ( .A1(\SB1_3_8/i0[10] ), .A2(
        \SB1_3_8/i0_4 ), .A3(\SB1_3_8/i0_3 ), .ZN(
        \SB1_3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_8/Component_Function_0/N2  ( .A1(\SB1_3_8/i0[8] ), .A2(
        \SB1_3_8/i0[7] ), .A3(\SB1_3_8/i0[6] ), .ZN(
        \SB1_3_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_8/Component_Function_0/N1  ( .A1(\SB1_3_8/i0[10] ), .A2(
        \SB1_3_8/i0[9] ), .ZN(\SB1_3_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_1/N3  ( .A1(\SB1_3_8/i1_5 ), .A2(
        \SB1_3_8/i0[6] ), .A3(\SB1_3_8/i0[9] ), .ZN(
        \SB1_3_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_8/Component_Function_1/N2  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i1_7 ), .A3(\SB1_3_8/i0[8] ), .ZN(
        \SB1_3_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_8/Component_Function_1/N1  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i1[9] ), .ZN(\SB1_3_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_5/N4  ( .A1(\SB1_3_8/i0[9] ), .A2(
        \SB1_3_8/i0[6] ), .A3(\SB1_3_8/i0_4 ), .ZN(
        \SB1_3_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_8/Component_Function_5/N2  ( .A1(\SB1_3_8/i0_0 ), .A2(
        \SB1_3_8/i0[6] ), .A3(\SB1_3_8/i0[10] ), .ZN(
        \SB1_3_8/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_8/Component_Function_5/N1  ( .A1(\SB1_3_8/i0_0 ), .A2(
        \SB1_3_8/i3[0] ), .ZN(\SB1_3_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N4  ( .A1(\SB1_3_9/i0[7] ), .A2(
        \SB1_3_9/i0_3 ), .A3(\SB1_3_9/i0_0 ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N3  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i0_4 ), .A3(\SB1_3_9/i0[10] ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N2  ( .A1(\SB1_3_9/i0[8] ), .A2(
        \SB1_3_9/i0[7] ), .A3(\SB1_3_9/i0[6] ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_9/Component_Function_0/N1  ( .A1(\SB1_3_9/i0[10] ), .A2(
        \SB1_3_9/i0[9] ), .ZN(\SB1_3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_1/N4  ( .A1(\SB1_3_9/i1_7 ), .A2(
        \SB1_3_9/i0[8] ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_1/N3  ( .A1(\SB1_3_9/i1_5 ), .A2(
        \SB1_3_9/i0[6] ), .A3(\SB1_3_9/i0[9] ), .ZN(
        \SB1_3_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_9/Component_Function_1/N2  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i1_7 ), .A3(\SB1_3_9/i0[8] ), .ZN(
        \SB1_3_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_9/Component_Function_1/N1  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i1[9] ), .ZN(\SB1_3_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_5/N4  ( .A1(\SB1_3_9/i0[9] ), .A2(
        \SB1_3_9/i0[6] ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_5/N2  ( .A1(\SB1_3_9/i0_0 ), .A2(
        \SB1_3_9/i0[6] ), .A3(\SB1_3_9/i0[10] ), .ZN(
        \SB1_3_9/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_9/Component_Function_5/N1  ( .A1(\SB1_3_9/i0_0 ), .A2(
        \SB1_3_9/i3[0] ), .ZN(\SB1_3_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_0/N4  ( .A1(\SB1_3_10/i0[7] ), .A2(
        \SB1_3_10/i0_3 ), .A3(\SB1_3_10/i0_0 ), .ZN(
        \SB1_3_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_10/Component_Function_0/N3  ( .A1(\SB1_3_10/i0[10] ), .A2(
        \SB1_3_10/i0_4 ), .A3(\SB1_3_10/i0_3 ), .ZN(
        \SB1_3_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_10/Component_Function_0/N2  ( .A1(\SB1_3_10/i0[8] ), .A2(
        \SB1_3_10/i0[7] ), .A3(\SB1_3_10/i0[6] ), .ZN(
        \SB1_3_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_10/Component_Function_0/N1  ( .A1(\SB1_3_10/i0[10] ), .A2(
        \SB1_3_10/i0[9] ), .ZN(\SB1_3_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_1/N4  ( .A1(\SB1_3_10/i1_7 ), .A2(
        \SB1_3_10/i0[8] ), .A3(\SB1_3_10/i0_4 ), .ZN(
        \SB1_3_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_10/Component_Function_1/N3  ( .A1(\SB1_3_10/i1_5 ), .A2(
        \SB1_3_10/i0[6] ), .A3(\SB1_3_10/i0[9] ), .ZN(
        \SB1_3_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_10/Component_Function_1/N2  ( .A1(\SB1_3_10/i0_3 ), .A2(
        \SB1_3_10/i1_7 ), .A3(\SB1_3_10/i0[8] ), .ZN(
        \SB1_3_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_10/Component_Function_1/N1  ( .A1(\SB1_3_10/i0_3 ), .A2(
        \SB1_3_10/i1[9] ), .ZN(\SB1_3_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_5/N4  ( .A1(\SB1_3_10/i0[9] ), .A2(
        \SB1_3_10/i0[6] ), .A3(\SB1_3_10/i0_4 ), .ZN(
        \SB1_3_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_10/Component_Function_5/N2  ( .A1(\SB1_3_10/i0_0 ), .A2(
        \SB1_3_10/i0[6] ), .A3(\SB1_3_10/i0[10] ), .ZN(
        \SB1_3_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_10/Component_Function_5/N1  ( .A1(\SB1_3_10/i0_0 ), .A2(
        \SB1_3_10/i3[0] ), .ZN(\SB1_3_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N4  ( .A1(\SB1_3_11/i0[7] ), .A2(
        \SB1_3_11/i0_3 ), .A3(\SB1_3_11/i0_0 ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N3  ( .A1(\SB1_3_11/i0[10] ), .A2(
        \SB1_3_11/i0_4 ), .A3(\SB1_3_11/i0_3 ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N2  ( .A1(\SB1_3_11/i0[8] ), .A2(
        \SB1_3_11/i0[7] ), .A3(\SB1_3_11/i0[6] ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_11/Component_Function_0/N1  ( .A1(\SB1_3_11/i0[10] ), .A2(
        \SB1_3_11/i0[9] ), .ZN(\SB1_3_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_1/N4  ( .A1(\SB1_3_11/i1_7 ), .A2(
        \SB1_3_11/i0[8] ), .A3(\SB1_3_11/i0_4 ), .ZN(
        \SB1_3_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_11/Component_Function_1/N3  ( .A1(\SB1_3_11/i1_5 ), .A2(
        \SB1_3_11/i0[6] ), .A3(\SB1_3_11/i0[9] ), .ZN(
        \SB1_3_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_11/Component_Function_1/N2  ( .A1(n831), .A2(\SB1_3_11/i1_7 ), .A3(\SB1_3_11/i0[8] ), .ZN(\SB1_3_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_11/Component_Function_1/N1  ( .A1(n831), .A2(
        \SB1_3_11/i1[9] ), .ZN(\SB1_3_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_5/N4  ( .A1(\SB1_3_11/i0_4 ), .A2(
        \SB1_3_11/i0[6] ), .A3(\SB1_3_11/i0[9] ), .ZN(
        \SB1_3_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_11/Component_Function_5/N3  ( .A1(\SB1_3_11/i1[9] ), .A2(
        \SB1_3_11/i0_4 ), .A3(\SB1_3_11/i0_3 ), .ZN(
        \SB1_3_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_11/Component_Function_5/N2  ( .A1(\SB1_3_11/i0_0 ), .A2(
        \SB1_3_11/i0[6] ), .A3(\SB1_3_11/i0[10] ), .ZN(
        \SB1_3_11/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_11/Component_Function_5/N1  ( .A1(\SB1_3_11/i0_0 ), .A2(
        \SB1_3_11/i3[0] ), .ZN(\SB1_3_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_12/Component_Function_0/N4  ( .A1(\SB1_3_12/i0[7] ), .A2(
        \SB1_3_12/i0_3 ), .A3(\SB1_3_12/i0_0 ), .ZN(
        \SB1_3_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_12/Component_Function_0/N3  ( .A1(\SB1_3_12/i0[10] ), .A2(
        \SB1_3_12/i0_4 ), .A3(\SB1_3_12/i0_3 ), .ZN(
        \SB1_3_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_12/Component_Function_0/N2  ( .A1(\SB1_3_12/i0[8] ), .A2(
        \SB1_3_12/i0[7] ), .A3(\SB1_3_12/i0[6] ), .ZN(
        \SB1_3_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_12/Component_Function_0/N1  ( .A1(\SB1_3_12/i0[10] ), .A2(
        \SB1_3_12/i0[9] ), .ZN(\SB1_3_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_12/Component_Function_1/N3  ( .A1(\SB1_3_12/i1_5 ), .A2(
        \SB1_3_12/i0[6] ), .A3(\SB1_3_12/i0[9] ), .ZN(
        \SB1_3_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_12/Component_Function_1/N2  ( .A1(\SB1_3_12/i0_3 ), .A2(
        \SB1_3_12/i1_7 ), .A3(\SB1_3_12/i0[8] ), .ZN(
        \SB1_3_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_12/Component_Function_1/N1  ( .A1(\SB1_3_12/i0_3 ), .A2(
        \SB1_3_12/i1[9] ), .ZN(\SB1_3_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_12/Component_Function_5/N4  ( .A1(\SB1_3_12/i0[9] ), .A2(
        \SB1_3_12/i0[6] ), .A3(\SB1_3_12/i0_4 ), .ZN(
        \SB1_3_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_12/Component_Function_5/N2  ( .A1(\SB1_3_12/i0_0 ), .A2(
        \SB1_3_12/i0[6] ), .A3(\SB1_3_12/i0[10] ), .ZN(
        \SB1_3_12/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_12/Component_Function_5/N1  ( .A1(\SB1_3_12/i0_0 ), .A2(
        \SB1_3_12/i3[0] ), .ZN(\SB1_3_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N4  ( .A1(\SB1_3_13/i0[7] ), .A2(
        \SB1_3_13/i0_3 ), .A3(\SB1_3_13/i0_0 ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N3  ( .A1(\SB1_3_13/i0[10] ), .A2(
        \SB1_3_13/i0_4 ), .A3(\SB1_3_13/i0_3 ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N2  ( .A1(\SB1_3_13/i0[8] ), .A2(
        \SB1_3_13/i0[7] ), .A3(\SB1_3_13/i0[6] ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_13/Component_Function_0/N1  ( .A1(\SB1_3_13/i0[10] ), .A2(
        \SB1_3_13/i0[9] ), .ZN(\SB1_3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_1/N4  ( .A1(\SB1_3_13/i1_7 ), .A2(
        \SB1_3_13/i0[8] ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_13/Component_Function_1/N3  ( .A1(\SB1_3_13/i1_5 ), .A2(
        \SB1_3_13/i0[6] ), .A3(\SB1_3_13/i0[9] ), .ZN(
        \SB1_3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_1/N2  ( .A1(\SB1_3_13/i0_3 ), .A2(
        \SB1_3_13/i1_7 ), .A3(\SB1_3_13/i0[8] ), .ZN(
        \SB1_3_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_13/Component_Function_1/N1  ( .A1(\SB1_3_13/i0_3 ), .A2(
        \SB1_3_13/i1[9] ), .ZN(\SB1_3_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_5/N4  ( .A1(\SB1_3_13/i0[9] ), .A2(
        \SB1_3_13/i0[6] ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_13/Component_Function_5/N2  ( .A1(\SB1_3_13/i0_0 ), .A2(
        \SB1_3_13/i0[6] ), .A3(\SB1_3_13/i0[10] ), .ZN(
        \SB1_3_13/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_13/Component_Function_5/N1  ( .A1(\SB1_3_13/i0_0 ), .A2(
        \SB1_3_13/i3[0] ), .ZN(\SB1_3_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_0/N4  ( .A1(\SB1_3_14/i0[7] ), .A2(
        \SB1_3_14/i0_3 ), .A3(\SB1_3_14/i0_0 ), .ZN(
        \SB1_3_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_0/N3  ( .A1(\SB1_3_14/i0[10] ), .A2(
        \SB1_3_14/i0_4 ), .A3(\SB1_3_14/i0_3 ), .ZN(
        \SB1_3_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_14/Component_Function_0/N2  ( .A1(\SB1_3_14/i0[8] ), .A2(
        \SB1_3_14/i0[7] ), .A3(\SB1_3_14/i0[6] ), .ZN(
        \SB1_3_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_14/Component_Function_0/N1  ( .A1(\SB1_3_14/i0[10] ), .A2(
        \SB1_3_14/i0[9] ), .ZN(\SB1_3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N4  ( .A1(\SB1_3_14/i1_7 ), .A2(
        \SB1_3_14/i0[8] ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N3  ( .A1(\SB1_3_14/i1_5 ), .A2(
        \SB1_3_14/i0[6] ), .A3(\SB1_3_14/i0[9] ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N2  ( .A1(\SB1_3_14/i0_3 ), .A2(
        \SB1_3_14/i1_7 ), .A3(\SB1_3_14/i0[8] ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_14/Component_Function_1/N1  ( .A1(\SB1_3_14/i0_3 ), .A2(
        \SB1_3_14/i1[9] ), .ZN(\SB1_3_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_5/N4  ( .A1(\SB1_3_14/i0[9] ), .A2(
        \SB1_3_14/i0[6] ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_5/N2  ( .A1(\SB1_3_14/i0_0 ), .A2(
        \SB1_3_14/i0[6] ), .A3(\SB1_3_14/i0[10] ), .ZN(
        \SB1_3_14/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_14/Component_Function_5/N1  ( .A1(\SB1_3_14/i0_0 ), .A2(
        \SB1_3_14/i3[0] ), .ZN(\SB1_3_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_0/N3  ( .A1(\SB1_3_15/i0[10] ), .A2(
        \SB1_3_15/i0_4 ), .A3(\SB1_3_15/i0_3 ), .ZN(
        \SB1_3_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_15/Component_Function_0/N2  ( .A1(\SB1_3_15/i0[8] ), .A2(
        \SB1_3_15/i0[7] ), .A3(\SB1_3_15/i0[6] ), .ZN(
        \SB1_3_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_15/Component_Function_0/N1  ( .A1(\SB1_3_15/i0[10] ), .A2(
        \SB1_3_15/i0[9] ), .ZN(\SB1_3_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_1/N4  ( .A1(\SB1_3_15/i1_7 ), .A2(
        \SB1_3_15/i0[8] ), .A3(\SB1_3_15/i0_4 ), .ZN(
        \SB1_3_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_15/Component_Function_1/N3  ( .A1(\SB1_3_15/i1_5 ), .A2(
        \SB1_3_15/i0[6] ), .A3(\SB1_3_15/i0[9] ), .ZN(
        \SB1_3_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_15/Component_Function_1/N2  ( .A1(n1647), .A2(
        \SB1_3_15/i1_7 ), .A3(\SB1_3_15/i0[8] ), .ZN(
        \SB1_3_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_15/Component_Function_1/N1  ( .A1(n1647), .A2(
        \SB1_3_15/i1[9] ), .ZN(\SB1_3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_5/N4  ( .A1(\SB1_3_15/i0[9] ), .A2(
        \SB1_3_15/i0[6] ), .A3(\SB1_3_15/i0_4 ), .ZN(
        \SB1_3_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_15/Component_Function_5/N2  ( .A1(\SB1_3_15/i0_0 ), .A2(
        \SB1_3_15/i0[6] ), .A3(\SB1_3_15/i0[10] ), .ZN(
        \SB1_3_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_15/Component_Function_5/N1  ( .A1(\SB1_3_15/i0_0 ), .A2(
        \SB1_3_15/i3[0] ), .ZN(\SB1_3_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N4  ( .A1(\SB1_3_16/i0[7] ), .A2(
        \SB1_3_16/i0_3 ), .A3(\SB1_3_16/i0_0 ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N3  ( .A1(\SB1_3_16/i0[10] ), .A2(
        \SB1_3_16/i0_4 ), .A3(\SB1_3_16/i0_3 ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N2  ( .A1(\SB1_3_16/i0[8] ), .A2(
        \SB1_3_16/i0[7] ), .A3(\SB1_3_16/i0[6] ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_16/Component_Function_0/N1  ( .A1(\SB1_3_16/i0[10] ), .A2(
        \SB1_3_16/i0[9] ), .ZN(\SB1_3_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_1/N4  ( .A1(\SB1_3_16/i1_7 ), .A2(
        \SB1_3_16/i0[8] ), .A3(\SB1_3_16/i0_4 ), .ZN(
        \SB1_3_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_1/N3  ( .A1(\SB1_3_16/i1_5 ), .A2(
        \SB1_3_16/i0[6] ), .A3(\SB1_3_16/i0[9] ), .ZN(
        \SB1_3_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_16/Component_Function_1/N2  ( .A1(\SB1_3_16/i0_3 ), .A2(
        \SB1_3_16/i1_7 ), .A3(\SB1_3_16/i0[8] ), .ZN(
        \SB1_3_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_16/Component_Function_1/N1  ( .A1(\SB1_3_16/i0_3 ), .A2(
        \SB1_3_16/i1[9] ), .ZN(\SB1_3_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_5/N2  ( .A1(\SB1_3_16/i0_0 ), .A2(
        \SB1_3_16/i0[6] ), .A3(\SB1_3_16/i0[10] ), .ZN(
        \SB1_3_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_16/Component_Function_5/N1  ( .A1(\SB1_3_16/i0_0 ), .A2(
        \SB1_3_16/i3[0] ), .ZN(\SB1_3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_17/Component_Function_0/N4  ( .A1(\SB1_3_17/i0[7] ), .A2(
        \SB1_3_17/i0_3 ), .A3(\SB1_3_17/i0_0 ), .ZN(
        \SB1_3_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_17/Component_Function_0/N3  ( .A1(\SB1_3_17/i0[10] ), .A2(
        \SB1_3_17/i0_4 ), .A3(\SB1_3_17/i0_3 ), .ZN(
        \SB1_3_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_17/Component_Function_0/N2  ( .A1(\SB1_3_17/i0[8] ), .A2(
        \SB1_3_17/i0[7] ), .A3(\SB1_3_17/i0[6] ), .ZN(
        \SB1_3_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_17/Component_Function_0/N1  ( .A1(\SB1_3_17/i0[10] ), .A2(
        \SB1_3_17/i0[9] ), .ZN(\SB1_3_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_17/Component_Function_1/N4  ( .A1(\SB1_3_17/i1_7 ), .A2(
        \SB1_3_17/i0[8] ), .A3(\SB1_3_17/i0_4 ), .ZN(
        \SB1_3_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_17/Component_Function_1/N3  ( .A1(\SB1_3_17/i1_5 ), .A2(
        \SB1_3_17/i0[6] ), .A3(\SB1_3_17/i0[9] ), .ZN(
        \SB1_3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_17/Component_Function_1/N2  ( .A1(\SB1_3_17/i0_3 ), .A2(
        \SB1_3_17/i1_7 ), .A3(\SB1_3_17/i0[8] ), .ZN(
        \SB1_3_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_17/Component_Function_1/N1  ( .A1(\SB1_3_17/i0_3 ), .A2(
        \SB1_3_17/i1[9] ), .ZN(\SB1_3_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_17/Component_Function_5/N1  ( .A1(\SB1_3_17/i0_0 ), .A2(
        \SB1_3_17/i3[0] ), .ZN(\SB1_3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_0/N4  ( .A1(\SB1_3_18/i0[7] ), .A2(
        \SB1_3_18/i0_3 ), .A3(\SB1_3_18/i0_0 ), .ZN(
        \SB1_3_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_18/Component_Function_0/N3  ( .A1(\SB1_3_18/i0[10] ), .A2(
        \SB1_3_18/i0_4 ), .A3(\SB1_3_18/i0_3 ), .ZN(
        \SB1_3_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_18/Component_Function_0/N2  ( .A1(\SB1_3_18/i0[8] ), .A2(
        \SB1_3_18/i0[7] ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_18/Component_Function_0/N1  ( .A1(\SB1_3_18/i0[10] ), .A2(
        \SB1_3_18/i0[9] ), .ZN(\SB1_3_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_1/N4  ( .A1(\SB1_3_18/i1_7 ), .A2(
        \SB1_3_18/i0[8] ), .A3(\SB1_3_18/i0_4 ), .ZN(
        \SB1_3_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_18/Component_Function_1/N3  ( .A1(\SB1_3_18/i1_5 ), .A2(
        \SB1_3_18/i0[6] ), .A3(\SB1_3_18/i0[9] ), .ZN(
        \SB1_3_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_18/Component_Function_1/N2  ( .A1(\SB1_3_18/i0_3 ), .A2(
        \SB1_3_18/i1_7 ), .A3(\SB1_3_18/i0[8] ), .ZN(
        \SB1_3_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_18/Component_Function_1/N1  ( .A1(\SB1_3_18/i0_3 ), .A2(
        \SB1_3_18/i1[9] ), .ZN(\SB1_3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_5/N2  ( .A1(\SB1_3_18/i0_0 ), .A2(
        \SB1_3_18/i0[6] ), .A3(\SB1_3_18/i0[10] ), .ZN(
        \SB1_3_18/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_18/Component_Function_5/N1  ( .A1(\SB1_3_18/i0_0 ), .A2(
        \SB1_3_18/i3[0] ), .ZN(\SB1_3_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_0/N4  ( .A1(\SB1_3_19/i0[7] ), .A2(
        \SB1_3_19/i0_3 ), .A3(\SB1_3_19/i0_0 ), .ZN(
        \SB1_3_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_19/Component_Function_0/N3  ( .A1(\SB1_3_19/i0[10] ), .A2(
        \SB1_3_19/i0_4 ), .A3(\SB1_3_19/i0_3 ), .ZN(
        \SB1_3_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_19/Component_Function_0/N2  ( .A1(\SB1_3_19/i0[8] ), .A2(
        \SB1_3_19/i0[7] ), .A3(\SB1_3_19/i0[6] ), .ZN(
        \SB1_3_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_19/Component_Function_0/N1  ( .A1(\SB1_3_19/i0[10] ), .A2(
        \SB1_3_19/i0[9] ), .ZN(\SB1_3_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_1/N4  ( .A1(\SB1_3_19/i1_7 ), .A2(
        \SB1_3_19/i0[8] ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_19/Component_Function_1/N3  ( .A1(\SB1_3_19/i1_5 ), .A2(
        \SB1_3_19/i0[6] ), .A3(\SB1_3_19/i0[9] ), .ZN(
        \SB1_3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_19/Component_Function_1/N2  ( .A1(\SB1_3_19/i0_3 ), .A2(
        \SB1_3_19/i1_7 ), .A3(\SB1_3_19/i0[8] ), .ZN(
        \SB1_3_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_19/Component_Function_1/N1  ( .A1(\SB1_3_19/i0_3 ), .A2(
        \SB1_3_19/i1[9] ), .ZN(\SB1_3_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_5/N4  ( .A1(\SB1_3_19/i0[9] ), .A2(
        \SB1_3_19/i0[6] ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_19/Component_Function_5/N2  ( .A1(\SB1_3_19/i0_0 ), .A2(
        \SB1_3_19/i0[6] ), .A3(\SB1_3_19/i0[10] ), .ZN(
        \SB1_3_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_19/Component_Function_5/N1  ( .A1(\SB1_3_19/i0_0 ), .A2(
        \SB1_3_19/i3[0] ), .ZN(\SB1_3_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_0/N4  ( .A1(\SB1_3_20/i0[7] ), .A2(
        \SB1_3_20/i0_3 ), .A3(\SB1_3_20/i0_0 ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_20/Component_Function_0/N3  ( .A1(\SB1_3_20/i0[10] ), .A2(
        \SB1_3_20/i0_4 ), .A3(\SB1_3_20/i0_3 ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_20/Component_Function_0/N2  ( .A1(\SB1_3_20/i0[8] ), .A2(
        \SB1_3_20/i0[7] ), .A3(\SB1_3_20/i0[6] ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_20/Component_Function_0/N1  ( .A1(\SB1_3_20/i0[10] ), .A2(
        \SB1_3_20/i0[9] ), .ZN(\SB1_3_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_1/N3  ( .A1(\SB1_3_20/i1_5 ), .A2(
        \SB1_3_20/i0[6] ), .A3(\SB1_3_20/i0[9] ), .ZN(
        \SB1_3_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_20/Component_Function_1/N2  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i1_7 ), .A3(\SB1_3_20/i0[8] ), .ZN(
        \SB1_3_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_20/Component_Function_1/N1  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i1[9] ), .ZN(\SB1_3_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_5/N4  ( .A1(\SB1_3_20/i0[9] ), .A2(
        \SB1_3_20/i0[6] ), .A3(\SB1_3_20/i0_4 ), .ZN(
        \SB1_3_20/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_3_20/Component_Function_5/N1  ( .A1(\SB1_3_20/i0_0 ), .A2(
        \SB1_3_20/i3[0] ), .ZN(\SB1_3_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_0/N4  ( .A1(\SB1_3_21/i0[7] ), .A2(
        \SB1_3_21/i0_3 ), .A3(\SB1_3_21/i0_0 ), .ZN(
        \SB1_3_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_21/Component_Function_0/N2  ( .A1(\SB1_3_21/i0[8] ), .A2(
        \SB1_3_21/i0[7] ), .A3(\SB1_3_21/i0[6] ), .ZN(
        \SB1_3_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_21/Component_Function_0/N1  ( .A1(\SB1_3_21/i0[10] ), .A2(
        \SB1_3_21/i0[9] ), .ZN(\SB1_3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_1/N4  ( .A1(\SB1_3_21/i1_7 ), .A2(
        \SB1_3_21/i0[8] ), .A3(\SB1_3_21/i0_4 ), .ZN(
        \SB1_3_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_21/Component_Function_1/N3  ( .A1(\SB1_3_21/i1_5 ), .A2(
        \SB1_3_21/i0[6] ), .A3(\SB1_3_21/i0[9] ), .ZN(
        \SB1_3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_21/Component_Function_1/N2  ( .A1(\SB1_3_21/i0_3 ), .A2(
        \SB1_3_21/i1_7 ), .A3(\SB1_3_21/i0[8] ), .ZN(
        \SB1_3_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_21/Component_Function_1/N1  ( .A1(\SB1_3_21/i0_3 ), .A2(
        \SB1_3_21/i1[9] ), .ZN(\SB1_3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_5/N4  ( .A1(\SB1_3_21/i0[9] ), .A2(
        \SB1_3_21/i0[6] ), .A3(\SB1_3_21/i0_4 ), .ZN(
        \SB1_3_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_21/Component_Function_5/N2  ( .A1(\SB1_3_21/i0_0 ), .A2(
        \SB1_3_21/i0[6] ), .A3(\SB1_3_21/i0[10] ), .ZN(
        \SB1_3_21/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_21/Component_Function_5/N1  ( .A1(\SB1_3_21/i0_0 ), .A2(
        \SB1_3_21/i3[0] ), .ZN(\SB1_3_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_0/N4  ( .A1(\SB1_3_22/i0[7] ), .A2(
        \SB1_3_22/i0_3 ), .A3(\SB1_3_22/i0_0 ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_22/Component_Function_0/N3  ( .A1(\SB1_3_22/i0[10] ), .A2(
        \SB1_3_22/i0_4 ), .A3(\SB1_3_22/i0_3 ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_22/Component_Function_0/N2  ( .A1(\SB1_3_22/i0[8] ), .A2(
        \SB1_3_22/i0[7] ), .A3(\SB1_3_22/i0[6] ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_22/Component_Function_0/N1  ( .A1(\SB1_3_22/i0[10] ), .A2(
        \SB1_3_22/i0[9] ), .ZN(\SB1_3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_1/N4  ( .A1(\SB1_3_22/i1_7 ), .A2(
        \SB1_3_22/i0[8] ), .A3(\SB1_3_22/i0_4 ), .ZN(
        \SB1_3_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_22/Component_Function_1/N3  ( .A1(\SB1_3_22/i1_5 ), .A2(
        \SB1_3_22/i0[6] ), .A3(\SB1_3_22/i0[9] ), .ZN(
        \SB1_3_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_22/Component_Function_1/N2  ( .A1(\SB1_3_22/i0_3 ), .A2(
        \SB1_3_22/i1_7 ), .A3(\SB1_3_22/i0[8] ), .ZN(
        \SB1_3_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_22/Component_Function_1/N1  ( .A1(\SB1_3_22/i0_3 ), .A2(
        \SB1_3_22/i1[9] ), .ZN(\SB1_3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_5/N4  ( .A1(\SB1_3_22/i0[9] ), .A2(
        \SB1_3_22/i0[6] ), .A3(\SB1_3_22/i0_4 ), .ZN(
        \SB1_3_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_22/Component_Function_5/N2  ( .A1(\SB1_3_22/i0_0 ), .A2(
        \SB1_3_22/i0[6] ), .A3(\SB1_3_22/i0[10] ), .ZN(
        \SB1_3_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_22/Component_Function_5/N1  ( .A1(\SB1_3_22/i0_0 ), .A2(
        \SB1_3_22/i3[0] ), .ZN(\SB1_3_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_0/N4  ( .A1(\SB1_3_23/i0[7] ), .A2(
        \SB1_3_23/i0_3 ), .A3(\SB1_3_23/i0_0 ), .ZN(
        \SB1_3_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_23/Component_Function_0/N3  ( .A1(\SB1_3_23/i0_3 ), .A2(
        \SB1_3_23/i0_4 ), .A3(\SB1_3_23/i0[10] ), .ZN(
        \SB1_3_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_23/Component_Function_0/N2  ( .A1(\SB1_3_23/i0[8] ), .A2(
        \SB1_3_23/i0[7] ), .A3(\SB1_3_23/i0[6] ), .ZN(
        \SB1_3_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_23/Component_Function_0/N1  ( .A1(\SB1_3_23/i0[10] ), .A2(
        \SB1_3_23/i0[9] ), .ZN(\SB1_3_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_1/N3  ( .A1(\SB1_3_23/i1_5 ), .A2(
        \SB1_3_23/i0[6] ), .A3(\SB1_3_23/i0[9] ), .ZN(
        \SB1_3_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_23/Component_Function_1/N2  ( .A1(\SB1_3_23/i0_3 ), .A2(
        \SB1_3_23/i1_7 ), .A3(\SB1_3_23/i0[8] ), .ZN(
        \SB1_3_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_23/Component_Function_1/N1  ( .A1(\SB1_3_23/i0_3 ), .A2(
        \SB1_3_23/i1[9] ), .ZN(\SB1_3_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_5/N4  ( .A1(\SB1_3_23/i0[9] ), .A2(
        \SB1_3_23/i0[6] ), .A3(\SB1_3_23/i0_4 ), .ZN(
        \SB1_3_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_23/Component_Function_5/N2  ( .A1(\SB1_3_23/i0_0 ), .A2(
        \SB1_3_23/i0[6] ), .A3(\SB1_3_23/i0[10] ), .ZN(
        \SB1_3_23/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_23/Component_Function_5/N1  ( .A1(\SB1_3_23/i0_0 ), .A2(
        \SB1_3_23/i3[0] ), .ZN(\SB1_3_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_0/N4  ( .A1(\SB1_3_24/i0[7] ), .A2(
        \SB1_3_24/i0_3 ), .A3(\SB1_3_24/i0_0 ), .ZN(
        \SB1_3_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_0/N3  ( .A1(\SB1_3_24/i0[10] ), .A2(
        \SB1_3_24/i0_4 ), .A3(\SB1_3_24/i0_3 ), .ZN(
        \SB1_3_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_24/Component_Function_0/N2  ( .A1(\SB1_3_24/i0[8] ), .A2(
        \SB1_3_24/i0[7] ), .A3(\SB1_3_24/i0[6] ), .ZN(
        \SB1_3_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_24/Component_Function_0/N1  ( .A1(\SB1_3_24/i0[10] ), .A2(
        \SB1_3_24/i0[9] ), .ZN(\SB1_3_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N4  ( .A1(\SB1_3_24/i1_7 ), .A2(
        \SB1_3_24/i0[8] ), .A3(\SB1_3_24/i0_4 ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N3  ( .A1(\SB1_3_24/i1_5 ), .A2(
        \SB1_3_24/i0[6] ), .A3(\SB1_3_24/i0[9] ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N2  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i1_7 ), .A3(\SB1_3_24/i0[8] ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_24/Component_Function_1/N1  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i1[9] ), .ZN(\SB1_3_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_5/N4  ( .A1(\SB1_3_24/i0[9] ), .A2(
        \SB1_3_24/i0[6] ), .A3(\SB1_3_24/i0_4 ), .ZN(
        \SB1_3_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_5/N2  ( .A1(\SB1_3_24/i0_0 ), .A2(
        \SB1_3_24/i0[6] ), .A3(\SB1_3_24/i0[10] ), .ZN(
        \SB1_3_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_24/Component_Function_5/N1  ( .A1(\SB1_3_24/i0_0 ), .A2(
        \SB1_3_24/i3[0] ), .ZN(\SB1_3_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N4  ( .A1(\SB1_3_25/i0[7] ), .A2(
        n804), .A3(\SB1_3_25/i0_0 ), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N3  ( .A1(\SB1_3_25/i0[10] ), .A2(
        \SB1_3_25/i0_4 ), .A3(n804), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N2  ( .A1(\SB1_3_25/i0[8] ), .A2(
        \SB1_3_25/i0[7] ), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_25/Component_Function_0/N1  ( .A1(\SB1_3_25/i0[10] ), .A2(
        \SB1_3_25/i0[9] ), .ZN(\SB1_3_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_1/N3  ( .A1(\SB1_3_25/i1_5 ), .A2(
        \SB1_3_25/i0[6] ), .A3(\SB1_3_25/i0[9] ), .ZN(
        \SB1_3_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_25/Component_Function_1/N2  ( .A1(n804), .A2(\SB1_3_25/i1_7 ), .A3(\SB1_3_25/i0[8] ), .ZN(\SB1_3_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_25/Component_Function_1/N1  ( .A1(\SB1_3_25/i0_3 ), .A2(
        \SB1_3_25/i1[9] ), .ZN(\SB1_3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_5/N4  ( .A1(\SB1_3_25/i0[9] ), .A2(
        \SB1_3_25/i0[6] ), .A3(\SB1_3_25/i0_4 ), .ZN(
        \SB1_3_25/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_3_25/Component_Function_5/N1  ( .A1(\SB1_3_25/i0_0 ), .A2(
        \SB1_3_25/i3[0] ), .ZN(\SB1_3_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_0/N4  ( .A1(\SB1_3_26/i0[7] ), .A2(
        \SB1_3_26/i0_3 ), .A3(\SB1_3_26/i0_0 ), .ZN(
        \SB1_3_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_26/Component_Function_0/N3  ( .A1(\SB1_3_26/i0[10] ), .A2(
        \SB1_3_26/i0_4 ), .A3(\SB1_3_26/i0_3 ), .ZN(
        \SB1_3_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_26/Component_Function_0/N2  ( .A1(\SB1_3_26/i0[8] ), .A2(
        \SB1_3_26/i0[7] ), .A3(\SB1_3_26/i0[6] ), .ZN(
        \SB1_3_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_26/Component_Function_0/N1  ( .A1(\SB1_3_26/i0[10] ), .A2(
        \SB1_3_26/i0[9] ), .ZN(\SB1_3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_1/N4  ( .A1(\SB1_3_26/i1_7 ), .A2(
        \SB1_3_26/i0[8] ), .A3(\SB1_3_26/i0_4 ), .ZN(
        \SB1_3_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_26/Component_Function_1/N3  ( .A1(\SB1_3_26/i1_5 ), .A2(
        \SB1_3_26/i0[6] ), .A3(\SB1_3_26/i0[9] ), .ZN(
        \SB1_3_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_26/Component_Function_1/N2  ( .A1(\SB1_3_26/i0_3 ), .A2(
        \SB1_3_26/i1_7 ), .A3(\SB1_3_26/i0[8] ), .ZN(
        \SB1_3_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_26/Component_Function_1/N1  ( .A1(\SB1_3_26/i0_3 ), .A2(
        \SB1_3_26/i1[9] ), .ZN(\SB1_3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_5/N4  ( .A1(\SB1_3_26/i0[9] ), .A2(
        \SB1_3_26/i0[6] ), .A3(\SB1_3_26/i0_4 ), .ZN(
        \SB1_3_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_26/Component_Function_5/N2  ( .A1(\SB1_3_26/i0_0 ), .A2(
        \SB1_3_26/i0[6] ), .A3(\SB1_3_26/i0[10] ), .ZN(
        \SB1_3_26/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_26/Component_Function_5/N1  ( .A1(\SB1_3_26/i0_0 ), .A2(
        \SB1_3_26/i3[0] ), .ZN(\SB1_3_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_0/N3  ( .A1(\SB1_3_27/i0[10] ), .A2(
        \SB1_3_27/i0_4 ), .A3(\SB1_3_27/i0_3 ), .ZN(
        \SB1_3_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_27/Component_Function_0/N2  ( .A1(\SB1_3_27/i0[8] ), .A2(
        \SB1_3_27/i0[7] ), .A3(\SB1_3_27/i0[6] ), .ZN(
        \SB1_3_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_27/Component_Function_0/N1  ( .A1(\SB1_3_27/i0[10] ), .A2(
        \SB1_3_27/i0[9] ), .ZN(\SB1_3_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_1/N4  ( .A1(\SB1_3_27/i1_7 ), .A2(
        \SB1_3_27/i0[8] ), .A3(\SB1_3_27/i0_4 ), .ZN(
        \SB1_3_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_27/Component_Function_1/N3  ( .A1(\SB1_3_27/i1_5 ), .A2(
        \SB1_3_27/i0[6] ), .A3(\SB1_3_27/i0[9] ), .ZN(
        \SB1_3_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_27/Component_Function_1/N2  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i1_7 ), .A3(\SB1_3_27/i0[8] ), .ZN(
        \SB1_3_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_27/Component_Function_1/N1  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i1[9] ), .ZN(\SB1_3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_5/N4  ( .A1(\SB1_3_27/i0[9] ), .A2(
        \SB1_3_27/i0[6] ), .A3(\SB1_3_27/i0_4 ), .ZN(
        \SB1_3_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_27/Component_Function_5/N2  ( .A1(\SB1_3_27/i0_0 ), .A2(
        \SB1_3_27/i0[6] ), .A3(\SB1_3_27/i0[10] ), .ZN(
        \SB1_3_27/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_27/Component_Function_5/N1  ( .A1(\SB1_3_27/i0_0 ), .A2(
        \SB1_3_27/i3[0] ), .ZN(\SB1_3_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_0/N4  ( .A1(\SB1_3_28/i0[7] ), .A2(
        \SB1_3_28/i0_3 ), .A3(\SB1_3_28/i0_0 ), .ZN(
        \SB1_3_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_28/Component_Function_0/N3  ( .A1(\SB1_3_28/i0[10] ), .A2(
        \SB1_3_28/i0_4 ), .A3(\SB1_3_28/i0_3 ), .ZN(
        \SB1_3_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_28/Component_Function_0/N2  ( .A1(\SB1_3_28/i0[8] ), .A2(
        \SB1_3_28/i0[7] ), .A3(\SB1_3_28/i0[6] ), .ZN(
        \SB1_3_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_28/Component_Function_0/N1  ( .A1(\SB1_3_28/i0[10] ), .A2(
        \SB1_3_28/i0[9] ), .ZN(\SB1_3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_1/N4  ( .A1(\SB1_3_28/i1_7 ), .A2(
        \SB1_3_28/i0[8] ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_28/Component_Function_1/N3  ( .A1(\SB1_3_28/i1_5 ), .A2(
        \SB1_3_28/i0[6] ), .A3(\SB1_3_28/i0[9] ), .ZN(
        \SB1_3_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_28/Component_Function_1/N2  ( .A1(\SB1_3_28/i0_3 ), .A2(
        \SB1_3_28/i1_7 ), .A3(\SB1_3_28/i0[8] ), .ZN(
        \SB1_3_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_28/Component_Function_1/N1  ( .A1(\SB1_3_28/i0_3 ), .A2(
        \SB1_3_28/i1[9] ), .ZN(\SB1_3_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_5/N4  ( .A1(\SB1_3_28/i0[9] ), .A2(
        \SB1_3_28/i0[6] ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_28/Component_Function_5/N2  ( .A1(\SB1_3_28/i0_0 ), .A2(
        \SB1_3_28/i0[6] ), .A3(\SB1_3_28/i0[10] ), .ZN(
        \SB1_3_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_28/Component_Function_5/N1  ( .A1(\SB1_3_28/i0_0 ), .A2(
        \SB1_3_28/i3[0] ), .ZN(\SB1_3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N4  ( .A1(\SB1_3_29/i0[7] ), .A2(
        \SB1_3_29/i0_3 ), .A3(\SB1_3_29/i0_0 ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N3  ( .A1(\SB1_3_29/i0[10] ), .A2(
        \SB1_3_29/i0_4 ), .A3(\SB1_3_29/i0_3 ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N2  ( .A1(\SB1_3_29/i0[8] ), .A2(
        \SB1_3_29/i0[7] ), .A3(\SB1_3_29/i0[6] ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_29/Component_Function_0/N1  ( .A1(\SB1_3_29/i0[10] ), .A2(
        \SB1_3_29/i0[9] ), .ZN(\SB1_3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_1/N4  ( .A1(\SB1_3_29/i1_7 ), .A2(
        \SB1_3_29/i0[8] ), .A3(\SB1_3_29/i0_4 ), .ZN(
        \SB1_3_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_29/Component_Function_1/N3  ( .A1(\SB1_3_29/i1_5 ), .A2(
        \SB1_3_29/i0[6] ), .A3(\SB1_3_29/i0[9] ), .ZN(
        \SB1_3_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_29/Component_Function_1/N2  ( .A1(\SB1_3_29/i0_3 ), .A2(
        \SB1_3_29/i1_7 ), .A3(\SB1_3_29/i0[8] ), .ZN(
        \SB1_3_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_29/Component_Function_1/N1  ( .A1(\SB1_3_29/i0_3 ), .A2(
        \SB1_3_29/i1[9] ), .ZN(\SB1_3_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_5/N4  ( .A1(\SB1_3_29/i0[9] ), .A2(
        \SB1_3_29/i0[6] ), .A3(\SB1_3_29/i0_4 ), .ZN(
        \SB1_3_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_29/Component_Function_5/N2  ( .A1(\SB1_3_29/i0_0 ), .A2(
        \SB1_3_29/i0[6] ), .A3(\SB1_3_29/i0[10] ), .ZN(
        \SB1_3_29/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_29/Component_Function_5/N1  ( .A1(\SB1_3_29/i0_0 ), .A2(
        \SB1_3_29/i3[0] ), .ZN(\SB1_3_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_0/N4  ( .A1(\SB1_3_30/i0[7] ), .A2(
        \SB1_3_30/i0_3 ), .A3(\SB1_3_30/i0_0 ), .ZN(
        \SB1_3_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_30/Component_Function_0/N3  ( .A1(\SB1_3_30/i0[10] ), .A2(
        \SB1_3_30/i0_4 ), .A3(\SB1_3_30/i0_3 ), .ZN(
        \SB1_3_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_30/Component_Function_0/N2  ( .A1(\SB1_3_30/i0[8] ), .A2(
        \SB1_3_30/i0[7] ), .A3(\SB1_3_30/i0[6] ), .ZN(
        \SB1_3_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_30/Component_Function_0/N1  ( .A1(\SB1_3_30/i0[10] ), .A2(
        \SB1_3_30/i0[9] ), .ZN(\SB1_3_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_1/N4  ( .A1(\SB1_3_30/i1_7 ), .A2(
        \SB1_3_30/i0[8] ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_30/Component_Function_1/N2  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i1_7 ), .A3(\SB1_3_30/i0[8] ), .ZN(
        \SB1_3_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_30/Component_Function_1/N1  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i1[9] ), .ZN(\SB1_3_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_5/N4  ( .A1(\SB1_3_30/i0[9] ), .A2(
        \SB1_3_30/i0[6] ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_30/Component_Function_5/N2  ( .A1(\SB1_3_30/i0_0 ), .A2(
        \SB1_3_30/i0[6] ), .A3(\SB1_3_30/i0[10] ), .ZN(
        \SB1_3_30/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_30/Component_Function_5/N1  ( .A1(\SB1_3_30/i0_0 ), .A2(
        \SB1_3_30/i3[0] ), .ZN(\SB1_3_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_31/Component_Function_0/N4  ( .A1(\SB1_3_31/i0[7] ), .A2(
        \SB1_3_31/i0_3 ), .A3(\SB1_3_31/i0_0 ), .ZN(
        \SB1_3_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_31/Component_Function_0/N3  ( .A1(\SB1_3_31/i0[10] ), .A2(
        \SB1_3_31/i0_4 ), .A3(\SB1_3_31/i0_3 ), .ZN(
        \SB1_3_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_31/Component_Function_0/N2  ( .A1(\SB1_3_31/i0[8] ), .A2(
        \SB1_3_31/i0[7] ), .A3(\SB1_3_31/i0[6] ), .ZN(
        \SB1_3_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_31/Component_Function_0/N1  ( .A1(\SB1_3_31/i0[10] ), .A2(
        \SB1_3_31/i0[9] ), .ZN(\SB1_3_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_31/Component_Function_1/N4  ( .A1(\SB1_3_31/i1_7 ), .A2(
        \SB1_3_31/i0[8] ), .A3(\SB1_3_31/i0_4 ), .ZN(
        \SB1_3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_31/Component_Function_1/N3  ( .A1(\SB1_3_31/i1_5 ), .A2(
        \SB1_3_31/i0[6] ), .A3(\SB1_3_31/i0[9] ), .ZN(
        \SB1_3_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_31/Component_Function_1/N2  ( .A1(\SB1_3_31/i0_3 ), .A2(
        \SB1_3_31/i1_7 ), .A3(\SB1_3_31/i0[8] ), .ZN(
        \SB1_3_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_31/Component_Function_1/N1  ( .A1(\SB1_3_31/i0_3 ), .A2(
        \SB1_3_31/i1[9] ), .ZN(\SB1_3_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_31/Component_Function_5/N4  ( .A1(\SB1_3_31/i0[9] ), .A2(
        \SB1_3_31/i0[6] ), .A3(\SB1_3_31/i0_4 ), .ZN(
        \SB1_3_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_31/Component_Function_5/N2  ( .A1(\SB1_3_31/i0_0 ), .A2(
        \SB1_3_31/i0[6] ), .A3(\SB1_3_31/i0[10] ), .ZN(
        \SB1_3_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_31/Component_Function_5/N1  ( .A1(\SB1_3_31/i0_0 ), .A2(
        \SB1_3_31/i3[0] ), .ZN(\SB1_3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_0/N4  ( .A1(\SB2_3_0/i0[7] ), .A2(
        \SB2_3_0/i0_3 ), .A3(\SB2_3_0/i0_0 ), .ZN(
        \SB2_3_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_0/Component_Function_0/N3  ( .A1(\SB2_3_0/i0[10] ), .A2(
        \SB2_3_0/i0_4 ), .A3(\SB2_3_0/i0_3 ), .ZN(
        \SB2_3_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_0/Component_Function_0/N2  ( .A1(\SB2_3_0/i0[8] ), .A2(
        \SB2_3_0/i0[7] ), .A3(\SB2_3_0/i0[6] ), .ZN(
        \SB2_3_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_0/Component_Function_0/N1  ( .A1(\SB2_3_0/i0[10] ), .A2(
        \SB2_3_0/i0[9] ), .ZN(\SB2_3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_1/N4  ( .A1(\SB2_3_0/i1_7 ), .A2(
        \SB2_3_0/i0[8] ), .A3(\SB2_3_0/i0_4 ), .ZN(
        \SB2_3_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_0/Component_Function_1/N3  ( .A1(\SB2_3_0/i1_5 ), .A2(
        \SB2_3_0/i0[6] ), .A3(\SB2_3_0/i0[9] ), .ZN(
        \SB2_3_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_0/Component_Function_1/N2  ( .A1(\SB2_3_0/i0_3 ), .A2(
        \SB2_3_0/i1_7 ), .A3(\SB2_3_0/i0[8] ), .ZN(
        \SB2_3_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_0/Component_Function_1/N1  ( .A1(\SB2_3_0/i0_3 ), .A2(
        \SB2_3_0/i1[9] ), .ZN(\SB2_3_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_5/N4  ( .A1(\SB2_3_0/i0[9] ), .A2(
        \SB2_3_0/i0[6] ), .A3(\SB2_3_0/i0_4 ), .ZN(
        \SB2_3_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_0/Component_Function_5/N2  ( .A1(\SB2_3_0/i0_0 ), .A2(
        \SB2_3_0/i0[6] ), .A3(\SB2_3_0/i0[10] ), .ZN(
        \SB2_3_0/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_0/Component_Function_5/N1  ( .A1(\SB2_3_0/i0_0 ), .A2(
        \SB2_3_0/i3[0] ), .ZN(\SB2_3_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_0/N4  ( .A1(\SB2_3_1/i0[7] ), .A2(
        \SB2_3_1/i0_3 ), .A3(\SB2_3_1/i0_0 ), .ZN(
        \SB2_3_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_1/Component_Function_0/N3  ( .A1(\SB2_3_1/i0[10] ), .A2(
        \SB2_3_1/i0_4 ), .A3(\SB2_3_1/i0_3 ), .ZN(
        \SB2_3_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_1/Component_Function_0/N2  ( .A1(\SB2_3_1/i0[8] ), .A2(
        \SB2_3_1/i0[7] ), .A3(n1637), .ZN(
        \SB2_3_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_1/Component_Function_0/N1  ( .A1(\SB2_3_1/i0[10] ), .A2(
        \SB2_3_1/i0[9] ), .ZN(\SB2_3_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_1/N4  ( .A1(\SB2_3_1/i1_7 ), .A2(
        \SB2_3_1/i0[8] ), .A3(\SB2_3_1/i0_4 ), .ZN(
        \SB2_3_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_1/Component_Function_1/N3  ( .A1(\SB2_3_1/i1_5 ), .A2(n1637), 
        .A3(\SB2_3_1/i0[9] ), .ZN(\SB2_3_1/Component_Function_1/NAND4_in[2] )
         );
  NAND3_X1 \SB2_3_1/Component_Function_1/N2  ( .A1(\SB2_3_1/i0_3 ), .A2(
        \SB2_3_1/i1_7 ), .A3(\SB2_3_1/i0[8] ), .ZN(
        \SB2_3_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_1/Component_Function_1/N1  ( .A1(\SB2_3_1/i0_3 ), .A2(
        \SB2_3_1/i1[9] ), .ZN(\SB2_3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_5/N2  ( .A1(\SB2_3_1/i0_0 ), .A2(n1637), 
        .A3(\SB2_3_1/i0[10] ), .ZN(\SB2_3_1/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X1 \SB2_3_1/Component_Function_5/N1  ( .A1(\SB2_3_1/i0_0 ), .A2(
        \SB2_3_1/i3[0] ), .ZN(\SB2_3_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_0/N4  ( .A1(\SB2_3_2/i0[7] ), .A2(
        \SB2_3_2/i0_3 ), .A3(\SB2_3_2/i0_0 ), .ZN(
        \SB2_3_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_2/Component_Function_0/N3  ( .A1(\SB2_3_2/i0[10] ), .A2(
        \SB2_3_2/i0_4 ), .A3(\SB2_3_2/i0_3 ), .ZN(
        \SB2_3_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_2/Component_Function_0/N2  ( .A1(\SB2_3_2/i0[8] ), .A2(
        \SB2_3_2/i0[7] ), .A3(\SB2_3_2/i0[6] ), .ZN(
        \SB2_3_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_2/Component_Function_0/N1  ( .A1(\SB2_3_2/i0[10] ), .A2(
        \SB2_3_2/i0[9] ), .ZN(\SB2_3_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_1/N4  ( .A1(\SB2_3_2/i1_7 ), .A2(
        \SB2_3_2/i0[8] ), .A3(\SB2_3_2/i0_4 ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_2/Component_Function_1/N3  ( .A1(\SB2_3_2/i1_5 ), .A2(
        \SB2_3_2/i0[6] ), .A3(\SB2_3_2/i0[9] ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_2/Component_Function_1/N2  ( .A1(\SB2_3_2/i0_3 ), .A2(
        \SB2_3_2/i1_7 ), .A3(\SB2_3_2/i0[8] ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_2/Component_Function_5/N4  ( .A1(\SB2_3_2/i0[9] ), .A2(
        \SB2_3_2/i0[6] ), .A3(\SB2_3_2/i0_4 ), .ZN(
        \SB2_3_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_2/Component_Function_5/N2  ( .A1(\SB2_3_2/i0_0 ), .A2(
        \SB2_3_2/i0[6] ), .A3(\SB2_3_2/i0[10] ), .ZN(
        \SB2_3_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_2/Component_Function_5/N1  ( .A1(\SB2_3_2/i0_0 ), .A2(
        \SB2_3_2/i3[0] ), .ZN(\SB2_3_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_0/N4  ( .A1(\SB2_3_3/i0[7] ), .A2(
        \SB2_3_3/i0_3 ), .A3(\SB2_3_3/i0_0 ), .ZN(
        \SB2_3_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_0/N3  ( .A1(\SB2_3_3/i0[10] ), .A2(
        \SB2_3_3/i0_4 ), .A3(\SB2_3_3/i0_3 ), .ZN(
        \SB2_3_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_3/Component_Function_0/N2  ( .A1(\SB2_3_3/i0[8] ), .A2(
        \SB2_3_3/i0[7] ), .A3(\SB2_3_3/i0[6] ), .ZN(
        \SB2_3_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_3/Component_Function_0/N1  ( .A1(\SB2_3_3/i0[10] ), .A2(
        \SB2_3_3/i0[9] ), .ZN(\SB2_3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_1/N4  ( .A1(\SB2_3_3/i1_7 ), .A2(
        \SB2_3_3/i0[8] ), .A3(\SB2_3_3/i0_4 ), .ZN(
        \SB2_3_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_1/N3  ( .A1(\SB2_3_3/i1_5 ), .A2(
        \SB2_3_3/i0[6] ), .A3(\SB2_3_3/i0[9] ), .ZN(
        \SB2_3_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_3/Component_Function_1/N2  ( .A1(\SB2_3_3/i0_3 ), .A2(
        \SB2_3_3/i1_7 ), .A3(\SB2_3_3/i0[8] ), .ZN(
        \SB2_3_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_3/Component_Function_1/N1  ( .A1(\SB2_3_3/i0_3 ), .A2(
        \SB2_3_3/i1[9] ), .ZN(\SB2_3_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_5/N2  ( .A1(\SB2_3_3/i0_0 ), .A2(
        \SB2_3_3/i0[6] ), .A3(\SB2_3_3/i0[10] ), .ZN(
        \SB2_3_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_3/Component_Function_5/N1  ( .A1(\SB2_3_3/i0_0 ), .A2(
        \SB2_3_3/i3[0] ), .ZN(\SB2_3_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_0/N4  ( .A1(\SB2_3_4/i0[7] ), .A2(
        \SB2_3_4/i0_3 ), .A3(\SB2_3_4/i0_0 ), .ZN(
        \SB2_3_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_0/N3  ( .A1(\SB2_3_4/i0[10] ), .A2(
        \SB2_3_4/i0_4 ), .A3(\SB2_3_4/i0_3 ), .ZN(
        \SB2_3_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_4/Component_Function_0/N2  ( .A1(\SB2_3_4/i0[8] ), .A2(
        \SB2_3_4/i0[7] ), .A3(\SB2_3_4/i0[6] ), .ZN(
        \SB2_3_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_4/Component_Function_0/N1  ( .A1(\SB2_3_4/i0[10] ), .A2(
        n2133), .ZN(\SB2_3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_1/N4  ( .A1(\SB2_3_4/i1_7 ), .A2(
        \SB2_3_4/i0[8] ), .A3(\SB2_3_4/i0_4 ), .ZN(
        \SB2_3_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_1/N3  ( .A1(\SB2_3_4/i1_5 ), .A2(
        \SB2_3_4/i0[6] ), .A3(\RI3[3][162] ), .ZN(
        \SB2_3_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_4/Component_Function_1/N2  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i1_7 ), .A3(\SB2_3_4/i0[8] ), .ZN(
        \SB2_3_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_4/Component_Function_1/N1  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i1[9] ), .ZN(\SB2_3_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_5/N4  ( .A1(n2133), .A2(\SB2_3_4/i0[6] ), .A3(\SB2_3_4/i0_4 ), .ZN(\SB2_3_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_5/N2  ( .A1(\SB2_3_4/i0_0 ), .A2(
        \SB2_3_4/i0[6] ), .A3(\SB2_3_4/i0[10] ), .ZN(
        \SB2_3_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_4/Component_Function_5/N1  ( .A1(\SB2_3_4/i0_0 ), .A2(
        \SB2_3_4/i3[0] ), .ZN(\SB2_3_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_0/N4  ( .A1(\SB2_3_5/i0[7] ), .A2(
        \SB2_3_5/i0_3 ), .A3(\SB2_3_5/i0_0 ), .ZN(
        \SB2_3_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_5/Component_Function_0/N3  ( .A1(\SB2_3_5/i0[10] ), .A2(
        \SB2_3_5/i0_4 ), .A3(\SB2_3_5/i0_3 ), .ZN(
        \SB2_3_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_5/Component_Function_0/N2  ( .A1(\SB2_3_5/i0[8] ), .A2(
        \SB2_3_5/i0[7] ), .A3(\SB2_3_5/i0[6] ), .ZN(
        \SB2_3_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_5/Component_Function_0/N1  ( .A1(\SB2_3_5/i0[10] ), .A2(
        n2110), .ZN(\SB2_3_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_1/N4  ( .A1(\SB2_3_5/i1_7 ), .A2(
        \SB2_3_5/i0[8] ), .A3(\SB2_3_5/i0_4 ), .ZN(
        \SB2_3_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_5/Component_Function_1/N3  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[6] ), .A3(n2110), .ZN(
        \SB2_3_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_5/Component_Function_1/N2  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i1_7 ), .A3(\SB2_3_5/i0[8] ), .ZN(
        \SB2_3_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_5/Component_Function_1/N1  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i1[9] ), .ZN(\SB2_3_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_5/N4  ( .A1(\RI3[3][156] ), .A2(
        \SB2_3_5/i0[6] ), .A3(\SB2_3_5/i0_4 ), .ZN(
        \SB2_3_5/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_5/Component_Function_5/N1  ( .A1(\SB2_3_5/i0_0 ), .A2(
        \SB2_3_5/i3[0] ), .ZN(\SB2_3_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_0/N4  ( .A1(\SB2_3_6/i0[7] ), .A2(
        \SB2_3_6/i0_3 ), .A3(\SB2_3_6/i0_0 ), .ZN(
        \SB2_3_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_6/Component_Function_0/N3  ( .A1(\SB2_3_6/i0[10] ), .A2(
        \RI3[3][154] ), .A3(\SB2_3_6/i0_3 ), .ZN(
        \SB2_3_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_6/Component_Function_0/N2  ( .A1(\SB2_3_6/i0[8] ), .A2(
        \SB2_3_6/i0[7] ), .A3(n2143), .ZN(
        \SB2_3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_6/Component_Function_0/N1  ( .A1(\SB2_3_6/i0[10] ), .A2(
        \SB2_3_6/i0[9] ), .ZN(\SB2_3_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_1/N4  ( .A1(\SB2_3_6/i1_7 ), .A2(
        \SB2_3_6/i0[8] ), .A3(\RI3[3][154] ), .ZN(
        \SB2_3_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_6/Component_Function_1/N3  ( .A1(\SB2_3_6/i1_5 ), .A2(n2143), 
        .A3(\SB2_3_6/i0[9] ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[2] )
         );
  NAND3_X1 \SB2_3_6/Component_Function_1/N2  ( .A1(\SB2_3_6/i0_3 ), .A2(
        \SB2_3_6/i1_7 ), .A3(\SB2_3_6/i0[8] ), .ZN(
        \SB2_3_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_6/Component_Function_1/N1  ( .A1(\SB2_3_6/i0_3 ), .A2(
        \SB2_3_6/i1[9] ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_5/N4  ( .A1(\RI3[3][150] ), .A2(
        \RI3[3][151] ), .A3(\RI3[3][154] ), .ZN(
        \SB2_3_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_6/Component_Function_5/N3  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \RI3[3][154] ), .A3(\SB2_3_6/i0_3 ), .ZN(
        \SB2_3_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_6/Component_Function_5/N2  ( .A1(\SB2_3_6/i0_0 ), .A2(
        \RI3[3][151] ), .A3(\SB2_3_6/i0[10] ), .ZN(
        \SB2_3_6/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_6/Component_Function_5/N1  ( .A1(\SB2_3_6/i0_0 ), .A2(
        \SB2_3_6/i3[0] ), .ZN(\SB2_3_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_0/N4  ( .A1(\SB2_3_7/i0[7] ), .A2(
        \SB2_3_7/i0_3 ), .A3(\SB2_3_7/i0_0 ), .ZN(
        \SB2_3_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_7/Component_Function_0/N3  ( .A1(\SB2_3_7/i0[10] ), .A2(
        \SB2_3_7/i0_4 ), .A3(\SB2_3_7/i0_3 ), .ZN(
        \SB2_3_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_7/Component_Function_0/N2  ( .A1(\SB2_3_7/i0[8] ), .A2(
        \SB2_3_7/i0[7] ), .A3(\SB2_3_7/i0[6] ), .ZN(
        \SB2_3_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_7/Component_Function_0/N1  ( .A1(\SB2_3_7/i0[10] ), .A2(
        \SB2_3_7/i0[9] ), .ZN(\SB2_3_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_1/N4  ( .A1(\SB2_3_7/i1_7 ), .A2(
        \SB2_3_7/i0[8] ), .A3(\SB2_3_7/i0_4 ), .ZN(
        \SB2_3_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_7/Component_Function_1/N3  ( .A1(\SB2_3_7/i1_5 ), .A2(
        \SB2_3_7/i0[6] ), .A3(\SB2_3_7/i0[9] ), .ZN(
        \SB2_3_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_7/Component_Function_1/N2  ( .A1(\SB2_3_7/i0_3 ), .A2(
        \SB2_3_7/i1_7 ), .A3(\SB2_3_7/i0[8] ), .ZN(
        \SB2_3_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_7/Component_Function_1/N1  ( .A1(\SB2_3_7/i0_3 ), .A2(
        \SB2_3_7/i1[9] ), .ZN(\SB2_3_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_5/N2  ( .A1(\SB2_3_7/i0_0 ), .A2(
        \SB2_3_7/i0[6] ), .A3(\SB2_3_7/i0[10] ), .ZN(
        \SB2_3_7/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_7/Component_Function_5/N1  ( .A1(\SB2_3_7/i0_0 ), .A2(
        \SB2_3_7/i3[0] ), .ZN(\SB2_3_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_0/N4  ( .A1(\SB2_3_8/i0[7] ), .A2(
        \SB2_3_8/i0_3 ), .A3(\SB2_3_8/i0_0 ), .ZN(
        \SB2_3_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_0/N3  ( .A1(\SB2_3_8/i0[10] ), .A2(
        \SB2_3_8/i0_4 ), .A3(\SB2_3_8/i0_3 ), .ZN(
        \SB2_3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_8/Component_Function_0/N2  ( .A1(\SB2_3_8/i0[8] ), .A2(
        \SB2_3_8/i0[7] ), .A3(\SB2_3_8/i0[6] ), .ZN(
        \SB2_3_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_8/Component_Function_0/N1  ( .A1(\SB2_3_8/i0[10] ), .A2(
        n1639), .ZN(\SB2_3_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_1/N4  ( .A1(\SB2_3_8/i1_7 ), .A2(
        \SB2_3_8/i0[8] ), .A3(\SB2_3_8/i0_4 ), .ZN(
        \SB2_3_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_1/N3  ( .A1(\SB2_3_8/i1_5 ), .A2(
        \SB2_3_8/i0[6] ), .A3(n1639), .ZN(
        \SB2_3_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_8/Component_Function_1/N2  ( .A1(\SB2_3_8/i0_3 ), .A2(
        \SB2_3_8/i1_7 ), .A3(\SB2_3_8/i0[8] ), .ZN(
        \SB2_3_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_8/Component_Function_1/N1  ( .A1(\SB2_3_8/i0_3 ), .A2(
        \SB2_3_8/i1[9] ), .ZN(\SB2_3_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_5/N4  ( .A1(\RI3[3][138] ), .A2(
        \SB2_3_8/i0[6] ), .A3(\SB2_3_8/i0_4 ), .ZN(
        \SB2_3_8/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_8/Component_Function_5/N1  ( .A1(\SB2_3_8/i0_0 ), .A2(
        \SB2_3_8/i3[0] ), .ZN(\SB2_3_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_0/N3  ( .A1(\SB2_3_9/i0[10] ), .A2(
        \SB2_3_9/i0_4 ), .A3(\SB2_3_9/i0_3 ), .ZN(
        \SB2_3_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_9/Component_Function_0/N2  ( .A1(\SB2_3_9/i0[8] ), .A2(
        \SB2_3_9/i0[7] ), .A3(\SB2_3_9/i0[6] ), .ZN(
        \SB2_3_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_9/Component_Function_0/N1  ( .A1(\SB2_3_9/i0[10] ), .A2(n546), .ZN(\SB2_3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_1/N4  ( .A1(\SB2_3_9/i1_7 ), .A2(
        \SB2_3_9/i0[8] ), .A3(\SB2_3_9/i0_4 ), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_9/Component_Function_1/N3  ( .A1(\SB2_3_9/i1_5 ), .A2(
        \SB2_3_9/i0[6] ), .A3(n546), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_9/Component_Function_1/N2  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i1_7 ), .A3(\SB2_3_9/i0[8] ), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_9/Component_Function_1/N1  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i1[9] ), .ZN(\SB2_3_9/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_9/Component_Function_5/N1  ( .A1(\SB2_3_9/i0_0 ), .A2(
        \SB2_3_9/i3[0] ), .ZN(\SB2_3_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_0/N4  ( .A1(\SB2_3_10/i0[7] ), .A2(
        \SB2_3_10/i0_3 ), .A3(\SB2_3_10/i0_0 ), .ZN(
        \SB2_3_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_10/Component_Function_0/N3  ( .A1(\SB2_3_10/i0[10] ), .A2(
        \SB2_3_10/i0_4 ), .A3(\SB2_3_10/i0_3 ), .ZN(
        \SB2_3_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_10/Component_Function_0/N2  ( .A1(\SB2_3_10/i0[8] ), .A2(
        \SB2_3_10/i0[7] ), .A3(\SB2_3_10/i0[6] ), .ZN(
        \SB2_3_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_10/Component_Function_0/N1  ( .A1(\SB2_3_10/i0[10] ), .A2(
        \SB2_3_10/i0[9] ), .ZN(\SB2_3_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_1/N4  ( .A1(\SB2_3_10/i1_7 ), .A2(
        \SB2_3_10/i0[8] ), .A3(\SB2_3_10/i0_4 ), .ZN(
        \SB2_3_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_10/Component_Function_1/N3  ( .A1(\SB2_3_10/i1_5 ), .A2(
        \SB2_3_10/i0[6] ), .A3(\SB2_3_10/i0[9] ), .ZN(
        \SB2_3_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_10/Component_Function_1/N2  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i1_7 ), .A3(\SB2_3_10/i0[8] ), .ZN(
        \SB2_3_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_10/Component_Function_1/N1  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i1[9] ), .ZN(\SB2_3_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_5/N4  ( .A1(\RI3[3][126] ), .A2(
        \SB2_3_10/i0[6] ), .A3(\SB2_3_10/i0_4 ), .ZN(
        \SB2_3_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_10/Component_Function_5/N2  ( .A1(\SB2_3_10/i0_0 ), .A2(
        \SB2_3_10/i0[6] ), .A3(\SB2_3_10/i0[10] ), .ZN(
        \SB2_3_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_10/Component_Function_5/N1  ( .A1(\SB2_3_10/i0_0 ), .A2(
        \SB2_3_10/i3[0] ), .ZN(\SB2_3_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_0/N4  ( .A1(\SB2_3_11/i0[7] ), .A2(
        \SB2_3_11/i0_3 ), .A3(\SB2_3_11/i0_0 ), .ZN(
        \SB2_3_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_0/N3  ( .A1(\SB2_3_11/i0[10] ), .A2(
        \RI3[3][124] ), .A3(\SB2_3_11/i0_3 ), .ZN(
        \SB2_3_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_11/Component_Function_0/N2  ( .A1(\SB2_3_11/i0[8] ), .A2(
        \SB2_3_11/i0[7] ), .A3(\SB2_3_11/i0[6] ), .ZN(
        \SB2_3_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_11/Component_Function_0/N1  ( .A1(\SB2_3_11/i0[10] ), .A2(
        \SB2_3_11/i0[9] ), .ZN(\SB2_3_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_1/N4  ( .A1(\SB2_3_11/i1_7 ), .A2(
        \SB2_3_11/i0[8] ), .A3(\RI3[3][124] ), .ZN(
        \SB2_3_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_1/N3  ( .A1(\SB2_3_11/i1_5 ), .A2(
        \SB2_3_11/i0[6] ), .A3(\SB2_3_11/i0[9] ), .ZN(
        \SB2_3_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_11/Component_Function_1/N2  ( .A1(\SB2_3_11/i0_3 ), .A2(
        \SB2_3_11/i1_7 ), .A3(\SB2_3_11/i0[8] ), .ZN(
        \SB2_3_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_11/Component_Function_1/N1  ( .A1(\SB2_3_11/i0_3 ), .A2(
        \SB2_3_11/i1[9] ), .ZN(\SB2_3_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_5/N4  ( .A1(\SB2_3_11/i0[9] ), .A2(
        \SB2_3_11/i0[6] ), .A3(\RI3[3][124] ), .ZN(
        \SB2_3_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_5/N3  ( .A1(\SB2_3_11/i1[9] ), .A2(
        \RI3[3][124] ), .A3(\SB2_3_11/i0_3 ), .ZN(
        \SB2_3_11/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_11/Component_Function_5/N1  ( .A1(\SB2_3_11/i0_0 ), .A2(
        \SB2_3_11/i3[0] ), .ZN(\SB2_3_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_0/N4  ( .A1(\SB2_3_12/i0[7] ), .A2(
        \SB2_3_12/i0_3 ), .A3(\SB2_3_12/i0_0 ), .ZN(
        \SB2_3_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_0/N3  ( .A1(\SB2_3_12/i0[10] ), .A2(
        \SB2_3_12/i0_4 ), .A3(\SB2_3_12/i0_3 ), .ZN(
        \SB2_3_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_12/Component_Function_0/N2  ( .A1(\SB2_3_12/i0[8] ), .A2(
        \SB2_3_12/i0[7] ), .A3(\SB2_3_12/i0[6] ), .ZN(
        \SB2_3_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_12/Component_Function_0/N1  ( .A1(\SB2_3_12/i0[10] ), .A2(
        \SB2_3_12/i0[9] ), .ZN(\SB2_3_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_1/N4  ( .A1(\SB2_3_12/i1_7 ), .A2(
        \SB2_3_12/i0[8] ), .A3(\SB2_3_12/i0_4 ), .ZN(
        \SB2_3_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_1/N3  ( .A1(\SB2_3_12/i1_5 ), .A2(
        \SB2_3_12/i0[6] ), .A3(\SB2_3_12/i0[9] ), .ZN(
        \SB2_3_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_12/Component_Function_1/N2  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i1_7 ), .A3(\SB2_3_12/i0[8] ), .ZN(
        \SB2_3_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_12/Component_Function_1/N1  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i1[9] ), .ZN(\SB2_3_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_5/N4  ( .A1(\SB2_3_12/i0[9] ), .A2(
        \SB2_3_12/i0[6] ), .A3(\SB2_3_12/i0_4 ), .ZN(
        \SB2_3_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_5/N2  ( .A1(\SB2_3_12/i0_0 ), .A2(
        \SB2_3_12/i0[6] ), .A3(\SB2_3_12/i0[10] ), .ZN(
        \SB2_3_12/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_12/Component_Function_5/N1  ( .A1(\SB2_3_12/i0_0 ), .A2(
        \SB2_3_12/i3[0] ), .ZN(\SB2_3_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_0/N4  ( .A1(\SB2_3_13/i0[7] ), .A2(
        \SB2_3_13/i0_3 ), .A3(\SB2_3_13/i0_0 ), .ZN(
        \SB2_3_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_13/Component_Function_0/N3  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i0_4 ), .A3(\SB2_3_13/i0[10] ), .ZN(
        \SB2_3_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_0/N2  ( .A1(\SB2_3_13/i0[8] ), .A2(
        \SB2_3_13/i0[7] ), .A3(\SB2_3_13/i0[6] ), .ZN(
        \SB2_3_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_13/Component_Function_0/N1  ( .A1(\SB2_3_13/i0[10] ), .A2(
        n2107), .ZN(\SB2_3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_1/N4  ( .A1(\SB2_3_13/i1_7 ), .A2(
        \SB2_3_13/i0[8] ), .A3(\SB2_3_13/i0_4 ), .ZN(
        \SB2_3_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_13/Component_Function_1/N3  ( .A1(\SB2_3_13/i1_5 ), .A2(
        \SB2_3_13/i0[6] ), .A3(n2107), .ZN(
        \SB2_3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_1/N2  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i1_7 ), .A3(\SB2_3_13/i0[8] ), .ZN(
        \SB2_3_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_13/Component_Function_1/N1  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i1[9] ), .ZN(\SB2_3_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_5/N3  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i0_4 ), .A3(\SB2_3_13/i1[9] ), .ZN(
        \SB2_3_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_5/N2  ( .A1(\SB2_3_13/i0_0 ), .A2(
        \SB2_3_13/i0[6] ), .A3(\SB2_3_13/i0[10] ), .ZN(
        \SB2_3_13/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_13/Component_Function_5/N1  ( .A1(\SB2_3_13/i0_0 ), .A2(
        \SB2_3_13/i3[0] ), .ZN(\SB2_3_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_0/N4  ( .A1(\SB2_3_14/i0[7] ), .A2(
        \SB2_3_14/i0_3 ), .A3(\SB2_3_14/i0_0 ), .ZN(
        \SB2_3_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_0/N3  ( .A1(\SB2_3_14/i0[10] ), .A2(
        n1945), .A3(\SB2_3_14/i0_3 ), .ZN(
        \SB2_3_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_14/Component_Function_0/N2  ( .A1(\SB2_3_14/i0[8] ), .A2(
        \SB2_3_14/i0[7] ), .A3(\SB2_3_14/i0[6] ), .ZN(
        \SB2_3_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_14/Component_Function_0/N1  ( .A1(\SB2_3_14/i0[10] ), .A2(
        \SB2_3_14/i0[9] ), .ZN(\SB2_3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_1/N4  ( .A1(\SB2_3_14/i1_7 ), .A2(
        \SB2_3_14/i0[8] ), .A3(n1945), .ZN(
        \SB2_3_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_1/N3  ( .A1(\SB2_3_14/i1_5 ), .A2(
        \SB2_3_14/i0[6] ), .A3(\SB2_3_14/i0[9] ), .ZN(
        \SB2_3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_14/Component_Function_1/N2  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i1_7 ), .A3(\SB2_3_14/i0[8] ), .ZN(
        \SB2_3_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_14/Component_Function_1/N1  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i1[9] ), .ZN(\SB2_3_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_5/N4  ( .A1(\SB2_3_14/i0[9] ), .A2(
        \SB2_3_14/i0[6] ), .A3(\RI3[3][106] ), .ZN(
        \SB2_3_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_5/N2  ( .A1(\SB2_3_14/i0_0 ), .A2(
        \SB2_3_14/i0[6] ), .A3(\SB2_3_14/i0[10] ), .ZN(
        \SB2_3_14/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_14/Component_Function_5/N1  ( .A1(\SB2_3_14/i0_0 ), .A2(
        \SB2_3_14/i3[0] ), .ZN(\SB2_3_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_0/N4  ( .A1(\SB2_3_15/i0[7] ), .A2(
        \SB2_3_15/i0_3 ), .A3(\SB2_3_15/i0_0 ), .ZN(
        \SB2_3_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_15/Component_Function_0/N3  ( .A1(\SB2_3_15/i0[10] ), .A2(
        \SB2_3_15/i0_4 ), .A3(\SB2_3_15/i0_3 ), .ZN(
        \SB2_3_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_15/Component_Function_0/N2  ( .A1(\SB2_3_15/i0[8] ), .A2(
        \SB2_3_15/i0[7] ), .A3(n2097), .ZN(
        \SB2_3_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_15/Component_Function_0/N1  ( .A1(\SB2_3_15/i0[10] ), .A2(
        \SB2_3_15/i0[9] ), .ZN(\SB2_3_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_1/N4  ( .A1(n1965), .A2(
        \SB2_3_15/i0[8] ), .A3(\SB2_3_15/i0_4 ), .ZN(
        \SB2_3_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_15/Component_Function_1/N3  ( .A1(\SB2_3_15/i1_5 ), .A2(
        n2097), .A3(\SB2_3_15/i0[9] ), .ZN(
        \SB2_3_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_15/Component_Function_1/N2  ( .A1(\SB2_3_15/i0_3 ), .A2(
        n1965), .A3(\SB2_3_15/i0[8] ), .ZN(
        \SB2_3_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_15/Component_Function_1/N1  ( .A1(\SB2_3_15/i0_3 ), .A2(
        \SB2_3_15/i1[9] ), .ZN(\SB2_3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_5/N4  ( .A1(\SB2_3_15/i0[9] ), .A2(
        n2097), .A3(\SB2_3_15/i0_4 ), .ZN(
        \SB2_3_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_15/Component_Function_5/N2  ( .A1(\SB2_3_15/i0_0 ), .A2(
        n2097), .A3(\SB2_3_15/i0[10] ), .ZN(
        \SB2_3_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_15/Component_Function_5/N1  ( .A1(\SB2_3_15/i0_0 ), .A2(
        \SB2_3_15/i3[0] ), .ZN(\SB2_3_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_0/N4  ( .A1(n2134), .A2(
        \SB2_3_16/i0_3 ), .A3(\SB2_3_16/i0_0 ), .ZN(
        \SB2_3_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_16/Component_Function_0/N3  ( .A1(\SB2_3_16/i0[10] ), .A2(
        \RI3[3][94] ), .A3(\SB2_3_16/i0_3 ), .ZN(
        \SB2_3_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_16/Component_Function_0/N2  ( .A1(\SB2_3_16/i0[8] ), .A2(
        n2134), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_16/Component_Function_0/N1  ( .A1(\SB2_3_16/i0[10] ), .A2(
        n2114), .ZN(\SB2_3_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_1/N4  ( .A1(\SB2_3_16/i1_7 ), .A2(
        \SB2_3_16/i0[8] ), .A3(\RI3[3][94] ), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_16/Component_Function_1/N3  ( .A1(\SB2_3_16/i1_5 ), .A2(
        \SB2_3_16/i0[6] ), .A3(n2114), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_16/Component_Function_1/N2  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i1_7 ), .A3(\SB2_3_16/i0[8] ), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_16/Component_Function_1/N1  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i1[9] ), .ZN(\SB2_3_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_5/N4  ( .A1(\RI3[3][90] ), .A2(
        \SB2_3_16/i0[6] ), .A3(\RI3[3][94] ), .ZN(
        \SB2_3_16/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_16/Component_Function_5/N1  ( .A1(\SB2_3_16/i0_0 ), .A2(
        \SB2_3_16/i3[0] ), .ZN(\SB2_3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_17/Component_Function_0/N3  ( .A1(\SB2_3_17/i0[10] ), .A2(
        \SB2_3_17/i0_4 ), .A3(\SB2_3_17/i0_3 ), .ZN(
        \SB2_3_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_17/Component_Function_0/N2  ( .A1(\SB2_3_17/i0[8] ), .A2(
        \SB2_3_17/i0[7] ), .A3(\SB2_3_17/i0[6] ), .ZN(
        \SB2_3_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_17/Component_Function_0/N1  ( .A1(\SB2_3_17/i0[10] ), .A2(
        \SB2_3_17/i0[9] ), .ZN(\SB2_3_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_17/Component_Function_1/N4  ( .A1(\SB2_3_17/i1_7 ), .A2(
        \SB2_3_17/i0[8] ), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_1/N3  ( .A1(\SB2_3_17/i1_5 ), .A2(
        \SB2_3_17/i0[6] ), .A3(\SB2_3_17/i0[9] ), .ZN(
        \SB2_3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_17/Component_Function_1/N2  ( .A1(\SB2_3_17/i0_3 ), .A2(
        \SB2_3_17/i1_7 ), .A3(\SB2_3_17/i0[8] ), .ZN(
        \SB2_3_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_17/Component_Function_1/N1  ( .A1(\SB2_3_17/i0_3 ), .A2(
        \SB2_3_17/i1[9] ), .ZN(\SB2_3_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_17/Component_Function_5/N1  ( .A1(\SB2_3_17/i0_0 ), .A2(
        \SB2_3_17/i3[0] ), .ZN(\SB2_3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_0/N4  ( .A1(\SB2_3_18/i0[7] ), .A2(
        \SB2_3_18/i0_3 ), .A3(\SB2_3_18/i0_0 ), .ZN(
        \SB2_3_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_18/Component_Function_0/N3  ( .A1(\SB2_3_18/i0[10] ), .A2(
        \SB2_3_18/i0_4 ), .A3(\SB2_3_18/i0_3 ), .ZN(
        \SB2_3_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_18/Component_Function_0/N2  ( .A1(\SB2_3_18/i0[8] ), .A2(
        \SB2_3_18/i0[7] ), .A3(\SB2_3_18/i0[6] ), .ZN(
        \SB2_3_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_18/Component_Function_0/N1  ( .A1(\SB2_3_18/i0[10] ), .A2(
        \SB2_3_18/i0[9] ), .ZN(\SB2_3_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_1/N4  ( .A1(\SB2_3_18/i1_7 ), .A2(
        \SB2_3_18/i0[8] ), .A3(\SB2_3_18/i0_4 ), .ZN(
        \SB2_3_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_18/Component_Function_1/N3  ( .A1(\SB2_3_18/i1_5 ), .A2(
        \SB2_3_18/i0[6] ), .A3(\SB2_3_18/i0[9] ), .ZN(
        \SB2_3_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_18/Component_Function_1/N2  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i1_7 ), .A3(\SB2_3_18/i0[8] ), .ZN(
        \SB2_3_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_18/Component_Function_1/N1  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i1[9] ), .ZN(\SB2_3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_5/N4  ( .A1(\SB2_3_18/i0[9] ), .A2(
        \SB2_3_18/i0[6] ), .A3(\SB2_3_18/i0_4 ), .ZN(
        \SB2_3_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_18/Component_Function_5/N3  ( .A1(\SB2_3_18/i1[9] ), .A2(
        \SB2_3_18/i0_4 ), .A3(\SB2_3_18/i0_3 ), .ZN(
        \SB2_3_18/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_18/Component_Function_5/N1  ( .A1(\SB2_3_18/i0_0 ), .A2(
        \SB2_3_18/i3[0] ), .ZN(\SB2_3_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_0/N4  ( .A1(\SB2_3_19/i0[7] ), .A2(
        \SB2_3_19/i0_3 ), .A3(\SB2_3_19/i0_0 ), .ZN(
        \SB2_3_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_19/Component_Function_0/N3  ( .A1(\SB2_3_19/i0[10] ), .A2(
        \SB2_3_19/i0_4 ), .A3(\SB2_3_19/i0_3 ), .ZN(
        \SB2_3_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_19/Component_Function_0/N2  ( .A1(\SB2_3_19/i0[8] ), .A2(
        \SB2_3_19/i0[7] ), .A3(\SB2_3_19/i0[6] ), .ZN(
        \SB2_3_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_19/Component_Function_0/N1  ( .A1(\SB2_3_19/i0[10] ), .A2(
        n1623), .ZN(\SB2_3_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_1/N4  ( .A1(\SB2_3_19/i1_7 ), .A2(
        \SB2_3_19/i0[8] ), .A3(\SB2_3_19/i0_4 ), .ZN(
        \SB2_3_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_19/Component_Function_1/N3  ( .A1(\SB2_3_19/i1_5 ), .A2(
        \SB2_3_19/i0[6] ), .A3(n1623), .ZN(
        \SB2_3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_19/Component_Function_1/N2  ( .A1(\SB2_3_19/i0_3 ), .A2(
        \SB2_3_19/i1_7 ), .A3(\SB2_3_19/i0[8] ), .ZN(
        \SB2_3_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_19/Component_Function_1/N1  ( .A1(\SB2_3_19/i0_3 ), .A2(
        \SB2_3_19/i1[9] ), .ZN(\SB2_3_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_19/Component_Function_5/N1  ( .A1(\SB2_3_19/i0_0 ), .A2(
        \SB2_3_19/i3[0] ), .ZN(\SB2_3_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_0/N4  ( .A1(\SB2_3_20/i0[7] ), .A2(
        \SB2_3_20/i0_3 ), .A3(\SB2_3_20/i0_0 ), .ZN(
        \SB2_3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_0/N3  ( .A1(\SB2_3_20/i0[10] ), .A2(
        \SB2_3_20/i0_3 ), .A3(\SB2_3_20/i0_4 ), .ZN(
        \SB2_3_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_20/Component_Function_0/N2  ( .A1(\SB2_3_20/i0[8] ), .A2(
        \SB2_3_20/i0[7] ), .A3(\SB2_3_20/i0[6] ), .ZN(
        \SB2_3_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_20/Component_Function_0/N1  ( .A1(\SB2_3_20/i0[10] ), .A2(
        \SB2_3_20/i0[9] ), .ZN(\SB2_3_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_1/N4  ( .A1(\SB2_3_20/i1_7 ), .A2(
        \SB2_3_20/i0[8] ), .A3(\SB2_3_20/i0_4 ), .ZN(
        \SB2_3_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_1/N3  ( .A1(\SB2_3_20/i1_5 ), .A2(
        \SB2_3_20/i0[6] ), .A3(\SB2_3_20/i0[9] ), .ZN(
        \SB2_3_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_20/Component_Function_1/N2  ( .A1(\SB2_3_20/i0_3 ), .A2(
        \SB2_3_20/i1_7 ), .A3(\SB2_3_20/i0[8] ), .ZN(
        \SB2_3_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_20/Component_Function_1/N1  ( .A1(\SB2_3_20/i0_3 ), .A2(
        \SB2_3_20/i1[9] ), .ZN(\SB2_3_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_5/N4  ( .A1(\SB2_3_20/i0[9] ), .A2(
        \SB2_3_20/i0[6] ), .A3(\SB2_3_20/i0_4 ), .ZN(
        \SB2_3_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_5/N2  ( .A1(\SB2_3_20/i0_0 ), .A2(
        \RI3[3][67] ), .A3(\SB2_3_20/i0[10] ), .ZN(
        \SB2_3_20/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_20/Component_Function_5/N1  ( .A1(\SB2_3_20/i0_0 ), .A2(
        \SB2_3_20/i3[0] ), .ZN(\SB2_3_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_0/N4  ( .A1(\SB2_3_21/i0[7] ), .A2(
        \SB2_3_21/i0_3 ), .A3(\SB2_3_21/i0_0 ), .ZN(
        \SB2_3_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_21/Component_Function_0/N3  ( .A1(\SB2_3_21/i0[10] ), .A2(
        \RI3[3][64] ), .A3(\SB2_3_21/i0_3 ), .ZN(
        \SB2_3_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_21/Component_Function_0/N2  ( .A1(\SB2_3_21/i0[8] ), .A2(
        \SB2_3_21/i0[7] ), .A3(\SB2_3_21/i0[6] ), .ZN(
        \SB2_3_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_21/Component_Function_0/N1  ( .A1(\SB2_3_21/i0[10] ), .A2(
        \SB2_3_21/i0[9] ), .ZN(\SB2_3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_1/N4  ( .A1(\SB2_3_21/i1_7 ), .A2(
        \SB2_3_21/i0[8] ), .A3(\RI3[3][64] ), .ZN(
        \SB2_3_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_21/Component_Function_1/N3  ( .A1(\SB2_3_21/i1_5 ), .A2(
        \SB2_3_21/i0[6] ), .A3(\SB2_3_21/i0[9] ), .ZN(
        \SB2_3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_21/Component_Function_1/N2  ( .A1(\SB2_3_21/i0_3 ), .A2(
        \SB2_3_21/i1_7 ), .A3(\SB2_3_21/i0[8] ), .ZN(
        \SB2_3_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_21/Component_Function_1/N1  ( .A1(\SB2_3_21/i0_3 ), .A2(
        \SB2_3_21/i1[9] ), .ZN(\SB2_3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_5/N4  ( .A1(\SB2_3_21/i0[9] ), .A2(
        \SB2_3_21/i0[6] ), .A3(\RI3[3][64] ), .ZN(
        \SB2_3_21/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_21/Component_Function_5/N1  ( .A1(\SB2_3_21/i0_0 ), .A2(
        \SB2_3_21/i3[0] ), .ZN(\SB2_3_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_0/N4  ( .A1(\SB2_3_22/i0[7] ), .A2(
        \SB2_3_22/i0_3 ), .A3(\SB2_3_22/i0_0 ), .ZN(
        \SB2_3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_22/Component_Function_0/N3  ( .A1(\SB2_3_22/i0[10] ), .A2(
        \SB2_3_22/i0_4 ), .A3(\SB2_3_22/i0_3 ), .ZN(
        \SB2_3_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_22/Component_Function_0/N2  ( .A1(\SB2_3_22/i0[8] ), .A2(
        \SB2_3_22/i0[7] ), .A3(\SB2_3_22/i0[6] ), .ZN(
        \SB2_3_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_22/Component_Function_0/N1  ( .A1(\SB2_3_22/i0[10] ), .A2(
        \SB2_3_22/i0[9] ), .ZN(\SB2_3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_1/N4  ( .A1(\SB2_3_22/i1_7 ), .A2(
        \SB2_3_22/i0[8] ), .A3(\SB2_3_22/i0_4 ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_22/Component_Function_1/N3  ( .A1(\SB2_3_22/i1_5 ), .A2(
        \SB2_3_22/i0[6] ), .A3(\SB2_3_22/i0[9] ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_22/Component_Function_1/N2  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i1_7 ), .A3(\SB2_3_22/i0[8] ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_22/Component_Function_1/N1  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i1[9] ), .ZN(\SB2_3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_5/N4  ( .A1(\SB2_3_22/i0[9] ), .A2(
        \RI3[3][55] ), .A3(\SB2_3_22/i0_4 ), .ZN(
        \SB2_3_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_22/Component_Function_5/N2  ( .A1(\SB2_3_22/i0_0 ), .A2(
        \SB2_3_22/i0[6] ), .A3(\SB2_3_22/i0[10] ), .ZN(
        \SB2_3_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_22/Component_Function_5/N1  ( .A1(\SB2_3_22/i0_0 ), .A2(
        \SB2_3_22/i3[0] ), .ZN(\SB2_3_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_0/N4  ( .A1(\SB2_3_23/i0[7] ), .A2(
        \SB2_3_23/i0_3 ), .A3(\SB2_3_23/i0_0 ), .ZN(
        \SB2_3_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_23/Component_Function_0/N3  ( .A1(\SB2_3_23/i0[10] ), .A2(
        \SB2_3_23/i0_4 ), .A3(\SB2_3_23/i0_3 ), .ZN(
        \SB2_3_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_23/Component_Function_0/N2  ( .A1(\SB2_3_23/i0[8] ), .A2(
        \SB2_3_23/i0[7] ), .A3(\SB2_3_23/i0[6] ), .ZN(
        \SB2_3_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_23/Component_Function_0/N1  ( .A1(\SB2_3_23/i0[10] ), .A2(
        \SB2_3_23/i0[9] ), .ZN(\SB2_3_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_1/N4  ( .A1(\SB2_3_23/i1_7 ), .A2(
        \SB2_3_23/i0[8] ), .A3(\SB2_3_23/i0_4 ), .ZN(
        \SB2_3_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_23/Component_Function_1/N3  ( .A1(\SB2_3_23/i1_5 ), .A2(
        \SB2_3_23/i0[6] ), .A3(\SB2_3_23/i0[9] ), .ZN(
        \SB2_3_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_23/Component_Function_1/N2  ( .A1(\SB2_3_23/i0_3 ), .A2(
        \SB2_3_23/i1_7 ), .A3(\SB2_3_23/i0[8] ), .ZN(
        \SB2_3_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_23/Component_Function_1/N1  ( .A1(\SB2_3_23/i0_3 ), .A2(
        \SB2_3_23/i1[9] ), .ZN(\SB2_3_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_5/N4  ( .A1(\SB2_3_23/i0[9] ), .A2(
        \SB2_3_23/i0[6] ), .A3(\SB2_3_23/i0_4 ), .ZN(
        \SB2_3_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_0/N4  ( .A1(\SB2_3_24/i0[7] ), .A2(
        \SB2_3_24/i0_3 ), .A3(\SB2_3_24/i0_0 ), .ZN(
        \SB2_3_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_0/N3  ( .A1(\SB2_3_24/i0[10] ), .A2(
        \SB2_3_24/i0_4 ), .A3(\SB2_3_24/i0_3 ), .ZN(
        \SB2_3_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_24/Component_Function_0/N2  ( .A1(\SB2_3_24/i0[8] ), .A2(
        \SB2_3_24/i0[7] ), .A3(\SB2_3_24/i0[6] ), .ZN(
        \SB2_3_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_24/Component_Function_0/N1  ( .A1(\SB2_3_24/i0[10] ), .A2(
        \SB2_3_24/i0[9] ), .ZN(\SB2_3_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_24/Component_Function_1/N4  ( .A1(\SB2_3_24/i1_7 ), .A2(
        \SB2_3_24/i0[8] ), .A3(\SB2_3_24/i0_4 ), .ZN(
        \SB2_3_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_1/N3  ( .A1(\SB2_3_24/i1_5 ), .A2(
        \SB2_3_24/i0[6] ), .A3(\SB2_3_24/i0[9] ), .ZN(
        \SB2_3_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_24/Component_Function_1/N2  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB2_3_24/i1_7 ), .A3(\SB2_3_24/i0[8] ), .ZN(
        \SB2_3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_24/Component_Function_1/N1  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB2_3_24/i1[9] ), .ZN(\SB2_3_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_24/Component_Function_5/N2  ( .A1(\SB2_3_24/i0_0 ), .A2(
        \SB2_3_24/i0[6] ), .A3(\SB2_3_24/i0[10] ), .ZN(
        \SB2_3_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_24/Component_Function_5/N1  ( .A1(\SB2_3_24/i0_0 ), .A2(
        \SB2_3_24/i3[0] ), .ZN(\SB2_3_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_25/Component_Function_0/N4  ( .A1(\SB2_3_25/i0[7] ), .A2(
        \SB2_3_25/i0_3 ), .A3(\SB2_3_25/i0_0 ), .ZN(
        \SB2_3_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_25/Component_Function_0/N3  ( .A1(\SB2_3_25/i0[10] ), .A2(
        \SB2_3_25/i0_4 ), .A3(\SB2_3_25/i0_3 ), .ZN(
        \SB2_3_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_25/Component_Function_0/N2  ( .A1(\SB2_3_25/i0[8] ), .A2(
        \SB2_3_25/i0[7] ), .A3(\SB2_3_25/i0[6] ), .ZN(
        \SB2_3_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_25/Component_Function_0/N1  ( .A1(\SB2_3_25/i0[10] ), .A2(
        \SB2_3_25/i0[9] ), .ZN(\SB2_3_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_25/Component_Function_1/N4  ( .A1(\SB2_3_25/i1_7 ), .A2(
        \SB2_3_25/i0[8] ), .A3(\SB2_3_25/i0_4 ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_25/Component_Function_1/N3  ( .A1(\SB2_3_25/i1_5 ), .A2(
        \SB2_3_25/i0[6] ), .A3(\SB2_3_25/i0[9] ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_25/Component_Function_1/N2  ( .A1(\SB2_3_25/i0_3 ), .A2(
        \SB2_3_25/i1_7 ), .A3(\SB2_3_25/i0[8] ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_25/Component_Function_1/N1  ( .A1(\SB2_3_25/i0_3 ), .A2(
        \SB2_3_25/i1[9] ), .ZN(\SB2_3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_25/Component_Function_5/N4  ( .A1(\SB2_3_25/i0[9] ), .A2(
        \RI3[3][37] ), .A3(\SB2_3_25/i0_4 ), .ZN(
        \SB2_3_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_25/Component_Function_5/N2  ( .A1(\SB2_3_25/i0_0 ), .A2(
        \SB2_3_25/i0[6] ), .A3(\SB2_3_25/i0[10] ), .ZN(
        \SB2_3_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_25/Component_Function_5/N1  ( .A1(\SB2_3_25/i0_0 ), .A2(
        \SB2_3_25/i3[0] ), .ZN(\SB2_3_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_0/N4  ( .A1(\SB2_3_26/i0[7] ), .A2(
        \SB2_3_26/i0_3 ), .A3(\SB2_3_26/i0_0 ), .ZN(
        \SB2_3_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_26/Component_Function_0/N3  ( .A1(\SB2_3_26/i0[10] ), .A2(
        \SB2_3_26/i0_4 ), .A3(\SB2_3_26/i0_3 ), .ZN(
        \SB2_3_26/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_26/Component_Function_0/N1  ( .A1(\SB2_3_26/i0[10] ), .A2(
        \SB2_3_26/i0[9] ), .ZN(\SB2_3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_1/N4  ( .A1(\SB2_3_26/i1_7 ), .A2(
        \SB2_3_26/i0[8] ), .A3(\SB2_3_26/i0_4 ), .ZN(
        \SB2_3_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_26/Component_Function_1/N3  ( .A1(\SB2_3_26/i1_5 ), .A2(
        \SB2_3_26/i0[6] ), .A3(\SB2_3_26/i0[9] ), .ZN(
        \SB2_3_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_26/Component_Function_1/N2  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i1_7 ), .A3(\SB2_3_26/i0[8] ), .ZN(
        \SB2_3_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_26/Component_Function_1/N1  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i1[9] ), .ZN(\SB2_3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_5/N4  ( .A1(\SB2_3_26/i0[9] ), .A2(
        \SB2_3_26/i0[6] ), .A3(\SB2_3_26/i0_4 ), .ZN(
        \SB2_3_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_27/Component_Function_0/N4  ( .A1(\SB2_3_27/i0[7] ), .A2(
        \SB2_3_27/i0_3 ), .A3(\SB2_3_27/i0_0 ), .ZN(
        \SB2_3_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_27/Component_Function_0/N3  ( .A1(\SB2_3_27/i0[10] ), .A2(
        \SB2_3_27/i0_4 ), .A3(\SB2_3_27/i0_3 ), .ZN(
        \SB2_3_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_27/Component_Function_0/N2  ( .A1(\SB2_3_27/i0[8] ), .A2(
        \SB2_3_27/i0[7] ), .A3(\SB2_3_27/i0[6] ), .ZN(
        \SB2_3_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_27/Component_Function_0/N1  ( .A1(\SB2_3_27/i0[10] ), .A2(
        \SB2_3_27/i0[9] ), .ZN(\SB2_3_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_1/N4  ( .A1(\SB2_3_27/i1_7 ), .A2(
        \SB2_3_27/i0[8] ), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_27/Component_Function_1/N2  ( .A1(\SB2_3_27/i0_3 ), .A2(
        \SB2_3_27/i1_7 ), .A3(\SB2_3_27/i0[8] ), .ZN(
        \SB2_3_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_27/Component_Function_1/N1  ( .A1(\SB2_3_27/i0_3 ), .A2(
        \SB2_3_27/i1[9] ), .ZN(\SB2_3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_5/N4  ( .A1(\RI3[3][24] ), .A2(
        \SB2_3_27/i0[6] ), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_27/Component_Function_5/N1  ( .A1(\SB2_3_27/i0_0 ), .A2(
        \SB2_3_27/i3[0] ), .ZN(\SB2_3_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_0/N4  ( .A1(\SB2_3_28/i0[7] ), .A2(
        \SB2_3_28/i0_3 ), .A3(\SB2_3_28/i0_0 ), .ZN(
        \SB2_3_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_28/Component_Function_0/N3  ( .A1(\SB2_3_28/i0[10] ), .A2(
        \SB2_3_28/i0_4 ), .A3(\SB2_3_28/i0_3 ), .ZN(
        \SB2_3_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_28/Component_Function_0/N2  ( .A1(\SB2_3_28/i0[8] ), .A2(
        \SB2_3_28/i0[7] ), .A3(\SB2_3_28/i0[6] ), .ZN(
        \SB2_3_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_28/Component_Function_0/N1  ( .A1(\SB2_3_28/i0[10] ), .A2(
        \SB2_3_28/i0[9] ), .ZN(\SB2_3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_1/N4  ( .A1(\SB2_3_28/i1_7 ), .A2(
        \SB2_3_28/i0[8] ), .A3(\SB2_3_28/i0_4 ), .ZN(
        \SB2_3_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_28/Component_Function_1/N3  ( .A1(\SB2_3_28/i1_5 ), .A2(
        \SB2_3_28/i0[6] ), .A3(\SB2_3_28/i0[9] ), .ZN(
        \SB2_3_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_28/Component_Function_1/N2  ( .A1(\SB2_3_28/i0_3 ), .A2(
        \SB2_3_28/i1_7 ), .A3(\SB2_3_28/i0[8] ), .ZN(
        \SB2_3_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_28/Component_Function_1/N1  ( .A1(\SB2_3_28/i0_3 ), .A2(
        \SB2_3_28/i1[9] ), .ZN(\SB2_3_28/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_28/Component_Function_5/N1  ( .A1(\SB2_3_28/i0_0 ), .A2(
        \SB2_3_28/i3[0] ), .ZN(\SB2_3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_29/Component_Function_0/N4  ( .A1(\SB2_3_29/i0[7] ), .A2(
        \SB2_3_29/i0_3 ), .A3(\SB2_3_29/i0_0 ), .ZN(
        \SB2_3_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_29/Component_Function_0/N3  ( .A1(\SB2_3_29/i0[10] ), .A2(
        \SB2_3_29/i0_4 ), .A3(\SB2_3_29/i0_3 ), .ZN(
        \SB2_3_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_29/Component_Function_0/N2  ( .A1(\SB2_3_29/i0[8] ), .A2(
        \SB2_3_29/i0[7] ), .A3(n2115), .ZN(
        \SB2_3_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_29/Component_Function_0/N1  ( .A1(\SB2_3_29/i0[10] ), .A2(
        \SB2_3_29/i0[9] ), .ZN(\SB2_3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_29/Component_Function_1/N4  ( .A1(\SB2_3_29/i1_7 ), .A2(
        \SB2_3_29/i0[8] ), .A3(\SB2_3_29/i0_4 ), .ZN(
        \SB2_3_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_29/Component_Function_1/N3  ( .A1(\SB2_3_29/i1_5 ), .A2(
        n2115), .A3(\SB2_3_29/i0[9] ), .ZN(
        \SB2_3_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_29/Component_Function_1/N2  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i1_7 ), .A3(\SB2_3_29/i0[8] ), .ZN(
        \SB2_3_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_29/Component_Function_1/N1  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_29/Component_Function_5/N1  ( .A1(\SB2_3_29/i0_0 ), .A2(
        \SB2_3_29/i3[0] ), .ZN(\SB2_3_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_0/N4  ( .A1(\SB2_3_30/i0[7] ), .A2(
        \SB2_3_30/i0_3 ), .A3(\SB2_3_30/i0_0 ), .ZN(
        \SB2_3_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_30/Component_Function_0/N3  ( .A1(\SB2_3_30/i0[10] ), .A2(
        \SB2_3_30/i0_4 ), .A3(\SB2_3_30/i0_3 ), .ZN(
        \SB2_3_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_30/Component_Function_0/N2  ( .A1(\SB2_3_30/i0[8] ), .A2(
        \SB2_3_30/i0[7] ), .A3(\SB2_3_30/i0[6] ), .ZN(
        \SB2_3_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_30/Component_Function_0/N1  ( .A1(\SB2_3_30/i0[10] ), .A2(
        \SB2_3_30/i0[9] ), .ZN(\SB2_3_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_1/N4  ( .A1(\SB2_3_30/i1_7 ), .A2(
        \SB2_3_30/i0[8] ), .A3(\SB2_3_30/i0_4 ), .ZN(
        \SB2_3_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_30/Component_Function_1/N3  ( .A1(\SB2_3_30/i1_5 ), .A2(
        \SB2_3_30/i0[6] ), .A3(\SB2_3_30/i0[9] ), .ZN(
        \SB2_3_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_30/Component_Function_1/N2  ( .A1(\SB2_3_30/i0_3 ), .A2(
        \SB2_3_30/i1_7 ), .A3(\SB2_3_30/i0[8] ), .ZN(
        \SB2_3_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_30/Component_Function_1/N1  ( .A1(\SB2_3_30/i0_3 ), .A2(
        \SB2_3_30/i1[9] ), .ZN(\SB2_3_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_5/N2  ( .A1(\SB2_3_30/i0_0 ), .A2(
        \SB2_3_30/i0[6] ), .A3(\SB2_3_30/i0[10] ), .ZN(
        \SB2_3_30/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_30/Component_Function_5/N1  ( .A1(\SB2_3_30/i0_0 ), .A2(
        \SB2_3_30/i3[0] ), .ZN(\SB2_3_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_0/N4  ( .A1(n1513), .A2(
        \SB2_3_31/i0_3 ), .A3(\SB2_3_31/i0_0 ), .ZN(
        \SB2_3_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_31/Component_Function_0/N3  ( .A1(\SB2_3_31/i0[10] ), .A2(
        n1651), .A3(\SB2_3_31/i0_3 ), .ZN(
        \SB2_3_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_31/Component_Function_0/N2  ( .A1(\SB2_3_31/i0[8] ), .A2(
        n1513), .A3(\SB2_3_31/i0[6] ), .ZN(
        \SB2_3_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_31/Component_Function_0/N1  ( .A1(\SB2_3_31/i0[10] ), .A2(
        \SB2_3_31/i0[9] ), .ZN(\SB2_3_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_1/N4  ( .A1(\SB2_3_31/i1_7 ), .A2(
        \SB2_3_31/i0[8] ), .A3(n1652), .ZN(
        \SB2_3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_31/Component_Function_1/N3  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0[6] ), .A3(\SB2_3_31/i0[9] ), .ZN(
        \SB2_3_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_31/Component_Function_1/N2  ( .A1(\SB2_3_31/i0_3 ), .A2(
        \SB2_3_31/i1_7 ), .A3(\SB2_3_31/i0[8] ), .ZN(
        \SB2_3_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_31/Component_Function_1/N1  ( .A1(\SB2_3_31/i0_3 ), .A2(
        n1662), .ZN(\SB2_3_31/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_31/Component_Function_5/N1  ( .A1(\SB2_3_31/i0_0 ), .A2(
        \SB2_3_31/i3[0] ), .ZN(\SB2_3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_0/N4  ( .A1(\SB3_0/i0[7] ), .A2(
        \SB3_0/i0_3 ), .A3(\SB3_0/i0_0 ), .ZN(
        \SB3_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_0/Component_Function_0/N3  ( .A1(\SB3_0/i0[10] ), .A2(
        \SB3_0/i0_4 ), .A3(\SB3_0/i0_3 ), .ZN(
        \SB3_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_0/Component_Function_0/N2  ( .A1(\SB3_0/i0[8] ), .A2(
        \SB3_0/i0[7] ), .A3(\SB3_0/i0[6] ), .ZN(
        \SB3_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_0/Component_Function_0/N1  ( .A1(\SB3_0/i0[10] ), .A2(
        \SB3_0/i0[9] ), .ZN(\SB3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_1/N4  ( .A1(\SB3_0/i1_7 ), .A2(
        \SB3_0/i0[8] ), .A3(\SB3_0/i0_4 ), .ZN(
        \SB3_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_0/Component_Function_1/N3  ( .A1(\SB3_0/i1_5 ), .A2(
        \SB3_0/i0[6] ), .A3(\SB3_0/i0[9] ), .ZN(
        \SB3_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_0/Component_Function_1/N2  ( .A1(\SB3_0/i0_3 ), .A2(
        \SB3_0/i1_7 ), .A3(\SB3_0/i0[8] ), .ZN(
        \SB3_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_0/Component_Function_1/N1  ( .A1(\SB3_0/i0_3 ), .A2(
        \SB3_0/i1[9] ), .ZN(\SB3_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_5/N4  ( .A1(\SB3_0/i0[9] ), .A2(
        \SB3_0/i0[6] ), .A3(\SB3_0/i0_4 ), .ZN(
        \SB3_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_0/Component_Function_5/N2  ( .A1(\SB3_0/i0_0 ), .A2(
        \SB3_0/i0[6] ), .A3(\SB3_0/i0[10] ), .ZN(
        \SB3_0/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_0/Component_Function_5/N1  ( .A1(\SB3_0/i0_0 ), .A2(
        \SB3_0/i3[0] ), .ZN(\SB3_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_0/N3  ( .A1(\SB3_1/i0[10] ), .A2(
        \SB3_1/i0_4 ), .A3(\SB3_1/i0_3 ), .ZN(
        \SB3_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_1/Component_Function_0/N2  ( .A1(\SB3_1/i0[8] ), .A2(
        \SB3_1/i0[7] ), .A3(\SB3_1/i0[6] ), .ZN(
        \SB3_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_1/Component_Function_0/N1  ( .A1(\SB3_1/i0[10] ), .A2(
        \SB3_1/i0[9] ), .ZN(\SB3_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_1/N4  ( .A1(\SB3_1/i1_7 ), .A2(
        \SB3_1/i0[8] ), .A3(\SB3_1/i0_4 ), .ZN(
        \SB3_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_1/Component_Function_1/N3  ( .A1(\SB3_1/i1_5 ), .A2(
        \SB3_1/i0[6] ), .A3(\SB3_1/i0[9] ), .ZN(
        \SB3_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_1/Component_Function_1/N2  ( .A1(n856), .A2(\SB3_1/i1_7 ), 
        .A3(\SB3_1/i0[8] ), .ZN(\SB3_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_1/Component_Function_1/N1  ( .A1(n856), .A2(\SB3_1/i1[9] ), 
        .ZN(\SB3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_5/N4  ( .A1(\SB3_1/i0[9] ), .A2(
        \SB3_1/i0_4 ), .A3(\SB3_1/i0[6] ), .ZN(
        \SB3_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_1/Component_Function_5/N2  ( .A1(\SB3_1/i0_0 ), .A2(
        \SB3_1/i0[6] ), .A3(\SB3_1/i0[10] ), .ZN(
        \SB3_1/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_1/Component_Function_5/N1  ( .A1(\SB3_1/i0_0 ), .A2(
        \SB3_1/i3[0] ), .ZN(\SB3_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_0/N2  ( .A1(\SB3_2/i0[8] ), .A2(
        \SB3_2/i0[7] ), .A3(\SB3_2/i0[6] ), .ZN(
        \SB3_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_2/Component_Function_0/N1  ( .A1(\SB3_2/i0[10] ), .A2(
        \SB3_2/i0[9] ), .ZN(\SB3_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_1/N3  ( .A1(\SB3_2/i1_5 ), .A2(
        \SB3_2/i0[6] ), .A3(\SB3_2/i0[9] ), .ZN(
        \SB3_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_2/Component_Function_1/N2  ( .A1(\SB3_2/i0_3 ), .A2(
        \SB3_2/i1_7 ), .A3(\SB3_2/i0[8] ), .ZN(
        \SB3_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_2/Component_Function_1/N1  ( .A1(\SB3_2/i0_3 ), .A2(
        \SB3_2/i1[9] ), .ZN(\SB3_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_5/N2  ( .A1(\SB3_2/i0_0 ), .A2(
        \SB3_2/i0[6] ), .A3(\SB3_2/i0[10] ), .ZN(
        \SB3_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_2/Component_Function_5/N1  ( .A1(\SB3_2/i0_0 ), .A2(
        \SB3_2/i3[0] ), .ZN(\SB3_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_0/N4  ( .A1(\SB3_3/i0[7] ), .A2(
        \SB3_3/i0_3 ), .A3(\SB3_3/i0_0 ), .ZN(
        \SB3_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_3/Component_Function_0/N2  ( .A1(\SB3_3/i0[8] ), .A2(
        \SB3_3/i0[7] ), .A3(\SB3_3/i0[6] ), .ZN(
        \SB3_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_3/Component_Function_0/N1  ( .A1(\SB3_3/i0[10] ), .A2(
        \SB3_3/i0[9] ), .ZN(\SB3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_1/N4  ( .A1(\SB3_3/i1_7 ), .A2(
        \SB3_3/i0[8] ), .A3(\SB3_3/i0_4 ), .ZN(
        \SB3_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_3/Component_Function_1/N3  ( .A1(\SB3_3/i1_5 ), .A2(
        \SB3_3/i0[6] ), .A3(\SB3_3/i0[9] ), .ZN(
        \SB3_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_3/Component_Function_1/N2  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i1_7 ), .A3(\SB3_3/i0[8] ), .ZN(
        \SB3_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_3/Component_Function_1/N1  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i1[9] ), .ZN(\SB3_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_5/N4  ( .A1(\SB3_3/i0[9] ), .A2(
        \SB3_3/i0[6] ), .A3(\SB3_3/i0_4 ), .ZN(
        \SB3_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_3/Component_Function_5/N2  ( .A1(\SB3_3/i0_0 ), .A2(
        \SB3_3/i0[6] ), .A3(\SB3_3/i0[10] ), .ZN(
        \SB3_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_3/Component_Function_5/N1  ( .A1(\SB3_3/i0_0 ), .A2(
        \SB3_3/i3[0] ), .ZN(\SB3_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_0/N4  ( .A1(\SB3_4/i0[7] ), .A2(
        \SB3_4/i0_3 ), .A3(\SB3_4/i0_0 ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_0/N3  ( .A1(\SB3_4/i0[10] ), .A2(
        \SB3_4/i0_4 ), .A3(\SB3_4/i0_3 ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_4/Component_Function_0/N2  ( .A1(\SB3_4/i0[8] ), .A2(
        \SB3_4/i0[7] ), .A3(\SB3_4/i0[6] ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_4/Component_Function_0/N1  ( .A1(\SB3_4/i0[10] ), .A2(
        \SB3_4/i0[9] ), .ZN(\SB3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_1/N4  ( .A1(\SB3_4/i1_7 ), .A2(
        \SB3_4/i0[8] ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_1/N3  ( .A1(\SB3_4/i1_5 ), .A2(
        \SB3_4/i0[6] ), .A3(\SB3_4/i0[9] ), .ZN(
        \SB3_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_4/Component_Function_1/N2  ( .A1(\SB3_4/i0_3 ), .A2(
        \SB3_4/i1_7 ), .A3(\SB3_4/i0[8] ), .ZN(
        \SB3_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_4/Component_Function_1/N1  ( .A1(\SB3_4/i0_3 ), .A2(
        \SB3_4/i1[9] ), .ZN(\SB3_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_5/N4  ( .A1(\SB3_4/i0[9] ), .A2(
        \SB3_4/i0[6] ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_5/N2  ( .A1(\SB3_4/i0_0 ), .A2(
        \SB3_4/i0[6] ), .A3(\SB3_4/i0[10] ), .ZN(
        \SB3_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_4/Component_Function_5/N1  ( .A1(\SB3_4/i0_0 ), .A2(
        \SB3_4/i3[0] ), .ZN(\SB3_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_0/N3  ( .A1(\SB3_5/i0[10] ), .A2(
        \SB3_5/i0_4 ), .A3(\SB3_5/i0_3 ), .ZN(
        \SB3_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_5/Component_Function_0/N2  ( .A1(\SB3_5/i0[8] ), .A2(
        \SB3_5/i0[7] ), .A3(\SB3_5/i0[6] ), .ZN(
        \SB3_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_5/Component_Function_0/N1  ( .A1(\SB3_5/i0[10] ), .A2(
        \SB3_5/i0[9] ), .ZN(\SB3_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_1/N4  ( .A1(\SB3_5/i1_7 ), .A2(
        \SB3_5/i0[8] ), .A3(\SB3_5/i0_4 ), .ZN(
        \SB3_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_5/Component_Function_1/N3  ( .A1(\SB3_5/i1_5 ), .A2(
        \SB3_5/i0[6] ), .A3(\SB3_5/i0[9] ), .ZN(
        \SB3_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_5/Component_Function_1/N2  ( .A1(\SB3_5/i0_3 ), .A2(
        \SB3_5/i1_7 ), .A3(\SB3_5/i0[8] ), .ZN(
        \SB3_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_5/Component_Function_1/N1  ( .A1(\SB3_5/i0_3 ), .A2(
        \SB3_5/i1[9] ), .ZN(\SB3_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_5/N4  ( .A1(\SB3_5/i0[9] ), .A2(
        \SB3_5/i0[6] ), .A3(\SB3_5/i0_4 ), .ZN(
        \SB3_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_5/Component_Function_5/N2  ( .A1(\SB3_5/i0_0 ), .A2(
        \SB3_5/i0[6] ), .A3(\SB3_5/i0[10] ), .ZN(
        \SB3_5/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_5/Component_Function_5/N1  ( .A1(\SB3_5/i0_0 ), .A2(
        \SB3_5/i3[0] ), .ZN(\SB3_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_0/N3  ( .A1(\SB3_6/i0[10] ), .A2(
        \SB3_6/i0_4 ), .A3(n833), .ZN(\SB3_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_6/Component_Function_0/N2  ( .A1(\SB3_6/i0[8] ), .A2(
        \SB3_6/i0[7] ), .A3(\SB3_6/i0[6] ), .ZN(
        \SB3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_6/Component_Function_0/N1  ( .A1(\SB3_6/i0[10] ), .A2(
        \SB3_6/i0[9] ), .ZN(\SB3_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_1/N4  ( .A1(\SB3_6/i1_7 ), .A2(
        \SB3_6/i0[8] ), .A3(\SB3_6/i0_4 ), .ZN(
        \SB3_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_1/N3  ( .A1(\SB3_6/i1_5 ), .A2(
        \SB3_6/i0[6] ), .A3(\SB3_6/i0[9] ), .ZN(
        \SB3_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_6/Component_Function_1/N2  ( .A1(\SB3_6/i0_3 ), .A2(
        \SB3_6/i1_7 ), .A3(\SB3_6/i0[8] ), .ZN(
        \SB3_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_6/Component_Function_1/N1  ( .A1(\SB3_6/i0_3 ), .A2(
        \SB3_6/i1[9] ), .ZN(\SB3_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_5/N4  ( .A1(\SB3_6/i0[9] ), .A2(
        \SB3_6/i0[6] ), .A3(\SB3_6/i0_4 ), .ZN(
        \SB3_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_5/N3  ( .A1(n833), .A2(\SB3_6/i0_4 ), 
        .A3(\SB3_6/i1[9] ), .ZN(\SB3_6/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB3_6/Component_Function_5/N1  ( .A1(\SB3_6/i0_0 ), .A2(
        \SB3_6/i3[0] ), .ZN(\SB3_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_0/N3  ( .A1(\SB3_7/i0[10] ), .A2(
        \SB3_7/i0_4 ), .A3(\SB3_7/i0_3 ), .ZN(
        \SB3_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_7/Component_Function_0/N2  ( .A1(n798), .A2(\SB3_7/i0[7] ), 
        .A3(\SB3_7/i0[6] ), .ZN(\SB3_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_7/Component_Function_0/N1  ( .A1(\SB3_7/i0[10] ), .A2(
        \SB3_7/i0[9] ), .ZN(\SB3_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_1/N4  ( .A1(\SB3_7/i1_7 ), .A2(n798), 
        .A3(\SB3_7/i0_4 ), .ZN(\SB3_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_7/Component_Function_1/N3  ( .A1(\SB3_7/i1_5 ), .A2(
        \SB3_7/i0[6] ), .A3(\SB3_7/i0[9] ), .ZN(
        \SB3_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_7/Component_Function_1/N2  ( .A1(\SB3_7/i0_3 ), .A2(
        \SB3_7/i1_7 ), .A3(n798), .ZN(\SB3_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_7/Component_Function_1/N1  ( .A1(\SB3_7/i0_3 ), .A2(
        \SB3_7/i1[9] ), .ZN(\SB3_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_5/N4  ( .A1(\SB3_7/i0[9] ), .A2(
        \SB3_7/i0[6] ), .A3(\SB3_7/i0_4 ), .ZN(
        \SB3_7/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB3_7/Component_Function_5/N1  ( .A1(\SB3_7/i0_0 ), .A2(
        \SB3_7/i3[0] ), .ZN(\SB3_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_0/N4  ( .A1(\SB3_8/i0[7] ), .A2(
        \SB3_8/i0_3 ), .A3(\SB3_8/i0_0 ), .ZN(
        \SB3_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_0/N2  ( .A1(\SB3_8/i0[8] ), .A2(
        \SB3_8/i0[7] ), .A3(\SB3_8/i0[6] ), .ZN(
        \SB3_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_8/Component_Function_0/N1  ( .A1(\SB3_8/i0[10] ), .A2(
        \SB3_8/i0[9] ), .ZN(\SB3_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_1/N4  ( .A1(\SB3_8/i1_7 ), .A2(
        \SB3_8/i0[8] ), .A3(\SB3_8/i0_4 ), .ZN(
        \SB3_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_1/N3  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[6] ), .A3(\SB3_8/i0[9] ), .ZN(
        \SB3_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_8/Component_Function_1/N2  ( .A1(\SB3_8/i0_3 ), .A2(
        \SB3_8/i1_7 ), .A3(\SB3_8/i0[8] ), .ZN(
        \SB3_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_8/Component_Function_1/N1  ( .A1(\SB3_8/i0_3 ), .A2(
        \SB3_8/i1[9] ), .ZN(\SB3_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_5/N4  ( .A1(\SB3_8/i0[9] ), .A2(
        \SB3_8/i0[6] ), .A3(\SB3_8/i0_4 ), .ZN(
        \SB3_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_5/N2  ( .A1(\SB3_8/i0_0 ), .A2(
        \SB3_8/i0[6] ), .A3(\SB3_8/i0[10] ), .ZN(
        \SB3_8/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_8/Component_Function_5/N1  ( .A1(\SB3_8/i0_0 ), .A2(
        \SB3_8/i3[0] ), .ZN(\SB3_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_0/N4  ( .A1(\SB3_9/i0[7] ), .A2(
        \SB3_9/i0_3 ), .A3(\SB3_9/i0_0 ), .ZN(
        \SB3_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_0/N3  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i0_4 ), .A3(\SB3_9/i0[10] ), .ZN(
        \SB3_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_9/Component_Function_0/N2  ( .A1(\SB3_9/i0[8] ), .A2(
        \SB3_9/i0[7] ), .A3(\SB3_9/i0[6] ), .ZN(
        \SB3_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_9/Component_Function_0/N1  ( .A1(\SB3_9/i0[10] ), .A2(
        \SB3_9/i0[9] ), .ZN(\SB3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_1/N4  ( .A1(\SB3_9/i1_7 ), .A2(
        \SB3_9/i0[8] ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_1/N3  ( .A1(\SB3_9/i1_5 ), .A2(
        \SB3_9/i0[6] ), .A3(\SB3_9/i0[9] ), .ZN(
        \SB3_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_9/Component_Function_1/N2  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i1_7 ), .A3(\SB3_9/i0[8] ), .ZN(
        \SB3_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_9/Component_Function_1/N1  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i1[9] ), .ZN(\SB3_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_5/N4  ( .A1(\SB3_9/i0[9] ), .A2(
        \SB3_9/i0[6] ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_5/N2  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i0[6] ), .A3(\SB3_9/i0[10] ), .ZN(
        \SB3_9/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_9/Component_Function_5/N1  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i3[0] ), .ZN(\SB3_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_0/N3  ( .A1(\SB3_10/i0[10] ), .A2(
        \SB3_10/i0_4 ), .A3(n835), .ZN(
        \SB3_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_10/Component_Function_0/N2  ( .A1(\SB3_10/i0[8] ), .A2(
        \SB3_10/i0[7] ), .A3(\SB3_10/i0[6] ), .ZN(
        \SB3_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_10/Component_Function_0/N1  ( .A1(\SB3_10/i0[10] ), .A2(
        \SB3_10/i0[9] ), .ZN(\SB3_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_1/N4  ( .A1(\SB3_10/i1_7 ), .A2(
        \SB3_10/i0[8] ), .A3(\SB3_10/i0_4 ), .ZN(
        \SB3_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_10/Component_Function_1/N3  ( .A1(\SB3_10/i1_5 ), .A2(
        \SB3_10/i0[6] ), .A3(\SB3_10/i0[9] ), .ZN(
        \SB3_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_10/Component_Function_1/N2  ( .A1(n835), .A2(\SB3_10/i1_7 ), 
        .A3(\SB3_10/i0[8] ), .ZN(\SB3_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_10/Component_Function_1/N1  ( .A1(n835), .A2(\SB3_10/i1[9] ), 
        .ZN(\SB3_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_5/N4  ( .A1(\SB3_10/i0[9] ), .A2(
        \SB3_10/i0[6] ), .A3(\SB3_10/i0_4 ), .ZN(
        \SB3_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_10/Component_Function_5/N2  ( .A1(\SB3_10/i0_0 ), .A2(
        \SB3_10/i0[6] ), .A3(\SB3_10/i0[10] ), .ZN(
        \SB3_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_10/Component_Function_5/N1  ( .A1(\SB3_10/i0_0 ), .A2(
        \SB3_10/i3[0] ), .ZN(\SB3_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_0/N3  ( .A1(\SB3_11/i0[10] ), .A2(
        \SB3_11/i0_4 ), .A3(\SB3_11/i0_3 ), .ZN(
        \SB3_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_11/Component_Function_0/N2  ( .A1(\SB3_11/i0[8] ), .A2(
        \SB3_11/i0[7] ), .A3(\SB3_11/i0[6] ), .ZN(
        \SB3_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_11/Component_Function_0/N1  ( .A1(\SB3_11/i0[10] ), .A2(
        \SB3_11/i0[9] ), .ZN(\SB3_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_1/N2  ( .A1(\SB3_11/i0_3 ), .A2(
        \SB3_11/i1_7 ), .A3(\SB3_11/i0[8] ), .ZN(
        \SB3_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_11/Component_Function_1/N1  ( .A1(n840), .A2(\SB3_11/i1[9] ), 
        .ZN(\SB3_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_5/N2  ( .A1(\SB3_11/i0_0 ), .A2(
        \SB3_11/i0[6] ), .A3(\SB3_11/i0[10] ), .ZN(
        \SB3_11/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_11/Component_Function_5/N1  ( .A1(\SB3_11/i0_0 ), .A2(
        \SB3_11/i3[0] ), .ZN(\SB3_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_0/N2  ( .A1(\SB3_12/i0[8] ), .A2(
        \SB3_12/i0[7] ), .A3(\SB3_12/i0[6] ), .ZN(
        \SB3_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_12/Component_Function_0/N1  ( .A1(\SB3_12/i0[10] ), .A2(
        \SB3_12/i0[9] ), .ZN(\SB3_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_1/N4  ( .A1(\SB3_12/i1_7 ), .A2(
        \SB3_12/i0[8] ), .A3(\SB3_12/i0_4 ), .ZN(
        \SB3_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_12/Component_Function_1/N3  ( .A1(\SB3_12/i1_5 ), .A2(
        \SB3_12/i0[6] ), .A3(\SB3_12/i0[9] ), .ZN(
        \SB3_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_12/Component_Function_1/N2  ( .A1(\SB3_12/i0_3 ), .A2(
        \SB3_12/i1_7 ), .A3(\SB3_12/i0[8] ), .ZN(
        \SB3_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_12/Component_Function_1/N1  ( .A1(\SB3_12/i0_3 ), .A2(
        \SB3_12/i1[9] ), .ZN(\SB3_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_5/N4  ( .A1(\SB3_12/i0[9] ), .A2(
        \SB3_12/i0[6] ), .A3(\SB3_12/i0_4 ), .ZN(
        \SB3_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_12/Component_Function_5/N2  ( .A1(\SB3_12/i0_0 ), .A2(
        \SB3_12/i0[6] ), .A3(\SB3_12/i0[10] ), .ZN(
        \SB3_12/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_12/Component_Function_5/N1  ( .A1(\SB3_12/i0_0 ), .A2(
        \SB3_12/i3[0] ), .ZN(\SB3_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_0/N4  ( .A1(\SB3_13/i0[7] ), .A2(
        \SB3_13/i0_3 ), .A3(\SB3_13/i0_0 ), .ZN(
        \SB3_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_0/N3  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i0_4 ), .A3(\SB3_13/i0[10] ), .ZN(
        \SB3_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_13/Component_Function_0/N2  ( .A1(\SB3_13/i0[8] ), .A2(
        \SB3_13/i0[7] ), .A3(\SB3_13/i0[6] ), .ZN(
        \SB3_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_13/Component_Function_0/N1  ( .A1(\SB3_13/i0[10] ), .A2(
        \SB3_13/i0[9] ), .ZN(\SB3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_1/N4  ( .A1(\SB3_13/i1_7 ), .A2(
        \SB3_13/i0[8] ), .A3(\SB3_13/i0_4 ), .ZN(
        \SB3_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_1/N3  ( .A1(\SB3_13/i1_5 ), .A2(
        \SB3_13/i0[6] ), .A3(\SB3_13/i0[9] ), .ZN(
        \SB3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_13/Component_Function_1/N2  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i1_7 ), .A3(\SB3_13/i0[8] ), .ZN(
        \SB3_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_13/Component_Function_1/N1  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i1[9] ), .ZN(\SB3_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_5/N4  ( .A1(\SB3_13/i0[9] ), .A2(
        \SB3_13/i0[6] ), .A3(\SB3_13/i0_4 ), .ZN(
        \SB3_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_5/N2  ( .A1(\SB3_13/i0_0 ), .A2(
        \SB3_13/i0[6] ), .A3(\SB3_13/i0[10] ), .ZN(
        \SB3_13/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_13/Component_Function_5/N1  ( .A1(\SB3_13/i0_0 ), .A2(
        \SB3_13/i3[0] ), .ZN(\SB3_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_0/N3  ( .A1(\SB3_14/i0[10] ), .A2(
        \SB3_14/i0_4 ), .A3(\SB3_14/i0_3 ), .ZN(
        \SB3_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_0/N2  ( .A1(\SB3_14/i0[8] ), .A2(
        \SB3_14/i0[7] ), .A3(\SB3_14/i0[6] ), .ZN(
        \SB3_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_14/Component_Function_0/N1  ( .A1(\SB3_14/i0[10] ), .A2(
        \SB3_14/i0[9] ), .ZN(\SB3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_1/N4  ( .A1(\SB3_14/i1_7 ), .A2(
        \SB3_14/i0[8] ), .A3(\SB3_14/i0_4 ), .ZN(
        \SB3_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_14/Component_Function_1/N3  ( .A1(\SB3_14/i1_5 ), .A2(
        \SB3_14/i0[6] ), .A3(\SB3_14/i0[9] ), .ZN(
        \SB3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_1/N2  ( .A1(n860), .A2(\SB3_14/i1_7 ), 
        .A3(\SB3_14/i0[8] ), .ZN(\SB3_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_14/Component_Function_1/N1  ( .A1(n860), .A2(\SB3_14/i1[9] ), 
        .ZN(\SB3_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_5/N4  ( .A1(\SB3_14/i0[9] ), .A2(
        \SB3_14/i0[6] ), .A3(\SB3_14/i0_4 ), .ZN(
        \SB3_14/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB3_14/Component_Function_5/N1  ( .A1(\SB3_14/i0_0 ), .A2(
        \SB3_14/i3[0] ), .ZN(\SB3_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_15/Component_Function_0/N3  ( .A1(\SB3_15/i0[10] ), .A2(
        \SB3_15/i0_4 ), .A3(\SB3_15/i0_3 ), .ZN(
        \SB3_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_0/N2  ( .A1(\SB3_15/i0[8] ), .A2(
        \SB3_15/i0[7] ), .A3(\SB3_15/i0[6] ), .ZN(
        \SB3_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_15/Component_Function_0/N1  ( .A1(\SB3_15/i0[10] ), .A2(
        \SB3_15/i0[9] ), .ZN(\SB3_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_15/Component_Function_1/N4  ( .A1(\SB3_15/i1_7 ), .A2(
        \SB3_15/i0[8] ), .A3(\SB3_15/i0_4 ), .ZN(
        \SB3_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_15/Component_Function_1/N3  ( .A1(\SB3_15/i1_5 ), .A2(
        \SB3_15/i0[6] ), .A3(\SB3_15/i0[9] ), .ZN(
        \SB3_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_1/N2  ( .A1(\SB3_15/i0_3 ), .A2(
        \SB3_15/i1_7 ), .A3(\SB3_15/i0[8] ), .ZN(
        \SB3_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_15/Component_Function_1/N1  ( .A1(\SB3_15/i0_3 ), .A2(
        \SB3_15/i1[9] ), .ZN(\SB3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_15/Component_Function_5/N4  ( .A1(\SB3_15/i0[9] ), .A2(
        \SB3_15/i0[6] ), .A3(\SB3_15/i0_4 ), .ZN(
        \SB3_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_15/Component_Function_5/N2  ( .A1(\SB3_15/i0_0 ), .A2(
        \SB3_15/i0[6] ), .A3(\SB3_15/i0[10] ), .ZN(
        \SB3_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_15/Component_Function_5/N1  ( .A1(\SB3_15/i0_0 ), .A2(
        \SB3_15/i3[0] ), .ZN(\SB3_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_0/N4  ( .A1(\SB3_16/i0[7] ), .A2(n876), 
        .A3(\SB3_16/i0_0 ), .ZN(\SB3_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_16/Component_Function_0/N3  ( .A1(\SB3_16/i0[10] ), .A2(
        \SB3_16/i0_4 ), .A3(\SB3_16/i0_3 ), .ZN(
        \SB3_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_16/Component_Function_0/N2  ( .A1(\SB3_16/i0[8] ), .A2(
        \SB3_16/i0[7] ), .A3(\SB3_16/i0[6] ), .ZN(
        \SB3_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_16/Component_Function_0/N1  ( .A1(\SB3_16/i0[10] ), .A2(
        \SB3_16/i0[9] ), .ZN(\SB3_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_1/N4  ( .A1(\SB3_16/i1_7 ), .A2(
        \SB3_16/i0[8] ), .A3(\SB3_16/i0_4 ), .ZN(
        \SB3_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_16/Component_Function_1/N3  ( .A1(\SB3_16/i1_5 ), .A2(
        \SB3_16/i0[6] ), .A3(\SB3_16/i0[9] ), .ZN(
        \SB3_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_16/Component_Function_1/N2  ( .A1(n876), .A2(\SB3_16/i1_7 ), 
        .A3(\SB3_16/i0[8] ), .ZN(\SB3_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_16/Component_Function_1/N1  ( .A1(n876), .A2(\SB3_16/i1[9] ), 
        .ZN(\SB3_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_5/N4  ( .A1(\SB3_16/i0[9] ), .A2(
        \SB3_16/i0[6] ), .A3(\SB3_16/i0_4 ), .ZN(
        \SB3_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_16/Component_Function_5/N2  ( .A1(\SB3_16/i0_0 ), .A2(
        \SB3_16/i0[6] ), .A3(\SB3_16/i0[10] ), .ZN(
        \SB3_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_16/Component_Function_5/N1  ( .A1(\SB3_16/i0_0 ), .A2(
        \SB3_16/i3[0] ), .ZN(\SB3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_0/N3  ( .A1(\SB3_17/i0[10] ), .A2(
        \SB3_17/i0_4 ), .A3(n867), .ZN(
        \SB3_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_17/Component_Function_0/N2  ( .A1(\SB3_17/i0[8] ), .A2(
        \SB3_17/i0[7] ), .A3(\SB3_17/i0[6] ), .ZN(
        \SB3_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_17/Component_Function_0/N1  ( .A1(\SB3_17/i0[10] ), .A2(
        \SB3_17/i0[9] ), .ZN(\SB3_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_1/N4  ( .A1(\SB3_17/i1_7 ), .A2(
        \SB3_17/i0[8] ), .A3(\SB3_17/i0_4 ), .ZN(
        \SB3_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_17/Component_Function_1/N3  ( .A1(\SB3_17/i1_5 ), .A2(
        \SB3_17/i0[6] ), .A3(\SB3_17/i0[9] ), .ZN(
        \SB3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_17/Component_Function_1/N2  ( .A1(n867), .A2(\SB3_17/i1_7 ), 
        .A3(\SB3_17/i0[8] ), .ZN(\SB3_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_17/Component_Function_1/N1  ( .A1(n867), .A2(\SB3_17/i1[9] ), 
        .ZN(\SB3_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_5/N4  ( .A1(\SB3_17/i0[9] ), .A2(
        \SB3_17/i0[6] ), .A3(\SB3_17/i0_4 ), .ZN(
        \SB3_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_17/Component_Function_5/N2  ( .A1(\SB3_17/i0_0 ), .A2(
        \SB3_17/i0[6] ), .A3(\SB3_17/i0[10] ), .ZN(
        \SB3_17/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_17/Component_Function_5/N1  ( .A1(\SB3_17/i0_0 ), .A2(
        \SB3_17/i3[0] ), .ZN(\SB3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_18/Component_Function_0/N3  ( .A1(\SB3_18/i0[10] ), .A2(
        \SB3_18/i0_4 ), .A3(n869), .ZN(
        \SB3_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_0/N2  ( .A1(\SB3_18/i0[8] ), .A2(
        \SB3_18/i0[7] ), .A3(\SB3_18/i0[6] ), .ZN(
        \SB3_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_18/Component_Function_0/N1  ( .A1(\SB3_18/i0[10] ), .A2(
        \SB3_18/i0[9] ), .ZN(\SB3_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_18/Component_Function_1/N4  ( .A1(\SB3_18/i1_7 ), .A2(
        \SB3_18/i0[8] ), .A3(\SB3_18/i0_4 ), .ZN(
        \SB3_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_18/Component_Function_1/N3  ( .A1(\SB3_18/i1_5 ), .A2(
        \SB3_18/i0[6] ), .A3(\SB3_18/i0[9] ), .ZN(
        \SB3_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_1/N2  ( .A1(\SB3_18/i0_3 ), .A2(
        \SB3_18/i1_7 ), .A3(\SB3_18/i0[8] ), .ZN(
        \SB3_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_18/Component_Function_1/N1  ( .A1(n869), .A2(\SB3_18/i1[9] ), 
        .ZN(\SB3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_18/Component_Function_5/N3  ( .A1(\SB3_18/i1[9] ), .A2(
        \SB3_18/i0_4 ), .A3(\SB3_18/i0_3 ), .ZN(
        \SB3_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_5/N2  ( .A1(\SB3_18/i0[10] ), .A2(
        \SB3_18/i0[6] ), .A3(\SB3_18/i0_0 ), .ZN(
        \SB3_18/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_18/Component_Function_5/N1  ( .A1(\SB3_18/i0_0 ), .A2(
        \SB3_18/i3[0] ), .ZN(\SB3_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_0/N4  ( .A1(\SB3_19/i0[7] ), .A2(
        \SB3_19/i0_3 ), .A3(\SB3_19/i0_0 ), .ZN(
        \SB3_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_19/Component_Function_0/N3  ( .A1(\SB3_19/i0[10] ), .A2(
        \SB3_19/i0_4 ), .A3(\SB3_19/i0_3 ), .ZN(
        \SB3_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_19/Component_Function_0/N2  ( .A1(\SB3_19/i0[8] ), .A2(
        \SB3_19/i0[7] ), .A3(\SB3_19/i0[6] ), .ZN(
        \SB3_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_19/Component_Function_0/N1  ( .A1(\SB3_19/i0[10] ), .A2(
        \SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_1/N4  ( .A1(\SB3_19/i1_7 ), .A2(
        \SB3_19/i0[8] ), .A3(\SB3_19/i0_4 ), .ZN(
        \SB3_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_19/Component_Function_1/N3  ( .A1(\SB3_19/i0[9] ), .A2(
        \SB3_19/i0[6] ), .A3(\SB3_19/i1_5 ), .ZN(
        \SB3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_19/Component_Function_1/N2  ( .A1(\SB3_19/i0_3 ), .A2(
        \SB3_19/i1_7 ), .A3(\SB3_19/i0[8] ), .ZN(
        \SB3_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_19/Component_Function_1/N1  ( .A1(\SB3_19/i0_3 ), .A2(
        \SB3_19/i1[9] ), .ZN(\SB3_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_19/Component_Function_5/N1  ( .A1(\SB3_19/i0_0 ), .A2(
        \SB3_19/i3[0] ), .ZN(\SB3_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_0/N3  ( .A1(\SB3_20/i0[10] ), .A2(
        \SB3_20/i0_4 ), .A3(n864), .ZN(
        \SB3_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_20/Component_Function_0/N2  ( .A1(\SB3_20/i0[8] ), .A2(
        \SB3_20/i0[7] ), .A3(\SB3_20/i0[6] ), .ZN(
        \SB3_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_20/Component_Function_0/N1  ( .A1(\SB3_20/i0[10] ), .A2(
        \SB3_20/i0[9] ), .ZN(\SB3_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_1/N4  ( .A1(\SB3_20/i1_7 ), .A2(
        \SB3_20/i0[8] ), .A3(\SB3_20/i0_4 ), .ZN(
        \SB3_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_20/Component_Function_1/N3  ( .A1(\SB3_20/i1_5 ), .A2(
        \SB3_20/i0[6] ), .A3(\SB3_20/i0[9] ), .ZN(
        \SB3_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_20/Component_Function_1/N2  ( .A1(n864), .A2(\SB3_20/i1_7 ), 
        .A3(\SB3_20/i0[8] ), .ZN(\SB3_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_20/Component_Function_1/N1  ( .A1(n864), .A2(\SB3_20/i1[9] ), 
        .ZN(\SB3_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_5/N4  ( .A1(\SB3_20/i0[9] ), .A2(
        \SB3_20/i0[6] ), .A3(\SB3_20/i0_4 ), .ZN(
        \SB3_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_20/Component_Function_5/N2  ( .A1(\SB3_20/i0_0 ), .A2(
        \SB3_20/i0[6] ), .A3(\SB3_20/i0[10] ), .ZN(
        \SB3_20/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_20/Component_Function_5/N1  ( .A1(\SB3_20/i0_0 ), .A2(
        \SB3_20/i3[0] ), .ZN(\SB3_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_0/N4  ( .A1(\SB3_21/i0[7] ), .A2(n843), 
        .A3(\SB3_21/i0_0 ), .ZN(\SB3_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_21/Component_Function_0/N2  ( .A1(\SB3_21/i0[8] ), .A2(
        \SB3_21/i0[7] ), .A3(\SB3_21/i0[6] ), .ZN(
        \SB3_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_21/Component_Function_0/N1  ( .A1(\SB3_21/i0[10] ), .A2(
        \SB3_21/i0[9] ), .ZN(\SB3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_1/N3  ( .A1(\SB3_21/i1_5 ), .A2(
        \SB3_21/i0[6] ), .A3(\SB3_21/i0[9] ), .ZN(
        \SB3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_21/Component_Function_1/N2  ( .A1(\SB3_21/i0_3 ), .A2(
        \SB3_21/i1_7 ), .A3(\SB3_21/i0[8] ), .ZN(
        \SB3_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_21/Component_Function_1/N1  ( .A1(\SB3_21/i0_3 ), .A2(
        \SB3_21/i1[9] ), .ZN(\SB3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_5/N4  ( .A1(\SB3_21/i0[9] ), .A2(
        \SB3_21/i0[6] ), .A3(\SB3_21/i0_4 ), .ZN(
        \SB3_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_21/Component_Function_5/N2  ( .A1(\SB3_21/i0[6] ), .A2(
        \SB3_21/i0_0 ), .A3(\SB3_21/i0[10] ), .ZN(
        \SB3_21/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_21/Component_Function_5/N1  ( .A1(\SB3_21/i0_0 ), .A2(
        \SB3_21/i3[0] ), .ZN(\SB3_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_0/N3  ( .A1(\SB3_22/i0[10] ), .A2(
        \SB3_22/i0_4 ), .A3(\SB3_22/i0_3 ), .ZN(
        \SB3_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_22/Component_Function_0/N2  ( .A1(\SB3_22/i0[8] ), .A2(
        \SB3_22/i0[7] ), .A3(\SB3_22/i0[6] ), .ZN(
        \SB3_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_22/Component_Function_0/N1  ( .A1(\SB3_22/i0[10] ), .A2(
        \SB3_22/i0[9] ), .ZN(\SB3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_1/N4  ( .A1(\SB3_22/i1_7 ), .A2(
        \SB3_22/i0[8] ), .A3(\SB3_22/i0_4 ), .ZN(
        \SB3_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_22/Component_Function_1/N3  ( .A1(\SB3_22/i1_5 ), .A2(
        \SB3_22/i0[6] ), .A3(\SB3_22/i0[9] ), .ZN(
        \SB3_22/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB3_22/Component_Function_1/N1  ( .A1(\SB3_22/i0_3 ), .A2(
        \SB3_22/i1[9] ), .ZN(\SB3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_5/N4  ( .A1(\SB3_22/i0[9] ), .A2(
        \SB3_22/i0[6] ), .A3(\SB3_22/i0_4 ), .ZN(
        \SB3_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_22/Component_Function_5/N2  ( .A1(\SB3_22/i0_0 ), .A2(
        \SB3_22/i0[6] ), .A3(\SB3_22/i0[10] ), .ZN(
        \SB3_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_22/Component_Function_5/N1  ( .A1(\SB3_22/i0_0 ), .A2(
        \SB3_22/i3[0] ), .ZN(\SB3_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_0/N4  ( .A1(\SB3_23/i0[7] ), .A2(n847), 
        .A3(\SB3_23/i0_0 ), .ZN(\SB3_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_0/N3  ( .A1(\SB3_23/i0[10] ), .A2(
        \SB3_23/i0_4 ), .A3(n847), .ZN(
        \SB3_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_23/Component_Function_0/N2  ( .A1(\SB3_23/i0[8] ), .A2(
        \SB3_23/i0[7] ), .A3(\SB3_23/i0[6] ), .ZN(
        \SB3_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_23/Component_Function_0/N1  ( .A1(\SB3_23/i0[10] ), .A2(
        \SB3_23/i0[9] ), .ZN(\SB3_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_1/N4  ( .A1(\SB3_23/i1_7 ), .A2(
        \SB3_23/i0[8] ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_1/N3  ( .A1(\SB3_23/i1_5 ), .A2(
        \SB3_23/i0[6] ), .A3(\SB3_23/i0[9] ), .ZN(
        \SB3_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_23/Component_Function_1/N2  ( .A1(n847), .A2(\SB3_23/i1_7 ), 
        .A3(\SB3_23/i0[8] ), .ZN(\SB3_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_23/Component_Function_1/N1  ( .A1(n847), .A2(\SB3_23/i1[9] ), 
        .ZN(\SB3_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_5/N4  ( .A1(\SB3_23/i0[9] ), .A2(
        \SB3_23/i0[6] ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_5/N2  ( .A1(\SB3_23/i0_0 ), .A2(
        \SB3_23/i0[6] ), .A3(\SB3_23/i0[10] ), .ZN(
        \SB3_23/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_23/Component_Function_5/N1  ( .A1(\SB3_23/i0_0 ), .A2(
        \SB3_23/i3[0] ), .ZN(\SB3_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_0/N3  ( .A1(\SB3_24/i0[10] ), .A2(
        \SB3_24/i0_4 ), .A3(n872), .ZN(
        \SB3_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_24/Component_Function_0/N2  ( .A1(\SB3_24/i0[8] ), .A2(
        \SB3_24/i0[7] ), .A3(\SB3_24/i0[6] ), .ZN(
        \SB3_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_24/Component_Function_0/N1  ( .A1(\SB3_24/i0[10] ), .A2(
        \SB3_24/i0[9] ), .ZN(\SB3_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_1/N4  ( .A1(\SB3_24/i1_7 ), .A2(
        \SB3_24/i0[8] ), .A3(\SB3_24/i0_4 ), .ZN(
        \SB3_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_24/Component_Function_1/N3  ( .A1(\SB3_24/i1_5 ), .A2(
        \SB3_24/i0[6] ), .A3(\SB3_24/i0[9] ), .ZN(
        \SB3_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_24/Component_Function_1/N2  ( .A1(n872), .A2(\SB3_24/i1_7 ), 
        .A3(\SB3_24/i0[8] ), .ZN(\SB3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_24/Component_Function_1/N1  ( .A1(n872), .A2(\SB3_24/i1[9] ), 
        .ZN(\SB3_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_5/N4  ( .A1(\SB3_24/i0[9] ), .A2(
        \SB3_24/i0[6] ), .A3(\SB3_24/i0_4 ), .ZN(
        \SB3_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_24/Component_Function_5/N2  ( .A1(\SB3_24/i0_0 ), .A2(
        \SB3_24/i0[6] ), .A3(\SB3_24/i0[10] ), .ZN(
        \SB3_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_24/Component_Function_5/N1  ( .A1(\SB3_24/i0_0 ), .A2(
        \SB3_24/i3[0] ), .ZN(\SB3_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_0/N4  ( .A1(\SB3_25/i0[7] ), .A2(
        \SB3_25/i0_3 ), .A3(\SB3_25/i0_0 ), .ZN(
        \SB3_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_25/Component_Function_0/N3  ( .A1(\SB3_25/i0[10] ), .A2(
        \SB3_25/i0_4 ), .A3(\SB3_25/i0_3 ), .ZN(
        \SB3_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_25/Component_Function_0/N2  ( .A1(\SB3_25/i0[8] ), .A2(
        \SB3_25/i0[7] ), .A3(\SB3_25/i0[6] ), .ZN(
        \SB3_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_25/Component_Function_0/N1  ( .A1(\SB3_25/i0[10] ), .A2(
        \SB3_25/i0[9] ), .ZN(\SB3_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_1/N4  ( .A1(\SB3_25/i1_7 ), .A2(
        \SB3_25/i0[8] ), .A3(\SB3_25/i0_4 ), .ZN(
        \SB3_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_25/Component_Function_1/N3  ( .A1(\SB3_25/i1_5 ), .A2(
        \SB3_25/i0[6] ), .A3(\SB3_25/i0[9] ), .ZN(
        \SB3_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_25/Component_Function_1/N2  ( .A1(n845), .A2(\SB3_25/i1_7 ), 
        .A3(\SB3_25/i0[8] ), .ZN(\SB3_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_25/Component_Function_1/N1  ( .A1(n845), .A2(\SB3_25/i1[9] ), 
        .ZN(\SB3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_5/N2  ( .A1(\SB3_25/i0_0 ), .A2(
        \SB3_25/i0[6] ), .A3(\SB3_25/i0[10] ), .ZN(
        \SB3_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_25/Component_Function_5/N1  ( .A1(\SB3_25/i0_0 ), .A2(
        \SB3_25/i3[0] ), .ZN(\SB3_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_0/N3  ( .A1(\SB3_26/i0[10] ), .A2(
        \SB3_26/i0_4 ), .A3(\SB3_26/i0_3 ), .ZN(
        \SB3_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_26/Component_Function_0/N2  ( .A1(\SB3_26/i0[8] ), .A2(
        \SB3_26/i0[7] ), .A3(\SB3_26/i0[6] ), .ZN(
        \SB3_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_26/Component_Function_0/N1  ( .A1(\SB3_26/i0[10] ), .A2(
        \SB3_26/i0[9] ), .ZN(\SB3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_1/N4  ( .A1(\SB3_26/i1_7 ), .A2(
        \SB3_26/i0[8] ), .A3(\SB3_26/i0_4 ), .ZN(
        \SB3_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_26/Component_Function_1/N3  ( .A1(\SB3_26/i1_5 ), .A2(
        \SB3_26/i0[6] ), .A3(\SB3_26/i0[9] ), .ZN(
        \SB3_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_26/Component_Function_1/N2  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i1_7 ), .A3(\SB3_26/i0[8] ), .ZN(
        \SB3_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_26/Component_Function_1/N1  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i1[9] ), .ZN(\SB3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_5/N4  ( .A1(\SB3_26/i0[9] ), .A2(
        \SB3_26/i0[6] ), .A3(\SB3_26/i0_4 ), .ZN(
        \SB3_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_26/Component_Function_5/N2  ( .A1(\SB3_26/i0_0 ), .A2(
        \SB3_26/i0[6] ), .A3(\SB3_26/i0[10] ), .ZN(
        \SB3_26/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_26/Component_Function_5/N1  ( .A1(\SB3_26/i0_0 ), .A2(
        \SB3_26/i3[0] ), .ZN(\SB3_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_0/N3  ( .A1(\SB3_27/i0[10] ), .A2(
        \SB3_27/i0_4 ), .A3(n819), .ZN(
        \SB3_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_27/Component_Function_0/N2  ( .A1(\SB3_27/i0[8] ), .A2(
        \SB3_27/i0[7] ), .A3(\SB3_27/i0[6] ), .ZN(
        \SB3_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_27/Component_Function_0/N1  ( .A1(\SB3_27/i0[10] ), .A2(
        \SB3_27/i0[9] ), .ZN(\SB3_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_1/N4  ( .A1(\SB3_27/i1_7 ), .A2(
        \SB3_27/i0[8] ), .A3(\SB3_27/i0_4 ), .ZN(
        \SB3_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_27/Component_Function_1/N3  ( .A1(\SB3_27/i1_5 ), .A2(
        \SB3_27/i0[6] ), .A3(\SB3_27/i0[9] ), .ZN(
        \SB3_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_27/Component_Function_1/N2  ( .A1(n819), .A2(\SB3_27/i1_7 ), 
        .A3(\SB3_27/i0[8] ), .ZN(\SB3_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_27/Component_Function_1/N1  ( .A1(n819), .A2(\SB3_27/i1[9] ), 
        .ZN(\SB3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_5/N4  ( .A1(\SB3_27/i0[9] ), .A2(
        \SB3_27/i0[6] ), .A3(\SB3_27/i0_4 ), .ZN(
        \SB3_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_27/Component_Function_5/N2  ( .A1(\SB3_27/i0_0 ), .A2(
        \SB3_27/i0[6] ), .A3(\SB3_27/i0[10] ), .ZN(
        \SB3_27/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_27/Component_Function_5/N1  ( .A1(\SB3_27/i0_0 ), .A2(
        \SB3_27/i3[0] ), .ZN(\SB3_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_0/N3  ( .A1(\SB3_28/i0[10] ), .A2(
        \SB3_28/i0_4 ), .A3(\SB3_28/i0_3 ), .ZN(
        \SB3_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_0/N2  ( .A1(\SB3_28/i0[8] ), .A2(
        \SB3_28/i0[7] ), .A3(\SB3_28/i0[6] ), .ZN(
        \SB3_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_28/Component_Function_0/N1  ( .A1(\SB3_28/i0[10] ), .A2(
        \SB3_28/i0[9] ), .ZN(\SB3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_1/N4  ( .A1(\SB3_28/i1_7 ), .A2(
        \SB3_28/i0[8] ), .A3(\SB3_28/i0_4 ), .ZN(
        \SB3_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_28/Component_Function_1/N3  ( .A1(\SB3_28/i1_5 ), .A2(
        \SB3_28/i0[6] ), .A3(\SB3_28/i0[9] ), .ZN(
        \SB3_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_1/N2  ( .A1(n865), .A2(\SB3_28/i1_7 ), 
        .A3(\SB3_28/i0[8] ), .ZN(\SB3_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_28/Component_Function_1/N1  ( .A1(n865), .A2(\SB3_28/i1[9] ), 
        .ZN(\SB3_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_5/N4  ( .A1(\SB3_28/i0[9] ), .A2(
        \SB3_28/i0[6] ), .A3(\SB3_28/i0_4 ), .ZN(
        \SB3_28/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB3_28/Component_Function_5/N1  ( .A1(\SB3_28/i0_0 ), .A2(
        \SB3_28/i3[0] ), .ZN(\SB3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_0/N3  ( .A1(\SB3_29/i0[10] ), .A2(
        \SB3_29/i0_4 ), .A3(\SB3_29/i0_3 ), .ZN(
        \SB3_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_0/N2  ( .A1(\SB3_29/i0[8] ), .A2(
        \SB3_29/i0[7] ), .A3(\SB3_29/i0[6] ), .ZN(
        \SB3_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_29/Component_Function_0/N1  ( .A1(\SB3_29/i0[10] ), .A2(
        \SB3_29/i0[9] ), .ZN(\SB3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N4  ( .A1(\SB3_29/i1_7 ), .A2(
        \SB3_29/i0[8] ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N3  ( .A1(\SB3_29/i1_5 ), .A2(
        \SB3_29/i0[6] ), .A3(\SB3_29/i0[9] ), .ZN(
        \SB3_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N2  ( .A1(n861), .A2(\SB3_29/i1_7 ), 
        .A3(\SB3_29/i0[8] ), .ZN(\SB3_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_29/Component_Function_1/N1  ( .A1(n861), .A2(\SB3_29/i1[9] ), 
        .ZN(\SB3_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_5/N4  ( .A1(\SB3_29/i0[9] ), .A2(
        \SB3_29/i0[6] ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_29/Component_Function_5/N2  ( .A1(\SB3_29/i0_0 ), .A2(
        \SB3_29/i0[6] ), .A3(\SB3_29/i0[10] ), .ZN(
        \SB3_29/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_29/Component_Function_5/N1  ( .A1(\SB3_29/i0_0 ), .A2(
        \SB3_29/i3[0] ), .ZN(\SB3_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_0/N3  ( .A1(\SB3_30/i0[10] ), .A2(
        \SB3_30/i0_4 ), .A3(\SB3_30/i0_3 ), .ZN(
        \SB3_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_30/Component_Function_0/N2  ( .A1(\SB3_30/i0[8] ), .A2(
        \SB3_30/i0[7] ), .A3(\SB3_30/i0[6] ), .ZN(
        \SB3_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_30/Component_Function_0/N1  ( .A1(\SB3_30/i0[10] ), .A2(
        \SB3_30/i0[9] ), .ZN(\SB3_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_1/N4  ( .A1(\SB3_30/i1_7 ), .A2(
        \SB3_30/i0[8] ), .A3(\SB3_30/i0_4 ), .ZN(
        \SB3_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_30/Component_Function_1/N3  ( .A1(\SB3_30/i1_5 ), .A2(
        \SB3_30/i0[6] ), .A3(\SB3_30/i0[9] ), .ZN(
        \SB3_30/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB3_30/Component_Function_1/N1  ( .A1(\SB3_30/i0_3 ), .A2(
        \SB3_30/i1[9] ), .ZN(\SB3_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_5/N4  ( .A1(\SB3_30/i0[9] ), .A2(
        \SB3_30/i0[6] ), .A3(\SB3_30/i0_4 ), .ZN(
        \SB3_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_30/Component_Function_5/N2  ( .A1(\SB3_30/i0_0 ), .A2(
        \SB3_30/i0[6] ), .A3(\SB3_30/i0[10] ), .ZN(
        \SB3_30/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_30/Component_Function_5/N1  ( .A1(\SB3_30/i0_0 ), .A2(
        \SB3_30/i3[0] ), .ZN(\SB3_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_0/N4  ( .A1(\SB3_31/i0[7] ), .A2(n1669), 
        .A3(\SB3_31/i0_0 ), .ZN(\SB3_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_31/Component_Function_0/N3  ( .A1(\SB3_31/i0[10] ), .A2(
        \SB3_31/i0_4 ), .A3(\SB3_31/i0_3 ), .ZN(
        \SB3_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_31/Component_Function_0/N2  ( .A1(\SB3_31/i0[8] ), .A2(
        \SB3_31/i0[7] ), .A3(\SB3_31/i0[6] ), .ZN(
        \SB3_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_31/Component_Function_0/N1  ( .A1(\SB3_31/i0[10] ), .A2(
        \SB3_31/i0[9] ), .ZN(\SB3_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_1/N4  ( .A1(\SB3_31/i1_7 ), .A2(
        \SB3_31/i0[8] ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_31/Component_Function_1/N3  ( .A1(\SB3_31/i1_5 ), .A2(
        \SB3_31/i0[6] ), .A3(\SB3_31/i0[9] ), .ZN(
        \SB3_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_31/Component_Function_1/N2  ( .A1(n1669), .A2(\SB3_31/i1_7 ), 
        .A3(\SB3_31/i0[8] ), .ZN(\SB3_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_31/Component_Function_1/N1  ( .A1(n1669), .A2(\SB3_31/i1[9] ), 
        .ZN(\SB3_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_5/N4  ( .A1(\SB3_31/i0[9] ), .A2(
        \SB3_31/i0[6] ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_31/Component_Function_5/N2  ( .A1(\SB3_31/i0_0 ), .A2(
        \SB3_31/i0[6] ), .A3(\SB3_31/i0[10] ), .ZN(
        \SB3_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_31/Component_Function_5/N1  ( .A1(\SB3_31/i0_0 ), .A2(
        \SB3_31/i3[0] ), .ZN(\SB3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_0/Component_Function_0/N3  ( .A1(\SB4_0/i0[10] ), .A2(
        \SB4_0/i0_4 ), .A3(\SB4_0/i0_3 ), .ZN(
        \SB4_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_0/Component_Function_0/N2  ( .A1(\SB4_0/i0[8] ), .A2(
        \SB4_0/i0[7] ), .A3(\SB4_0/i0[6] ), .ZN(
        \SB4_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_0/Component_Function_0/N1  ( .A1(\SB4_0/i0[10] ), .A2(
        \SB4_0/i0[9] ), .ZN(\SB4_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_0/Component_Function_1/N4  ( .A1(\SB4_0/i1_7 ), .A2(
        \SB4_0/i0[8] ), .A3(\SB4_0/i0_4 ), .ZN(
        \SB4_0/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB4_0/Component_Function_1/N1  ( .A1(\SB4_0/i0_3 ), .A2(
        \SB4_0/i1[9] ), .ZN(\SB4_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_0/Component_Function_5/N4  ( .A1(\SB4_0/i0[9] ), .A2(
        \SB4_0/i0[6] ), .A3(\SB4_0/i0_4 ), .ZN(
        \SB4_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_0/Component_Function_5/N2  ( .A1(\SB4_0/i0_0 ), .A2(
        \SB4_0/i0[6] ), .A3(\SB4_0/i0[10] ), .ZN(
        \SB4_0/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_0/Component_Function_5/N1  ( .A1(\SB4_0/i0_0 ), .A2(
        \SB4_0/i3[0] ), .ZN(\SB4_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_1/Component_Function_0/N3  ( .A1(\SB4_1/i0[10] ), .A2(
        \SB4_1/i0_4 ), .A3(\SB4_1/i0_3 ), .ZN(
        \SB4_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_1/Component_Function_0/N2  ( .A1(\SB4_1/i0[8] ), .A2(
        \SB4_1/i0[7] ), .A3(\SB4_1/i0[6] ), .ZN(
        \SB4_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_1/Component_Function_0/N1  ( .A1(\SB4_1/i0[10] ), .A2(
        \SB4_1/i0[9] ), .ZN(\SB4_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_1/Component_Function_1/N3  ( .A1(\SB4_1/i1_5 ), .A2(
        \SB4_1/i0[6] ), .A3(\SB4_1/i0[9] ), .ZN(
        \SB4_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_1/Component_Function_1/N2  ( .A1(n857), .A2(\SB4_1/i1_7 ), 
        .A3(\SB4_1/i0[8] ), .ZN(\SB4_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_1/Component_Function_1/N1  ( .A1(\SB4_1/i0_3 ), .A2(
        \SB4_1/i1[9] ), .ZN(\SB4_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_1/Component_Function_5/N4  ( .A1(\SB4_1/i0[9] ), .A2(
        \SB4_1/i0[6] ), .A3(\SB4_1/i0_4 ), .ZN(
        \SB4_1/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_1/Component_Function_5/N1  ( .A1(\SB4_1/i0_0 ), .A2(
        \SB4_1/i3[0] ), .ZN(\SB4_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_0/N3  ( .A1(\SB4_2/i0[10] ), .A2(
        \SB4_2/i0_4 ), .A3(\SB4_2/i0_3 ), .ZN(
        \SB4_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_2/Component_Function_0/N2  ( .A1(\SB4_2/i0[8] ), .A2(
        \SB4_2/i0[7] ), .A3(\SB4_2/i0[6] ), .ZN(
        \SB4_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_2/Component_Function_0/N1  ( .A1(\SB4_2/i0[10] ), .A2(n785), 
        .ZN(\SB4_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_1/N3  ( .A1(\SB4_2/i1_5 ), .A2(
        \SB4_2/i0[6] ), .A3(n785), .ZN(
        \SB4_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_2/Component_Function_1/N2  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i1_7 ), .A3(\SB4_2/i0[8] ), .ZN(
        \SB4_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_2/Component_Function_1/N1  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i1[9] ), .ZN(\SB4_2/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB4_2/Component_Function_5/N1  ( .A1(\SB4_2/i0_0 ), .A2(n556), 
        .ZN(\SB4_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_3/Component_Function_0/N3  ( .A1(\SB4_3/i0[10] ), .A2(
        \SB4_3/i0_4 ), .A3(\SB4_3/i0_3 ), .ZN(
        \SB4_3/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB4_3/Component_Function_0/N1  ( .A1(\SB4_3/i0[10] ), .A2(
        \SB4_3/i0[9] ), .ZN(\SB4_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_3/Component_Function_1/N2  ( .A1(n859), .A2(\SB4_3/i1_7 ), 
        .A3(\SB4_3/i0[8] ), .ZN(\SB4_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_3/Component_Function_1/N1  ( .A1(n859), .A2(\SB4_3/i1[9] ), 
        .ZN(\SB4_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_3/Component_Function_5/N4  ( .A1(\SB4_3/i0[9] ), .A2(
        \SB4_3/i0[6] ), .A3(\SB4_3/i0_4 ), .ZN(
        \SB4_3/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_3/Component_Function_5/N1  ( .A1(\SB4_3/i0_0 ), .A2(
        \SB4_3/i3[0] ), .ZN(\SB4_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_4/Component_Function_0/N4  ( .A1(\SB4_4/i0[7] ), .A2(n1667), 
        .A3(\SB4_4/i0_0 ), .ZN(\SB4_4/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB4_4/Component_Function_0/N1  ( .A1(\SB4_4/i0[10] ), .A2(
        \SB4_4/i0[9] ), .ZN(\SB4_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_4/Component_Function_1/N4  ( .A1(\SB4_4/i1_7 ), .A2(
        \SB4_4/i0[8] ), .A3(\SB4_4/i0_4 ), .ZN(
        \SB4_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_4/Component_Function_1/N2  ( .A1(n1667), .A2(\SB4_4/i1_7 ), 
        .A3(\SB4_4/i0[8] ), .ZN(\SB4_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_4/Component_Function_1/N1  ( .A1(\SB4_4/i0_3 ), .A2(
        \SB4_4/i1[9] ), .ZN(\SB4_4/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB4_4/Component_Function_5/N1  ( .A1(\SB4_4/i0_0 ), .A2(
        \SB4_4/i3[0] ), .ZN(\SB4_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_0/N3  ( .A1(\SB4_5/i0[10] ), .A2(n834), 
        .A3(\SB4_5/i0_3 ), .ZN(\SB4_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_5/Component_Function_0/N2  ( .A1(\SB4_5/i0[8] ), .A2(n549), 
        .A3(\RI3[4][157] ), .ZN(\SB4_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_5/Component_Function_0/N1  ( .A1(\SB4_5/i0[10] ), .A2(
        \SB4_5/i0[9] ), .ZN(\SB4_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_1/N3  ( .A1(\SB4_5/i1_5 ), .A2(n810), 
        .A3(\SB4_5/i0[9] ), .ZN(\SB4_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_5/Component_Function_1/N2  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i1_7 ), .A3(\SB4_5/i0[8] ), .ZN(
        \SB4_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_5/Component_Function_1/N1  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i1[9] ), .ZN(\SB4_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_5/N4  ( .A1(\SB4_5/i0[9] ), .A2(n810), 
        .A3(n834), .ZN(\SB4_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_5/Component_Function_5/N2  ( .A1(\SB4_5/i0[10] ), .A2(n810), 
        .A3(\SB4_5/i0_0 ), .ZN(\SB4_5/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_5/Component_Function_5/N1  ( .A1(\SB4_5/i0_0 ), .A2(
        \SB4_5/i3[0] ), .ZN(\SB4_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_6/Component_Function_0/N3  ( .A1(\SB4_6/i0[10] ), .A2(
        \SB4_6/i0_4 ), .A3(n858), .ZN(\SB4_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_6/Component_Function_0/N2  ( .A1(\SB4_6/i0[8] ), .A2(
        \SB4_6/i0[7] ), .A3(\SB4_6/i0[6] ), .ZN(
        \SB4_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_6/Component_Function_0/N1  ( .A1(\SB4_6/i0[10] ), .A2(
        \SB4_6/i0[9] ), .ZN(\SB4_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_6/Component_Function_1/N3  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0[6] ), .A3(\SB4_6/i0[9] ), .ZN(
        \SB4_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB4_6/Component_Function_1/N1  ( .A1(n858), .A2(\SB4_6/i1[9] ), 
        .ZN(\SB4_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_6/Component_Function_5/N4  ( .A1(\SB4_6/i0[9] ), .A2(
        \SB4_6/i0[6] ), .A3(\SB4_6/i0_4 ), .ZN(
        \SB4_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_5/N2  ( .A1(\SB4_6/i0_0 ), .A2(
        \SB4_6/i0[6] ), .A3(\SB4_6/i0[10] ), .ZN(
        \SB4_6/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_6/Component_Function_5/N1  ( .A1(\SB4_6/i0_0 ), .A2(
        \SB4_6/i3[0] ), .ZN(\SB4_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_0/N2  ( .A1(\SB4_7/i0[8] ), .A2(
        \SB4_7/i0[7] ), .A3(\RI3[4][145] ), .ZN(
        \SB4_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_7/Component_Function_0/N1  ( .A1(\SB4_7/i0[10] ), .A2(
        \SB4_7/i0[9] ), .ZN(\SB4_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_1/N2  ( .A1(n877), .A2(\SB4_7/i1_7 ), 
        .A3(\SB4_7/i0[8] ), .ZN(\SB4_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_7/Component_Function_1/N1  ( .A1(\SB4_7/i0_3 ), .A2(
        \SB4_7/i1[9] ), .ZN(\SB4_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_5/N4  ( .A1(\SB4_7/i0[9] ), .A2(
        \SB4_7/i0[6] ), .A3(\SB4_7/i0_4 ), .ZN(
        \SB4_7/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_7/Component_Function_5/N1  ( .A1(\SB4_7/i0_0 ), .A2(
        \SB4_7/i3[0] ), .ZN(\SB4_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_0/N3  ( .A1(\SB4_8/i0[10] ), .A2(n1638), 
        .A3(\SB4_8/i0_3 ), .ZN(\SB4_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_8/Component_Function_0/N2  ( .A1(\SB4_8/i0[8] ), .A2(n1512), 
        .A3(\SB4_8/i0[6] ), .ZN(\SB4_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_8/Component_Function_0/N1  ( .A1(\SB4_8/i0[10] ), .A2(
        \SB4_8/i0[9] ), .ZN(\SB4_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_1/N2  ( .A1(n863), .A2(\SB4_8/i1_7 ), 
        .A3(\SB4_8/i0[8] ), .ZN(\SB4_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_8/Component_Function_1/N1  ( .A1(n863), .A2(\SB4_8/i1[9] ), 
        .ZN(\SB4_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_5/N4  ( .A1(\SB4_8/i0[9] ), .A2(
        \SB4_8/i0[6] ), .A3(n1638), .ZN(
        \SB4_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_8/Component_Function_5/N2  ( .A1(\SB4_8/i0_0 ), .A2(
        \SB4_8/i0[6] ), .A3(\SB4_8/i0[10] ), .ZN(
        \SB4_8/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_8/Component_Function_5/N1  ( .A1(\SB4_8/i0_0 ), .A2(
        \SB4_8/i3[0] ), .ZN(\SB4_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_9/Component_Function_0/N4  ( .A1(n836), .A2(n1663), .A3(
        \SB4_9/i0_0 ), .ZN(\SB4_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_0/N2  ( .A1(\SB4_9/i0[8] ), .A2(n836), 
        .A3(\SB4_9/i0[6] ), .ZN(\SB4_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_9/Component_Function_0/N1  ( .A1(\SB4_9/i0[10] ), .A2(
        \SB4_9/i0[9] ), .ZN(\SB4_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_9/Component_Function_1/N3  ( .A1(\SB4_9/i1_5 ), .A2(
        \SB4_9/i0[6] ), .A3(\SB4_9/i0[9] ), .ZN(
        \SB4_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_9/Component_Function_1/N2  ( .A1(n1663), .A2(\SB4_9/i1_7 ), 
        .A3(\SB4_9/i0[8] ), .ZN(\SB4_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_9/Component_Function_1/N1  ( .A1(\SB4_9/i0_3 ), .A2(
        \SB4_9/i1[9] ), .ZN(\SB4_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_9/Component_Function_5/N4  ( .A1(\SB4_9/i0[9] ), .A2(
        \SB4_9/i0[6] ), .A3(\RI3[4][136] ), .ZN(
        \SB4_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_5/N2  ( .A1(\SB4_9/i0_0 ), .A2(
        \SB4_9/i0[6] ), .A3(\SB4_9/i0[10] ), .ZN(
        \SB4_9/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_9/Component_Function_5/N1  ( .A1(\SB4_9/i0_0 ), .A2(
        \SB4_9/i3[0] ), .ZN(\SB4_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_10/Component_Function_0/N4  ( .A1(\SB4_10/i0[7] ), .A2(
        \SB4_10/i0_3 ), .A3(\SB4_10/i0_0 ), .ZN(
        \SB4_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_10/Component_Function_0/N2  ( .A1(\SB4_10/i0[8] ), .A2(
        \SB4_10/i0[7] ), .A3(\SB4_10/i0[6] ), .ZN(
        \SB4_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_10/Component_Function_0/N1  ( .A1(\SB4_10/i0[10] ), .A2(
        \SB4_10/i0[9] ), .ZN(\SB4_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_10/Component_Function_1/N3  ( .A1(\SB4_10/i1_5 ), .A2(
        \SB4_10/i0[6] ), .A3(\SB4_10/i0[9] ), .ZN(
        \SB4_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_10/Component_Function_1/N2  ( .A1(\SB4_10/i0_3 ), .A2(
        \SB4_10/i1_7 ), .A3(\SB4_10/i0[8] ), .ZN(
        \SB4_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_10/Component_Function_1/N1  ( .A1(\SB4_10/i0_3 ), .A2(
        \SB4_10/i1[9] ), .ZN(\SB4_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_10/Component_Function_5/N4  ( .A1(\SB4_10/i0[9] ), .A2(
        \SB4_10/i0[6] ), .A3(\SB4_10/i0_4 ), .ZN(
        \SB4_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_10/Component_Function_5/N2  ( .A1(\SB4_10/i0_0 ), .A2(
        \SB4_10/i0[6] ), .A3(\SB4_10/i0[10] ), .ZN(
        \SB4_10/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_10/Component_Function_5/N1  ( .A1(\SB4_10/i0_0 ), .A2(
        \SB4_10/i3[0] ), .ZN(\SB4_10/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB4_11/Component_Function_0/N1  ( .A1(\SB4_11/i0[10] ), .A2(
        \SB4_11/i0[9] ), .ZN(\SB4_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_11/Component_Function_1/N3  ( .A1(\SB4_11/i1_5 ), .A2(
        \SB4_11/i0[6] ), .A3(\SB4_11/i0[9] ), .ZN(
        \SB4_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_11/Component_Function_1/N2  ( .A1(\SB4_11/i0_3 ), .A2(
        \SB4_11/i1_7 ), .A3(\SB4_11/i0[8] ), .ZN(
        \SB4_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_11/Component_Function_1/N1  ( .A1(n841), .A2(\SB4_11/i1[9] ), 
        .ZN(\SB4_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_11/Component_Function_5/N2  ( .A1(\SB4_11/i0_0 ), .A2(
        \SB4_11/i0[6] ), .A3(\SB4_11/i0[10] ), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_11/Component_Function_5/N1  ( .A1(\SB4_11/i0_0 ), .A2(
        \SB4_11/i3[0] ), .ZN(\SB4_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_12/Component_Function_0/N2  ( .A1(\SB4_12/i0[8] ), .A2(
        \SB4_12/i0[7] ), .A3(\SB4_12/i0[6] ), .ZN(
        \SB4_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_12/Component_Function_0/N1  ( .A1(\SB4_12/i0[10] ), .A2(
        \SB4_12/i0[9] ), .ZN(\SB4_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_12/Component_Function_1/N3  ( .A1(\SB4_12/i1_5 ), .A2(
        \SB4_12/i0[6] ), .A3(\SB4_12/i0[9] ), .ZN(
        \SB4_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_12/Component_Function_1/N2  ( .A1(\SB4_12/i0_3 ), .A2(
        \SB4_12/i1_7 ), .A3(\SB4_12/i0[8] ), .ZN(
        \SB4_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_12/Component_Function_1/N1  ( .A1(\SB4_12/i0_3 ), .A2(
        \SB4_12/i1[9] ), .ZN(\SB4_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_12/Component_Function_5/N4  ( .A1(\SB4_12/i0[9] ), .A2(
        \SB4_12/i0[6] ), .A3(\SB4_12/i0_4 ), .ZN(
        \SB4_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_12/Component_Function_5/N2  ( .A1(\SB4_12/i0_0 ), .A2(
        \SB4_12/i0[6] ), .A3(\SB4_12/i0[10] ), .ZN(
        \SB4_12/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_12/Component_Function_5/N1  ( .A1(\SB4_12/i0_0 ), .A2(
        \SB4_12/i3[0] ), .ZN(\SB4_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_13/Component_Function_0/N4  ( .A1(\SB4_13/i0[7] ), .A2(n2148), 
        .A3(\SB4_13/i0_0 ), .ZN(\SB4_13/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB4_13/Component_Function_0/N1  ( .A1(\SB4_13/i0[10] ), .A2(
        \SB4_13/i0[9] ), .ZN(\SB4_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_13/Component_Function_1/N4  ( .A1(\SB4_13/i1_7 ), .A2(
        \SB4_13/i0[8] ), .A3(\SB4_13/i0_4 ), .ZN(
        \SB4_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_13/Component_Function_1/N3  ( .A1(\SB4_13/i1_5 ), .A2(
        \SB4_13/i0[6] ), .A3(\SB4_13/i0[9] ), .ZN(
        \SB4_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_13/Component_Function_1/N2  ( .A1(n2148), .A2(\SB4_13/i1_7 ), 
        .A3(\SB4_13/i0[8] ), .ZN(\SB4_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_13/Component_Function_1/N1  ( .A1(\SB4_13/i0_3 ), .A2(
        \SB4_13/i1[9] ), .ZN(\SB4_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_13/Component_Function_5/N2  ( .A1(\SB4_13/i0_0 ), .A2(
        \SB4_13/i0[6] ), .A3(\SB4_13/i0[10] ), .ZN(
        \SB4_13/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_13/Component_Function_5/N1  ( .A1(\SB4_13/i0_0 ), .A2(
        \SB4_13/i3[0] ), .ZN(\SB4_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_0/N4  ( .A1(n553), .A2(\SB4_14/i0_3 ), 
        .A3(\SB4_14/i0_0 ), .ZN(\SB4_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_14/Component_Function_0/N2  ( .A1(\SB4_14/i0[8] ), .A2(n553), 
        .A3(\RI3[4][103] ), .ZN(\SB4_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_14/Component_Function_0/N1  ( .A1(\SB4_14/i0[10] ), .A2(
        \SB4_14/i0[9] ), .ZN(\SB4_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_1/N2  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i1_7 ), .A3(\SB4_14/i0[8] ), .ZN(
        \SB4_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_14/Component_Function_1/N1  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i1[9] ), .ZN(\SB4_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_5/N4  ( .A1(\SB4_14/i0[9] ), .A2(n806), 
        .A3(n799), .ZN(\SB4_14/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_14/Component_Function_5/N1  ( .A1(\SB4_14/i0_0 ), .A2(
        \SB4_14/i3[0] ), .ZN(\SB4_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_15/Component_Function_0/N2  ( .A1(\SB4_15/i0[8] ), .A2(
        \SB4_15/i0[7] ), .A3(\SB4_15/i0[6] ), .ZN(
        \SB4_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_15/Component_Function_0/N1  ( .A1(\SB4_15/i0[10] ), .A2(
        \SB4_15/i0[9] ), .ZN(\SB4_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_15/Component_Function_1/N4  ( .A1(\SB4_15/i1_7 ), .A2(
        \SB4_15/i0[8] ), .A3(\SB4_15/i0_4 ), .ZN(
        \SB4_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_15/Component_Function_1/N2  ( .A1(n871), .A2(\SB4_15/i1_7 ), 
        .A3(\SB4_15/i0[8] ), .ZN(\SB4_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_15/Component_Function_1/N1  ( .A1(\SB4_15/i0_3 ), .A2(
        \SB4_15/i1[9] ), .ZN(\SB4_15/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB4_15/Component_Function_5/N1  ( .A1(\SB4_15/i0_0 ), .A2(
        \SB4_15/i3[0] ), .ZN(\SB4_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_16/Component_Function_0/N3  ( .A1(\SB4_16/i0[10] ), .A2(
        \SB4_16/i0_4 ), .A3(\SB4_16/i0_3 ), .ZN(
        \SB4_16/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB4_16/Component_Function_0/N1  ( .A1(\SB4_16/i0[10] ), .A2(
        \SB4_16/i0[9] ), .ZN(\SB4_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_16/Component_Function_1/N3  ( .A1(\SB4_16/i1_5 ), .A2(
        \SB4_16/i0[6] ), .A3(\SB4_16/i0[9] ), .ZN(
        \SB4_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_16/Component_Function_1/N2  ( .A1(\SB4_16/i0_3 ), .A2(
        \SB4_16/i1_7 ), .A3(\SB4_16/i0[8] ), .ZN(
        \SB4_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_16/Component_Function_1/N1  ( .A1(\SB4_16/i0_3 ), .A2(
        \SB4_16/i1[9] ), .ZN(\SB4_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_16/Component_Function_5/N4  ( .A1(\SB4_16/i0[9] ), .A2(
        \SB4_16/i0[6] ), .A3(\SB4_16/i0_4 ), .ZN(
        \SB4_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_16/Component_Function_5/N2  ( .A1(\SB4_16/i0_0 ), .A2(
        \SB4_16/i0[6] ), .A3(\SB4_16/i0[10] ), .ZN(
        \SB4_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_16/Component_Function_5/N1  ( .A1(\SB4_16/i0_0 ), .A2(
        \SB4_16/i3[0] ), .ZN(\SB4_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_17/Component_Function_0/N4  ( .A1(\SB4_17/i0[7] ), .A2(n868), 
        .A3(\SB4_17/i0_0 ), .ZN(\SB4_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_0/N2  ( .A1(\SB4_17/i0[8] ), .A2(
        \SB4_17/i0[7] ), .A3(\RI3[4][85] ), .ZN(
        \SB4_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_17/Component_Function_0/N1  ( .A1(\SB4_17/i0[10] ), .A2(
        \SB4_17/i0[9] ), .ZN(\SB4_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N4  ( .A1(\SB4_17/i1_7 ), .A2(
        \SB4_17/i0[8] ), .A3(\SB4_17/i0_4 ), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N3  ( .A1(\SB4_17/i1_5 ), .A2(
        \SB4_17/i0[6] ), .A3(\SB4_17/i0[9] ), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N2  ( .A1(n868), .A2(\SB4_17/i1_7 ), 
        .A3(\SB4_17/i0[8] ), .ZN(\SB4_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_17/Component_Function_1/N1  ( .A1(\SB4_17/i0_3 ), .A2(
        \SB4_17/i1[9] ), .ZN(\SB4_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_17/Component_Function_5/N4  ( .A1(\SB4_17/i0[9] ), .A2(
        \SB4_17/i0[6] ), .A3(\SB4_17/i0_4 ), .ZN(
        \SB4_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_5/N2  ( .A1(\SB4_17/i0_0 ), .A2(
        \SB4_17/i0[6] ), .A3(\SB4_17/i0[10] ), .ZN(
        \SB4_17/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_17/Component_Function_5/N1  ( .A1(\SB4_17/i0_0 ), .A2(
        \SB4_17/i3[0] ), .ZN(\SB4_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_0/N3  ( .A1(\SB4_18/i0[10] ), .A2(
        \SB4_18/i0_4 ), .A3(n870), .ZN(
        \SB4_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_0/N2  ( .A1(\SB4_18/i0[8] ), .A2(
        \SB4_18/i0[7] ), .A3(\SB4_18/i0[6] ), .ZN(
        \SB4_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_18/Component_Function_0/N1  ( .A1(\SB4_18/i0[10] ), .A2(
        \SB4_18/i0[9] ), .ZN(\SB4_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_1/N3  ( .A1(\SB4_18/i1_5 ), .A2(
        \SB4_18/i0[6] ), .A3(\SB4_18/i0[9] ), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_1/N2  ( .A1(\SB4_18/i0_3 ), .A2(
        \SB4_18/i1_7 ), .A3(\SB4_18/i0[8] ), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_18/Component_Function_1/N1  ( .A1(\SB4_18/i0_3 ), .A2(n2113), 
        .ZN(\SB4_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_5/N4  ( .A1(\SB4_18/i0[9] ), .A2(
        \SB4_18/i0[6] ), .A3(\SB4_18/i0_4 ), .ZN(
        \SB4_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_18/Component_Function_5/N3  ( .A1(n2113), .A2(\SB4_18/i0_4 ), 
        .A3(n870), .ZN(\SB4_18/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB4_18/Component_Function_5/N1  ( .A1(\SB4_18/i0_0 ), .A2(
        \SB4_18/i3[0] ), .ZN(\SB4_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_0/N4  ( .A1(\SB4_19/i0[7] ), .A2(
        \SB4_19/i0_3 ), .A3(\SB4_19/i0_0 ), .ZN(
        \SB4_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_0/N3  ( .A1(\SB4_19/i0[10] ), .A2(
        \SB4_19/i0_4 ), .A3(\SB4_19/i0_3 ), .ZN(
        \SB4_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_0/N2  ( .A1(\SB4_19/i0[8] ), .A2(
        \SB4_19/i0[7] ), .A3(\SB4_19/i0[6] ), .ZN(
        \SB4_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_19/Component_Function_0/N1  ( .A1(\SB4_19/i0[10] ), .A2(
        \SB4_19/i0[9] ), .ZN(\SB4_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_1/N4  ( .A1(\SB4_19/i1_7 ), .A2(
        \SB4_19/i0[8] ), .A3(\SB4_19/i0_4 ), .ZN(
        \SB4_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_1/N3  ( .A1(\SB4_19/i1_5 ), .A2(
        \SB4_19/i0[6] ), .A3(\SB4_19/i0[9] ), .ZN(
        \SB4_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_1/N2  ( .A1(\SB4_19/i0_3 ), .A2(
        \SB4_19/i1_7 ), .A3(\SB4_19/i0[8] ), .ZN(
        \SB4_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_19/Component_Function_1/N1  ( .A1(\SB4_19/i0_3 ), .A2(
        \SB4_19/i1[9] ), .ZN(\SB4_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_5/N4  ( .A1(\SB4_19/i0[9] ), .A2(
        \SB4_19/i0[6] ), .A3(\SB4_19/i0_4 ), .ZN(
        \SB4_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_5/N3  ( .A1(\SB4_19/i1[9] ), .A2(
        \SB4_19/i0_4 ), .A3(\SB4_19/i0_3 ), .ZN(
        \SB4_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_5/N2  ( .A1(\SB4_19/i0_0 ), .A2(
        \SB4_19/i0[6] ), .A3(\SB4_19/i0[10] ), .ZN(
        \SB4_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_19/Component_Function_5/N1  ( .A1(\SB4_19/i0_0 ), .A2(
        \SB4_19/i3[0] ), .ZN(\SB4_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_20/Component_Function_0/N3  ( .A1(\SB4_20/i0[10] ), .A2(n844), 
        .A3(\SB4_20/i0_3 ), .ZN(\SB4_20/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB4_20/Component_Function_0/N1  ( .A1(\SB4_20/i0[10] ), .A2(
        \SB4_20/i0[9] ), .ZN(\SB4_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_20/Component_Function_1/N4  ( .A1(\SB4_20/i1_7 ), .A2(
        \SB4_20/i0[8] ), .A3(n844), .ZN(
        \SB4_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_1/N2  ( .A1(\SB4_20/i0_3 ), .A2(
        \SB4_20/i1_7 ), .A3(\SB4_20/i0[8] ), .ZN(
        \SB4_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_20/Component_Function_1/N1  ( .A1(\SB4_20/i0_3 ), .A2(
        \SB4_20/i1[9] ), .ZN(\SB4_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_20/Component_Function_5/N4  ( .A1(\SB4_20/i0[9] ), .A2(
        \SB4_20/i0[6] ), .A3(n844), .ZN(
        \SB4_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_5/N2  ( .A1(\SB4_20/i0_0 ), .A2(
        \SB4_20/i0[6] ), .A3(\SB4_20/i0[10] ), .ZN(
        \SB4_20/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_20/Component_Function_5/N1  ( .A1(\SB4_20/i0_0 ), .A2(
        \SB4_20/i3[0] ), .ZN(\SB4_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_0/N4  ( .A1(\SB4_21/i0[7] ), .A2(n854), 
        .A3(\SB4_21/i0_0 ), .ZN(\SB4_21/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB4_21/Component_Function_0/N1  ( .A1(\SB4_21/i0[10] ), .A2(
        \SB4_21/i0[9] ), .ZN(\SB4_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_1/N2  ( .A1(n854), .A2(\SB4_21/i1_7 ), 
        .A3(\SB4_21/i0[8] ), .ZN(\SB4_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_21/Component_Function_1/N1  ( .A1(\SB4_21/i0_3 ), .A2(
        \SB4_21/i1[9] ), .ZN(\SB4_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_5/N2  ( .A1(\SB4_21/i0_0 ), .A2(
        \SB4_21/i0[6] ), .A3(\SB4_21/i0[10] ), .ZN(
        \SB4_21/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_21/Component_Function_5/N1  ( .A1(\SB4_21/i0_0 ), .A2(
        \SB4_21/i3[0] ), .ZN(\SB4_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_22/Component_Function_0/N2  ( .A1(\SB4_22/i0[8] ), .A2(
        \SB4_22/i0[7] ), .A3(\SB4_22/i0[6] ), .ZN(
        \SB4_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_22/Component_Function_0/N1  ( .A1(\SB4_22/i0[10] ), .A2(n779), 
        .ZN(\SB4_22/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB4_22/Component_Function_1/N1  ( .A1(\SB4_22/i0_3 ), .A2(
        \SB4_22/i1[9] ), .ZN(\SB4_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_22/Component_Function_5/N2  ( .A1(\SB4_22/i0_0 ), .A2(
        \SB4_22/i0[6] ), .A3(\SB4_22/i0[10] ), .ZN(
        \SB4_22/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_22/Component_Function_5/N1  ( .A1(\SB4_22/i0_0 ), .A2(n550), 
        .ZN(\SB4_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_23/Component_Function_0/N4  ( .A1(\SB4_23/i0[7] ), .A2(n848), 
        .A3(\SB4_23/i0_0 ), .ZN(\SB4_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_0/N2  ( .A1(\SB4_23/i0[8] ), .A2(
        \SB4_23/i0[7] ), .A3(\SB4_23/i0[6] ), .ZN(
        \SB4_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_23/Component_Function_0/N1  ( .A1(\SB4_23/i0[10] ), .A2(
        \SB4_23/i0[9] ), .ZN(\SB4_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_23/Component_Function_1/N4  ( .A1(\SB4_23/i1_7 ), .A2(
        \SB4_23/i0[8] ), .A3(\SB4_23/i0_4 ), .ZN(
        \SB4_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_1/N3  ( .A1(\SB4_23/i1_5 ), .A2(
        \SB4_23/i0[6] ), .A3(\SB4_23/i0[9] ), .ZN(
        \SB4_23/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB4_23/Component_Function_1/N1  ( .A1(n2100), .A2(\SB4_23/i1[9] ), 
        .ZN(\SB4_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_23/Component_Function_5/N4  ( .A1(\SB4_23/i0[9] ), .A2(
        \SB4_23/i0[6] ), .A3(\SB4_23/i0_4 ), .ZN(
        \SB4_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_5/N2  ( .A1(\SB4_23/i0_0 ), .A2(
        \SB4_23/i0[6] ), .A3(\SB4_23/i0[10] ), .ZN(
        \SB4_23/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_23/Component_Function_5/N1  ( .A1(\SB4_23/i0_0 ), .A2(
        \SB4_23/i3[0] ), .ZN(\SB4_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_0/N3  ( .A1(\SB4_24/i0[10] ), .A2(
        \SB4_24/i0_4 ), .A3(n2135), .ZN(
        \SB4_24/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB4_24/Component_Function_0/N1  ( .A1(\SB4_24/i0[10] ), .A2(
        \SB4_24/i0[9] ), .ZN(\SB4_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_1/N4  ( .A1(\SB4_24/i1_7 ), .A2(
        \SB4_24/i0[8] ), .A3(\SB4_24/i0_4 ), .ZN(
        \SB4_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_1/N2  ( .A1(n2135), .A2(\SB4_24/i1_7 ), 
        .A3(\SB4_24/i0[8] ), .ZN(\SB4_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_24/Component_Function_1/N1  ( .A1(\SB4_24/i0_3 ), .A2(
        \SB4_24/i1[9] ), .ZN(\SB4_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_5/N4  ( .A1(\SB4_24/i0[9] ), .A2(
        \SB4_24/i0[6] ), .A3(\SB4_24/i0_4 ), .ZN(
        \SB4_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_5/N2  ( .A1(\SB4_24/i0_0 ), .A2(
        \SB4_24/i0[6] ), .A3(\SB4_24/i0[10] ), .ZN(
        \SB4_24/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_24/Component_Function_5/N1  ( .A1(\SB4_24/i0_0 ), .A2(
        \SB4_24/i3[0] ), .ZN(\SB4_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_0/N3  ( .A1(\SB4_25/i0[10] ), .A2(
        \SB4_25/i0_4 ), .A3(\SB4_25/i0_3 ), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_25/Component_Function_0/N2  ( .A1(\SB4_25/i0[8] ), .A2(n821), 
        .A3(\SB4_25/i0[6] ), .ZN(\SB4_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_25/Component_Function_0/N1  ( .A1(\SB4_25/i0[10] ), .A2(
        \SB4_25/i0[9] ), .ZN(\SB4_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_1/N2  ( .A1(\SB4_25/i0_3 ), .A2(
        \SB4_25/i1_7 ), .A3(\SB4_25/i0[8] ), .ZN(
        \SB4_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_25/Component_Function_1/N1  ( .A1(\SB4_25/i0_3 ), .A2(
        \SB4_25/i1[9] ), .ZN(\SB4_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_5/N4  ( .A1(\SB4_25/i0[9] ), .A2(
        \SB4_25/i0[6] ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_5/N2  ( .A1(\SB4_25/i0_0 ), .A2(
        \SB4_25/i0[6] ), .A3(\SB4_25/i0[10] ), .ZN(
        \SB4_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_25/Component_Function_5/N1  ( .A1(\SB4_25/i0_0 ), .A2(
        \SB4_25/i3[0] ), .ZN(\SB4_25/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB4_26/Component_Function_0/N1  ( .A1(\SB4_26/i0[10] ), .A2(
        \SB4_26/i0[9] ), .ZN(\SB4_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_1/N3  ( .A1(\SB4_26/i1_5 ), .A2(
        \SB4_26/i0[6] ), .A3(\SB4_26/i0[9] ), .ZN(
        \SB4_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_26/Component_Function_1/N2  ( .A1(n1671), .A2(\SB4_26/i1_7 ), 
        .A3(\SB4_26/i0[8] ), .ZN(\SB4_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_26/Component_Function_1/N1  ( .A1(\SB4_26/i0_3 ), .A2(
        \SB4_26/i1[9] ), .ZN(\SB4_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_5/N4  ( .A1(\SB4_26/i0[9] ), .A2(
        \SB4_26/i0[6] ), .A3(\SB4_26/i0_4 ), .ZN(
        \SB4_26/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_26/Component_Function_5/N1  ( .A1(\SB4_26/i0_0 ), .A2(
        \SB4_26/i3[0] ), .ZN(\SB4_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_0/N4  ( .A1(n552), .A2(n1949), .A3(
        \SB4_27/i0_0 ), .ZN(\SB4_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_27/Component_Function_0/N2  ( .A1(\SB4_27/i0[8] ), .A2(n552), 
        .A3(\SB4_27/i0[6] ), .ZN(\SB4_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_27/Component_Function_0/N1  ( .A1(\SB4_27/i0[10] ), .A2(
        \SB4_27/i0[9] ), .ZN(\SB4_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_1/N3  ( .A1(\SB4_27/i1_5 ), .A2(
        \SB4_27/i0[6] ), .A3(\SB4_27/i0[9] ), .ZN(
        \SB4_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_27/Component_Function_1/N2  ( .A1(n1949), .A2(\SB4_27/i1_7 ), 
        .A3(\SB4_27/i0[8] ), .ZN(\SB4_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_27/Component_Function_1/N1  ( .A1(n1949), .A2(\SB4_27/i1[9] ), 
        .ZN(\SB4_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_5/N4  ( .A1(\SB4_27/i0[9] ), .A2(
        \SB4_27/i0[6] ), .A3(n780), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_27/Component_Function_5/N2  ( .A1(\SB4_27/i0_0 ), .A2(
        \SB4_27/i0[6] ), .A3(\SB4_27/i0[10] ), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_27/Component_Function_5/N1  ( .A1(\SB4_27/i0_0 ), .A2(
        \SB4_27/i3[0] ), .ZN(\SB4_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_28/Component_Function_0/N2  ( .A1(\SB4_28/i0[8] ), .A2(
        \SB4_28/i0[7] ), .A3(\SB4_28/i0[6] ), .ZN(
        \SB4_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_28/Component_Function_0/N1  ( .A1(\SB4_28/i0[10] ), .A2(
        \SB4_28/i0[9] ), .ZN(\SB4_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_28/Component_Function_1/N3  ( .A1(\SB4_28/i1_5 ), .A2(
        \SB4_28/i0[6] ), .A3(\SB4_28/i0[9] ), .ZN(
        \SB4_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_28/Component_Function_1/N2  ( .A1(n866), .A2(\SB4_28/i1_7 ), 
        .A3(\SB4_28/i0[8] ), .ZN(\SB4_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_28/Component_Function_1/N1  ( .A1(\SB4_28/i0_3 ), .A2(
        \SB4_28/i1[9] ), .ZN(\SB4_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_28/Component_Function_5/N4  ( .A1(\SB4_28/i0[9] ), .A2(
        \SB4_28/i0[6] ), .A3(\SB4_28/i0_4 ), .ZN(
        \SB4_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_28/Component_Function_5/N2  ( .A1(\SB4_28/i0_0 ), .A2(
        \SB4_28/i0[6] ), .A3(\SB4_28/i0[10] ), .ZN(
        \SB4_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_28/Component_Function_5/N1  ( .A1(\SB4_28/i0_0 ), .A2(
        \SB4_28/i3[0] ), .ZN(\SB4_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_29/Component_Function_0/N4  ( .A1(n1963), .A2(\SB4_29/i0_3 ), 
        .A3(\SB4_29/i0_0 ), .ZN(\SB4_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_29/Component_Function_0/N2  ( .A1(\SB4_29/i0[8] ), .A2(n1963), 
        .A3(n791), .ZN(\SB4_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_29/Component_Function_0/N1  ( .A1(\SB4_29/i0[10] ), .A2(n790), 
        .ZN(\SB4_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_29/Component_Function_1/N4  ( .A1(n554), .A2(\SB4_29/i0[8] ), 
        .A3(n2131), .ZN(\SB4_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_29/Component_Function_1/N2  ( .A1(\SB4_29/i0_3 ), .A2(n554), 
        .A3(\SB4_29/i0[8] ), .ZN(\SB4_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_29/Component_Function_1/N1  ( .A1(\SB4_29/i0_3 ), .A2(
        \SB4_29/i1[9] ), .ZN(\SB4_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_29/Component_Function_5/N2  ( .A1(\SB4_29/i0_0 ), .A2(n791), 
        .A3(\SB4_29/i0[10] ), .ZN(\SB4_29/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X1 \SB4_29/Component_Function_5/N1  ( .A1(\SB4_29/i0_0 ), .A2(n555), 
        .ZN(\SB4_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_30/Component_Function_0/N3  ( .A1(\SB4_30/i0[10] ), .A2(
        \SB4_30/i0_4 ), .A3(n1668), .ZN(
        \SB4_30/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB4_30/Component_Function_0/N1  ( .A1(\SB4_30/i0[10] ), .A2(
        \SB4_30/i0[9] ), .ZN(\SB4_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_30/Component_Function_1/N4  ( .A1(\SB4_30/i1_7 ), .A2(
        \SB4_30/i0[8] ), .A3(\SB4_30/i0_4 ), .ZN(
        \SB4_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_30/Component_Function_1/N2  ( .A1(n1668), .A2(\SB4_30/i1_7 ), 
        .A3(\SB4_30/i0[8] ), .ZN(\SB4_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_30/Component_Function_1/N1  ( .A1(\SB4_30/i0_3 ), .A2(
        \SB4_30/i1[9] ), .ZN(\SB4_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_30/Component_Function_5/N2  ( .A1(\SB4_30/i0_0 ), .A2(
        \SB4_30/i0[6] ), .A3(\SB4_30/i0[10] ), .ZN(
        \SB4_30/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_30/Component_Function_5/N1  ( .A1(\SB4_30/i0_0 ), .A2(
        \SB4_30/i3[0] ), .ZN(\SB4_30/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB4_31/Component_Function_0/N1  ( .A1(\SB4_31/i0[10] ), .A2(
        \SB4_31/i0[9] ), .ZN(\SB4_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N3  ( .A1(n1964), .A2(\SB4_31/i0[6] ), 
        .A3(\SB4_31/i0[9] ), .ZN(\SB4_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N2  ( .A1(n2106), .A2(\SB4_31/i1_7 ), 
        .A3(\SB4_31/i0[8] ), .ZN(\SB4_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_31/Component_Function_1/N1  ( .A1(n1670), .A2(\SB4_31/i1[9] ), 
        .ZN(\SB4_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_31/Component_Function_5/N4  ( .A1(\SB4_31/i0[9] ), .A2(
        \SB4_31/i0[6] ), .A3(\SB4_31/i0_4 ), .ZN(
        \SB4_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_31/Component_Function_5/N2  ( .A1(\SB4_31/i0_0 ), .A2(
        \SB4_31/i0[6] ), .A3(\SB4_31/i0[10] ), .ZN(
        \SB4_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_31/Component_Function_5/N1  ( .A1(\SB4_31/i0_0 ), .A2(
        \SB4_31/i3[0] ), .ZN(\SB4_31/Component_Function_5/NAND4_in[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_31_5  ( .A(\MC_ARK_ARC_1_0/temp6[0] ), .B(
        \MC_ARK_ARC_1_0/temp5[0] ), .ZN(\RI1[1][0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_31_5  ( .A(\MC_ARK_ARC_1_0/temp3[0] ), .B(
        \MC_ARK_ARC_1_0/temp4[0] ), .ZN(\MC_ARK_ARC_1_0/temp6[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_31_5  ( .A(\MC_ARK_ARC_1_0/temp1[0] ), .B(
        \MC_ARK_ARC_1_0/temp2[0] ), .ZN(\MC_ARK_ARC_1_0/temp5[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_31_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[36] ), 
        .B(n389), .ZN(\MC_ARK_ARC_1_0/temp4[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_31_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[66] ), .ZN(\MC_ARK_ARC_1_0/temp3[0] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_31_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[162] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[138] ), .ZN(\MC_ARK_ARC_1_0/temp2[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_31_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[186] ), .ZN(\MC_ARK_ARC_1_0/temp1[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_31_4  ( .A(\MC_ARK_ARC_1_0/temp5[1] ), .B(
        \MC_ARK_ARC_1_0/temp6[1] ), .ZN(\RI1[1][1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_31_4  ( .A(\MC_ARK_ARC_1_0/temp3[1] ), .B(
        \MC_ARK_ARC_1_0/temp4[1] ), .ZN(\MC_ARK_ARC_1_0/temp6[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_31_4  ( .A(\MC_ARK_ARC_1_0/temp1[1] ), .B(
        \MC_ARK_ARC_1_0/temp2[1] ), .ZN(\MC_ARK_ARC_1_0/temp5[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_31_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[37] ), 
        .B(n427), .ZN(\MC_ARK_ARC_1_0/temp4[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_31_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[67] ), .ZN(\MC_ARK_ARC_1_0/temp3[1] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_31_4  ( .A(\RI5[0][163] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[139] ), .ZN(\MC_ARK_ARC_1_0/temp2[1] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_31_4  ( .A(\RI5[0][1] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[187] ), .ZN(\MC_ARK_ARC_1_0/temp1[1] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_31_3  ( .A(\MC_ARK_ARC_1_0/temp5[2] ), .B(
        \MC_ARK_ARC_1_0/temp6[2] ), .ZN(\RI1[1][2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_31_3  ( .A(\MC_ARK_ARC_1_0/temp3[2] ), .B(
        \MC_ARK_ARC_1_0/temp4[2] ), .ZN(\MC_ARK_ARC_1_0/temp6[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_31_3  ( .A(\MC_ARK_ARC_1_0/temp2[2] ), .B(
        \MC_ARK_ARC_1_0/temp1[2] ), .ZN(\MC_ARK_ARC_1_0/temp5[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_31_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[38] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[27] ), .ZN(\MC_ARK_ARC_1_0/temp4[2] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_31_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[104] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_0/temp3[2] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_31_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[164] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[140] ), .ZN(\MC_ARK_ARC_1_0/temp2[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_31_3  ( .A(\RI5[0][2] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[188] ), .ZN(\MC_ARK_ARC_1_0/temp1[2] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_31_2  ( .A(\MC_ARK_ARC_1_0/temp5[3] ), .B(
        \MC_ARK_ARC_1_0/temp6[3] ), .ZN(\RI1[1][3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_31_2  ( .A(\MC_ARK_ARC_1_0/temp3[3] ), .B(
        \MC_ARK_ARC_1_0/temp4[3] ), .ZN(\MC_ARK_ARC_1_0/temp6[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_31_2  ( .A(\MC_ARK_ARC_1_0/temp2[3] ), .B(
        \MC_ARK_ARC_1_0/temp1[3] ), .ZN(\MC_ARK_ARC_1_0/temp5[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_31_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[39] ), 
        .B(n466), .ZN(\MC_ARK_ARC_1_0/temp4[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_31_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[69] ), .ZN(\MC_ARK_ARC_1_0/temp3[3] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_31_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .B(\RI5[0][165] ), .ZN(\MC_ARK_ARC_1_0/temp2[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_31_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[3] ), 
        .B(n1959), .ZN(\MC_ARK_ARC_1_0/temp1[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_31_1  ( .A(\MC_ARK_ARC_1_0/temp6[4] ), .B(
        \MC_ARK_ARC_1_0/temp5[4] ), .ZN(\RI1[1][4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_31_1  ( .A(\MC_ARK_ARC_1_0/temp3[4] ), .B(
        \MC_ARK_ARC_1_0/temp4[4] ), .ZN(\MC_ARK_ARC_1_0/temp6[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_31_1  ( .A(\MC_ARK_ARC_1_0/temp2[4] ), .B(
        \MC_ARK_ARC_1_0/temp1[4] ), .ZN(\MC_ARK_ARC_1_0/temp5[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_31_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[40] ), 
        .B(n342), .ZN(\MC_ARK_ARC_1_0/temp4[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_31_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_0/temp3[4] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_31_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[142] ), .ZN(\MC_ARK_ARC_1_0/temp2[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_31_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[190] ), .ZN(\MC_ARK_ARC_1_0/temp1[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_31_0  ( .A(n1961), .B(n469), .ZN(
        \MC_ARK_ARC_1_0/temp4[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_31_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .B(n1962), .ZN(\MC_ARK_ARC_1_0/temp3[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_31_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[143] ), .ZN(\MC_ARK_ARC_1_0/temp2[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_31_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[5] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[191] ), .ZN(\MC_ARK_ARC_1_0/temp1[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_30_5  ( .A(\MC_ARK_ARC_1_0/temp5[6] ), .B(
        \MC_ARK_ARC_1_0/temp6[6] ), .ZN(\RI1[1][6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_30_5  ( .A(\MC_ARK_ARC_1_0/temp3[6] ), .B(
        \MC_ARK_ARC_1_0/temp4[6] ), .ZN(\MC_ARK_ARC_1_0/temp6[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_30_5  ( .A(\MC_ARK_ARC_1_0/temp1[6] ), .B(
        \MC_ARK_ARC_1_0/temp2[6] ), .ZN(\MC_ARK_ARC_1_0/temp5[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_30_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .B(n330), .ZN(\MC_ARK_ARC_1_0/temp4[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_30_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[108] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[72] ), .ZN(\MC_ARK_ARC_1_0/temp3[6] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_30_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[144] ), .ZN(\MC_ARK_ARC_1_0/temp2[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_30_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_0/temp1[6] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_30_4  ( .A(\MC_ARK_ARC_1_0/temp5[7] ), .B(
        \MC_ARK_ARC_1_0/temp6[7] ), .ZN(\RI1[1][7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_30_4  ( .A(\MC_ARK_ARC_1_0/temp3[7] ), .B(
        \MC_ARK_ARC_1_0/temp4[7] ), .ZN(\MC_ARK_ARC_1_0/temp6[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_30_4  ( .A(\MC_ARK_ARC_1_0/temp1[7] ), .B(
        \MC_ARK_ARC_1_0/temp2[7] ), .ZN(\MC_ARK_ARC_1_0/temp5[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_30_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .B(n323), .ZN(\MC_ARK_ARC_1_0/temp4[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_30_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[73] ), .ZN(\MC_ARK_ARC_1_0/temp3[7] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_30_4  ( .A(\RI5[0][169] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[145] ), .ZN(\MC_ARK_ARC_1_0/temp2[7] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_30_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .B(\RI5[0][1] ), .ZN(\MC_ARK_ARC_1_0/temp1[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_30_3  ( .A(\MC_ARK_ARC_1_0/temp6[8] ), .B(
        \MC_ARK_ARC_1_0/temp5[8] ), .ZN(\RI1[1][8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_30_3  ( .A(\MC_ARK_ARC_1_0/temp3[8] ), .B(
        \MC_ARK_ARC_1_0/temp4[8] ), .ZN(\MC_ARK_ARC_1_0/temp6[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_30_3  ( .A(\MC_ARK_ARC_1_0/temp2[8] ), .B(
        \MC_ARK_ARC_1_0/temp1[8] ), .ZN(\MC_ARK_ARC_1_0/temp5[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_30_3  ( .A(n1475), .B(n317), .ZN(
        \MC_ARK_ARC_1_0/temp4[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_30_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[74] ), .ZN(\MC_ARK_ARC_1_0/temp3[8] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_30_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[146] ), 
        .B(\RI5[0][170] ), .ZN(\MC_ARK_ARC_1_0/temp2[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_30_3  ( .A(\RI5[0][2] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_0/temp1[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_30_2  ( .A(\MC_ARK_ARC_1_0/temp5[9] ), .B(
        \MC_ARK_ARC_1_0/temp6[9] ), .ZN(\RI1[1][9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_30_2  ( .A(\MC_ARK_ARC_1_0/temp3[9] ), .B(
        \MC_ARK_ARC_1_0/temp4[9] ), .ZN(\MC_ARK_ARC_1_0/temp6[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_30_2  ( .A(\MC_ARK_ARC_1_0/temp1[9] ), .B(
        \MC_ARK_ARC_1_0/temp2[9] ), .ZN(\MC_ARK_ARC_1_0/temp5[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_30_2  ( .A(\RI5[0][45] ), .B(n486), .ZN(
        \MC_ARK_ARC_1_0/temp4[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_30_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[111] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[75] ), .ZN(\MC_ARK_ARC_1_0/temp3[9] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_30_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[171] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[147] ), .ZN(\MC_ARK_ARC_1_0/temp2[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_30_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[3] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_0/temp1[9] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_30_1  ( .A(\MC_ARK_ARC_1_0/temp5[10] ), .B(
        \MC_ARK_ARC_1_0/temp6[10] ), .ZN(\RI1[1][10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_30_1  ( .A(\MC_ARK_ARC_1_0/temp3[10] ), .B(
        \MC_ARK_ARC_1_0/temp4[10] ), .ZN(\MC_ARK_ARC_1_0/temp6[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_30_1  ( .A(\MC_ARK_ARC_1_0/temp2[10] ), .B(
        \MC_ARK_ARC_1_0/temp1[10] ), .ZN(\MC_ARK_ARC_1_0/temp5[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_30_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .B(n502), .ZN(\MC_ARK_ARC_1_0/temp4[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_30_1  ( .A(\RI5[0][76] ), .B(\RI5[0][112] ), 
        .ZN(\MC_ARK_ARC_1_0/temp3[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_30_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[148] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_30_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_0/temp1[10] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_30_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[47] ), 
        .B(\MC_ARK_ARC_1_0/buf_keyinput[11] ), .ZN(\MC_ARK_ARC_1_0/temp4[11] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_30_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[113] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_30_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[149] ), 
        .B(n2150), .ZN(\MC_ARK_ARC_1_0/temp2[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_30_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[5] ), 
        .B(n2146), .ZN(\MC_ARK_ARC_1_0/temp1[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_29_5  ( .A(\MC_ARK_ARC_1_0/temp6[12] ), .B(
        \MC_ARK_ARC_1_0/temp5[12] ), .ZN(\RI1[1][12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_29_5  ( .A(\MC_ARK_ARC_1_0/temp3[12] ), .B(
        \MC_ARK_ARC_1_0/temp4[12] ), .ZN(\MC_ARK_ARC_1_0/temp6[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_29_5  ( .A(\MC_ARK_ARC_1_0/temp1[12] ), .B(
        \MC_ARK_ARC_1_0/temp2[12] ), .ZN(\MC_ARK_ARC_1_0/temp5[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_29_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .B(n290), .ZN(\MC_ARK_ARC_1_0/temp4[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_29_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[78] ), .ZN(\MC_ARK_ARC_1_0/temp3[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_29_5  ( .A(\RI5[0][174] ), .B(\RI5[0][150] ), 
        .ZN(\MC_ARK_ARC_1_0/temp2[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_29_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_0/temp1[12] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_29_4  ( .A(\MC_ARK_ARC_1_0/temp5[13] ), .B(
        \MC_ARK_ARC_1_0/temp6[13] ), .ZN(\RI1[1][13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_29_4  ( .A(\MC_ARK_ARC_1_0/temp3[13] ), .B(
        \MC_ARK_ARC_1_0/temp4[13] ), .ZN(\MC_ARK_ARC_1_0/temp6[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_29_4  ( .A(\MC_ARK_ARC_1_0/temp1[13] ), .B(
        \MC_ARK_ARC_1_0/temp2[13] ), .ZN(\MC_ARK_ARC_1_0/temp5[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_29_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[49] ), 
        .B(n283), .ZN(\MC_ARK_ARC_1_0/temp4[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_29_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[79] ), .ZN(\MC_ARK_ARC_1_0/temp3[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_29_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[151] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_29_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_0/temp1[13] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_29_3  ( .A(\MC_ARK_ARC_1_0/temp6[14] ), .B(
        \MC_ARK_ARC_1_0/temp5[14] ), .ZN(\RI1[1][14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_29_3  ( .A(\MC_ARK_ARC_1_0/temp3[14] ), .B(
        \MC_ARK_ARC_1_0/temp4[14] ), .ZN(\MC_ARK_ARC_1_0/temp6[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_29_3  ( .A(\MC_ARK_ARC_1_0/temp2[14] ), .B(
        \MC_ARK_ARC_1_0/temp1[14] ), .ZN(\MC_ARK_ARC_1_0/temp5[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_29_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[50] ), 
        .B(n378), .ZN(\MC_ARK_ARC_1_0/temp4[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_29_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[80] ), 
        .B(n1941), .ZN(\MC_ARK_ARC_1_0/temp3[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_29_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[176] ), 
        .B(\RI5[0][152] ), .ZN(\MC_ARK_ARC_1_0/temp2[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_29_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_0/temp1[14] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_29_2  ( .A(\MC_ARK_ARC_1_0/temp5[15] ), .B(
        \MC_ARK_ARC_1_0/temp6[15] ), .ZN(\RI1[1][15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_29_2  ( .A(\MC_ARK_ARC_1_0/temp3[15] ), .B(
        \MC_ARK_ARC_1_0/temp4[15] ), .ZN(\MC_ARK_ARC_1_0/temp6[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_29_2  ( .A(\MC_ARK_ARC_1_0/temp2[15] ), .B(
        \MC_ARK_ARC_1_0/temp1[15] ), .ZN(\MC_ARK_ARC_1_0/temp5[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_29_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .B(n501), .ZN(\MC_ARK_ARC_1_0/temp4[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_29_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[117] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[81] ), .ZN(\MC_ARK_ARC_1_0/temp3[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_29_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[177] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[153] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_29_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[15] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_0/temp1[15] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_29_1  ( .A(\MC_ARK_ARC_1_0/temp5[16] ), .B(
        \MC_ARK_ARC_1_0/temp6[16] ), .ZN(\RI1[1][16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_29_1  ( .A(\MC_ARK_ARC_1_0/temp3[16] ), .B(
        \MC_ARK_ARC_1_0/temp4[16] ), .ZN(\MC_ARK_ARC_1_0/temp6[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_29_1  ( .A(\MC_ARK_ARC_1_0/temp2[16] ), .B(
        \MC_ARK_ARC_1_0/temp1[16] ), .ZN(\MC_ARK_ARC_1_0/temp5[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_29_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[52] ), 
        .B(n263), .ZN(\MC_ARK_ARC_1_0/temp4[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_29_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[118] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[82] ), .ZN(\MC_ARK_ARC_1_0/temp3[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_29_1  ( .A(\RI5[0][178] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[154] ), .ZN(\MC_ARK_ARC_1_0/temp2[16] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_29_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_0/temp1[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_29_0  ( .A(n1631), .B(n256), .ZN(
        \MC_ARK_ARC_1_0/temp4[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_29_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[83] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[119] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_29_0  ( .A(n2116), .B(n1660), .ZN(
        \MC_ARK_ARC_1_0/temp2[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_29_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[17] ), 
        .B(n2146), .ZN(\MC_ARK_ARC_1_0/temp1[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_28_5  ( .A(\MC_ARK_ARC_1_0/temp5[18] ), .B(
        \MC_ARK_ARC_1_0/temp6[18] ), .ZN(\RI1[1][18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_28_5  ( .A(\MC_ARK_ARC_1_0/temp3[18] ), .B(
        \MC_ARK_ARC_1_0/temp4[18] ), .ZN(\MC_ARK_ARC_1_0/temp6[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_28_5  ( .A(\MC_ARK_ARC_1_0/temp1[18] ), .B(
        \MC_ARK_ARC_1_0/temp2[18] ), .ZN(\MC_ARK_ARC_1_0/temp5[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_28_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[54] ), 
        .B(n250), .ZN(\MC_ARK_ARC_1_0/temp4[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_28_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[84] ), .ZN(\MC_ARK_ARC_1_0/temp3[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_28_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .B(\RI5[0][156] ), .ZN(\MC_ARK_ARC_1_0/temp2[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_28_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_0/temp1[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_28_4  ( .A(\MC_ARK_ARC_1_0/temp5[19] ), .B(
        \MC_ARK_ARC_1_0/temp6[19] ), .ZN(\RI1[1][19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_28_4  ( .A(\MC_ARK_ARC_1_0/temp3[19] ), .B(
        \MC_ARK_ARC_1_0/temp4[19] ), .ZN(\MC_ARK_ARC_1_0/temp6[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_28_4  ( .A(\MC_ARK_ARC_1_0/temp1[19] ), .B(
        \MC_ARK_ARC_1_0/temp2[19] ), .ZN(\MC_ARK_ARC_1_0/temp5[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_28_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[55] ), 
        .B(n244), .ZN(\MC_ARK_ARC_1_0/temp4[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_28_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[85] ), .ZN(\MC_ARK_ARC_1_0/temp3[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_28_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[181] ), 
        .B(\RI5[0][157] ), .ZN(\MC_ARK_ARC_1_0/temp2[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_28_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[13] ), .ZN(\MC_ARK_ARC_1_0/temp1[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_28_3  ( .A(\MC_ARK_ARC_1_0/temp5[20] ), .B(
        \MC_ARK_ARC_1_0/temp6[20] ), .ZN(\RI1[1][20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_28_3  ( .A(\MC_ARK_ARC_1_0/temp3[20] ), .B(
        \MC_ARK_ARC_1_0/temp4[20] ), .ZN(\MC_ARK_ARC_1_0/temp6[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_28_3  ( .A(\MC_ARK_ARC_1_0/temp1[20] ), .B(
        \MC_ARK_ARC_1_0/temp2[20] ), .ZN(\MC_ARK_ARC_1_0/temp5[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_28_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[56] ), 
        .B(n238), .ZN(\MC_ARK_ARC_1_0/temp4[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_28_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[86] ), .ZN(\MC_ARK_ARC_1_0/temp3[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_28_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[158] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_28_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_0/temp1[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_28_2  ( .A(\MC_ARK_ARC_1_0/temp5[21] ), .B(
        \MC_ARK_ARC_1_0/temp6[21] ), .ZN(\RI1[1][21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_28_2  ( .A(\MC_ARK_ARC_1_0/temp3[21] ), .B(
        \MC_ARK_ARC_1_0/temp4[21] ), .ZN(\MC_ARK_ARC_1_0/temp6[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_28_2  ( .A(\MC_ARK_ARC_1_0/temp2[21] ), .B(
        \MC_ARK_ARC_1_0/temp1[21] ), .ZN(\MC_ARK_ARC_1_0/temp5[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_28_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[57] ), 
        .B(n485), .ZN(\MC_ARK_ARC_1_0/temp4[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_28_2  ( .A(\RI5[0][123] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[87] ), .ZN(\MC_ARK_ARC_1_0/temp3[21] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_28_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[159] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[183] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_28_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[15] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_0/temp1[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_28_1  ( .A(\MC_ARK_ARC_1_0/temp5[22] ), .B(
        \MC_ARK_ARC_1_0/temp6[22] ), .ZN(\RI1[1][22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_28_1  ( .A(\MC_ARK_ARC_1_0/temp3[22] ), .B(
        \MC_ARK_ARC_1_0/temp4[22] ), .ZN(\MC_ARK_ARC_1_0/temp6[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_28_1  ( .A(\MC_ARK_ARC_1_0/temp1[22] ), .B(
        \MC_ARK_ARC_1_0/temp2[22] ), .ZN(\MC_ARK_ARC_1_0/temp5[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_28_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[58] ), 
        .B(n511), .ZN(\MC_ARK_ARC_1_0/temp4[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_28_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_0/temp3[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_28_1  ( .A(\RI5[0][184] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[160] ), .ZN(\MC_ARK_ARC_1_0/temp2[22] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_28_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_0/temp1[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_28_0  ( .A(n787), .B(n217), .ZN(
        \MC_ARK_ARC_1_0/temp4[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_28_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[89] ), 
        .B(n1939), .ZN(\MC_ARK_ARC_1_0/temp3[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_28_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[161] ), 
        .B(n795), .ZN(\MC_ARK_ARC_1_0/temp2[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_28_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[17] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[23] ), .ZN(\MC_ARK_ARC_1_0/temp1[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_27_5  ( .A(\MC_ARK_ARC_1_0/temp5[24] ), .B(
        \MC_ARK_ARC_1_0/temp6[24] ), .ZN(\RI1[1][24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_27_5  ( .A(\MC_ARK_ARC_1_0/temp3[24] ), .B(
        \MC_ARK_ARC_1_0/temp4[24] ), .ZN(\MC_ARK_ARC_1_0/temp6[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_27_5  ( .A(\MC_ARK_ARC_1_0/temp1[24] ), .B(
        \MC_ARK_ARC_1_0/temp2[24] ), .ZN(\MC_ARK_ARC_1_0/temp5[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_27_5  ( .A(\RI5[0][60] ), .B(n210), .ZN(
        \MC_ARK_ARC_1_0/temp4[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_27_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[90] ), .ZN(\MC_ARK_ARC_1_0/temp3[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_27_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_27_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[18] ), .ZN(\MC_ARK_ARC_1_0/temp1[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_27_4  ( .A(\MC_ARK_ARC_1_0/temp5[25] ), .B(
        \MC_ARK_ARC_1_0/temp6[25] ), .ZN(\RI1[1][25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_27_4  ( .A(\MC_ARK_ARC_1_0/temp3[25] ), .B(
        \MC_ARK_ARC_1_0/temp4[25] ), .ZN(\MC_ARK_ARC_1_0/temp6[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_27_4  ( .A(\MC_ARK_ARC_1_0/temp1[25] ), .B(
        \MC_ARK_ARC_1_0/temp2[25] ), .ZN(\MC_ARK_ARC_1_0/temp5[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_27_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[129] ), .ZN(\MC_ARK_ARC_1_0/temp4[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_27_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_0/temp3[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_27_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[187] ), 
        .B(\RI5[0][163] ), .ZN(\MC_ARK_ARC_1_0/temp2[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_27_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[19] ), .ZN(\MC_ARK_ARC_1_0/temp1[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_27_3  ( .A(\MC_ARK_ARC_1_0/temp5[26] ), .B(
        \MC_ARK_ARC_1_0/temp6[26] ), .ZN(\RI1[1][26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_27_3  ( .A(\MC_ARK_ARC_1_0/temp3[26] ), .B(
        \MC_ARK_ARC_1_0/temp4[26] ), .ZN(\MC_ARK_ARC_1_0/temp6[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_27_3  ( .A(\MC_ARK_ARC_1_0/temp1[26] ), .B(
        \MC_ARK_ARC_1_0/temp2[26] ), .ZN(\MC_ARK_ARC_1_0/temp5[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_27_3  ( .A(\RI5[0][62] ), .B(Key[187]), .ZN(
        \MC_ARK_ARC_1_0/temp4[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_27_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_27_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[164] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_27_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_0/temp1[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_27_2  ( .A(\RI5[0][63] ), .B(n372), .ZN(
        \MC_ARK_ARC_1_0/temp4[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_27_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[93] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[129] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_27_2  ( .A(\RI5[0][165] ), .B(n1495), .ZN(
        \MC_ARK_ARC_1_0/temp2[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_27_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[21] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[27] ), .ZN(\MC_ARK_ARC_1_0/temp1[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_27_1  ( .A(\MC_ARK_ARC_1_0/temp5[28] ), .B(
        \MC_ARK_ARC_1_0/temp6[28] ), .ZN(\RI1[1][28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_27_1  ( .A(\MC_ARK_ARC_1_0/temp3[28] ), .B(
        \MC_ARK_ARC_1_0/temp4[28] ), .ZN(\MC_ARK_ARC_1_0/temp6[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_27_1  ( .A(\MC_ARK_ARC_1_0/temp2[28] ), .B(
        \MC_ARK_ARC_1_0/temp1[28] ), .ZN(\MC_ARK_ARC_1_0/temp5[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_27_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .B(n503), .ZN(\MC_ARK_ARC_1_0/temp4[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_27_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[130] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[94] ), .ZN(\MC_ARK_ARC_1_0/temp3[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_27_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_27_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[28] ), .ZN(\MC_ARK_ARC_1_0/temp1[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_27_0  ( .A(\MC_ARK_ARC_1_0/temp5[29] ), .B(
        \MC_ARK_ARC_1_0/temp6[29] ), .ZN(\RI1[1][29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_27_0  ( .A(\MC_ARK_ARC_1_0/temp3[29] ), .B(
        \MC_ARK_ARC_1_0/temp4[29] ), .ZN(\MC_ARK_ARC_1_0/temp6[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_27_0  ( .A(\MC_ARK_ARC_1_0/temp1[29] ), .B(
        \MC_ARK_ARC_1_0/temp2[29] ), .ZN(\MC_ARK_ARC_1_0/temp5[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_27_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[65] ), 
        .B(n359), .ZN(\MC_ARK_ARC_1_0/temp4[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_27_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[191] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_27_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[23] ), 
        .B(n1960), .ZN(\MC_ARK_ARC_1_0/temp1[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_26_5  ( .A(\MC_ARK_ARC_1_0/temp5[30] ), .B(
        \MC_ARK_ARC_1_0/temp6[30] ), .ZN(\RI1[1][30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_26_5  ( .A(\MC_ARK_ARC_1_0/temp3[30] ), .B(
        \MC_ARK_ARC_1_0/temp4[30] ), .ZN(\MC_ARK_ARC_1_0/temp6[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_26_5  ( .A(\MC_ARK_ARC_1_0/temp1[30] ), .B(
        \MC_ARK_ARC_1_0/temp2[30] ), .ZN(\MC_ARK_ARC_1_0/temp5[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_26_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[66] ), 
        .B(n465), .ZN(\MC_ARK_ARC_1_0/temp4[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_26_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[96] ), .ZN(\MC_ARK_ARC_1_0/temp3[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_26_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_26_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[24] ), .ZN(\MC_ARK_ARC_1_0/temp1[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_26_4  ( .A(\MC_ARK_ARC_1_0/temp5[31] ), .B(
        \MC_ARK_ARC_1_0/temp6[31] ), .ZN(\RI1[1][31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_26_4  ( .A(\MC_ARK_ARC_1_0/temp3[31] ), .B(
        \MC_ARK_ARC_1_0/temp4[31] ), .ZN(\MC_ARK_ARC_1_0/temp6[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_26_4  ( .A(\MC_ARK_ARC_1_0/temp1[31] ), .B(
        \MC_ARK_ARC_1_0/temp2[31] ), .ZN(\MC_ARK_ARC_1_0/temp5[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_26_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[142] ), .ZN(\MC_ARK_ARC_1_0/temp4[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_26_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[133] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[97] ), .ZN(\MC_ARK_ARC_1_0/temp3[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_26_4  ( .A(\RI5[0][1] ), .B(\RI5[0][169] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_26_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[25] ), .ZN(\MC_ARK_ARC_1_0/temp1[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_26_3  ( .A(\MC_ARK_ARC_1_0/temp5[32] ), .B(
        \MC_ARK_ARC_1_0/temp6[32] ), .ZN(\RI1[1][32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_26_3  ( .A(\MC_ARK_ARC_1_0/temp3[32] ), .B(
        \MC_ARK_ARC_1_0/temp4[32] ), .ZN(\MC_ARK_ARC_1_0/temp6[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_26_3  ( .A(\MC_ARK_ARC_1_0/temp2[32] ), .B(
        \MC_ARK_ARC_1_0/temp1[32] ), .ZN(\MC_ARK_ARC_1_0/temp5[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_26_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[68] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[184] ), .ZN(\MC_ARK_ARC_1_0/temp4[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_26_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[98] ), .ZN(\MC_ARK_ARC_1_0/temp3[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_26_3  ( .A(\RI5[0][170] ), .B(\RI5[0][2] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_26_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[32] ), .ZN(\MC_ARK_ARC_1_0/temp1[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_26_2  ( .A(\MC_ARK_ARC_1_0/temp6[33] ), .B(
        \MC_ARK_ARC_1_0/temp5[33] ), .ZN(\RI1[1][33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_26_2  ( .A(\MC_ARK_ARC_1_0/temp3[33] ), .B(
        \MC_ARK_ARC_1_0/temp4[33] ), .ZN(\MC_ARK_ARC_1_0/temp6[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_26_2  ( .A(\MC_ARK_ARC_1_0/temp2[33] ), .B(
        \MC_ARK_ARC_1_0/temp1[33] ), .ZN(\MC_ARK_ARC_1_0/temp5[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_26_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[69] ), 
        .B(n333), .ZN(\MC_ARK_ARC_1_0/temp4[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_26_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[135] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[99] ), .ZN(\MC_ARK_ARC_1_0/temp3[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_26_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[171] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[3] ), .ZN(\MC_ARK_ARC_1_0/temp2[33] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_26_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[27] ), .ZN(\MC_ARK_ARC_1_0/temp1[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_26_1  ( .A(\MC_ARK_ARC_1_0/temp5[34] ), .B(
        \MC_ARK_ARC_1_0/temp6[34] ), .ZN(\RI1[1][34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_26_1  ( .A(\MC_ARK_ARC_1_0/temp3[34] ), .B(
        \MC_ARK_ARC_1_0/temp4[34] ), .ZN(\MC_ARK_ARC_1_0/temp6[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_26_1  ( .A(\MC_ARK_ARC_1_0/temp1[34] ), .B(
        \MC_ARK_ARC_1_0/temp2[34] ), .ZN(\MC_ARK_ARC_1_0/temp5[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_26_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .B(n496), .ZN(\MC_ARK_ARC_1_0/temp4[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_26_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_26_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_26_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[28] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[34] ), .ZN(\MC_ARK_ARC_1_0/temp1[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_26_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .B(n482), .ZN(\MC_ARK_ARC_1_0/temp4[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_26_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[101] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[137] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_26_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[5] ), 
        .B(n2151), .ZN(\MC_ARK_ARC_1_0/temp2[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_26_0  ( .A(n1508), .B(n1470), .ZN(
        \MC_ARK_ARC_1_0/temp1[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_25_5  ( .A(\MC_ARK_ARC_1_0/temp5[36] ), .B(
        \MC_ARK_ARC_1_0/temp6[36] ), .ZN(\RI1[1][36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_25_5  ( .A(\MC_ARK_ARC_1_0/temp3[36] ), .B(
        \MC_ARK_ARC_1_0/temp4[36] ), .ZN(\MC_ARK_ARC_1_0/temp6[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_25_5  ( .A(\MC_ARK_ARC_1_0/temp1[36] ), .B(
        \MC_ARK_ARC_1_0/temp2[36] ), .ZN(\MC_ARK_ARC_1_0/temp5[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_25_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[72] ), 
        .B(n404), .ZN(\MC_ARK_ARC_1_0/temp4[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_25_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[102] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_25_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[6] ), 
        .B(\RI5[0][174] ), .ZN(\MC_ARK_ARC_1_0/temp2[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_25_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[30] ), .ZN(\MC_ARK_ARC_1_0/temp1[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_25_4  ( .A(\MC_ARK_ARC_1_0/temp5[37] ), .B(
        \MC_ARK_ARC_1_0/temp6[37] ), .ZN(\RI1[1][37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_25_4  ( .A(\MC_ARK_ARC_1_0/temp3[37] ), .B(
        \MC_ARK_ARC_1_0/temp4[37] ), .ZN(\MC_ARK_ARC_1_0/temp6[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_25_4  ( .A(\MC_ARK_ARC_1_0/temp1[37] ), .B(
        \MC_ARK_ARC_1_0/temp2[37] ), .ZN(\MC_ARK_ARC_1_0/temp5[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_25_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .B(n306), .ZN(\MC_ARK_ARC_1_0/temp4[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_25_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_25_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_25_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[37] ), .ZN(\MC_ARK_ARC_1_0/temp1[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_25_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[94] ), .ZN(\MC_ARK_ARC_1_0/temp4[38] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_25_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_25_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_0/temp2[38] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_25_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_0/temp1[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_25_2  ( .A(\MC_ARK_ARC_1_0/temp5[39] ), .B(
        \MC_ARK_ARC_1_0/temp6[39] ), .ZN(\RI1[1][39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_25_2  ( .A(\MC_ARK_ARC_1_0/temp3[39] ), .B(
        \MC_ARK_ARC_1_0/temp4[39] ), .ZN(\MC_ARK_ARC_1_0/temp6[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_25_2  ( .A(\MC_ARK_ARC_1_0/temp1[39] ), .B(
        \MC_ARK_ARC_1_0/temp2[39] ), .ZN(\MC_ARK_ARC_1_0/temp5[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_25_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .B(n438), .ZN(\MC_ARK_ARC_1_0/temp4[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_25_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[141] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_25_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[177] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_0/temp2[39] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_25_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[39] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_0/temp1[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_25_1  ( .A(\MC_ARK_ARC_1_0/temp5[40] ), .B(
        \MC_ARK_ARC_1_0/temp6[40] ), .ZN(\RI1[1][40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_25_1  ( .A(\MC_ARK_ARC_1_0/temp3[40] ), .B(
        \MC_ARK_ARC_1_0/temp4[40] ), .ZN(\MC_ARK_ARC_1_0/temp6[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_25_1  ( .A(\MC_ARK_ARC_1_0/temp2[40] ), .B(
        \MC_ARK_ARC_1_0/temp1[40] ), .ZN(\MC_ARK_ARC_1_0/temp5[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_25_1  ( .A(\RI5[0][76] ), .B(
        \MC_ARK_ARC_1_0/buf_keyinput[40] ), .ZN(\MC_ARK_ARC_1_0/temp4[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_25_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[106] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_25_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[10] ), 
        .B(\RI5[0][178] ), .ZN(\MC_ARK_ARC_1_0/temp2[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_25_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[34] ), .ZN(\MC_ARK_ARC_1_0/temp1[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_25_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .B(n463), .ZN(\MC_ARK_ARC_1_0/temp4[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_25_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[143] ), 
        .B(n1962), .ZN(\MC_ARK_ARC_1_0/temp3[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_25_0  ( .A(n2146), .B(n1660), .ZN(
        \MC_ARK_ARC_1_0/temp2[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_25_0  ( .A(n1483), .B(n1507), .ZN(
        \MC_ARK_ARC_1_0/temp1[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_24_5  ( .A(\MC_ARK_ARC_1_0/temp5[42] ), .B(
        \MC_ARK_ARC_1_0/temp6[42] ), .ZN(\RI1[1][42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_24_5  ( .A(\MC_ARK_ARC_1_0/temp4[42] ), .B(
        \MC_ARK_ARC_1_0/temp3[42] ), .ZN(\MC_ARK_ARC_1_0/temp6[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_24_5  ( .A(\MC_ARK_ARC_1_0/temp1[42] ), .B(
        \MC_ARK_ARC_1_0/temp2[42] ), .ZN(\MC_ARK_ARC_1_0/temp5[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_24_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[78] ), 
        .B(n388), .ZN(\MC_ARK_ARC_1_0/temp4[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_24_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[144] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[108] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_24_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_24_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[36] ), .ZN(\MC_ARK_ARC_1_0/temp1[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_24_4  ( .A(\MC_ARK_ARC_1_0/temp5[43] ), .B(
        \MC_ARK_ARC_1_0/temp6[43] ), .ZN(\RI1[1][43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_24_4  ( .A(\MC_ARK_ARC_1_0/temp3[43] ), .B(
        \MC_ARK_ARC_1_0/temp4[43] ), .ZN(\MC_ARK_ARC_1_0/temp6[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_24_4  ( .A(\MC_ARK_ARC_1_0/temp1[43] ), .B(
        \MC_ARK_ARC_1_0/temp2[43] ), .ZN(\MC_ARK_ARC_1_0/temp5[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_24_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .B(n266), .ZN(\MC_ARK_ARC_1_0/temp4[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_24_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_24_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_24_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[37] ), .ZN(\MC_ARK_ARC_1_0/temp1[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_24_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[80] ), 
        .B(n259), .ZN(\MC_ARK_ARC_1_0/temp4[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_24_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[146] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_24_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[14] ), .ZN(\MC_ARK_ARC_1_0/temp2[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_24_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[38] ), 
        .B(n1475), .ZN(\MC_ARK_ARC_1_0/temp1[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_24_2  ( .A(\MC_ARK_ARC_1_0/temp5[45] ), .B(
        \MC_ARK_ARC_1_0/temp6[45] ), .ZN(\RI1[1][45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_24_2  ( .A(\MC_ARK_ARC_1_0/temp3[45] ), .B(
        \MC_ARK_ARC_1_0/temp4[45] ), .ZN(\MC_ARK_ARC_1_0/temp6[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_24_2  ( .A(\MC_ARK_ARC_1_0/temp2[45] ), .B(
        \MC_ARK_ARC_1_0/temp1[45] ), .ZN(\MC_ARK_ARC_1_0/temp5[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_24_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[81] ), 
        .B(n252), .ZN(\MC_ARK_ARC_1_0/temp4[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_24_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[147] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[111] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_24_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[15] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[183] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_24_2  ( .A(\RI5[0][45] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[39] ), .ZN(\MC_ARK_ARC_1_0/temp1[45] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_24_1  ( .A(\MC_ARK_ARC_1_0/temp5[46] ), .B(
        \MC_ARK_ARC_1_0/temp6[46] ), .ZN(\RI1[1][46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_24_1  ( .A(\MC_ARK_ARC_1_0/temp3[46] ), .B(
        \MC_ARK_ARC_1_0/temp4[46] ), .ZN(\MC_ARK_ARC_1_0/temp6[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_24_1  ( .A(\MC_ARK_ARC_1_0/temp1[46] ), .B(
        \MC_ARK_ARC_1_0/temp2[46] ), .ZN(\MC_ARK_ARC_1_0/temp5[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_24_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[82] ), 
        .B(n510), .ZN(\MC_ARK_ARC_1_0/temp4[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_24_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[148] ), 
        .B(\RI5[0][112] ), .ZN(\MC_ARK_ARC_1_0/temp3[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_24_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[16] ), 
        .B(\RI5[0][184] ), .ZN(\MC_ARK_ARC_1_0/temp2[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_24_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[46] ), .ZN(\MC_ARK_ARC_1_0/temp1[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_24_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[83] ), 
        .B(n461), .ZN(\MC_ARK_ARC_1_0/temp4[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_24_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[149] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_24_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[17] ), 
        .B(n795), .ZN(\MC_ARK_ARC_1_0/temp2[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_24_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[47] ), 
        .B(n1483), .ZN(\MC_ARK_ARC_1_0/temp1[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_23_5  ( .A(\MC_ARK_ARC_1_0/temp5[48] ), .B(
        \MC_ARK_ARC_1_0/temp6[48] ), .ZN(\RI1[1][48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_23_5  ( .A(\MC_ARK_ARC_1_0/temp3[48] ), .B(
        \MC_ARK_ARC_1_0/temp4[48] ), .ZN(\MC_ARK_ARC_1_0/temp6[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_23_5  ( .A(\MC_ARK_ARC_1_0/temp1[48] ), .B(
        \MC_ARK_ARC_1_0/temp2[48] ), .ZN(\MC_ARK_ARC_1_0/temp5[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_23_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .B(n234), .ZN(\MC_ARK_ARC_1_0/temp4[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_23_5  ( .A(\RI5[0][150] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[114] ), .ZN(\MC_ARK_ARC_1_0/temp3[48] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_23_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[186] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_23_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_0/temp1[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_23_4  ( .A(\MC_ARK_ARC_1_0/temp5[49] ), .B(
        \MC_ARK_ARC_1_0/temp6[49] ), .ZN(\RI1[1][49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_23_4  ( .A(\MC_ARK_ARC_1_0/temp3[49] ), .B(
        \MC_ARK_ARC_1_0/temp4[49] ), .ZN(\MC_ARK_ARC_1_0/temp6[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_23_4  ( .A(\MC_ARK_ARC_1_0/temp1[49] ), .B(
        \MC_ARK_ARC_1_0/temp2[49] ), .ZN(\MC_ARK_ARC_1_0/temp5[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_23_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[85] ), 
        .B(n377), .ZN(\MC_ARK_ARC_1_0/temp4[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_23_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_23_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[187] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_23_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[43] ), .ZN(\MC_ARK_ARC_1_0/temp1[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_23_3  ( .A(\MC_ARK_ARC_1_0/temp5[50] ), .B(
        \MC_ARK_ARC_1_0/temp6[50] ), .ZN(\RI1[1][50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_23_3  ( .A(\MC_ARK_ARC_1_0/temp3[50] ), .B(
        \MC_ARK_ARC_1_0/temp4[50] ), .ZN(\MC_ARK_ARC_1_0/temp6[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_23_3  ( .A(\MC_ARK_ARC_1_0/temp2[50] ), .B(
        \MC_ARK_ARC_1_0/temp1[50] ), .ZN(\MC_ARK_ARC_1_0/temp5[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_23_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[179] ), .ZN(\MC_ARK_ARC_1_0/temp4[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_23_3  ( .A(\RI5[0][152] ), .B(n1940), .ZN(
        \MC_ARK_ARC_1_0/temp3[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_23_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_0/temp2[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_23_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[50] ), 
        .B(n1474), .ZN(\MC_ARK_ARC_1_0/temp1[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_23_2  ( .A(\MC_ARK_ARC_1_0/temp5[51] ), .B(
        \MC_ARK_ARC_1_0/temp6[51] ), .ZN(\RI1[1][51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_23_2  ( .A(\MC_ARK_ARC_1_0/temp3[51] ), .B(
        \MC_ARK_ARC_1_0/temp4[51] ), .ZN(\MC_ARK_ARC_1_0/temp6[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_23_2  ( .A(\MC_ARK_ARC_1_0/temp1[51] ), .B(
        \MC_ARK_ARC_1_0/temp2[51] ), .ZN(\MC_ARK_ARC_1_0/temp5[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_23_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[87] ), 
        .B(n213), .ZN(\MC_ARK_ARC_1_0/temp4[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_23_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[153] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[117] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_23_2  ( .A(n1959), .B(
        \MC_ARK_ARC_1_0/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_0/temp2[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_23_2  ( .A(\RI5[0][45] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[51] ), .ZN(\MC_ARK_ARC_1_0/temp1[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_23_1  ( .A(\MC_ARK_ARC_1_0/temp5[52] ), .B(
        \MC_ARK_ARC_1_0/temp6[52] ), .ZN(\RI1[1][52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_23_1  ( .A(\MC_ARK_ARC_1_0/temp3[52] ), .B(
        \MC_ARK_ARC_1_0/temp4[52] ), .ZN(\MC_ARK_ARC_1_0/temp6[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_23_1  ( .A(\MC_ARK_ARC_1_0/temp1[52] ), .B(
        \MC_ARK_ARC_1_0/temp2[52] ), .ZN(\MC_ARK_ARC_1_0/temp5[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_23_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .B(n484), .ZN(\MC_ARK_ARC_1_0/temp4[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_23_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[118] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_23_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_23_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[46] ), .ZN(\MC_ARK_ARC_1_0/temp1[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_23_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[89] ), 
        .B(n474), .ZN(\MC_ARK_ARC_1_0/temp4[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_23_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[119] ), 
        .B(n2117), .ZN(\MC_ARK_ARC_1_0/temp3[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_23_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[191] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[23] ), .ZN(\MC_ARK_ARC_1_0/temp2[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_23_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[47] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[53] ), .ZN(\MC_ARK_ARC_1_0/temp1[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_22_5  ( .A(\MC_ARK_ARC_1_0/temp5[54] ), .B(
        \MC_ARK_ARC_1_0/temp6[54] ), .ZN(\RI1[1][54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_22_5  ( .A(\MC_ARK_ARC_1_0/temp3[54] ), .B(
        \MC_ARK_ARC_1_0/temp4[54] ), .ZN(\MC_ARK_ARC_1_0/temp6[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_22_5  ( .A(\MC_ARK_ARC_1_0/temp1[54] ), .B(
        \MC_ARK_ARC_1_0/temp2[54] ), .ZN(\MC_ARK_ARC_1_0/temp5[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_22_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[90] ), 
        .B(n406), .ZN(\MC_ARK_ARC_1_0/temp4[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_22_5  ( .A(\RI5[0][156] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[120] ), .ZN(\MC_ARK_ARC_1_0/temp3[54] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_22_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_0/temp2[54] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_22_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[48] ), .ZN(\MC_ARK_ARC_1_0/temp1[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_22_4  ( .A(\MC_ARK_ARC_1_0/temp5[55] ), .B(
        \MC_ARK_ARC_1_0/temp6[55] ), .ZN(\RI1[1][55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_22_4  ( .A(\MC_ARK_ARC_1_0/temp3[55] ), .B(
        \MC_ARK_ARC_1_0/temp4[55] ), .ZN(\MC_ARK_ARC_1_0/temp6[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_22_4  ( .A(\MC_ARK_ARC_1_0/temp1[55] ), .B(
        \MC_ARK_ARC_1_0/temp2[55] ), .ZN(\MC_ARK_ARC_1_0/temp5[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_22_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[62] ), .ZN(\MC_ARK_ARC_1_0/temp4[55] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_22_4  ( .A(\RI5[0][157] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[121] ), .ZN(\MC_ARK_ARC_1_0/temp3[55] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_22_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[25] ), 
        .B(\RI5[0][1] ), .ZN(\MC_ARK_ARC_1_0/temp2[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_22_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[49] ), .ZN(\MC_ARK_ARC_1_0/temp1[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_22_3  ( .A(\MC_ARK_ARC_1_0/temp5[56] ), .B(
        \MC_ARK_ARC_1_0/temp6[56] ), .ZN(\RI1[1][56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_22_3  ( .A(\MC_ARK_ARC_1_0/temp3[56] ), .B(
        \MC_ARK_ARC_1_0/temp4[56] ), .ZN(\MC_ARK_ARC_1_0/temp6[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_22_3  ( .A(\MC_ARK_ARC_1_0/temp2[56] ), .B(
        \MC_ARK_ARC_1_0/temp1[56] ), .ZN(\MC_ARK_ARC_1_0/temp5[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_22_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[92] ), 
        .B(Key[13]), .ZN(\MC_ARK_ARC_1_0/temp4[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_22_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[122] ), 
        .B(n2137), .ZN(\MC_ARK_ARC_1_0/temp3[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_22_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[26] ), 
        .B(\RI5[0][2] ), .ZN(\MC_ARK_ARC_1_0/temp2[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_22_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[56] ), .ZN(\MC_ARK_ARC_1_0/temp1[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_22_2  ( .A(\MC_ARK_ARC_1_0/temp5[57] ), .B(
        \MC_ARK_ARC_1_0/temp6[57] ), .ZN(\RI1[1][57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_22_2  ( .A(\MC_ARK_ARC_1_0/temp3[57] ), .B(
        \MC_ARK_ARC_1_0/temp4[57] ), .ZN(\MC_ARK_ARC_1_0/temp6[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_22_2  ( .A(\MC_ARK_ARC_1_0/temp1[57] ), .B(
        \MC_ARK_ARC_1_0/temp2[57] ), .ZN(\MC_ARK_ARC_1_0/temp5[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_22_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[93] ), 
        .B(n478), .ZN(\MC_ARK_ARC_1_0/temp4[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_22_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[159] ), 
        .B(\RI5[0][123] ), .ZN(\MC_ARK_ARC_1_0/temp3[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_22_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[3] ), .ZN(\MC_ARK_ARC_1_0/temp2[57] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_22_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[57] ), .ZN(\MC_ARK_ARC_1_0/temp1[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_22_1  ( .A(\MC_ARK_ARC_1_0/temp5[58] ), .B(
        \MC_ARK_ARC_1_0/temp6[58] ), .ZN(\RI1[1][58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_22_1  ( .A(\MC_ARK_ARC_1_0/temp3[58] ), .B(
        \MC_ARK_ARC_1_0/temp4[58] ), .ZN(\MC_ARK_ARC_1_0/temp6[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_22_1  ( .A(\MC_ARK_ARC_1_0/temp2[58] ), .B(
        \MC_ARK_ARC_1_0/temp1[58] ), .ZN(\MC_ARK_ARC_1_0/temp5[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_22_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[94] ), 
        .B(n348), .ZN(\MC_ARK_ARC_1_0/temp4[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_22_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_22_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[28] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_0/temp2[58] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_22_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[58] ), .ZN(\MC_ARK_ARC_1_0/temp1[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_22_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[95] ), 
        .B(n464), .ZN(\MC_ARK_ARC_1_0/temp4[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_22_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[161] ), 
        .B(n1938), .ZN(\MC_ARK_ARC_1_0/temp3[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_22_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[5] ), 
        .B(n1960), .ZN(\MC_ARK_ARC_1_0/temp2[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_22_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[53] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[59] ), .ZN(\MC_ARK_ARC_1_0/temp1[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_21_5  ( .A(\MC_ARK_ARC_1_0/temp5[60] ), .B(
        \MC_ARK_ARC_1_0/temp6[60] ), .ZN(\RI1[1][60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_21_5  ( .A(\MC_ARK_ARC_1_0/temp3[60] ), .B(
        \MC_ARK_ARC_1_0/temp4[60] ), .ZN(\MC_ARK_ARC_1_0/temp6[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_21_5  ( .A(\MC_ARK_ARC_1_0/temp1[60] ), .B(
        \MC_ARK_ARC_1_0/temp2[60] ), .ZN(\MC_ARK_ARC_1_0/temp5[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_21_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .B(n400), .ZN(\MC_ARK_ARC_1_0/temp4[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_21_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[162] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[126] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_21_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_0/temp2[60] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_21_5  ( .A(\RI5[0][60] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[54] ), .ZN(\MC_ARK_ARC_1_0/temp1[60] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_21_4  ( .A(\MC_ARK_ARC_1_0/temp5[61] ), .B(
        \MC_ARK_ARC_1_0/temp6[61] ), .ZN(\RI1[1][61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_21_4  ( .A(\MC_ARK_ARC_1_0/temp3[61] ), .B(
        \MC_ARK_ARC_1_0/temp4[61] ), .ZN(\MC_ARK_ARC_1_0/temp6[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_21_4  ( .A(\MC_ARK_ARC_1_0/temp1[61] ), .B(
        \MC_ARK_ARC_1_0/temp2[61] ), .ZN(\MC_ARK_ARC_1_0/temp5[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_21_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .B(n329), .ZN(\MC_ARK_ARC_1_0/temp4[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_21_4  ( .A(\RI5[0][163] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[127] ), .ZN(\MC_ARK_ARC_1_0/temp3[61] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_21_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_0/temp2[61] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_21_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[55] ), .ZN(\MC_ARK_ARC_1_0/temp1[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_21_3  ( .A(\MC_ARK_ARC_1_0/temp6[62] ), .B(
        \MC_ARK_ARC_1_0/temp5[62] ), .ZN(\RI1[1][62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_21_3  ( .A(\MC_ARK_ARC_1_0/temp3[62] ), .B(
        \MC_ARK_ARC_1_0/temp4[62] ), .ZN(\MC_ARK_ARC_1_0/temp6[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_21_3  ( .A(\MC_ARK_ARC_1_0/temp1[62] ), .B(
        \MC_ARK_ARC_1_0/temp2[62] ), .ZN(\MC_ARK_ARC_1_0/temp5[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_21_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[98] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[118] ), .ZN(\MC_ARK_ARC_1_0/temp4[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_21_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[164] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_21_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[8] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[32] ), .ZN(\MC_ARK_ARC_1_0/temp2[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_21_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[56] ), 
        .B(\RI5[0][62] ), .ZN(\MC_ARK_ARC_1_0/temp1[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_21_2  ( .A(\MC_ARK_ARC_1_0/temp5[63] ), .B(
        \MC_ARK_ARC_1_0/temp6[63] ), .ZN(\RI1[1][63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_21_2  ( .A(\MC_ARK_ARC_1_0/temp3[63] ), .B(
        \MC_ARK_ARC_1_0/temp4[63] ), .ZN(\MC_ARK_ARC_1_0/temp6[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_21_2  ( .A(\MC_ARK_ARC_1_0/temp2[63] ), .B(
        \MC_ARK_ARC_1_0/temp1[63] ), .ZN(\MC_ARK_ARC_1_0/temp5[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_21_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[99] ), 
        .B(n316), .ZN(\MC_ARK_ARC_1_0/temp4[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_21_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[129] ), 
        .B(\RI5[0][165] ), .ZN(\MC_ARK_ARC_1_0/temp3[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_21_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[9] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_0/temp2[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_21_2  ( .A(\RI5[0][63] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[57] ), .ZN(\MC_ARK_ARC_1_0/temp1[63] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_21_1  ( .A(\MC_ARK_ARC_1_0/temp5[64] ), .B(
        \MC_ARK_ARC_1_0/temp6[64] ), .ZN(\RI1[1][64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_21_1  ( .A(\MC_ARK_ARC_1_0/temp3[64] ), .B(
        \MC_ARK_ARC_1_0/temp4[64] ), .ZN(\MC_ARK_ARC_1_0/temp6[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_21_1  ( .A(\MC_ARK_ARC_1_0/temp2[64] ), .B(
        \MC_ARK_ARC_1_0/temp1[64] ), .ZN(\MC_ARK_ARC_1_0/temp5[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_21_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[100] ), 
        .B(n449), .ZN(\MC_ARK_ARC_1_0/temp4[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_21_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_21_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_0/temp2[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_21_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[58] ), .ZN(\MC_ARK_ARC_1_0/temp1[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_21_0  ( .A(\MC_ARK_ARC_1_0/temp3[65] ), .B(
        \MC_ARK_ARC_1_0/temp4[65] ), .ZN(\MC_ARK_ARC_1_0/temp6[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_21_0  ( .A(\MC_ARK_ARC_1_0/temp1[65] ), .B(
        \MC_ARK_ARC_1_0/temp2[65] ), .ZN(\MC_ARK_ARC_1_0/temp5[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_21_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[101] ), 
        .B(n458), .ZN(\MC_ARK_ARC_1_0/temp4[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_21_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[131] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[167] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_21_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[11] ), 
        .B(n1509), .ZN(\MC_ARK_ARC_1_0/temp2[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_21_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[65] ), 
        .B(n787), .ZN(\MC_ARK_ARC_1_0/temp1[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_20_5  ( .A(\MC_ARK_ARC_1_0/temp3[66] ), .B(
        \MC_ARK_ARC_1_0/temp4[66] ), .ZN(\MC_ARK_ARC_1_0/temp6[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_20_5  ( .A(\MC_ARK_ARC_1_0/temp1[66] ), .B(
        \MC_ARK_ARC_1_0/temp2[66] ), .ZN(\MC_ARK_ARC_1_0/temp5[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_20_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .B(n296), .ZN(\MC_ARK_ARC_1_0/temp4[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_20_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[132] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_20_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_0/temp2[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_20_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[66] ), 
        .B(\RI5[0][60] ), .ZN(\MC_ARK_ARC_1_0/temp1[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_20_4  ( .A(\MC_ARK_ARC_1_0/temp5[67] ), .B(
        \MC_ARK_ARC_1_0/temp6[67] ), .ZN(\RI1[1][67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_20_4  ( .A(\MC_ARK_ARC_1_0/temp3[67] ), .B(
        \MC_ARK_ARC_1_0/temp4[67] ), .ZN(\MC_ARK_ARC_1_0/temp6[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_20_4  ( .A(\MC_ARK_ARC_1_0/temp1[67] ), .B(
        \MC_ARK_ARC_1_0/temp2[67] ), .ZN(\MC_ARK_ARC_1_0/temp5[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_20_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[103] ), 
        .B(Key[90]), .ZN(\MC_ARK_ARC_1_0/temp4[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_20_4  ( .A(\RI5[0][169] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[133] ), .ZN(\MC_ARK_ARC_1_0/temp3[67] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_20_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[37] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[13] ), .ZN(\MC_ARK_ARC_1_0/temp2[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_20_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[61] ), .ZN(\MC_ARK_ARC_1_0/temp1[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_20_3  ( .A(\MC_ARK_ARC_1_0/temp6[68] ), .B(
        \MC_ARK_ARC_1_0/temp5[68] ), .ZN(\RI1[1][68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_20_3  ( .A(\MC_ARK_ARC_1_0/temp3[68] ), .B(
        \MC_ARK_ARC_1_0/temp4[68] ), .ZN(\MC_ARK_ARC_1_0/temp6[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_20_3  ( .A(\MC_ARK_ARC_1_0/temp2[68] ), .B(
        \MC_ARK_ARC_1_0/temp1[68] ), .ZN(\MC_ARK_ARC_1_0/temp5[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_20_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[104] ), 
        .B(n457), .ZN(\MC_ARK_ARC_1_0/temp4[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_20_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[134] ), 
        .B(\RI5[0][170] ), .ZN(\MC_ARK_ARC_1_0/temp3[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_20_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[38] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[14] ), .ZN(\MC_ARK_ARC_1_0/temp2[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_20_3  ( .A(\RI5[0][62] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_0/temp1[68] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_20_2  ( .A(\MC_ARK_ARC_1_0/temp5[69] ), .B(
        \MC_ARK_ARC_1_0/temp6[69] ), .ZN(\RI1[1][69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_20_2  ( .A(\MC_ARK_ARC_1_0/temp3[69] ), .B(
        \MC_ARK_ARC_1_0/temp4[69] ), .ZN(\MC_ARK_ARC_1_0/temp6[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_20_2  ( .A(\MC_ARK_ARC_1_0/temp2[69] ), .B(
        \MC_ARK_ARC_1_0/temp1[69] ), .ZN(\MC_ARK_ARC_1_0/temp5[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_20_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[105] ), 
        .B(n477), .ZN(\MC_ARK_ARC_1_0/temp4[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_20_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[171] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[135] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_20_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[39] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[15] ), .ZN(\MC_ARK_ARC_1_0/temp2[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_20_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[69] ), 
        .B(\RI5[0][63] ), .ZN(\MC_ARK_ARC_1_0/temp1[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_20_1  ( .A(\MC_ARK_ARC_1_0/temp5[70] ), .B(
        \MC_ARK_ARC_1_0/temp6[70] ), .ZN(\RI1[1][70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_20_1  ( .A(\MC_ARK_ARC_1_0/temp3[70] ), .B(
        \MC_ARK_ARC_1_0/temp4[70] ), .ZN(\MC_ARK_ARC_1_0/temp6[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_20_1  ( .A(\MC_ARK_ARC_1_0/temp2[70] ), .B(
        \MC_ARK_ARC_1_0/temp1[70] ), .ZN(\MC_ARK_ARC_1_0/temp5[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_20_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[106] ), 
        .B(n269), .ZN(\MC_ARK_ARC_1_0/temp4[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_20_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[136] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_20_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_0/temp2[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_20_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[64] ), .ZN(\MC_ARK_ARC_1_0/temp1[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_20_0  ( .A(n1962), .B(n439), .ZN(
        \MC_ARK_ARC_1_0/temp4[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_20_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[137] ), 
        .B(n2150), .ZN(\MC_ARK_ARC_1_0/temp3[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_20_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[17] ), 
        .B(n1961), .ZN(\MC_ARK_ARC_1_0/temp2[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_20_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[65] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[71] ), .ZN(\MC_ARK_ARC_1_0/temp1[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_19_5  ( .A(\MC_ARK_ARC_1_0/temp5[72] ), .B(
        \MC_ARK_ARC_1_0/temp6[72] ), .ZN(\RI1[1][72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_19_5  ( .A(\MC_ARK_ARC_1_0/temp3[72] ), .B(
        \MC_ARK_ARC_1_0/temp4[72] ), .ZN(\MC_ARK_ARC_1_0/temp6[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_19_5  ( .A(\MC_ARK_ARC_1_0/temp1[72] ), .B(
        \MC_ARK_ARC_1_0/temp2[72] ), .ZN(\MC_ARK_ARC_1_0/temp5[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_19_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[108] ), 
        .B(n255), .ZN(\MC_ARK_ARC_1_0/temp4[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_19_5  ( .A(\RI5[0][174] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[138] ), .ZN(\MC_ARK_ARC_1_0/temp3[72] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_19_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[18] ), .ZN(\MC_ARK_ARC_1_0/temp2[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_19_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[66] ), .ZN(\MC_ARK_ARC_1_0/temp1[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_19_4  ( .A(\MC_ARK_ARC_1_0/temp5[73] ), .B(
        \MC_ARK_ARC_1_0/temp6[73] ), .ZN(\RI1[1][73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_19_4  ( .A(\MC_ARK_ARC_1_0/temp3[73] ), .B(
        \MC_ARK_ARC_1_0/temp4[73] ), .ZN(\MC_ARK_ARC_1_0/temp6[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_19_4  ( .A(\MC_ARK_ARC_1_0/temp1[73] ), .B(
        \MC_ARK_ARC_1_0/temp2[73] ), .ZN(\MC_ARK_ARC_1_0/temp5[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_19_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[109] ), 
        .B(n249), .ZN(\MC_ARK_ARC_1_0/temp4[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_19_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[139] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_19_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[19] ), .ZN(\MC_ARK_ARC_1_0/temp2[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_19_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[67] ), .ZN(\MC_ARK_ARC_1_0/temp1[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_19_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[110] ), 
        .B(Key[139]), .ZN(\MC_ARK_ARC_1_0/temp4[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_19_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[140] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_19_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[20] ), 
        .B(n1474), .ZN(\MC_ARK_ARC_1_0/temp2[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_19_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_0/temp1[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_19_2  ( .A(\MC_ARK_ARC_1_0/temp5[75] ), .B(
        \MC_ARK_ARC_1_0/temp6[75] ), .ZN(\RI1[1][75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_19_2  ( .A(\MC_ARK_ARC_1_0/temp3[75] ), .B(
        \MC_ARK_ARC_1_0/temp4[75] ), .ZN(\MC_ARK_ARC_1_0/temp6[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_19_2  ( .A(\MC_ARK_ARC_1_0/temp1[75] ), .B(
        \MC_ARK_ARC_1_0/temp2[75] ), .ZN(\MC_ARK_ARC_1_0/temp5[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_19_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[111] ), 
        .B(n476), .ZN(\MC_ARK_ARC_1_0/temp4[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_19_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[177] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_19_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[21] ), 
        .B(\RI5[0][45] ), .ZN(\MC_ARK_ARC_1_0/temp2[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_19_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[69] ), .ZN(\MC_ARK_ARC_1_0/temp1[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_19_1  ( .A(\MC_ARK_ARC_1_0/temp5[76] ), .B(
        \MC_ARK_ARC_1_0/temp6[76] ), .ZN(\RI1[1][76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_19_1  ( .A(\MC_ARK_ARC_1_0/temp3[76] ), .B(
        \MC_ARK_ARC_1_0/temp4[76] ), .ZN(\MC_ARK_ARC_1_0/temp6[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_19_1  ( .A(\MC_ARK_ARC_1_0/temp1[76] ), .B(
        \MC_ARK_ARC_1_0/temp2[76] ), .ZN(\MC_ARK_ARC_1_0/temp5[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_19_1  ( .A(\RI5[0][112] ), .B(n230), .ZN(
        \MC_ARK_ARC_1_0/temp4[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_19_1  ( .A(\RI5[0][178] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[142] ), .ZN(\MC_ARK_ARC_1_0/temp3[76] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_19_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[22] ), .ZN(\MC_ARK_ARC_1_0/temp2[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_19_1  ( .A(\RI5[0][76] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_0/temp1[76] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_19_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .B(n223), .ZN(\MC_ARK_ARC_1_0/temp4[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_19_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[143] ), 
        .B(n1659), .ZN(\MC_ARK_ARC_1_0/temp3[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_19_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[47] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[23] ), .ZN(\MC_ARK_ARC_1_0/temp2[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_19_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[77] ), .ZN(\MC_ARK_ARC_1_0/temp1[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_18_5  ( .A(\MC_ARK_ARC_1_0/temp5[78] ), .B(
        \MC_ARK_ARC_1_0/temp6[78] ), .ZN(\RI1[1][78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_18_5  ( .A(\MC_ARK_ARC_1_0/temp3[78] ), .B(
        \MC_ARK_ARC_1_0/temp4[78] ), .ZN(\MC_ARK_ARC_1_0/temp6[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_18_5  ( .A(\MC_ARK_ARC_1_0/temp1[78] ), .B(
        \MC_ARK_ARC_1_0/temp2[78] ), .ZN(\MC_ARK_ARC_1_0/temp5[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_18_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[114] ), 
        .B(n216), .ZN(\MC_ARK_ARC_1_0/temp4[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_18_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[144] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_18_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[24] ), .ZN(\MC_ARK_ARC_1_0/temp2[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_18_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[72] ), .ZN(\MC_ARK_ARC_1_0/temp1[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_18_4  ( .A(\MC_ARK_ARC_1_0/temp6[79] ), .B(
        \MC_ARK_ARC_1_0/temp5[79] ), .ZN(\RI1[1][79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_18_4  ( .A(\MC_ARK_ARC_1_0/temp4[79] ), .B(
        \MC_ARK_ARC_1_0/temp3[79] ), .ZN(\MC_ARK_ARC_1_0/temp6[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_18_4  ( .A(\MC_ARK_ARC_1_0/temp1[79] ), .B(
        \MC_ARK_ARC_1_0/temp2[79] ), .ZN(\MC_ARK_ARC_1_0/temp5[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_18_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[87] ), .ZN(\MC_ARK_ARC_1_0/temp4[79] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_18_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[145] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_18_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[25] ), .ZN(\MC_ARK_ARC_1_0/temp2[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_18_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[73] ), .ZN(\MC_ARK_ARC_1_0/temp1[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_18_3  ( .A(\MC_ARK_ARC_1_0/temp5[80] ), .B(
        \MC_ARK_ARC_1_0/temp6[80] ), .ZN(\RI1[1][80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_18_3  ( .A(\MC_ARK_ARC_1_0/temp3[80] ), .B(
        \MC_ARK_ARC_1_0/temp4[80] ), .ZN(\MC_ARK_ARC_1_0/temp6[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_18_3  ( .A(\MC_ARK_ARC_1_0/temp2[80] ), .B(
        \MC_ARK_ARC_1_0/temp1[80] ), .ZN(\MC_ARK_ARC_1_0/temp5[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_18_3  ( .A(n1940), .B(
        \MC_ARK_ARC_1_0/buf_keyinput[80] ), .ZN(\MC_ARK_ARC_1_0/temp4[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_18_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[146] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_18_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[50] ), .ZN(\MC_ARK_ARC_1_0/temp2[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_18_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[80] ), .ZN(\MC_ARK_ARC_1_0/temp1[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_18_2  ( .A(\MC_ARK_ARC_1_0/temp6[81] ), .B(
        \MC_ARK_ARC_1_0/temp5[81] ), .ZN(\RI1[1][81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_18_2  ( .A(\MC_ARK_ARC_1_0/temp3[81] ), .B(
        \MC_ARK_ARC_1_0/temp4[81] ), .ZN(\MC_ARK_ARC_1_0/temp6[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_18_2  ( .A(\MC_ARK_ARC_1_0/temp1[81] ), .B(
        \MC_ARK_ARC_1_0/temp2[81] ), .ZN(\MC_ARK_ARC_1_0/temp5[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_18_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[117] ), 
        .B(n498), .ZN(\MC_ARK_ARC_1_0/temp4[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_18_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[183] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[147] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_18_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[27] ), .ZN(\MC_ARK_ARC_1_0/temp2[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_18_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[81] ), .ZN(\MC_ARK_ARC_1_0/temp1[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_18_1  ( .A(\MC_ARK_ARC_1_0/temp5[82] ), .B(
        \MC_ARK_ARC_1_0/temp6[82] ), .ZN(\RI1[1][82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_18_1  ( .A(\MC_ARK_ARC_1_0/temp3[82] ), .B(
        \MC_ARK_ARC_1_0/temp4[82] ), .ZN(\MC_ARK_ARC_1_0/temp6[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_18_1  ( .A(\MC_ARK_ARC_1_0/temp1[82] ), .B(
        \MC_ARK_ARC_1_0/temp2[82] ), .ZN(\MC_ARK_ARC_1_0/temp5[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_18_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[118] ), 
        .B(n473), .ZN(\MC_ARK_ARC_1_0/temp4[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_18_1  ( .A(\RI5[0][184] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[148] ), .ZN(\MC_ARK_ARC_1_0/temp3[82] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_18_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[28] ), .ZN(\MC_ARK_ARC_1_0/temp2[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_18_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[82] ), 
        .B(\RI5[0][76] ), .ZN(\MC_ARK_ARC_1_0/temp1[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_18_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[119] ), 
        .B(n456), .ZN(\MC_ARK_ARC_1_0/temp4[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_18_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[149] ), 
        .B(n794), .ZN(\MC_ARK_ARC_1_0/temp3[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_18_0  ( .A(n1960), .B(n1632), .ZN(
        \MC_ARK_ARC_1_0/temp2[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_18_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[83] ), .ZN(\MC_ARK_ARC_1_0/temp1[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_17_5  ( .A(\MC_ARK_ARC_1_0/temp5[84] ), .B(
        \MC_ARK_ARC_1_0/temp6[84] ), .ZN(\RI1[1][84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_17_5  ( .A(\MC_ARK_ARC_1_0/temp3[84] ), .B(
        \MC_ARK_ARC_1_0/temp4[84] ), .ZN(\MC_ARK_ARC_1_0/temp6[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_17_5  ( .A(\MC_ARK_ARC_1_0/temp1[84] ), .B(
        \MC_ARK_ARC_1_0/temp2[84] ), .ZN(\MC_ARK_ARC_1_0/temp5[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_17_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[120] ), 
        .B(n358), .ZN(\MC_ARK_ARC_1_0/temp4[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_17_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[186] ), 
        .B(\RI5[0][150] ), .ZN(\MC_ARK_ARC_1_0/temp3[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_17_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[30] ), .ZN(\MC_ARK_ARC_1_0/temp2[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_17_4  ( .A(\MC_ARK_ARC_1_0/temp5[85] ), .B(
        \MC_ARK_ARC_1_0/temp6[85] ), .ZN(\RI1[1][85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_17_4  ( .A(\MC_ARK_ARC_1_0/temp3[85] ), .B(
        \MC_ARK_ARC_1_0/temp4[85] ), .ZN(\MC_ARK_ARC_1_0/temp6[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_17_4  ( .A(\MC_ARK_ARC_1_0/temp1[85] ), .B(
        \MC_ARK_ARC_1_0/temp2[85] ), .ZN(\MC_ARK_ARC_1_0/temp5[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_17_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[121] ), 
        .B(n351), .ZN(\MC_ARK_ARC_1_0/temp4[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_17_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[187] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[151] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_17_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[31] ), .ZN(\MC_ARK_ARC_1_0/temp2[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_17_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[79] ), .ZN(\MC_ARK_ARC_1_0/temp1[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_17_3  ( .A(\MC_ARK_ARC_1_0/temp5[86] ), .B(
        \MC_ARK_ARC_1_0/temp6[86] ), .ZN(\RI1[1][86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_17_3  ( .A(\MC_ARK_ARC_1_0/temp3[86] ), .B(
        \MC_ARK_ARC_1_0/temp4[86] ), .ZN(\MC_ARK_ARC_1_0/temp6[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_17_3  ( .A(\MC_ARK_ARC_1_0/temp2[86] ), .B(
        \MC_ARK_ARC_1_0/temp1[86] ), .ZN(\MC_ARK_ARC_1_0/temp5[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_17_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[122] ), 
        .B(n344), .ZN(\MC_ARK_ARC_1_0/temp4[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_17_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[188] ), 
        .B(\RI5[0][152] ), .ZN(\MC_ARK_ARC_1_0/temp3[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_17_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[56] ), .ZN(\MC_ARK_ARC_1_0/temp2[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_17_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[80] ), .ZN(\MC_ARK_ARC_1_0/temp1[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_17_2  ( .A(\MC_ARK_ARC_1_0/temp5[87] ), .B(
        \MC_ARK_ARC_1_0/temp6[87] ), .ZN(\RI1[1][87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_17_2  ( .A(\MC_ARK_ARC_1_0/temp3[87] ), .B(
        \MC_ARK_ARC_1_0/temp4[87] ), .ZN(\MC_ARK_ARC_1_0/temp6[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_17_2  ( .A(\MC_ARK_ARC_1_0/temp2[87] ), .B(
        \MC_ARK_ARC_1_0/temp1[87] ), .ZN(\MC_ARK_ARC_1_0/temp5[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_17_2  ( .A(\RI5[0][123] ), .B(n480), .ZN(
        \MC_ARK_ARC_1_0/temp4[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_17_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[153] ), 
        .B(n1495), .ZN(\MC_ARK_ARC_1_0/temp3[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_17_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[57] ), .ZN(\MC_ARK_ARC_1_0/temp2[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_17_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[87] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[81] ), .ZN(\MC_ARK_ARC_1_0/temp1[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_17_1  ( .A(\MC_ARK_ARC_1_0/temp5[88] ), .B(
        \MC_ARK_ARC_1_0/temp6[88] ), .ZN(\RI1[1][88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_17_1  ( .A(\MC_ARK_ARC_1_0/temp3[88] ), .B(
        \MC_ARK_ARC_1_0/temp4[88] ), .ZN(\MC_ARK_ARC_1_0/temp6[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_17_1  ( .A(\MC_ARK_ARC_1_0/temp2[88] ), .B(
        \MC_ARK_ARC_1_0/temp1[88] ), .ZN(\MC_ARK_ARC_1_0/temp5[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_17_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[124] ), 
        .B(n332), .ZN(\MC_ARK_ARC_1_0/temp4[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_17_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_17_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[34] ), .ZN(\MC_ARK_ARC_1_0/temp2[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_17_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[82] ), .ZN(\MC_ARK_ARC_1_0/temp1[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_17_0  ( .A(n1939), .B(n325), .ZN(
        \MC_ARK_ARC_1_0/temp4[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_17_0  ( .A(n2116), .B(
        \MC_ARK_ARC_1_0/buf_datainput[191] ), .ZN(\MC_ARK_ARC_1_0/temp3[89] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_17_0  ( .A(n1508), .B(
        \MC_ARK_ARC_1_0/buf_datainput[59] ), .ZN(\MC_ARK_ARC_1_0/temp2[89] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_17_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[89] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[83] ), .ZN(\MC_ARK_ARC_1_0/temp1[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_16_5  ( .A(\MC_ARK_ARC_1_0/temp6[90] ), .B(
        \MC_ARK_ARC_1_0/temp5[90] ), .ZN(\RI1[1][90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_16_5  ( .A(\MC_ARK_ARC_1_0/temp3[90] ), .B(
        \MC_ARK_ARC_1_0/temp4[90] ), .ZN(\MC_ARK_ARC_1_0/temp6[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_16_5  ( .A(\MC_ARK_ARC_1_0/temp1[90] ), .B(
        \MC_ARK_ARC_1_0/temp2[90] ), .ZN(\MC_ARK_ARC_1_0/temp5[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_16_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[126] ), 
        .B(n394), .ZN(\MC_ARK_ARC_1_0/temp4[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_16_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[0] ), 
        .B(\RI5[0][156] ), .ZN(\MC_ARK_ARC_1_0/temp3[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_16_5  ( .A(\RI5[0][60] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[36] ), .ZN(\MC_ARK_ARC_1_0/temp2[90] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_16_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[84] ), .ZN(\MC_ARK_ARC_1_0/temp1[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_16_4  ( .A(\MC_ARK_ARC_1_0/temp5[91] ), .B(
        \MC_ARK_ARC_1_0/temp6[91] ), .ZN(\RI1[1][91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_16_4  ( .A(\MC_ARK_ARC_1_0/temp3[91] ), .B(
        \MC_ARK_ARC_1_0/temp4[91] ), .ZN(\MC_ARK_ARC_1_0/temp6[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_16_4  ( .A(\MC_ARK_ARC_1_0/temp1[91] ), .B(
        \MC_ARK_ARC_1_0/temp2[91] ), .ZN(\MC_ARK_ARC_1_0/temp5[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_16_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[127] ), 
        .B(n428), .ZN(\MC_ARK_ARC_1_0/temp4[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_16_4  ( .A(\RI5[0][1] ), .B(\RI5[0][157] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_16_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[37] ), .ZN(\MC_ARK_ARC_1_0/temp2[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_16_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_0/temp1[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_16_3  ( .A(\MC_ARK_ARC_1_0/temp3[92] ), .B(
        \MC_ARK_ARC_1_0/temp4[92] ), .ZN(\MC_ARK_ARC_1_0/temp6[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_16_3  ( .A(\MC_ARK_ARC_1_0/temp1[92] ), .B(
        \MC_ARK_ARC_1_0/temp2[92] ), .ZN(\MC_ARK_ARC_1_0/temp5[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_16_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[89] ), .ZN(\MC_ARK_ARC_1_0/temp4[92] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_16_3  ( .A(n2137), .B(\RI5[0][2] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_16_3  ( .A(\RI5[0][62] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_0/temp2[92] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_16_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[92] ), .ZN(\MC_ARK_ARC_1_0/temp1[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_16_2  ( .A(\MC_ARK_ARC_1_0/temp5[93] ), .B(
        \MC_ARK_ARC_1_0/temp6[93] ), .ZN(\RI1[1][93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_16_2  ( .A(\MC_ARK_ARC_1_0/temp3[93] ), .B(
        \MC_ARK_ARC_1_0/temp4[93] ), .ZN(\MC_ARK_ARC_1_0/temp6[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_16_2  ( .A(\MC_ARK_ARC_1_0/temp2[93] ), .B(
        \MC_ARK_ARC_1_0/temp1[93] ), .ZN(\MC_ARK_ARC_1_0/temp5[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_16_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[129] ), 
        .B(n512), .ZN(\MC_ARK_ARC_1_0/temp4[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_16_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[159] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[3] ), .ZN(\MC_ARK_ARC_1_0/temp3[93] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_16_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[39] ), 
        .B(\RI5[0][63] ), .ZN(\MC_ARK_ARC_1_0/temp2[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_16_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[93] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[87] ), .ZN(\MC_ARK_ARC_1_0/temp1[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_16_1  ( .A(\MC_ARK_ARC_1_0/temp5[94] ), .B(
        \MC_ARK_ARC_1_0/temp6[94] ), .ZN(\RI1[1][94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_16_1  ( .A(\MC_ARK_ARC_1_0/temp3[94] ), .B(
        \MC_ARK_ARC_1_0/temp4[94] ), .ZN(\MC_ARK_ARC_1_0/temp6[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_16_1  ( .A(\MC_ARK_ARC_1_0/temp2[94] ), .B(
        \MC_ARK_ARC_1_0/temp1[94] ), .ZN(\MC_ARK_ARC_1_0/temp5[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_16_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[130] ), 
        .B(n450), .ZN(\MC_ARK_ARC_1_0/temp4[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_16_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_16_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[64] ), .ZN(\MC_ARK_ARC_1_0/temp2[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_16_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_0/temp1[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_16_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[131] ), 
        .B(\MC_ARK_ARC_1_0/buf_keyinput[95] ), .ZN(\MC_ARK_ARC_1_0/temp4[95] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_16_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[5] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[161] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_16_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[65] ), 
        .B(n1961), .ZN(\MC_ARK_ARC_1_0/temp2[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_16_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[89] ), 
        .B(n875), .ZN(\MC_ARK_ARC_1_0/temp1[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_15_5  ( .A(\MC_ARK_ARC_1_0/temp5[96] ), .B(
        \MC_ARK_ARC_1_0/temp6[96] ), .ZN(\RI1[1][96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_15_5  ( .A(\MC_ARK_ARC_1_0/temp3[96] ), .B(
        \MC_ARK_ARC_1_0/temp4[96] ), .ZN(\MC_ARK_ARC_1_0/temp6[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_15_5  ( .A(\MC_ARK_ARC_1_0/temp1[96] ), .B(
        \MC_ARK_ARC_1_0/temp2[96] ), .ZN(\MC_ARK_ARC_1_0/temp5[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_15_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .B(n494), .ZN(\MC_ARK_ARC_1_0/temp4[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_15_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_15_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_0/temp2[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_15_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[90] ), .ZN(\MC_ARK_ARC_1_0/temp1[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_15_4  ( .A(\MC_ARK_ARC_1_0/temp5[97] ), .B(
        \MC_ARK_ARC_1_0/temp6[97] ), .ZN(\RI1[1][97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_15_4  ( .A(\MC_ARK_ARC_1_0/temp3[97] ), .B(
        \MC_ARK_ARC_1_0/temp4[97] ), .ZN(\MC_ARK_ARC_1_0/temp6[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_15_4  ( .A(\MC_ARK_ARC_1_0/temp1[97] ), .B(
        \MC_ARK_ARC_1_0/temp2[97] ), .ZN(\MC_ARK_ARC_1_0/temp5[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_15_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[133] ), 
        .B(n272), .ZN(\MC_ARK_ARC_1_0/temp4[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_15_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .B(\RI5[0][163] ), .ZN(\MC_ARK_ARC_1_0/temp3[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_15_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[43] ), .ZN(\MC_ARK_ARC_1_0/temp2[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_15_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_0/temp1[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_15_3  ( .A(\MC_ARK_ARC_1_0/temp6[98] ), .B(
        \MC_ARK_ARC_1_0/temp5[98] ), .ZN(\RI1[1][98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_15_3  ( .A(\MC_ARK_ARC_1_0/temp3[98] ), .B(
        \MC_ARK_ARC_1_0/temp4[98] ), .ZN(\MC_ARK_ARC_1_0/temp6[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_15_3  ( .A(\MC_ARK_ARC_1_0/temp2[98] ), .B(
        \MC_ARK_ARC_1_0/temp1[98] ), .ZN(\MC_ARK_ARC_1_0/temp5[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_15_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[134] ), 
        .B(n265), .ZN(\MC_ARK_ARC_1_0/temp4[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_15_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[164] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_0/temp3[98] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_15_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[68] ), 
        .B(n1474), .ZN(\MC_ARK_ARC_1_0/temp2[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_15_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[98] ), .ZN(\MC_ARK_ARC_1_0/temp1[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_15_2  ( .A(\MC_ARK_ARC_1_0/temp5[99] ), .B(
        \MC_ARK_ARC_1_0/temp6[99] ), .ZN(\RI1[1][99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_15_2  ( .A(\MC_ARK_ARC_1_0/temp3[99] ), .B(
        \MC_ARK_ARC_1_0/temp4[99] ), .ZN(\MC_ARK_ARC_1_0/temp6[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_15_2  ( .A(\MC_ARK_ARC_1_0/temp2[99] ), .B(
        \MC_ARK_ARC_1_0/temp1[99] ), .ZN(\MC_ARK_ARC_1_0/temp5[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_15_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[135] ), 
        .B(n258), .ZN(\MC_ARK_ARC_1_0/temp4[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_15_2  ( .A(\RI5[0][165] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_0/temp3[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_15_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[69] ), 
        .B(\RI5[0][45] ), .ZN(\MC_ARK_ARC_1_0/temp2[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_15_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[93] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[99] ), .ZN(\MC_ARK_ARC_1_0/temp1[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_15_1  ( .A(\MC_ARK_ARC_1_0/temp5[100] ), .B(
        \MC_ARK_ARC_1_0/temp6[100] ), .ZN(\RI1[1][100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_15_1  ( .A(\MC_ARK_ARC_1_0/temp3[100] ), .B(
        \MC_ARK_ARC_1_0/temp4[100] ), .ZN(\MC_ARK_ARC_1_0/temp6[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_15_1  ( .A(\MC_ARK_ARC_1_0/temp2[100] ), .B(
        \MC_ARK_ARC_1_0/temp1[100] ), .ZN(\MC_ARK_ARC_1_0/temp5[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_15_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[136] ), 
        .B(n419), .ZN(\MC_ARK_ARC_1_0/temp4[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_15_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_15_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[46] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_15_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[94] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_15_0  ( .A(\MC_ARK_ARC_1_0/temp3[101] ), .B(
        \MC_ARK_ARC_1_0/temp4[101] ), .ZN(\MC_ARK_ARC_1_0/temp6[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_15_0  ( .A(\MC_ARK_ARC_1_0/temp2[101] ), .B(
        \MC_ARK_ARC_1_0/temp1[101] ), .ZN(\MC_ARK_ARC_1_0/temp5[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_15_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[137] ), 
        .B(n245), .ZN(\MC_ARK_ARC_1_0/temp4[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_15_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .B(n2147), .ZN(\MC_ARK_ARC_1_0/temp3[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_15_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[47] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_15_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[101] ), 
        .B(n874), .ZN(\MC_ARK_ARC_1_0/temp1[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_14_5  ( .A(\MC_ARK_ARC_1_0/temp5[102] ), .B(
        \MC_ARK_ARC_1_0/temp6[102] ), .ZN(\RI1[1][102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_14_5  ( .A(\MC_ARK_ARC_1_0/temp3[102] ), .B(
        \MC_ARK_ARC_1_0/temp4[102] ), .ZN(\MC_ARK_ARC_1_0/temp6[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_14_5  ( .A(\MC_ARK_ARC_1_0/temp1[102] ), .B(
        \MC_ARK_ARC_1_0/temp2[102] ), .ZN(\MC_ARK_ARC_1_0/temp5[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_14_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .B(n395), .ZN(\MC_ARK_ARC_1_0/temp4[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_14_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_14_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[48] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_14_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[96] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_14_4  ( .A(\MC_ARK_ARC_1_0/temp5[103] ), .B(
        \MC_ARK_ARC_1_0/temp6[103] ), .ZN(\RI1[1][103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_14_4  ( .A(\MC_ARK_ARC_1_0/temp3[103] ), .B(
        \MC_ARK_ARC_1_0/temp4[103] ), .ZN(\MC_ARK_ARC_1_0/temp6[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_14_4  ( .A(\MC_ARK_ARC_1_0/temp1[103] ), .B(
        \MC_ARK_ARC_1_0/temp2[103] ), .ZN(\MC_ARK_ARC_1_0/temp5[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_14_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[70] ), .ZN(\MC_ARK_ARC_1_0/temp4[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_14_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[13] ), 
        .B(\RI5[0][169] ), .ZN(\MC_ARK_ARC_1_0/temp3[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_14_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[49] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_14_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[97] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_14_3  ( .A(\MC_ARK_ARC_1_0/temp6[104] ), .B(
        \MC_ARK_ARC_1_0/temp5[104] ), .ZN(\RI1[1][104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_14_3  ( .A(\MC_ARK_ARC_1_0/temp3[104] ), .B(
        \MC_ARK_ARC_1_0/temp4[104] ), .ZN(\MC_ARK_ARC_1_0/temp6[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_14_3  ( .A(\MC_ARK_ARC_1_0/temp2[104] ), .B(
        \MC_ARK_ARC_1_0/temp1[104] ), .ZN(\MC_ARK_ARC_1_0/temp5[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_14_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[173] ), .ZN(
        \MC_ARK_ARC_1_0/temp4[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_14_3  ( .A(\RI5[0][170] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[14] ), .ZN(\MC_ARK_ARC_1_0/temp3[104] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_14_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[50] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_14_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[104] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[98] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_14_2  ( .A(\MC_ARK_ARC_1_0/temp5[105] ), .B(
        \MC_ARK_ARC_1_0/temp6[105] ), .ZN(\RI1[1][105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_14_2  ( .A(\MC_ARK_ARC_1_0/temp3[105] ), .B(
        \MC_ARK_ARC_1_0/temp4[105] ), .ZN(\MC_ARK_ARC_1_0/temp6[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_14_2  ( .A(\MC_ARK_ARC_1_0/temp2[105] ), .B(
        \MC_ARK_ARC_1_0/temp1[105] ), .ZN(\MC_ARK_ARC_1_0/temp5[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_14_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .B(n219), .ZN(\MC_ARK_ARC_1_0/temp4[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_14_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[171] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[15] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_14_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[51] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_14_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[99] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_14_1  ( .A(\MC_ARK_ARC_1_0/temp5[106] ), .B(
        \MC_ARK_ARC_1_0/temp6[106] ), .ZN(\RI1[1][106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_14_1  ( .A(\MC_ARK_ARC_1_0/temp3[106] ), .B(
        \MC_ARK_ARC_1_0/temp4[106] ), .ZN(\MC_ARK_ARC_1_0/temp6[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_14_1  ( .A(\MC_ARK_ARC_1_0/temp1[106] ), .B(
        \MC_ARK_ARC_1_0/temp2[106] ), .ZN(\MC_ARK_ARC_1_0/temp5[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_14_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[142] ), 
        .B(n483), .ZN(\MC_ARK_ARC_1_0/temp4[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_14_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_14_1  ( .A(\RI5[0][76] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[52] ), .ZN(\MC_ARK_ARC_1_0/temp2[106] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_14_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_14_0  ( .A(\MC_ARK_ARC_1_0/temp3[107] ), .B(
        \MC_ARK_ARC_1_0/temp4[107] ), .ZN(\MC_ARK_ARC_1_0/temp6[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_14_0  ( .A(\MC_ARK_ARC_1_0/temp1[107] ), .B(
        \MC_ARK_ARC_1_0/temp2[107] ), .ZN(\MC_ARK_ARC_1_0/temp5[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_14_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[143] ), 
        .B(n205), .ZN(\MC_ARK_ARC_1_0/temp4[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_14_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[17] ), 
        .B(n2151), .ZN(\MC_ARK_ARC_1_0/temp3[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_14_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .B(n1631), .ZN(\MC_ARK_ARC_1_0/temp2[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_14_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[101] ), 
        .B(n1480), .ZN(\MC_ARK_ARC_1_0/temp1[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_13_5  ( .A(\MC_ARK_ARC_1_0/temp5[108] ), .B(
        \MC_ARK_ARC_1_0/temp6[108] ), .ZN(\RI1[1][108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_13_5  ( .A(\MC_ARK_ARC_1_0/temp3[108] ), .B(
        \MC_ARK_ARC_1_0/temp4[108] ), .ZN(\MC_ARK_ARC_1_0/temp6[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_13_5  ( .A(\MC_ARK_ARC_1_0/temp1[108] ), .B(
        \MC_ARK_ARC_1_0/temp2[108] ), .ZN(\MC_ARK_ARC_1_0/temp5[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_13_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[144] ), 
        .B(n454), .ZN(\MC_ARK_ARC_1_0/temp4[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_13_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[18] ), 
        .B(\RI5[0][174] ), .ZN(\MC_ARK_ARC_1_0/temp3[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_13_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[54] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_13_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[108] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[102] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_13_4  ( .A(\MC_ARK_ARC_1_0/temp5[109] ), .B(
        \MC_ARK_ARC_1_0/temp6[109] ), .ZN(\RI1[1][109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_13_4  ( .A(\MC_ARK_ARC_1_0/temp3[109] ), .B(
        \MC_ARK_ARC_1_0/temp4[109] ), .ZN(\MC_ARK_ARC_1_0/temp6[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_13_4  ( .A(\MC_ARK_ARC_1_0/temp1[109] ), .B(
        \MC_ARK_ARC_1_0/temp2[109] ), .ZN(\MC_ARK_ARC_1_0/temp5[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_13_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[152] ), .ZN(
        \MC_ARK_ARC_1_0/temp4[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_13_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_13_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[55] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_13_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_13_3  ( .A(\MC_ARK_ARC_1_0/temp6[110] ), .B(
        \MC_ARK_ARC_1_0/temp5[110] ), .ZN(\RI1[1][110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_13_3  ( .A(\MC_ARK_ARC_1_0/temp3[110] ), .B(
        \MC_ARK_ARC_1_0/temp4[110] ), .ZN(\MC_ARK_ARC_1_0/temp6[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_13_3  ( .A(\MC_ARK_ARC_1_0/temp1[110] ), .B(
        \MC_ARK_ARC_1_0/temp2[110] ), .ZN(\MC_ARK_ARC_1_0/temp5[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_13_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[146] ), 
        .B(n468), .ZN(\MC_ARK_ARC_1_0/temp4[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_13_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[20] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_13_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[56] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[80] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_13_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_13_2  ( .A(\MC_ARK_ARC_1_0/temp6[111] ), .B(
        \MC_ARK_ARC_1_0/temp5[111] ), .ZN(\RI1[1][111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_13_2  ( .A(\MC_ARK_ARC_1_0/temp3[111] ), .B(
        \MC_ARK_ARC_1_0/temp4[111] ), .ZN(\MC_ARK_ARC_1_0/temp6[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_13_2  ( .A(\MC_ARK_ARC_1_0/temp1[111] ), .B(
        \MC_ARK_ARC_1_0/temp2[111] ), .ZN(\MC_ARK_ARC_1_0/temp5[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_13_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[147] ), 
        .B(n361), .ZN(\MC_ARK_ARC_1_0/temp4[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_13_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[177] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[21] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_13_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[81] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[57] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_13_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[111] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[105] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_13_1  ( .A(\MC_ARK_ARC_1_0/temp5[112] ), .B(
        \MC_ARK_ARC_1_0/temp6[112] ), .ZN(\RI1[1][112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_13_1  ( .A(\MC_ARK_ARC_1_0/temp3[112] ), .B(
        \MC_ARK_ARC_1_0/temp4[112] ), .ZN(\MC_ARK_ARC_1_0/temp6[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_13_1  ( .A(\MC_ARK_ARC_1_0/temp2[112] ), .B(
        \MC_ARK_ARC_1_0/temp1[112] ), .ZN(\MC_ARK_ARC_1_0/temp5[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_13_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[148] ), 
        .B(n354), .ZN(\MC_ARK_ARC_1_0/temp4[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_13_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .B(\RI5[0][178] ), .ZN(\MC_ARK_ARC_1_0/temp3[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_13_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[58] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_13_1  ( .A(\RI5[0][112] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[106] ), .ZN(\MC_ARK_ARC_1_0/temp1[112] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_13_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[149] ), 
        .B(n448), .ZN(\MC_ARK_ARC_1_0/temp4[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_13_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[23] ), 
        .B(n1659), .ZN(\MC_ARK_ARC_1_0/temp3[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_13_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[83] ), 
        .B(n788), .ZN(\MC_ARK_ARC_1_0/temp2[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_13_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .B(n1480), .ZN(\MC_ARK_ARC_1_0/temp1[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_12_5  ( .A(\MC_ARK_ARC_1_0/temp5[114] ), .B(
        \MC_ARK_ARC_1_0/temp6[114] ), .ZN(\RI1[1][114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_12_5  ( .A(\MC_ARK_ARC_1_0/temp3[114] ), .B(
        \MC_ARK_ARC_1_0/temp4[114] ), .ZN(\MC_ARK_ARC_1_0/temp6[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_12_5  ( .A(\MC_ARK_ARC_1_0/temp1[114] ), .B(
        \MC_ARK_ARC_1_0/temp2[114] ), .ZN(\MC_ARK_ARC_1_0/temp5[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_12_5  ( .A(\RI5[0][150] ), .B(n407), .ZN(
        \MC_ARK_ARC_1_0/temp4[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_12_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_12_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .B(\RI5[0][60] ), .ZN(\MC_ARK_ARC_1_0/temp2[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_12_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[108] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_12_4  ( .A(\MC_ARK_ARC_1_0/temp5[115] ), .B(
        \MC_ARK_ARC_1_0/temp6[115] ), .ZN(\RI1[1][115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_12_4  ( .A(\MC_ARK_ARC_1_0/temp3[115] ), .B(
        \MC_ARK_ARC_1_0/temp4[115] ), .ZN(\MC_ARK_ARC_1_0/temp6[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_12_4  ( .A(\MC_ARK_ARC_1_0/temp1[115] ), .B(
        \MC_ARK_ARC_1_0/temp2[115] ), .ZN(\MC_ARK_ARC_1_0/temp5[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_12_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[151] ), 
        .B(n335), .ZN(\MC_ARK_ARC_1_0/temp4[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_12_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_12_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[61] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_12_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_12_3  ( .A(\MC_ARK_ARC_1_0/temp5[116] ), .B(
        \MC_ARK_ARC_1_0/temp6[116] ), .ZN(\RI1[1][116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_12_3  ( .A(\MC_ARK_ARC_1_0/temp3[116] ), .B(
        \MC_ARK_ARC_1_0/temp4[116] ), .ZN(\MC_ARK_ARC_1_0/temp6[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_12_3  ( .A(\MC_ARK_ARC_1_0/temp1[116] ), .B(
        \MC_ARK_ARC_1_0/temp2[116] ), .ZN(\MC_ARK_ARC_1_0/temp5[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_12_3  ( .A(\RI5[0][152] ), .B(n328), .ZN(
        \MC_ARK_ARC_1_0/temp4[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_12_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[26] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_12_3  ( .A(\RI5[0][62] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[86] ), .ZN(\MC_ARK_ARC_1_0/temp2[116] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_12_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[110] ), 
        .B(n1941), .ZN(\MC_ARK_ARC_1_0/temp1[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_12_2  ( .A(\MC_ARK_ARC_1_0/temp3[117] ), .B(
        \MC_ARK_ARC_1_0/temp4[117] ), .ZN(\MC_ARK_ARC_1_0/temp6[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_12_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[153] ), 
        .B(n437), .ZN(\MC_ARK_ARC_1_0/temp4[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_12_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[183] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_12_2  ( .A(\RI5[0][63] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[87] ), .ZN(\MC_ARK_ARC_1_0/temp2[117] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_12_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[117] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[111] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_12_1  ( .A(\MC_ARK_ARC_1_0/temp3[118] ), .B(
        \MC_ARK_ARC_1_0/temp4[118] ), .ZN(\MC_ARK_ARC_1_0/temp6[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_12_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[154] ), 
        .B(n505), .ZN(\MC_ARK_ARC_1_0/temp4[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_12_1  ( .A(\RI5[0][184] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[28] ), .ZN(\MC_ARK_ARC_1_0/temp3[118] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_12_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[64] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_12_1  ( .A(\RI5[0][112] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[118] ), .ZN(\MC_ARK_ARC_1_0/temp1[118] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_12_0  ( .A(\MC_ARK_ARC_1_0/temp1[119] ), .B(
        \MC_ARK_ARC_1_0/temp2[119] ), .ZN(\MC_ARK_ARC_1_0/temp5[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_12_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[155] ), 
        .B(n459), .ZN(\MC_ARK_ARC_1_0/temp4[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_12_0  ( .A(n1470), .B(
        \MC_ARK_ARC_1_0/buf_datainput[185] ), .ZN(\MC_ARK_ARC_1_0/temp3[119] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_12_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[65] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[89] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_12_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[119] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[113] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_11_5  ( .A(\MC_ARK_ARC_1_0/temp6[120] ), .B(
        \MC_ARK_ARC_1_0/temp5[120] ), .ZN(\RI1[1][120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_11_5  ( .A(\MC_ARK_ARC_1_0/temp3[120] ), .B(
        \MC_ARK_ARC_1_0/temp4[120] ), .ZN(\MC_ARK_ARC_1_0/temp6[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_11_5  ( .A(\MC_ARK_ARC_1_0/temp1[120] ), .B(
        \MC_ARK_ARC_1_0/temp2[120] ), .ZN(\MC_ARK_ARC_1_0/temp5[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_11_5  ( .A(\RI5[0][156] ), .B(n301), .ZN(
        \MC_ARK_ARC_1_0/temp4[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_11_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[186] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_11_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[66] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_11_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[114] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_11_4  ( .A(\MC_ARK_ARC_1_0/temp6[121] ), .B(
        \MC_ARK_ARC_1_0/temp5[121] ), .ZN(\RI1[1][121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_11_4  ( .A(\MC_ARK_ARC_1_0/temp3[121] ), .B(
        \MC_ARK_ARC_1_0/temp4[121] ), .ZN(\MC_ARK_ARC_1_0/temp6[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_11_4  ( .A(\MC_ARK_ARC_1_0/temp1[121] ), .B(
        \MC_ARK_ARC_1_0/temp2[121] ), .ZN(\MC_ARK_ARC_1_0/temp5[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_11_4  ( .A(\RI5[0][157] ), .B(n295), .ZN(
        \MC_ARK_ARC_1_0/temp4[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_11_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[187] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_11_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[67] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_11_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_11_3  ( .A(\MC_ARK_ARC_1_0/temp5[122] ), .B(
        \MC_ARK_ARC_1_0/temp6[122] ), .ZN(\RI1[1][122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_11_3  ( .A(\MC_ARK_ARC_1_0/temp3[122] ), .B(
        \MC_ARK_ARC_1_0/temp4[122] ), .ZN(\MC_ARK_ARC_1_0/temp6[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_11_3  ( .A(\MC_ARK_ARC_1_0/temp1[122] ), .B(
        \MC_ARK_ARC_1_0/temp2[122] ), .ZN(\MC_ARK_ARC_1_0/temp5[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_11_3  ( .A(n2138), .B(n423), .ZN(
        \MC_ARK_ARC_1_0/temp4[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_11_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[188] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_11_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[68] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_11_3  ( .A(n1941), .B(
        \MC_ARK_ARC_1_0/buf_datainput[122] ), .ZN(\MC_ARK_ARC_1_0/temp1[122] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_11_2  ( .A(\MC_ARK_ARC_1_0/temp5[123] ), .B(
        \MC_ARK_ARC_1_0/temp6[123] ), .ZN(\RI1[1][123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_11_2  ( .A(\MC_ARK_ARC_1_0/temp3[123] ), .B(
        \MC_ARK_ARC_1_0/temp4[123] ), .ZN(\MC_ARK_ARC_1_0/temp6[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_11_2  ( .A(\MC_ARK_ARC_1_0/temp1[123] ), .B(
        \MC_ARK_ARC_1_0/temp2[123] ), .ZN(\MC_ARK_ARC_1_0/temp5[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_11_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[159] ), 
        .B(n440), .ZN(\MC_ARK_ARC_1_0/temp4[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_11_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[33] ), 
        .B(n1959), .ZN(\MC_ARK_ARC_1_0/temp3[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_11_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[69] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[93] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_11_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[117] ), 
        .B(\RI5[0][123] ), .ZN(\MC_ARK_ARC_1_0/temp1[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_11_1  ( .A(\MC_ARK_ARC_1_0/temp5[124] ), .B(
        \MC_ARK_ARC_1_0/temp6[124] ), .ZN(\RI1[1][124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_11_1  ( .A(\MC_ARK_ARC_1_0/temp3[124] ), .B(
        \MC_ARK_ARC_1_0/temp4[124] ), .ZN(\MC_ARK_ARC_1_0/temp6[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_11_1  ( .A(\MC_ARK_ARC_1_0/temp2[124] ), .B(
        \MC_ARK_ARC_1_0/temp1[124] ), .ZN(\MC_ARK_ARC_1_0/temp5[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_11_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[160] ), 
        .B(n275), .ZN(\MC_ARK_ARC_1_0/temp4[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_11_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_11_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[70] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_11_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[118] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_11_0  ( .A(\MC_ARK_ARC_1_0/temp1[125] ), .B(
        \MC_ARK_ARC_1_0/temp2[125] ), .ZN(\MC_ARK_ARC_1_0/temp5[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_11_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[161] ), 
        .B(n435), .ZN(\MC_ARK_ARC_1_0/temp4[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_11_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[191] ), 
        .B(n1509), .ZN(\MC_ARK_ARC_1_0/temp3[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_11_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .B(n874), .ZN(\MC_ARK_ARC_1_0/temp2[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_11_0  ( .A(n1939), .B(
        \MC_ARK_ARC_1_0/buf_datainput[119] ), .ZN(\MC_ARK_ARC_1_0/temp1[125] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_10_5  ( .A(\MC_ARK_ARC_1_0/temp5[126] ), .B(
        \MC_ARK_ARC_1_0/temp6[126] ), .ZN(\RI1[1][126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_10_5  ( .A(\MC_ARK_ARC_1_0/temp3[126] ), .B(
        \MC_ARK_ARC_1_0/temp4[126] ), .ZN(\MC_ARK_ARC_1_0/temp6[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_10_5  ( .A(\MC_ARK_ARC_1_0/temp1[126] ), .B(
        \MC_ARK_ARC_1_0/temp2[126] ), .ZN(\MC_ARK_ARC_1_0/temp5[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_10_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[162] ), 
        .B(n402), .ZN(\MC_ARK_ARC_1_0/temp4[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_10_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_0/temp3[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_10_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[72] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_10_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_10_4  ( .A(\MC_ARK_ARC_1_0/temp6[127] ), .B(
        \MC_ARK_ARC_1_0/temp5[127] ), .ZN(\RI1[1][127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_10_4  ( .A(\MC_ARK_ARC_1_0/temp3[127] ), .B(
        \MC_ARK_ARC_1_0/temp4[127] ), .ZN(\MC_ARK_ARC_1_0/temp6[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_10_4  ( .A(\MC_ARK_ARC_1_0/temp1[127] ), .B(
        \MC_ARK_ARC_1_0/temp2[127] ), .ZN(\MC_ARK_ARC_1_0/temp5[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_10_4  ( .A(\RI5[0][163] ), .B(n383), .ZN(
        \MC_ARK_ARC_1_0/temp4[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_10_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[37] ), 
        .B(\RI5[0][1] ), .ZN(\MC_ARK_ARC_1_0/temp3[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_10_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[73] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_10_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_10_3  ( .A(\MC_ARK_ARC_1_0/temp6[128] ), .B(
        \MC_ARK_ARC_1_0/temp5[128] ), .ZN(\RI1[1][128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_10_3  ( .A(\MC_ARK_ARC_1_0/temp3[128] ), .B(
        \MC_ARK_ARC_1_0/temp4[128] ), .ZN(\MC_ARK_ARC_1_0/temp6[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_10_3  ( .A(\MC_ARK_ARC_1_0/temp1[128] ), .B(
        \MC_ARK_ARC_1_0/temp2[128] ), .ZN(\MC_ARK_ARC_1_0/temp5[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_10_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[164] ), 
        .B(n248), .ZN(\MC_ARK_ARC_1_0/temp4[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_10_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[38] ), 
        .B(\RI5[0][2] ), .ZN(\MC_ARK_ARC_1_0/temp3[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_10_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[98] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_10_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_10_2  ( .A(\MC_ARK_ARC_1_0/temp5[129] ), .B(
        \MC_ARK_ARC_1_0/temp6[129] ), .ZN(\RI1[1][129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_10_2  ( .A(\MC_ARK_ARC_1_0/temp3[129] ), .B(
        \MC_ARK_ARC_1_0/temp4[129] ), .ZN(\MC_ARK_ARC_1_0/temp6[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_10_2  ( .A(\MC_ARK_ARC_1_0/temp2[129] ), .B(
        \MC_ARK_ARC_1_0/temp1[129] ), .ZN(\MC_ARK_ARC_1_0/temp5[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_10_2  ( .A(\RI5[0][165] ), .B(n242), .ZN(
        \MC_ARK_ARC_1_0/temp4[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_10_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[3] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[39] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_10_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[99] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_10_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[129] ), 
        .B(\RI5[0][123] ), .ZN(\MC_ARK_ARC_1_0/temp1[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_10_1  ( .A(\MC_ARK_ARC_1_0/temp6[130] ), .B(
        \MC_ARK_ARC_1_0/temp5[130] ), .ZN(\RI1[1][130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_10_1  ( .A(\MC_ARK_ARC_1_0/temp3[130] ), .B(
        \MC_ARK_ARC_1_0/temp4[130] ), .ZN(\MC_ARK_ARC_1_0/temp6[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_10_1  ( .A(\MC_ARK_ARC_1_0/temp1[130] ), .B(
        \MC_ARK_ARC_1_0/temp2[130] ), .ZN(\MC_ARK_ARC_1_0/temp5[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_10_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .B(n507), .ZN(\MC_ARK_ARC_1_0/temp4[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_10_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[40] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_10_1  ( .A(\RI5[0][76] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[100] ), .ZN(\MC_ARK_ARC_1_0/temp2[130] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_10_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[130] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_10_0  ( .A(\MC_ARK_ARC_1_0/temp4[131] ), .B(
        \MC_ARK_ARC_1_0/temp3[131] ), .ZN(\MC_ARK_ARC_1_0/temp6[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_10_0  ( .A(\MC_ARK_ARC_1_0/temp1[131] ), .B(
        \MC_ARK_ARC_1_0/temp2[131] ), .ZN(\MC_ARK_ARC_1_0/temp5[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_10_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .B(n489), .ZN(\MC_ARK_ARC_1_0/temp4[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_10_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[5] ), 
        .B(n1483), .ZN(\MC_ARK_ARC_1_0/temp3[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_10_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[101] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[77] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_10_0  ( .A(n1939), .B(
        \MC_ARK_ARC_1_0/buf_datainput[131] ), .ZN(\MC_ARK_ARC_1_0/temp1[131] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_9_5  ( .A(\MC_ARK_ARC_1_0/temp5[132] ), .B(
        \MC_ARK_ARC_1_0/temp6[132] ), .ZN(\RI1[1][132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_9_5  ( .A(\MC_ARK_ARC_1_0/temp3[132] ), .B(
        \MC_ARK_ARC_1_0/temp4[132] ), .ZN(\MC_ARK_ARC_1_0/temp6[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_9_5  ( .A(\MC_ARK_ARC_1_0/temp2[132] ), .B(
        \MC_ARK_ARC_1_0/temp1[132] ), .ZN(\MC_ARK_ARC_1_0/temp5[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_9_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[168] ), 
        .B(n222), .ZN(\MC_ARK_ARC_1_0/temp4[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_9_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_0/temp3[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_9_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[78] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_9_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[126] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_9_4  ( .A(\MC_ARK_ARC_1_0/temp5[133] ), .B(
        \MC_ARK_ARC_1_0/temp6[133] ), .ZN(\RI1[1][133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_9_4  ( .A(\MC_ARK_ARC_1_0/temp3[133] ), .B(
        \MC_ARK_ARC_1_0/temp4[133] ), .ZN(\MC_ARK_ARC_1_0/temp6[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_9_4  ( .A(\MC_ARK_ARC_1_0/temp1[133] ), .B(
        \MC_ARK_ARC_1_0/temp2[133] ), .ZN(\MC_ARK_ARC_1_0/temp5[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_9_4  ( .A(\RI5[0][169] ), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[45] ), .ZN(\MC_ARK_ARC_1_0/temp4[133] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_9_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_0/temp3[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_9_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[79] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_9_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[133] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[127] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_9_3  ( .A(\MC_ARK_ARC_1_0/temp5[134] ), .B(
        \MC_ARK_ARC_1_0/temp6[134] ), .ZN(\RI1[1][134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_9_3  ( .A(\MC_ARK_ARC_1_0/temp4[134] ), .B(
        \MC_ARK_ARC_1_0/temp3[134] ), .ZN(\MC_ARK_ARC_1_0/temp6[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_9_3  ( .A(\MC_ARK_ARC_1_0/temp2[134] ), .B(
        \MC_ARK_ARC_1_0/temp1[134] ), .ZN(\MC_ARK_ARC_1_0/temp5[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_9_3  ( .A(\RI5[0][170] ), .B(n208), .ZN(
        \MC_ARK_ARC_1_0/temp4[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_9_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[8] ), 
        .B(n1473), .ZN(\MC_ARK_ARC_1_0/temp3[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_9_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[104] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[80] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_9_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_9_2  ( .A(\MC_ARK_ARC_1_0/temp5[135] ), .B(
        \MC_ARK_ARC_1_0/temp6[135] ), .ZN(\RI1[1][135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_9_2  ( .A(\MC_ARK_ARC_1_0/temp3[135] ), .B(
        \MC_ARK_ARC_1_0/temp4[135] ), .ZN(\MC_ARK_ARC_1_0/temp6[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_9_2  ( .A(\MC_ARK_ARC_1_0/temp2[135] ), .B(
        \MC_ARK_ARC_1_0/temp1[135] ), .ZN(\MC_ARK_ARC_1_0/temp5[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_9_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[171] ), 
        .B(n201), .ZN(\MC_ARK_ARC_1_0/temp4[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_9_2  ( .A(\RI5[0][45] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_0/temp3[135] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_9_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[81] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_9_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[135] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[129] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_9_1  ( .A(\MC_ARK_ARC_1_0/temp6[136] ), .B(
        \MC_ARK_ARC_1_0/temp5[136] ), .ZN(\RI1[1][136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_9_1  ( .A(\MC_ARK_ARC_1_0/temp3[136] ), .B(
        \MC_ARK_ARC_1_0/temp4[136] ), .ZN(\MC_ARK_ARC_1_0/temp6[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_9_1  ( .A(\MC_ARK_ARC_1_0/temp1[136] ), .B(
        \MC_ARK_ARC_1_0/temp2[136] ), .ZN(\MC_ARK_ARC_1_0/temp5[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_9_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_0/buf_keyinput[136] ), .ZN(
        \MC_ARK_ARC_1_0/temp4[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_9_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[10] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_9_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[82] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_9_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_9_0  ( .A(\MC_ARK_ARC_1_0/temp5[137] ), .B(
        \MC_ARK_ARC_1_0/temp6[137] ), .ZN(\RI1[1][137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_9_0  ( .A(\MC_ARK_ARC_1_0/temp3[137] ), .B(
        \MC_ARK_ARC_1_0/temp4[137] ), .ZN(\MC_ARK_ARC_1_0/temp6[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_9_0  ( .A(\MC_ARK_ARC_1_0/temp1[137] ), .B(
        \MC_ARK_ARC_1_0/temp2[137] ), .ZN(\MC_ARK_ARC_1_0/temp5[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_9_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[173] ), 
        .B(n432), .ZN(\MC_ARK_ARC_1_0/temp4[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_9_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[47] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[11] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_9_0  ( .A(n1480), .B(
        \MC_ARK_ARC_1_0/buf_datainput[83] ), .ZN(\MC_ARK_ARC_1_0/temp2[137] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_9_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[131] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_8_5  ( .A(\MC_ARK_ARC_1_0/temp6[138] ), .B(
        \MC_ARK_ARC_1_0/temp5[138] ), .ZN(\RI1[1][138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_8_5  ( .A(\MC_ARK_ARC_1_0/temp3[138] ), .B(
        \MC_ARK_ARC_1_0/temp4[138] ), .ZN(\MC_ARK_ARC_1_0/temp6[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_8_5  ( .A(\MC_ARK_ARC_1_0/temp1[138] ), .B(
        \MC_ARK_ARC_1_0/temp2[138] ), .ZN(\MC_ARK_ARC_1_0/temp5[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_8_5  ( .A(\RI5[0][174] ), .B(n398), .ZN(
        \MC_ARK_ARC_1_0/temp4[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_8_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[12] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_8_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[108] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[84] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_8_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[132] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_8_4  ( .A(\MC_ARK_ARC_1_0/temp5[139] ), .B(
        \MC_ARK_ARC_1_0/temp6[139] ), .ZN(\RI1[1][139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_8_4  ( .A(\MC_ARK_ARC_1_0/temp3[139] ), .B(
        \MC_ARK_ARC_1_0/temp4[139] ), .ZN(\MC_ARK_ARC_1_0/temp6[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_8_4  ( .A(\MC_ARK_ARC_1_0/temp2[139] ), .B(
        \MC_ARK_ARC_1_0/temp1[139] ), .ZN(\MC_ARK_ARC_1_0/temp5[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_8_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[175] ), 
        .B(n357), .ZN(\MC_ARK_ARC_1_0/temp4[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_8_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[13] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_8_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[85] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_8_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[133] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_8_3  ( .A(\MC_ARK_ARC_1_0/temp5[140] ), .B(
        \MC_ARK_ARC_1_0/temp6[140] ), .ZN(\RI1[1][140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_8_3  ( .A(\MC_ARK_ARC_1_0/temp3[140] ), .B(
        \MC_ARK_ARC_1_0/temp4[140] ), .ZN(\MC_ARK_ARC_1_0/temp6[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_8_3  ( .A(\MC_ARK_ARC_1_0/temp2[140] ), .B(
        \MC_ARK_ARC_1_0/temp1[140] ), .ZN(\MC_ARK_ARC_1_0/temp5[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_8_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[129] ), .ZN(
        \MC_ARK_ARC_1_0/temp4[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_8_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[14] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_8_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[86] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_8_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[134] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_8_2  ( .A(\MC_ARK_ARC_1_0/temp6[141] ), .B(
        \MC_ARK_ARC_1_0/temp5[141] ), .ZN(\RI1[1][141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_8_2  ( .A(\MC_ARK_ARC_1_0/temp3[141] ), .B(
        \MC_ARK_ARC_1_0/temp4[141] ), .ZN(\MC_ARK_ARC_1_0/temp6[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_8_2  ( .A(\MC_ARK_ARC_1_0/temp1[141] ), .B(
        \MC_ARK_ARC_1_0/temp2[141] ), .ZN(\MC_ARK_ARC_1_0/temp5[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_8_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[177] ), 
        .B(n460), .ZN(\MC_ARK_ARC_1_0/temp4[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_8_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[15] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[51] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_8_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[111] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[87] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_8_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[135] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_8_1  ( .A(\MC_ARK_ARC_1_0/temp5[142] ), .B(
        \MC_ARK_ARC_1_0/temp6[142] ), .ZN(\RI1[1][142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_8_1  ( .A(\MC_ARK_ARC_1_0/temp3[142] ), .B(
        \MC_ARK_ARC_1_0/temp4[142] ), .ZN(\MC_ARK_ARC_1_0/temp6[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_8_1  ( .A(\MC_ARK_ARC_1_0/temp2[142] ), .B(
        \MC_ARK_ARC_1_0/temp1[142] ), .ZN(\MC_ARK_ARC_1_0/temp5[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_8_1  ( .A(\RI5[0][178] ), .B(n472), .ZN(
        \MC_ARK_ARC_1_0/temp4[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_8_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[52] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_8_1  ( .A(\RI5[0][112] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_0/temp2[142] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_8_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[142] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_8_0  ( .A(\MC_ARK_ARC_1_0/temp3[143] ), .B(
        \MC_ARK_ARC_1_0/temp4[143] ), .ZN(\MC_ARK_ARC_1_0/temp6[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_8_0  ( .A(\MC_ARK_ARC_1_0/temp1[143] ), .B(
        \MC_ARK_ARC_1_0/temp2[143] ), .ZN(\MC_ARK_ARC_1_0/temp5[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_8_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[179] ), 
        .B(n462), .ZN(\MC_ARK_ARC_1_0/temp4[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_8_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[17] ), 
        .B(n1631), .ZN(\MC_ARK_ARC_1_0/temp3[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_8_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[89] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[113] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_8_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[143] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_7_5  ( .A(\MC_ARK_ARC_1_0/temp5[144] ), .B(
        \MC_ARK_ARC_1_0/temp6[144] ), .ZN(\RI1[1][144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_7_5  ( .A(\MC_ARK_ARC_1_0/temp3[144] ), .B(
        \MC_ARK_ARC_1_0/temp4[144] ), .ZN(\MC_ARK_ARC_1_0/temp6[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_7_5  ( .A(\MC_ARK_ARC_1_0/temp1[144] ), .B(
        \MC_ARK_ARC_1_0/temp2[144] ), .ZN(\MC_ARK_ARC_1_0/temp5[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_7_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .B(n324), .ZN(\MC_ARK_ARC_1_0/temp4[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_7_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[18] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_7_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[90] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_7_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[144] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[138] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_7_4  ( .A(\MC_ARK_ARC_1_0/temp5[145] ), .B(
        \MC_ARK_ARC_1_0/temp6[145] ), .ZN(\RI1[1][145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_7_4  ( .A(\MC_ARK_ARC_1_0/temp3[145] ), .B(
        \MC_ARK_ARC_1_0/temp4[145] ), .ZN(\MC_ARK_ARC_1_0/temp6[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_7_4  ( .A(\MC_ARK_ARC_1_0/temp1[145] ), .B(
        \MC_ARK_ARC_1_0/temp2[145] ), .ZN(\MC_ARK_ARC_1_0/temp5[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_7_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[181] ), 
        .B(n318), .ZN(\MC_ARK_ARC_1_0/temp4[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_7_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[19] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_7_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[91] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_7_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[139] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_7_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[182] ), 
        .B(n443), .ZN(\MC_ARK_ARC_1_0/temp4[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_7_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[56] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[20] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_7_3  ( .A(n1941), .B(
        \MC_ARK_ARC_1_0/buf_datainput[92] ), .ZN(\MC_ARK_ARC_1_0/temp2[146] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_7_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[140] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_7_2  ( .A(\MC_ARK_ARC_1_0/temp5[147] ), .B(
        \MC_ARK_ARC_1_0/temp6[147] ), .ZN(\RI1[1][147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_7_2  ( .A(\MC_ARK_ARC_1_0/temp3[147] ), .B(
        \MC_ARK_ARC_1_0/temp4[147] ), .ZN(\MC_ARK_ARC_1_0/temp6[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_7_2  ( .A(\MC_ARK_ARC_1_0/temp2[147] ), .B(
        \MC_ARK_ARC_1_0/temp1[147] ), .ZN(\MC_ARK_ARC_1_0/temp5[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_7_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[183] ), 
        .B(n497), .ZN(\MC_ARK_ARC_1_0/temp4[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_7_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[57] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[21] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_7_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[93] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[117] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_7_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[147] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_7_1  ( .A(\MC_ARK_ARC_1_0/temp6[148] ), .B(
        \MC_ARK_ARC_1_0/temp5[148] ), .ZN(\RI1[1][148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_7_1  ( .A(\MC_ARK_ARC_1_0/temp4[148] ), .B(
        \MC_ARK_ARC_1_0/temp3[148] ), .ZN(\MC_ARK_ARC_1_0/temp6[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_7_1  ( .A(\MC_ARK_ARC_1_0/temp1[148] ), .B(
        \MC_ARK_ARC_1_0/temp2[148] ), .ZN(\MC_ARK_ARC_1_0/temp5[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_7_1  ( .A(\RI5[0][184] ), .B(n488), .ZN(
        \MC_ARK_ARC_1_0/temp4[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_7_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[22] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_7_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[118] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[94] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_7_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[142] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_7_0  ( .A(\MC_ARK_ARC_1_0/temp1[149] ), .B(
        \MC_ARK_ARC_1_0/temp2[149] ), .ZN(\MC_ARK_ARC_1_0/temp5[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_7_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[185] ), 
        .B(n291), .ZN(\MC_ARK_ARC_1_0/temp4[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_7_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[23] ), 
        .B(n788), .ZN(\MC_ARK_ARC_1_0/temp3[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_7_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[119] ), 
        .B(n875), .ZN(\MC_ARK_ARC_1_0/temp2[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_7_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[143] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[149] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_6_5  ( .A(\MC_ARK_ARC_1_0/temp5[150] ), .B(
        \MC_ARK_ARC_1_0/temp6[150] ), .ZN(\RI1[1][150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_6_5  ( .A(\MC_ARK_ARC_1_0/temp3[150] ), .B(
        \MC_ARK_ARC_1_0/temp4[150] ), .ZN(\MC_ARK_ARC_1_0/temp6[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_6_5  ( .A(\MC_ARK_ARC_1_0/temp1[150] ), .B(
        \MC_ARK_ARC_1_0/temp2[150] ), .ZN(\MC_ARK_ARC_1_0/temp5[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_6_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[186] ), 
        .B(n479), .ZN(\MC_ARK_ARC_1_0/temp4[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_6_5  ( .A(\RI5[0][60] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[24] ), .ZN(\MC_ARK_ARC_1_0/temp3[150] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_6_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[96] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_6_5  ( .A(\RI5[0][150] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[144] ), .ZN(\MC_ARK_ARC_1_0/temp1[150] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_6_4  ( .A(\MC_ARK_ARC_1_0/temp5[151] ), .B(
        \MC_ARK_ARC_1_0/temp6[151] ), .ZN(\RI1[1][151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_6_4  ( .A(\MC_ARK_ARC_1_0/temp3[151] ), .B(
        \MC_ARK_ARC_1_0/temp4[151] ), .ZN(\MC_ARK_ARC_1_0/temp6[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_6_4  ( .A(\MC_ARK_ARC_1_0/temp1[151] ), .B(
        \MC_ARK_ARC_1_0/temp2[151] ), .ZN(\MC_ARK_ARC_1_0/temp5[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_6_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[187] ), 
        .B(n278), .ZN(\MC_ARK_ARC_1_0/temp4[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_6_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[25] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_6_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[97] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_6_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[145] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_6_3  ( .A(\MC_ARK_ARC_1_0/temp3[152] ), .B(
        \MC_ARK_ARC_1_0/temp4[152] ), .ZN(\MC_ARK_ARC_1_0/temp6[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_6_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[188] ), 
        .B(n271), .ZN(\MC_ARK_ARC_1_0/temp4[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_6_3  ( .A(\RI5[0][62] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_0/temp3[152] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_6_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[98] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_6_3  ( .A(\RI5[0][152] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[146] ), .ZN(\MC_ARK_ARC_1_0/temp1[152] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_6_2  ( .A(\MC_ARK_ARC_1_0/temp5[153] ), .B(
        \MC_ARK_ARC_1_0/temp6[153] ), .ZN(\RI1[1][153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_6_2  ( .A(\MC_ARK_ARC_1_0/temp3[153] ), .B(
        \MC_ARK_ARC_1_0/temp4[153] ), .ZN(\MC_ARK_ARC_1_0/temp6[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_6_2  ( .A(\MC_ARK_ARC_1_0/temp1[153] ), .B(
        \MC_ARK_ARC_1_0/temp2[153] ), .ZN(\MC_ARK_ARC_1_0/temp5[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_6_2  ( .A(n1959), .B(n467), .ZN(
        \MC_ARK_ARC_1_0/temp4[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_6_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[27] ), 
        .B(\RI5[0][63] ), .ZN(\MC_ARK_ARC_1_0/temp3[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_6_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[99] ), 
        .B(\RI5[0][123] ), .ZN(\MC_ARK_ARC_1_0/temp2[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_6_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[153] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[147] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_6_1  ( .A(\MC_ARK_ARC_1_0/temp5[154] ), .B(
        \MC_ARK_ARC_1_0/temp6[154] ), .ZN(\RI1[1][154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_6_1  ( .A(\MC_ARK_ARC_1_0/temp3[154] ), .B(
        \MC_ARK_ARC_1_0/temp4[154] ), .ZN(\MC_ARK_ARC_1_0/temp6[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_6_1  ( .A(\MC_ARK_ARC_1_0/temp1[154] ), .B(
        \MC_ARK_ARC_1_0/temp2[154] ), .ZN(\MC_ARK_ARC_1_0/temp5[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_6_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[190] ), 
        .B(n257), .ZN(\MC_ARK_ARC_1_0/temp4[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_6_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[28] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_6_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_6_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[148] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_6_0  ( .A(\MC_ARK_ARC_1_0/temp3[155] ), .B(
        \MC_ARK_ARC_1_0/temp4[155] ), .ZN(\MC_ARK_ARC_1_0/temp6[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_6_0  ( .A(\MC_ARK_ARC_1_0/temp2[155] ), .B(
        \MC_ARK_ARC_1_0/temp1[155] ), .ZN(\MC_ARK_ARC_1_0/temp5[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_6_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[191] ), 
        .B(n471), .ZN(\MC_ARK_ARC_1_0/temp4[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_6_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[65] ), 
        .B(n1960), .ZN(\MC_ARK_ARC_1_0/temp3[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_6_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[101] ), 
        .B(n1939), .ZN(\MC_ARK_ARC_1_0/temp2[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_6_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[149] ), 
        .B(n2116), .ZN(\MC_ARK_ARC_1_0/temp1[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_5_5  ( .A(\MC_ARK_ARC_1_0/temp5[156] ), .B(
        \MC_ARK_ARC_1_0/temp6[156] ), .ZN(\RI1[1][156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_5_5  ( .A(\MC_ARK_ARC_1_0/temp3[156] ), .B(
        \MC_ARK_ARC_1_0/temp4[156] ), .ZN(\MC_ARK_ARC_1_0/temp6[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_5_5  ( .A(\MC_ARK_ARC_1_0/temp1[156] ), .B(
        \MC_ARK_ARC_1_0/temp2[156] ), .ZN(\MC_ARK_ARC_1_0/temp5[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_5_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[0] ), 
        .B(n408), .ZN(\MC_ARK_ARC_1_0/temp4[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_5_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[30] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_5_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[102] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_5_5  ( .A(\RI5[0][156] ), .B(\RI5[0][150] ), 
        .ZN(\MC_ARK_ARC_1_0/temp1[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_5_4  ( .A(\MC_ARK_ARC_1_0/temp6[157] ), .B(
        \MC_ARK_ARC_1_0/temp5[157] ), .ZN(\RI1[1][157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_5_4  ( .A(\MC_ARK_ARC_1_0/temp3[157] ), .B(
        \MC_ARK_ARC_1_0/temp4[157] ), .ZN(\MC_ARK_ARC_1_0/temp6[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_5_4  ( .A(\MC_ARK_ARC_1_0/temp1[157] ), .B(
        \MC_ARK_ARC_1_0/temp2[157] ), .ZN(\MC_ARK_ARC_1_0/temp5[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_5_4  ( .A(\RI5[0][1] ), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[69] ), .ZN(\MC_ARK_ARC_1_0/temp4[157] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_5_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[31] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_5_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_5_4  ( .A(\RI5[0][157] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[151] ), .ZN(\MC_ARK_ARC_1_0/temp1[157] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_5_3  ( .A(\MC_ARK_ARC_1_0/temp2[158] ), .B(
        \MC_ARK_ARC_1_0/temp1[158] ), .ZN(\MC_ARK_ARC_1_0/temp5[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_5_3  ( .A(\RI5[0][2] ), .B(
        \MC_ARK_ARC_1_0/buf_keyinput[158] ), .ZN(\MC_ARK_ARC_1_0/temp4[158] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_5_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[68] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_5_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_5_3  ( .A(\RI5[0][152] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[158] ), .ZN(\MC_ARK_ARC_1_0/temp1[158] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_5_2  ( .A(\MC_ARK_ARC_1_0/temp5[159] ), .B(
        \MC_ARK_ARC_1_0/temp6[159] ), .ZN(\RI1[1][159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_5_2  ( .A(\MC_ARK_ARC_1_0/temp3[159] ), .B(
        \MC_ARK_ARC_1_0/temp4[159] ), .ZN(\MC_ARK_ARC_1_0/temp6[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_5_2  ( .A(\MC_ARK_ARC_1_0/temp1[159] ), .B(
        \MC_ARK_ARC_1_0/temp2[159] ), .ZN(\MC_ARK_ARC_1_0/temp5[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_5_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[3] ), 
        .B(n225), .ZN(\MC_ARK_ARC_1_0/temp4[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_5_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[69] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_5_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[129] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[105] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_5_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[159] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[153] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_5_1  ( .A(\MC_ARK_ARC_1_0/temp5[160] ), .B(
        \MC_ARK_ARC_1_0/temp6[160] ), .ZN(\RI1[1][160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_5_1  ( .A(\MC_ARK_ARC_1_0/temp3[160] ), .B(
        \MC_ARK_ARC_1_0/temp4[160] ), .ZN(\MC_ARK_ARC_1_0/temp6[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_5_1  ( .A(\MC_ARK_ARC_1_0/temp1[160] ), .B(
        \MC_ARK_ARC_1_0/temp2[160] ), .ZN(\MC_ARK_ARC_1_0/temp5[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_5_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[4] ), 
        .B(n493), .ZN(\MC_ARK_ARC_1_0/temp4[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_5_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[34] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_5_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_5_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_5_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[5] ), 
        .B(n470), .ZN(\MC_ARK_ARC_1_0/temp4[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_5_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .B(n1507), .ZN(\MC_ARK_ARC_1_0/temp3[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_5_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[131] ), 
        .B(n1962), .ZN(\MC_ARK_ARC_1_0/temp2[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_5_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[161] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[155] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_4_5  ( .A(\MC_ARK_ARC_1_0/temp6[162] ), .B(
        \MC_ARK_ARC_1_0/temp5[162] ), .ZN(\RI1[1][162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_4_5  ( .A(\MC_ARK_ARC_1_0/temp3[162] ), .B(
        \MC_ARK_ARC_1_0/temp4[162] ), .ZN(\MC_ARK_ARC_1_0/temp6[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_4_5  ( .A(\MC_ARK_ARC_1_0/temp1[162] ), .B(
        \MC_ARK_ARC_1_0/temp2[162] ), .ZN(\MC_ARK_ARC_1_0/temp5[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_4_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[6] ), 
        .B(n401), .ZN(\MC_ARK_ARC_1_0/temp4[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_4_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[36] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_4_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[108] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_4_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[162] ), 
        .B(\RI5[0][156] ), .ZN(\MC_ARK_ARC_1_0/temp1[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_4_4  ( .A(\MC_ARK_ARC_1_0/temp5[163] ), .B(
        \MC_ARK_ARC_1_0/temp6[163] ), .ZN(\RI1[1][163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_4_4  ( .A(\MC_ARK_ARC_1_0/temp3[163] ), .B(
        \MC_ARK_ARC_1_0/temp4[163] ), .ZN(\MC_ARK_ARC_1_0/temp6[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_4_4  ( .A(\MC_ARK_ARC_1_0/temp1[163] ), .B(
        \MC_ARK_ARC_1_0/temp2[163] ), .ZN(\MC_ARK_ARC_1_0/temp5[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_4_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .B(n198), .ZN(\MC_ARK_ARC_1_0/temp4[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_4_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[37] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_4_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[133] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_4_4  ( .A(\RI5[0][163] ), .B(\RI5[0][157] ), 
        .ZN(\MC_ARK_ARC_1_0/temp1[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_4_3  ( .A(\MC_ARK_ARC_1_0/temp5[164] ), .B(
        \MC_ARK_ARC_1_0/temp6[164] ), .ZN(\RI1[1][164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_4_3  ( .A(\MC_ARK_ARC_1_0/temp3[164] ), .B(
        \MC_ARK_ARC_1_0/temp4[164] ), .ZN(\MC_ARK_ARC_1_0/temp6[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_4_3  ( .A(\MC_ARK_ARC_1_0/temp2[164] ), .B(
        \MC_ARK_ARC_1_0/temp1[164] ), .ZN(\MC_ARK_ARC_1_0/temp5[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_4_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[8] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[105] ), .ZN(
        \MC_ARK_ARC_1_0/temp4[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_4_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[38] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_4_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[134] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_4_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[164] ), 
        .B(n2138), .ZN(\MC_ARK_ARC_1_0/temp1[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_4_2  ( .A(\MC_ARK_ARC_1_0/temp5[165] ), .B(
        \MC_ARK_ARC_1_0/temp6[165] ), .ZN(\RI1[1][165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_4_2  ( .A(\MC_ARK_ARC_1_0/temp3[165] ), .B(
        \MC_ARK_ARC_1_0/temp4[165] ), .ZN(\MC_ARK_ARC_1_0/temp6[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_4_2  ( .A(\MC_ARK_ARC_1_0/temp2[165] ), .B(
        \MC_ARK_ARC_1_0/temp1[165] ), .ZN(\MC_ARK_ARC_1_0/temp5[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_4_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[9] ), 
        .B(n499), .ZN(\MC_ARK_ARC_1_0/temp4[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_4_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[39] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_4_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[135] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[111] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_4_2  ( .A(\RI5[0][165] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[159] ), .ZN(\MC_ARK_ARC_1_0/temp1[165] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_4_1  ( .A(\MC_ARK_ARC_1_0/temp6[166] ), .B(
        \MC_ARK_ARC_1_0/temp5[166] ), .ZN(\RI1[1][166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_4_1  ( .A(\MC_ARK_ARC_1_0/temp3[166] ), .B(
        \MC_ARK_ARC_1_0/temp4[166] ), .ZN(\MC_ARK_ARC_1_0/temp6[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_4_1  ( .A(\MC_ARK_ARC_1_0/temp2[166] ), .B(
        \MC_ARK_ARC_1_0/temp1[166] ), .ZN(\MC_ARK_ARC_1_0/temp5[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_4_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[10] ), 
        .B(n506), .ZN(\MC_ARK_ARC_1_0/temp4[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_4_1  ( .A(\RI5[0][76] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[40] ), .ZN(\MC_ARK_ARC_1_0/temp3[166] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_4_1  ( .A(\RI5[0][112] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[136] ), .ZN(\MC_ARK_ARC_1_0/temp2[166] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_4_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_4_0  ( .A(n2147), .B(n353), .ZN(
        \MC_ARK_ARC_1_0/temp4[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_4_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .B(n1961), .ZN(\MC_ARK_ARC_1_0/temp3[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_4_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[137] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_4_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[161] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_3_5  ( .A(\MC_ARK_ARC_1_0/temp6[168] ), .B(
        \MC_ARK_ARC_1_0/temp5[168] ), .ZN(\RI1[1][168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_3_5  ( .A(\MC_ARK_ARC_1_0/temp3[168] ), .B(
        \MC_ARK_ARC_1_0/temp4[168] ), .ZN(\MC_ARK_ARC_1_0/temp6[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_3_5  ( .A(\MC_ARK_ARC_1_0/temp1[168] ), .B(
        \MC_ARK_ARC_1_0/temp2[168] ), .ZN(\MC_ARK_ARC_1_0/temp5[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_3_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[12] ), 
        .B(n403), .ZN(\MC_ARK_ARC_1_0/temp4[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_3_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[42] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_3_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[114] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_3_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_3_4  ( .A(\MC_ARK_ARC_1_0/temp5[169] ), .B(
        \MC_ARK_ARC_1_0/temp6[169] ), .ZN(\RI1[1][169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_3_4  ( .A(\MC_ARK_ARC_1_0/temp3[169] ), .B(
        \MC_ARK_ARC_1_0/temp4[169] ), .ZN(\MC_ARK_ARC_1_0/temp6[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_3_4  ( .A(\MC_ARK_ARC_1_0/temp1[169] ), .B(
        \MC_ARK_ARC_1_0/temp2[169] ), .ZN(\MC_ARK_ARC_1_0/temp5[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_3_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[13] ), 
        .B(n340), .ZN(\MC_ARK_ARC_1_0/temp4[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_3_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[43] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_3_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_3_4  ( .A(\RI5[0][169] ), .B(\RI5[0][163] ), 
        .ZN(\MC_ARK_ARC_1_0/temp1[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_3_3  ( .A(\MC_ARK_ARC_1_0/temp5[170] ), .B(
        \MC_ARK_ARC_1_0/temp6[170] ), .ZN(\RI1[1][170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_3_3  ( .A(\MC_ARK_ARC_1_0/temp3[170] ), .B(
        \MC_ARK_ARC_1_0/temp4[170] ), .ZN(\MC_ARK_ARC_1_0/temp6[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_3_3  ( .A(\MC_ARK_ARC_1_0/temp2[170] ), .B(
        \MC_ARK_ARC_1_0/temp1[170] ), .ZN(\MC_ARK_ARC_1_0/temp5[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_3_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[14] ), 
        .B(n384), .ZN(\MC_ARK_ARC_1_0/temp4[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_3_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[80] ), 
        .B(n1475), .ZN(\MC_ARK_ARC_1_0/temp3[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_3_3  ( .A(n1941), .B(
        \MC_ARK_ARC_1_0/buf_datainput[140] ), .ZN(\MC_ARK_ARC_1_0/temp2[170] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_3_3  ( .A(\RI5[0][170] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[164] ), .ZN(\MC_ARK_ARC_1_0/temp1[170] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_3_2  ( .A(\MC_ARK_ARC_1_0/temp5[171] ), .B(
        \MC_ARK_ARC_1_0/temp6[171] ), .ZN(\RI1[1][171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_3_2  ( .A(\MC_ARK_ARC_1_0/temp3[171] ), .B(
        \MC_ARK_ARC_1_0/temp4[171] ), .ZN(\MC_ARK_ARC_1_0/temp6[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_3_2  ( .A(\MC_ARK_ARC_1_0/temp1[171] ), .B(
        \MC_ARK_ARC_1_0/temp2[171] ), .ZN(\MC_ARK_ARC_1_0/temp5[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_3_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[15] ), 
        .B(n327), .ZN(\MC_ARK_ARC_1_0/temp4[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_3_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[81] ), 
        .B(\RI5[0][45] ), .ZN(\MC_ARK_ARC_1_0/temp3[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_3_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[117] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_3_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[171] ), 
        .B(\RI5[0][165] ), .ZN(\MC_ARK_ARC_1_0/temp1[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_3_1  ( .A(\MC_ARK_ARC_1_0/temp6[172] ), .B(
        \MC_ARK_ARC_1_0/temp5[172] ), .ZN(\RI1[1][172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_3_1  ( .A(\MC_ARK_ARC_1_0/temp4[172] ), .B(
        \MC_ARK_ARC_1_0/temp3[172] ), .ZN(\MC_ARK_ARC_1_0/temp6[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_3_1  ( .A(\MC_ARK_ARC_1_0/temp2[172] ), .B(
        \MC_ARK_ARC_1_0/temp1[172] ), .ZN(\MC_ARK_ARC_1_0/temp5[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_3_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[16] ), 
        .B(n444), .ZN(\MC_ARK_ARC_1_0/temp4[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_3_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[46] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_3_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[118] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_3_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_3_0  ( .A(\MC_ARK_ARC_1_0/temp1[173] ), .B(
        \MC_ARK_ARC_1_0/temp2[173] ), .ZN(\MC_ARK_ARC_1_0/temp5[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_3_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[17] ), 
        .B(n314), .ZN(\MC_ARK_ARC_1_0/temp4[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_3_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[83] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[47] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_3_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[143] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[119] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_3_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .B(n2150), .ZN(\MC_ARK_ARC_1_0/temp1[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_2_5  ( .A(\MC_ARK_ARC_1_0/temp5[174] ), .B(
        \MC_ARK_ARC_1_0/temp6[174] ), .ZN(\RI1[1][174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_2_5  ( .A(\MC_ARK_ARC_1_0/temp3[174] ), .B(
        \MC_ARK_ARC_1_0/temp4[174] ), .ZN(\MC_ARK_ARC_1_0/temp6[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_2_5  ( .A(\MC_ARK_ARC_1_0/temp1[174] ), .B(
        \MC_ARK_ARC_1_0/temp2[174] ), .ZN(\MC_ARK_ARC_1_0/temp5[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_2_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[18] ), 
        .B(n307), .ZN(\MC_ARK_ARC_1_0/temp4[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_2_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[48] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_2_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[144] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_2_5  ( .A(\RI5[0][174] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[168] ), .ZN(\MC_ARK_ARC_1_0/temp1[174] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_2_4  ( .A(\MC_ARK_ARC_1_0/temp5[175] ), .B(
        \MC_ARK_ARC_1_0/temp6[175] ), .ZN(\RI1[1][175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_2_4  ( .A(\MC_ARK_ARC_1_0/temp3[175] ), .B(
        \MC_ARK_ARC_1_0/temp4[175] ), .ZN(\MC_ARK_ARC_1_0/temp6[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_2_4  ( .A(\MC_ARK_ARC_1_0/temp1[175] ), .B(
        \MC_ARK_ARC_1_0/temp2[175] ), .ZN(\MC_ARK_ARC_1_0/temp5[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_2_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[134] ), .ZN(
        \MC_ARK_ARC_1_0/temp4[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_2_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[49] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_2_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_2_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[175] ), 
        .B(\RI5[0][169] ), .ZN(\MC_ARK_ARC_1_0/temp1[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_2_3  ( .A(\MC_ARK_ARC_1_0/temp5[176] ), .B(
        \MC_ARK_ARC_1_0/temp6[176] ), .ZN(\RI1[1][176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_2_3  ( .A(\MC_ARK_ARC_1_0/temp3[176] ), .B(
        \MC_ARK_ARC_1_0/temp4[176] ), .ZN(\MC_ARK_ARC_1_0/temp6[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_2_3  ( .A(\MC_ARK_ARC_1_0/temp1[176] ), .B(
        \MC_ARK_ARC_1_0/temp2[176] ), .ZN(\MC_ARK_ARC_1_0/temp5[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_2_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[20] ), 
        .B(n294), .ZN(\MC_ARK_ARC_1_0/temp4[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_2_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[50] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_2_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[122] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_2_3  ( .A(\RI5[0][170] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[176] ), .ZN(\MC_ARK_ARC_1_0/temp1[176] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_2_2  ( .A(\MC_ARK_ARC_1_0/temp1[177] ), .B(
        \MC_ARK_ARC_1_0/temp2[177] ), .ZN(\MC_ARK_ARC_1_0/temp5[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_2_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[21] ), 
        .B(n287), .ZN(\MC_ARK_ARC_1_0/temp4[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_2_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[87] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_2_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[147] ), 
        .B(\RI5[0][123] ), .ZN(\MC_ARK_ARC_1_0/temp2[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_2_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[171] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[177] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_2_1  ( .A(\MC_ARK_ARC_1_0/temp5[178] ), .B(
        \MC_ARK_ARC_1_0/temp6[178] ), .ZN(\RI1[1][178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_2_1  ( .A(\MC_ARK_ARC_1_0/temp3[178] ), .B(
        \MC_ARK_ARC_1_0/temp4[178] ), .ZN(\MC_ARK_ARC_1_0/temp6[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_2_1  ( .A(\MC_ARK_ARC_1_0/temp1[178] ), .B(
        \MC_ARK_ARC_1_0/temp2[178] ), .ZN(\MC_ARK_ARC_1_0/temp5[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_2_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .B(n281), .ZN(\MC_ARK_ARC_1_0/temp4[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_2_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[52] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_2_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_2_1  ( .A(\RI5[0][178] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[172] ), .ZN(\MC_ARK_ARC_1_0/temp1[178] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_2_0  ( .A(\MC_ARK_ARC_1_0/temp2[179] ), .B(
        \MC_ARK_ARC_1_0/temp1[179] ), .ZN(\MC_ARK_ARC_1_0/temp5[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_2_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[23] ), 
        .B(n274), .ZN(\MC_ARK_ARC_1_0/temp4[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_2_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[89] ), 
        .B(n1632), .ZN(\MC_ARK_ARC_1_0/temp3[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_2_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[149] ), 
        .B(n1938), .ZN(\MC_ARK_ARC_1_0/temp2[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_2_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[173] ), 
        .B(n1659), .ZN(\MC_ARK_ARC_1_0/temp1[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_1_5  ( .A(\MC_ARK_ARC_1_0/temp5[180] ), .B(
        \MC_ARK_ARC_1_0/temp6[180] ), .ZN(\RI1[1][180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_1_5  ( .A(\MC_ARK_ARC_1_0/temp3[180] ), .B(
        \MC_ARK_ARC_1_0/temp4[180] ), .ZN(\MC_ARK_ARC_1_0/temp6[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_1_5  ( .A(\MC_ARK_ARC_1_0/temp1[180] ), .B(
        \MC_ARK_ARC_1_0/temp2[180] ), .ZN(\MC_ARK_ARC_1_0/temp5[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_1_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[24] ), 
        .B(n267), .ZN(\MC_ARK_ARC_1_0/temp4[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_1_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[54] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_1_5  ( .A(\RI5[0][150] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[126] ), .ZN(\MC_ARK_ARC_1_0/temp2[180] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_1_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .B(\RI5[0][174] ), .ZN(\MC_ARK_ARC_1_0/temp1[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_1_4  ( .A(\MC_ARK_ARC_1_0/temp6[181] ), .B(
        \MC_ARK_ARC_1_0/temp5[181] ), .ZN(\RI1[1][181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_1_4  ( .A(\MC_ARK_ARC_1_0/temp3[181] ), .B(
        \MC_ARK_ARC_1_0/temp4[181] ), .ZN(\MC_ARK_ARC_1_0/temp6[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_1_4  ( .A(\MC_ARK_ARC_1_0/temp1[181] ), .B(
        \MC_ARK_ARC_1_0/temp2[181] ), .ZN(\MC_ARK_ARC_1_0/temp5[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_1_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[25] ), 
        .B(n260), .ZN(\MC_ARK_ARC_1_0/temp4[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_1_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[55] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_1_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[127] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_1_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_1_3  ( .A(\MC_ARK_ARC_1_0/temp5[182] ), .B(
        \MC_ARK_ARC_1_0/temp6[182] ), .ZN(\RI1[1][182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_1_3  ( .A(\MC_ARK_ARC_1_0/temp3[182] ), .B(
        \MC_ARK_ARC_1_0/temp4[182] ), .ZN(\MC_ARK_ARC_1_0/temp6[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_1_3  ( .A(\MC_ARK_ARC_1_0/temp1[182] ), .B(
        \MC_ARK_ARC_1_0/temp2[182] ), .ZN(\MC_ARK_ARC_1_0/temp5[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_1_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[26] ), 
        .B(Key[127]), .ZN(\MC_ARK_ARC_1_0/temp4[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_1_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[56] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[92] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_1_3  ( .A(\RI5[0][152] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[128] ), .ZN(\MC_ARK_ARC_1_0/temp2[182] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_1_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_1_2  ( .A(\MC_ARK_ARC_1_0/temp5[183] ), .B(
        \MC_ARK_ARC_1_0/temp6[183] ), .ZN(\RI1[1][183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_1_2  ( .A(\MC_ARK_ARC_1_0/temp3[183] ), .B(
        \MC_ARK_ARC_1_0/temp4[183] ), .ZN(\MC_ARK_ARC_1_0/temp6[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_1_2  ( .A(\MC_ARK_ARC_1_0/temp1[183] ), .B(
        \MC_ARK_ARC_1_0/temp2[183] ), .ZN(\MC_ARK_ARC_1_0/temp5[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_1_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[27] ), 
        .B(n451), .ZN(\MC_ARK_ARC_1_0/temp4[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_1_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[93] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[57] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_1_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[153] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[129] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_1_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[177] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[183] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_1_1  ( .A(\MC_ARK_ARC_1_0/temp5[184] ), .B(
        \MC_ARK_ARC_1_0/temp6[184] ), .ZN(\RI1[1][184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_1_1  ( .A(\MC_ARK_ARC_1_0/temp3[184] ), .B(
        \MC_ARK_ARC_1_0/temp4[184] ), .ZN(\MC_ARK_ARC_1_0/temp6[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_1_1  ( .A(\MC_ARK_ARC_1_0/temp1[184] ), .B(
        \MC_ARK_ARC_1_0/temp2[184] ), .ZN(\MC_ARK_ARC_1_0/temp5[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_1_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[28] ), 
        .B(n513), .ZN(\MC_ARK_ARC_1_0/temp4[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_1_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[58] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_1_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_1_1  ( .A(\RI5[0][184] ), .B(\RI5[0][178] ), 
        .ZN(\MC_ARK_ARC_1_0/temp1[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_1_0  ( .A(\MC_ARK_ARC_1_0/temp2[185] ), .B(
        \MC_ARK_ARC_1_0/temp1[185] ), .ZN(\MC_ARK_ARC_1_0/temp5[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_1_0  ( .A(n1470), .B(n491), .ZN(
        \MC_ARK_ARC_1_0/temp4[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_1_0  ( .A(n787), .B(
        \MC_ARK_ARC_1_0/buf_datainput[95] ), .ZN(\MC_ARK_ARC_1_0/temp3[185] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_1_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[131] ), 
        .B(n2117), .ZN(\MC_ARK_ARC_1_0/temp2[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_1_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[179] ), 
        .B(n794), .ZN(\MC_ARK_ARC_1_0/temp1[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_0_5  ( .A(\MC_ARK_ARC_1_0/temp5[186] ), .B(
        \MC_ARK_ARC_1_0/temp6[186] ), .ZN(\RI1[1][186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_0_5  ( .A(\MC_ARK_ARC_1_0/temp3[186] ), .B(
        \MC_ARK_ARC_1_0/temp4[186] ), .ZN(\MC_ARK_ARC_1_0/temp6[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_0_5  ( .A(\MC_ARK_ARC_1_0/temp1[186] ), .B(
        \MC_ARK_ARC_1_0/temp2[186] ), .ZN(\MC_ARK_ARC_1_0/temp5[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_0_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[30] ), 
        .B(n228), .ZN(\MC_ARK_ARC_1_0/temp4[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_0_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .B(\RI5[0][60] ), .ZN(\MC_ARK_ARC_1_0/temp3[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_0_5  ( .A(\RI5[0][156] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[132] ), .ZN(\MC_ARK_ARC_1_0/temp2[186] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_0_5  ( .A(\MC_ARK_ARC_1_0/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_0_4  ( .A(\MC_ARK_ARC_1_0/temp5[187] ), .B(
        \MC_ARK_ARC_1_0/temp6[187] ), .ZN(\RI1[1][187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_0_4  ( .A(\MC_ARK_ARC_1_0/temp3[187] ), .B(
        \MC_ARK_ARC_1_0/temp4[187] ), .ZN(\MC_ARK_ARC_1_0/temp6[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_0_4  ( .A(\MC_ARK_ARC_1_0/temp1[187] ), .B(
        \MC_ARK_ARC_1_0/temp2[187] ), .ZN(\MC_ARK_ARC_1_0/temp5[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_0_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_0/buf_keyinput[187] ), .ZN(
        \MC_ARK_ARC_1_0/temp4[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_0_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[61] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_0_4  ( .A(\RI5[0][157] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[133] ), .ZN(\MC_ARK_ARC_1_0/temp2[187] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_0_4  ( .A(\MC_ARK_ARC_1_0/buf_datainput[187] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_0_3  ( .A(\MC_ARK_ARC_1_0/temp5[188] ), .B(
        \MC_ARK_ARC_1_0/temp6[188] ), .ZN(\RI1[1][188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_0_3  ( .A(\MC_ARK_ARC_1_0/temp3[188] ), .B(
        \MC_ARK_ARC_1_0/temp4[188] ), .ZN(\MC_ARK_ARC_1_0/temp6[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_0_3  ( .A(\MC_ARK_ARC_1_0/temp1[188] ), .B(
        \MC_ARK_ARC_1_0/temp2[188] ), .ZN(\MC_ARK_ARC_1_0/temp5[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_0_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[32] ), 
        .B(n433), .ZN(\MC_ARK_ARC_1_0/temp4[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_0_3  ( .A(\RI5[0][62] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[98] ), .ZN(\MC_ARK_ARC_1_0/temp3[188] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_0_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[134] ), 
        .B(n2137), .ZN(\MC_ARK_ARC_1_0/temp2[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_0_3  ( .A(\MC_ARK_ARC_1_0/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[188] ), .ZN(
        \MC_ARK_ARC_1_0/temp1[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_0_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[33] ), 
        .B(n207), .ZN(\MC_ARK_ARC_1_0/temp4[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_0_2  ( .A(\RI5[0][63] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[99] ), .ZN(\MC_ARK_ARC_1_0/temp3[189] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_0_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[159] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[135] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_0_2  ( .A(\MC_ARK_ARC_1_0/buf_datainput[183] ), 
        .B(n1495), .ZN(\MC_ARK_ARC_1_0/temp1[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X7_0_1  ( .A(\MC_ARK_ARC_1_0/temp5[190] ), .B(
        \MC_ARK_ARC_1_0/temp6[190] ), .ZN(\RI1[1][190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X6_0_1  ( .A(\MC_ARK_ARC_1_0/temp3[190] ), .B(
        \MC_ARK_ARC_1_0/temp4[190] ), .ZN(\MC_ARK_ARC_1_0/temp6[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X5_0_1  ( .A(\MC_ARK_ARC_1_0/temp1[190] ), .B(
        \MC_ARK_ARC_1_0/temp2[190] ), .ZN(\MC_ARK_ARC_1_0/temp5[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_0_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[34] ), 
        .B(n508), .ZN(\MC_ARK_ARC_1_0/temp4[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_0_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_0_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[136] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_0_1  ( .A(\MC_ARK_ARC_1_0/buf_datainput[190] ), 
        .B(\RI5[0][184] ), .ZN(\MC_ARK_ARC_1_0/temp1[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X4_0_0  ( .A(n1508), .B(n430), .ZN(
        \MC_ARK_ARC_1_0/temp4[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X3_0_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[101] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[65] ), .ZN(
        \MC_ARK_ARC_1_0/temp3[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X2_0_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_0/buf_datainput[161] ), .ZN(
        \MC_ARK_ARC_1_0/temp2[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_0/X1_0_0  ( .A(\MC_ARK_ARC_1_0/buf_datainput[191] ), 
        .B(n794), .ZN(\MC_ARK_ARC_1_0/temp1[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_31_5  ( .A(\MC_ARK_ARC_1_1/temp5[0] ), .B(
        \MC_ARK_ARC_1_1/temp6[0] ), .ZN(\RI1[2][0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_31_5  ( .A(\MC_ARK_ARC_1_1/temp3[0] ), .B(
        \MC_ARK_ARC_1_1/temp4[0] ), .ZN(\MC_ARK_ARC_1_1/temp6[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_31_5  ( .A(\MC_ARK_ARC_1_1/temp1[0] ), .B(
        \MC_ARK_ARC_1_1/temp2[0] ), .ZN(\MC_ARK_ARC_1_1/temp5[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_31_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[36] ), 
        .B(n469), .ZN(\MC_ARK_ARC_1_1/temp4[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_31_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[66] ), .ZN(\MC_ARK_ARC_1_1/temp3[0] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_31_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[162] ), 
        .B(\RI5[1][138] ), .ZN(\MC_ARK_ARC_1_1/temp2[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_31_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[186] ), .ZN(\MC_ARK_ARC_1_1/temp1[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_31_4  ( .A(\MC_ARK_ARC_1_1/temp5[1] ), .B(
        \MC_ARK_ARC_1_1/temp6[1] ), .ZN(\RI1[2][1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_31_4  ( .A(\MC_ARK_ARC_1_1/temp3[1] ), .B(
        \MC_ARK_ARC_1_1/temp4[1] ), .ZN(\MC_ARK_ARC_1_1/temp6[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_31_4  ( .A(\MC_ARK_ARC_1_1/temp1[1] ), .B(
        \MC_ARK_ARC_1_1/temp2[1] ), .ZN(\MC_ARK_ARC_1_1/temp5[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_31_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[37] ), 
        .B(n390), .ZN(\MC_ARK_ARC_1_1/temp4[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_31_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[67] ), .ZN(\MC_ARK_ARC_1_1/temp3[1] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_31_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[139] ), .ZN(\MC_ARK_ARC_1_1/temp2[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_31_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[187] ), .ZN(\MC_ARK_ARC_1_1/temp1[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_31_3  ( .A(\MC_ARK_ARC_1_1/temp5[2] ), .B(
        \MC_ARK_ARC_1_1/temp6[2] ), .ZN(\RI1[2][2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_31_3  ( .A(\MC_ARK_ARC_1_1/temp3[2] ), .B(
        \MC_ARK_ARC_1_1/temp4[2] ), .ZN(\MC_ARK_ARC_1_1/temp6[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_31_3  ( .A(\MC_ARK_ARC_1_1/temp1[2] ), .B(
        \MC_ARK_ARC_1_1/temp2[2] ), .ZN(\MC_ARK_ARC_1_1/temp5[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_31_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .B(n244), .ZN(\MC_ARK_ARC_1_1/temp4[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_31_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[68] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[104] ), .ZN(\MC_ARK_ARC_1_1/temp3[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_31_3  ( .A(n1624), .B(
        \MC_ARK_ARC_1_1/buf_datainput[140] ), .ZN(\MC_ARK_ARC_1_1/temp2[2] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_31_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_1/temp1[2] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_31_2  ( .A(\MC_ARK_ARC_1_1/temp5[3] ), .B(
        \MC_ARK_ARC_1_1/temp6[3] ), .ZN(\RI1[2][3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_31_2  ( .A(\MC_ARK_ARC_1_1/temp3[3] ), .B(
        \MC_ARK_ARC_1_1/temp4[3] ), .ZN(\MC_ARK_ARC_1_1/temp6[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_31_2  ( .A(\MC_ARK_ARC_1_1/temp2[3] ), .B(
        \MC_ARK_ARC_1_1/temp1[3] ), .ZN(\MC_ARK_ARC_1_1/temp5[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_31_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[39] ), 
        .B(n197), .ZN(\MC_ARK_ARC_1_1/temp4[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_31_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[69] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[105] ), .ZN(\MC_ARK_ARC_1_1/temp3[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_31_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[165] ), 
        .B(\RI5[1][141] ), .ZN(\MC_ARK_ARC_1_1/temp2[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_31_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[3] ), 
        .B(n1935), .ZN(\MC_ARK_ARC_1_1/temp1[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_31_1  ( .A(\MC_ARK_ARC_1_1/temp5[4] ), .B(
        \MC_ARK_ARC_1_1/temp6[4] ), .ZN(\RI1[2][4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_31_1  ( .A(\MC_ARK_ARC_1_1/temp3[4] ), .B(
        \MC_ARK_ARC_1_1/temp4[4] ), .ZN(\MC_ARK_ARC_1_1/temp6[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_31_1  ( .A(\MC_ARK_ARC_1_1/temp2[4] ), .B(
        \MC_ARK_ARC_1_1/temp1[4] ), .ZN(\MC_ARK_ARC_1_1/temp5[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_31_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[40] ), 
        .B(n475), .ZN(\MC_ARK_ARC_1_1/temp4[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_31_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[106] ), .ZN(\MC_ARK_ARC_1_1/temp3[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_31_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[142] ), .ZN(\MC_ARK_ARC_1_1/temp2[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_31_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[190] ), .ZN(\MC_ARK_ARC_1_1/temp1[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_31_0  ( .A(\MC_ARK_ARC_1_1/temp5[5] ), .B(
        \MC_ARK_ARC_1_1/temp6[5] ), .ZN(\RI1[2][5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_31_0  ( .A(\MC_ARK_ARC_1_1/temp3[5] ), .B(
        \MC_ARK_ARC_1_1/temp4[5] ), .ZN(\MC_ARK_ARC_1_1/temp6[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_31_0  ( .A(\MC_ARK_ARC_1_1/temp2[5] ), .B(
        \MC_ARK_ARC_1_1/temp1[5] ), .ZN(\MC_ARK_ARC_1_1/temp5[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_31_0  ( .A(n1497), .B(n286), .ZN(
        \MC_ARK_ARC_1_1/temp4[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_31_0  ( .A(n1952), .B(
        \MC_ARK_ARC_1_1/buf_datainput[107] ), .ZN(\MC_ARK_ARC_1_1/temp3[5] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_31_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[167] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[143] ), .ZN(\MC_ARK_ARC_1_1/temp2[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_31_0  ( .A(n1641), .B(n515), .ZN(
        \MC_ARK_ARC_1_1/temp1[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_30_5  ( .A(\MC_ARK_ARC_1_1/temp5[6] ), .B(
        \MC_ARK_ARC_1_1/temp6[6] ), .ZN(\RI1[2][6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_30_5  ( .A(\MC_ARK_ARC_1_1/temp3[6] ), .B(
        \MC_ARK_ARC_1_1/temp4[6] ), .ZN(\MC_ARK_ARC_1_1/temp6[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_30_5  ( .A(\MC_ARK_ARC_1_1/temp1[6] ), .B(
        \MC_ARK_ARC_1_1/temp2[6] ), .ZN(\MC_ARK_ARC_1_1/temp5[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_30_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[42] ), 
        .B(n241), .ZN(\MC_ARK_ARC_1_1/temp4[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_30_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[108] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[72] ), .ZN(\MC_ARK_ARC_1_1/temp3[6] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_30_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[144] ), .ZN(\MC_ARK_ARC_1_1/temp2[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_30_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_1/temp1[6] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_30_4  ( .A(\MC_ARK_ARC_1_1/temp5[7] ), .B(
        \MC_ARK_ARC_1_1/temp6[7] ), .ZN(\RI1[2][7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_30_4  ( .A(\MC_ARK_ARC_1_1/temp3[7] ), .B(
        \MC_ARK_ARC_1_1/temp4[7] ), .ZN(\MC_ARK_ARC_1_1/temp6[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_30_4  ( .A(\MC_ARK_ARC_1_1/temp1[7] ), .B(
        \MC_ARK_ARC_1_1/temp2[7] ), .ZN(\MC_ARK_ARC_1_1/temp5[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_30_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[43] ), 
        .B(n406), .ZN(\MC_ARK_ARC_1_1/temp4[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_30_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[73] ), .ZN(\MC_ARK_ARC_1_1/temp3[7] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_30_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[169] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[145] ), .ZN(\MC_ARK_ARC_1_1/temp2[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_30_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[7] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[1] ), .ZN(\MC_ARK_ARC_1_1/temp1[7] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_30_3  ( .A(\MC_ARK_ARC_1_1/temp5[8] ), .B(
        \MC_ARK_ARC_1_1/temp6[8] ), .ZN(\RI1[2][8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_30_3  ( .A(\MC_ARK_ARC_1_1/temp3[8] ), .B(
        \MC_ARK_ARC_1_1/temp4[8] ), .ZN(\MC_ARK_ARC_1_1/temp6[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_30_3  ( .A(\MC_ARK_ARC_1_1/temp2[8] ), .B(
        \MC_ARK_ARC_1_1/temp1[8] ), .ZN(\MC_ARK_ARC_1_1/temp5[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_30_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[44] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[8] ), .ZN(\MC_ARK_ARC_1_1/temp4[8] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_30_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[110] ), .ZN(\MC_ARK_ARC_1_1/temp3[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_30_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[170] ), .ZN(\MC_ARK_ARC_1_1/temp2[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_30_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[8] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_1/temp1[8] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_30_2  ( .A(\MC_ARK_ARC_1_1/temp6[9] ), .B(
        \MC_ARK_ARC_1_1/temp5[9] ), .ZN(\RI1[2][9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_30_2  ( .A(\MC_ARK_ARC_1_1/temp3[9] ), .B(
        \MC_ARK_ARC_1_1/temp4[9] ), .ZN(\MC_ARK_ARC_1_1/temp6[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_30_2  ( .A(\MC_ARK_ARC_1_1/temp1[9] ), .B(
        \MC_ARK_ARC_1_1/temp2[9] ), .ZN(\MC_ARK_ARC_1_1/temp5[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_30_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[45] ), 
        .B(n457), .ZN(\MC_ARK_ARC_1_1/temp4[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_30_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[111] ), 
        .B(\RI5[1][75] ), .ZN(\MC_ARK_ARC_1_1/temp3[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_30_2  ( .A(\RI5[1][147] ), .B(n1954), .ZN(
        \MC_ARK_ARC_1_1/temp2[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_30_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[3] ), 
        .B(\RI5[1][9] ), .ZN(\MC_ARK_ARC_1_1/temp1[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_30_1  ( .A(\MC_ARK_ARC_1_1/temp5[10] ), .B(
        \MC_ARK_ARC_1_1/temp6[10] ), .ZN(\RI1[2][10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_30_1  ( .A(\MC_ARK_ARC_1_1/temp3[10] ), .B(
        \MC_ARK_ARC_1_1/temp4[10] ), .ZN(\MC_ARK_ARC_1_1/temp6[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_30_1  ( .A(\MC_ARK_ARC_1_1/temp2[10] ), .B(
        \MC_ARK_ARC_1_1/temp1[10] ), .ZN(\MC_ARK_ARC_1_1/temp5[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_30_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[46] ), 
        .B(n237), .ZN(\MC_ARK_ARC_1_1/temp4[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_30_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[76] ), .ZN(\MC_ARK_ARC_1_1/temp3[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_30_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[148] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_30_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_1/temp1[10] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_30_0  ( .A(\MC_ARK_ARC_1_1/temp5[11] ), .B(
        \MC_ARK_ARC_1_1/temp6[11] ), .ZN(\RI1[2][11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_30_0  ( .A(\MC_ARK_ARC_1_1/temp2[11] ), .B(
        \MC_ARK_ARC_1_1/temp1[11] ), .ZN(\MC_ARK_ARC_1_1/temp5[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_30_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[47] ), 
        .B(n371), .ZN(\MC_ARK_ARC_1_1/temp4[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_30_0  ( .A(n1937), .B(
        \MC_ARK_ARC_1_1/buf_datainput[149] ), .ZN(\MC_ARK_ARC_1_1/temp2[11] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_30_0  ( .A(n1641), .B(n2105), .ZN(
        \MC_ARK_ARC_1_1/temp1[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_29_5  ( .A(\MC_ARK_ARC_1_1/temp5[12] ), .B(
        \MC_ARK_ARC_1_1/temp6[12] ), .ZN(\RI1[2][12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_29_5  ( .A(\MC_ARK_ARC_1_1/temp3[12] ), .B(
        \MC_ARK_ARC_1_1/temp4[12] ), .ZN(\MC_ARK_ARC_1_1/temp6[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_29_5  ( .A(\MC_ARK_ARC_1_1/temp1[12] ), .B(
        \MC_ARK_ARC_1_1/temp2[12] ), .ZN(\MC_ARK_ARC_1_1/temp5[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_29_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[48] ), 
        .B(n375), .ZN(\MC_ARK_ARC_1_1/temp4[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_29_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[78] ), .ZN(\MC_ARK_ARC_1_1/temp3[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_29_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[174] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[150] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_29_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_1/temp1[12] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_29_4  ( .A(\MC_ARK_ARC_1_1/temp5[13] ), .B(
        \MC_ARK_ARC_1_1/temp6[13] ), .ZN(\RI1[2][13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_29_4  ( .A(\MC_ARK_ARC_1_1/temp3[13] ), .B(
        \MC_ARK_ARC_1_1/temp4[13] ), .ZN(\MC_ARK_ARC_1_1/temp6[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_29_4  ( .A(\MC_ARK_ARC_1_1/temp1[13] ), .B(
        \MC_ARK_ARC_1_1/temp2[13] ), .ZN(\MC_ARK_ARC_1_1/temp5[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_29_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[49] ), 
        .B(n494), .ZN(\MC_ARK_ARC_1_1/temp4[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_29_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[79] ), .ZN(\MC_ARK_ARC_1_1/temp3[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_29_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[151] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_29_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_1/temp1[13] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_29_3  ( .A(\MC_ARK_ARC_1_1/temp5[14] ), .B(
        \MC_ARK_ARC_1_1/temp6[14] ), .ZN(\RI1[2][14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_29_3  ( .A(\MC_ARK_ARC_1_1/temp3[14] ), .B(
        \MC_ARK_ARC_1_1/temp4[14] ), .ZN(\MC_ARK_ARC_1_1/temp6[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_29_3  ( .A(\MC_ARK_ARC_1_1/temp1[14] ), .B(
        \MC_ARK_ARC_1_1/temp2[14] ), .ZN(\MC_ARK_ARC_1_1/temp5[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_29_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[70] ), .ZN(\MC_ARK_ARC_1_1/temp4[14] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_29_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[80] ), .ZN(\MC_ARK_ARC_1_1/temp3[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_29_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_29_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_1/temp1[14] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_29_2  ( .A(\MC_ARK_ARC_1_1/temp5[15] ), .B(
        \MC_ARK_ARC_1_1/temp6[15] ), .ZN(\RI1[2][15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_29_2  ( .A(\MC_ARK_ARC_1_1/temp3[15] ), .B(
        \MC_ARK_ARC_1_1/temp4[15] ), .ZN(\MC_ARK_ARC_1_1/temp6[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_29_2  ( .A(\MC_ARK_ARC_1_1/temp1[15] ), .B(
        \MC_ARK_ARC_1_1/temp2[15] ), .ZN(\MC_ARK_ARC_1_1/temp5[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_29_2  ( .A(\RI5[1][51] ), .B(n468), .ZN(
        \MC_ARK_ARC_1_1/temp4[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_29_2  ( .A(\RI5[1][117] ), .B(\RI5[1][81] ), 
        .ZN(\MC_ARK_ARC_1_1/temp3[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_29_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .B(\RI5[1][177] ), .ZN(\MC_ARK_ARC_1_1/temp2[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_29_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .B(\RI5[1][9] ), .ZN(\MC_ARK_ARC_1_1/temp1[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_29_1  ( .A(\MC_ARK_ARC_1_1/temp6[16] ), .B(
        \MC_ARK_ARC_1_1/temp5[16] ), .ZN(\RI1[2][16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_29_1  ( .A(\MC_ARK_ARC_1_1/temp4[16] ), .B(
        \MC_ARK_ARC_1_1/temp3[16] ), .ZN(\MC_ARK_ARC_1_1/temp6[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_29_1  ( .A(\MC_ARK_ARC_1_1/temp1[16] ), .B(
        \MC_ARK_ARC_1_1/temp2[16] ), .ZN(\MC_ARK_ARC_1_1/temp5[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_29_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[52] ), 
        .B(n321), .ZN(\MC_ARK_ARC_1_1/temp4[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_29_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[118] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[82] ), .ZN(\MC_ARK_ARC_1_1/temp3[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_29_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[154] ), 
        .B(n1953), .ZN(\MC_ARK_ARC_1_1/temp2[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_29_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_1/temp1[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_29_0  ( .A(n838), .B(n495), .ZN(
        \MC_ARK_ARC_1_1/temp4[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_29_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[119] ), 
        .B(n813), .ZN(\MC_ARK_ARC_1_1/temp3[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_29_0  ( .A(n2153), .B(
        \MC_ARK_ARC_1_1/buf_datainput[179] ), .ZN(\MC_ARK_ARC_1_1/temp2[17] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_29_0  ( .A(n2105), .B(n1642), .ZN(
        \MC_ARK_ARC_1_1/temp1[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_28_5  ( .A(\MC_ARK_ARC_1_1/temp5[18] ), .B(
        \MC_ARK_ARC_1_1/temp6[18] ), .ZN(\RI1[2][18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_28_5  ( .A(\MC_ARK_ARC_1_1/temp3[18] ), .B(
        \MC_ARK_ARC_1_1/temp4[18] ), .ZN(\MC_ARK_ARC_1_1/temp6[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_28_5  ( .A(\MC_ARK_ARC_1_1/temp1[18] ), .B(
        \MC_ARK_ARC_1_1/temp2[18] ), .ZN(\MC_ARK_ARC_1_1/temp5[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_28_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[54] ), 
        .B(n489), .ZN(\MC_ARK_ARC_1_1/temp4[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_28_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[84] ), .ZN(\MC_ARK_ARC_1_1/temp3[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_28_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[180] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[156] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_28_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_1/temp1[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_28_4  ( .A(\MC_ARK_ARC_1_1/temp5[19] ), .B(
        \MC_ARK_ARC_1_1/temp6[19] ), .ZN(\RI1[2][19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_28_4  ( .A(\MC_ARK_ARC_1_1/temp4[19] ), .B(
        \MC_ARK_ARC_1_1/temp3[19] ), .ZN(\MC_ARK_ARC_1_1/temp6[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_28_4  ( .A(\MC_ARK_ARC_1_1/temp1[19] ), .B(
        \MC_ARK_ARC_1_1/temp2[19] ), .ZN(\MC_ARK_ARC_1_1/temp5[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_28_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[55] ), 
        .B(n364), .ZN(\MC_ARK_ARC_1_1/temp4[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_28_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[85] ), .ZN(\MC_ARK_ARC_1_1/temp3[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_28_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[157] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_28_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[13] ), .ZN(\MC_ARK_ARC_1_1/temp1[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_28_3  ( .A(\MC_ARK_ARC_1_1/temp5[20] ), .B(
        \MC_ARK_ARC_1_1/temp6[20] ), .ZN(\RI1[2][20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_28_3  ( .A(\MC_ARK_ARC_1_1/temp3[20] ), .B(
        \MC_ARK_ARC_1_1/temp4[20] ), .ZN(\MC_ARK_ARC_1_1/temp6[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_28_3  ( .A(\MC_ARK_ARC_1_1/temp1[20] ), .B(
        \MC_ARK_ARC_1_1/temp2[20] ), .ZN(\MC_ARK_ARC_1_1/temp5[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_28_3  ( .A(\RI5[1][56] ), .B(
        \MC_ARK_ARC_1_3/buf_keyinput[172] ), .ZN(\MC_ARK_ARC_1_1/temp4[20] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_28_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[86] ), .ZN(\MC_ARK_ARC_1_1/temp3[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_28_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[158] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_28_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_1/temp1[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_28_2  ( .A(\MC_ARK_ARC_1_1/temp2[21] ), .B(
        \MC_ARK_ARC_1_1/temp1[21] ), .ZN(\MC_ARK_ARC_1_1/temp5[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_28_2  ( .A(\RI5[1][57] ), .B(n271), .ZN(
        \MC_ARK_ARC_1_1/temp4[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_28_2  ( .A(\RI5[1][123] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[87] ), .ZN(\MC_ARK_ARC_1_1/temp3[21] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_28_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[159] ), 
        .B(n1486), .ZN(\MC_ARK_ARC_1_1/temp2[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_28_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_1/temp1[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_28_1  ( .A(\MC_ARK_ARC_1_1/temp6[22] ), .B(
        \MC_ARK_ARC_1_1/temp5[22] ), .ZN(\RI1[2][22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_28_1  ( .A(\MC_ARK_ARC_1_1/temp3[22] ), .B(
        \MC_ARK_ARC_1_1/temp4[22] ), .ZN(\MC_ARK_ARC_1_1/temp6[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_28_1  ( .A(\MC_ARK_ARC_1_1/temp2[22] ), .B(
        \MC_ARK_ARC_1_1/temp1[22] ), .ZN(\MC_ARK_ARC_1_1/temp5[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_28_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .B(n225), .ZN(\MC_ARK_ARC_1_1/temp4[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_28_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_28_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[184] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_28_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_1/temp1[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_28_0  ( .A(\MC_ARK_ARC_1_1/temp3[23] ), .B(
        \MC_ARK_ARC_1_1/temp4[23] ), .ZN(\MC_ARK_ARC_1_1/temp6[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_28_0  ( .A(\MC_ARK_ARC_1_1/temp2[23] ), .B(
        \MC_ARK_ARC_1_1/temp1[23] ), .ZN(\MC_ARK_ARC_1_1/temp5[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_28_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[59] ), 
        .B(n360), .ZN(\MC_ARK_ARC_1_1/temp4[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_28_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[125] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[89] ), .ZN(\MC_ARK_ARC_1_1/temp3[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_28_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[161] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[185] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_28_0  ( .A(n1926), .B(n1643), .ZN(
        \MC_ARK_ARC_1_1/temp1[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_27_5  ( .A(\MC_ARK_ARC_1_1/temp5[24] ), .B(
        \MC_ARK_ARC_1_1/temp6[24] ), .ZN(\RI1[2][24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_27_5  ( .A(\MC_ARK_ARC_1_1/temp3[24] ), .B(
        \MC_ARK_ARC_1_1/temp4[24] ), .ZN(\MC_ARK_ARC_1_1/temp6[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_27_5  ( .A(\MC_ARK_ARC_1_1/temp1[24] ), .B(
        \MC_ARK_ARC_1_1/temp2[24] ), .ZN(\MC_ARK_ARC_1_1/temp5[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_27_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[60] ), 
        .B(n455), .ZN(\MC_ARK_ARC_1_1/temp4[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_27_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[90] ), .ZN(\MC_ARK_ARC_1_1/temp3[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_27_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_27_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[18] ), .ZN(\MC_ARK_ARC_1_1/temp1[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_27_4  ( .A(\MC_ARK_ARC_1_1/temp5[25] ), .B(
        \MC_ARK_ARC_1_1/temp6[25] ), .ZN(\RI1[2][25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_27_4  ( .A(\MC_ARK_ARC_1_1/temp3[25] ), .B(
        \MC_ARK_ARC_1_1/temp4[25] ), .ZN(\MC_ARK_ARC_1_1/temp6[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_27_4  ( .A(\MC_ARK_ARC_1_1/temp1[25] ), .B(
        \MC_ARK_ARC_1_1/temp2[25] ), .ZN(\MC_ARK_ARC_1_1/temp5[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_27_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[61] ), 
        .B(n396), .ZN(\MC_ARK_ARC_1_1/temp4[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_27_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_1/temp3[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_27_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[163] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_27_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[19] ), .ZN(\MC_ARK_ARC_1_1/temp1[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_27_3  ( .A(\MC_ARK_ARC_1_1/temp5[26] ), .B(
        \MC_ARK_ARC_1_1/temp6[26] ), .ZN(\RI1[2][26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_27_3  ( .A(\MC_ARK_ARC_1_1/temp3[26] ), .B(
        \MC_ARK_ARC_1_1/temp4[26] ), .ZN(\MC_ARK_ARC_1_1/temp6[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_27_3  ( .A(\MC_ARK_ARC_1_1/temp1[26] ), .B(
        \MC_ARK_ARC_1_1/temp2[26] ), .ZN(\MC_ARK_ARC_1_1/temp5[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_27_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .B(n221), .ZN(\MC_ARK_ARC_1_1/temp4[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_27_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_27_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .B(n1625), .ZN(\MC_ARK_ARC_1_1/temp2[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_27_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_1/temp1[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_27_2  ( .A(\MC_ARK_ARC_1_1/temp6[27] ), .B(
        \MC_ARK_ARC_1_1/temp5[27] ), .ZN(\RI1[2][27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_27_2  ( .A(\MC_ARK_ARC_1_1/temp3[27] ), .B(
        \MC_ARK_ARC_1_1/temp4[27] ), .ZN(\MC_ARK_ARC_1_1/temp6[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_27_2  ( .A(\MC_ARK_ARC_1_1/temp2[27] ), .B(
        \MC_ARK_ARC_1_1/temp1[27] ), .ZN(\MC_ARK_ARC_1_1/temp5[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_27_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[27] ), .ZN(\MC_ARK_ARC_1_1/temp4[27] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_27_2  ( .A(\RI5[1][93] ), .B(\RI5[1][129] ), 
        .ZN(\MC_ARK_ARC_1_1/temp3[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_27_2  ( .A(n1935), .B(
        \MC_ARK_ARC_1_1/buf_datainput[165] ), .ZN(\MC_ARK_ARC_1_1/temp2[27] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_27_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_1/temp1[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_27_1  ( .A(\MC_ARK_ARC_1_1/temp5[28] ), .B(
        \MC_ARK_ARC_1_1/temp6[28] ), .ZN(\RI1[2][28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_27_1  ( .A(\MC_ARK_ARC_1_1/temp3[28] ), .B(
        \MC_ARK_ARC_1_1/temp4[28] ), .ZN(\MC_ARK_ARC_1_1/temp6[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_27_1  ( .A(\MC_ARK_ARC_1_1/temp1[28] ), .B(
        \MC_ARK_ARC_1_1/temp2[28] ), .ZN(\MC_ARK_ARC_1_1/temp5[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_27_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[64] ), 
        .B(n310), .ZN(\MC_ARK_ARC_1_1/temp4[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_27_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[130] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[94] ), .ZN(\MC_ARK_ARC_1_1/temp3[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_27_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[190] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_27_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[28] ), .ZN(\MC_ARK_ARC_1_1/temp1[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_27_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[65] ), 
        .B(n263), .ZN(\MC_ARK_ARC_1_1/temp4[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_27_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[131] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_27_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[167] ), 
        .B(n515), .ZN(\MC_ARK_ARC_1_1/temp2[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_27_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .B(n1927), .ZN(\MC_ARK_ARC_1_1/temp1[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_26_5  ( .A(\MC_ARK_ARC_1_1/temp6[30] ), .B(
        \MC_ARK_ARC_1_1/temp5[30] ), .ZN(\RI1[2][30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_26_5  ( .A(\MC_ARK_ARC_1_1/temp3[30] ), .B(
        \MC_ARK_ARC_1_1/temp4[30] ), .ZN(\MC_ARK_ARC_1_1/temp6[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_26_5  ( .A(\MC_ARK_ARC_1_1/temp1[30] ), .B(
        \MC_ARK_ARC_1_1/temp2[30] ), .ZN(\MC_ARK_ARC_1_1/temp5[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_26_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[66] ), 
        .B(n431), .ZN(\MC_ARK_ARC_1_1/temp4[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_26_5  ( .A(\RI5[1][132] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[96] ), .ZN(\MC_ARK_ARC_1_1/temp3[30] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_26_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_26_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[24] ), .ZN(\MC_ARK_ARC_1_1/temp1[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_26_4  ( .A(\MC_ARK_ARC_1_1/temp5[31] ), .B(
        \MC_ARK_ARC_1_1/temp6[31] ), .ZN(\RI1[2][31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_26_4  ( .A(\MC_ARK_ARC_1_1/temp3[31] ), .B(
        \MC_ARK_ARC_1_1/temp4[31] ), .ZN(\MC_ARK_ARC_1_1/temp6[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_26_4  ( .A(\MC_ARK_ARC_1_1/temp1[31] ), .B(
        \MC_ARK_ARC_1_1/temp2[31] ), .ZN(\MC_ARK_ARC_1_1/temp5[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_26_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[67] ), 
        .B(n465), .ZN(\MC_ARK_ARC_1_1/temp4[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_26_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[133] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[97] ), .ZN(\MC_ARK_ARC_1_1/temp3[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_26_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[169] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_26_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[25] ), .ZN(\MC_ARK_ARC_1_1/temp1[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_26_3  ( .A(\MC_ARK_ARC_1_1/temp5[32] ), .B(
        \MC_ARK_ARC_1_1/temp6[32] ), .ZN(\RI1[2][32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_26_3  ( .A(\MC_ARK_ARC_1_1/temp3[32] ), .B(
        \MC_ARK_ARC_1_1/temp4[32] ), .ZN(\MC_ARK_ARC_1_1/temp6[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_26_3  ( .A(\MC_ARK_ARC_1_1/temp1[32] ), .B(
        \MC_ARK_ARC_1_1/temp2[32] ), .ZN(\MC_ARK_ARC_1_1/temp5[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_26_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[68] ), 
        .B(n306), .ZN(\MC_ARK_ARC_1_1/temp4[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_26_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[98] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[134] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_26_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[170] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_1/temp2[32] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_26_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[32] ), .ZN(\MC_ARK_ARC_1_1/temp1[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_26_2  ( .A(\MC_ARK_ARC_1_1/temp5[33] ), .B(
        \MC_ARK_ARC_1_1/temp6[33] ), .ZN(\RI1[2][33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_26_2  ( .A(\MC_ARK_ARC_1_1/temp3[33] ), .B(
        \MC_ARK_ARC_1_1/temp4[33] ), .ZN(\MC_ARK_ARC_1_1/temp6[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_26_2  ( .A(\MC_ARK_ARC_1_1/temp1[33] ), .B(
        \MC_ARK_ARC_1_1/temp2[33] ), .ZN(\MC_ARK_ARC_1_1/temp5[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_26_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[69] ), 
        .B(n259), .ZN(\MC_ARK_ARC_1_1/temp4[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_26_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .B(\RI5[1][135] ), .ZN(\MC_ARK_ARC_1_1/temp3[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_26_2  ( .A(n1954), .B(
        \MC_ARK_ARC_1_1/buf_datainput[3] ), .ZN(\MC_ARK_ARC_1_1/temp2[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_26_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_1/temp1[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_26_1  ( .A(\MC_ARK_ARC_1_1/temp5[34] ), .B(
        \MC_ARK_ARC_1_1/temp6[34] ), .ZN(\RI1[2][34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_26_1  ( .A(\MC_ARK_ARC_1_1/temp3[34] ), .B(
        \MC_ARK_ARC_1_1/temp4[34] ), .ZN(\MC_ARK_ARC_1_1/temp6[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_26_1  ( .A(\MC_ARK_ARC_1_1/temp1[34] ), .B(
        \MC_ARK_ARC_1_1/temp2[34] ), .ZN(\MC_ARK_ARC_1_1/temp5[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_26_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[70] ), 
        .B(n213), .ZN(\MC_ARK_ARC_1_1/temp4[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_26_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[136] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_26_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_26_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[28] ), .ZN(\MC_ARK_ARC_1_1/temp1[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_26_0  ( .A(n1952), .B(n348), .ZN(
        \MC_ARK_ARC_1_1/temp4[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_26_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[137] ), 
        .B(n2125), .ZN(\MC_ARK_ARC_1_1/temp3[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_26_0  ( .A(n1937), .B(n1640), .ZN(
        \MC_ARK_ARC_1_1/temp2[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_26_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .B(n519), .ZN(\MC_ARK_ARC_1_1/temp1[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_25_5  ( .A(\MC_ARK_ARC_1_1/temp5[36] ), .B(
        \MC_ARK_ARC_1_1/temp6[36] ), .ZN(\RI1[2][36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_25_5  ( .A(\MC_ARK_ARC_1_1/temp3[36] ), .B(
        \MC_ARK_ARC_1_1/temp4[36] ), .ZN(\MC_ARK_ARC_1_1/temp6[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_25_5  ( .A(\MC_ARK_ARC_1_1/temp1[36] ), .B(
        \MC_ARK_ARC_1_1/temp2[36] ), .ZN(\MC_ARK_ARC_1_1/temp5[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_25_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[72] ), 
        .B(n458), .ZN(\MC_ARK_ARC_1_1/temp4[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_25_5  ( .A(\RI5[1][138] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[102] ), .ZN(\MC_ARK_ARC_1_1/temp3[36] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_25_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[174] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_25_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[30] ), .ZN(\MC_ARK_ARC_1_1/temp1[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_25_4  ( .A(\MC_ARK_ARC_1_1/temp5[37] ), .B(
        \MC_ARK_ARC_1_1/temp6[37] ), .ZN(\RI1[2][37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_25_4  ( .A(\MC_ARK_ARC_1_1/temp3[37] ), .B(
        \MC_ARK_ARC_1_1/temp4[37] ), .ZN(\MC_ARK_ARC_1_1/temp6[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_25_4  ( .A(\MC_ARK_ARC_1_1/temp1[37] ), .B(
        \MC_ARK_ARC_1_1/temp2[37] ), .ZN(\MC_ARK_ARC_1_1/temp5[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_25_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .B(n445), .ZN(\MC_ARK_ARC_1_1/temp4[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_25_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_25_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[7] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_25_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[37] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[31] ), .ZN(\MC_ARK_ARC_1_1/temp1[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_25_3  ( .A(\MC_ARK_ARC_1_1/temp5[38] ), .B(
        \MC_ARK_ARC_1_1/temp6[38] ), .ZN(\RI1[2][38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_25_3  ( .A(\MC_ARK_ARC_1_1/temp3[38] ), .B(
        \MC_ARK_ARC_1_1/temp4[38] ), .ZN(\MC_ARK_ARC_1_1/temp6[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_25_3  ( .A(\MC_ARK_ARC_1_1/temp2[38] ), .B(
        \MC_ARK_ARC_1_1/temp1[38] ), .ZN(\MC_ARK_ARC_1_1/temp5[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_25_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[74] ), 
        .B(n209), .ZN(\MC_ARK_ARC_1_1/temp4[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_25_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_25_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[8] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_25_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_1/temp1[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_25_2  ( .A(\MC_ARK_ARC_1_1/temp1[39] ), .B(
        \MC_ARK_ARC_1_1/temp2[39] ), .ZN(\MC_ARK_ARC_1_1/temp5[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_25_2  ( .A(\RI5[1][75] ), .B(n344), .ZN(
        \MC_ARK_ARC_1_1/temp4[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_25_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[105] ), 
        .B(\RI5[1][141] ), .ZN(\MC_ARK_ARC_1_1/temp3[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_25_2  ( .A(\RI5[1][177] ), .B(\RI5[1][9] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_25_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[39] ), .ZN(\MC_ARK_ARC_1_1/temp1[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_25_1  ( .A(\MC_ARK_ARC_1_1/temp5[40] ), .B(
        \MC_ARK_ARC_1_1/temp6[40] ), .ZN(\RI1[2][40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_25_1  ( .A(\MC_ARK_ARC_1_1/temp3[40] ), .B(
        \MC_ARK_ARC_1_1/temp4[40] ), .ZN(\MC_ARK_ARC_1_1/temp6[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_25_1  ( .A(\MC_ARK_ARC_1_1/temp1[40] ), .B(
        \MC_ARK_ARC_1_1/temp2[40] ), .ZN(\MC_ARK_ARC_1_1/temp5[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_25_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[76] ), 
        .B(n512), .ZN(\MC_ARK_ARC_1_1/temp4[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_25_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[142] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_25_1  ( .A(n1953), .B(
        \MC_ARK_ARC_1_1/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_1/temp2[40] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_25_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[34] ), .ZN(\MC_ARK_ARC_1_1/temp1[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_25_0  ( .A(\MC_ARK_ARC_1_1/temp6[41] ), .B(
        \MC_ARK_ARC_1_1/temp5[41] ), .ZN(\RI1[2][41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_25_0  ( .A(\MC_ARK_ARC_1_1/temp4[41] ), .B(
        \MC_ARK_ARC_1_1/temp3[41] ), .ZN(\MC_ARK_ARC_1_1/temp6[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_25_0  ( .A(\MC_ARK_ARC_1_1/temp2[41] ), .B(
        \MC_ARK_ARC_1_1/temp1[41] ), .ZN(\MC_ARK_ARC_1_1/temp5[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_25_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[77] ), 
        .B(n251), .ZN(\MC_ARK_ARC_1_1/temp4[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_25_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[143] ), 
        .B(n852), .ZN(\MC_ARK_ARC_1_1/temp3[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_25_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[179] ), 
        .B(n2104), .ZN(\MC_ARK_ARC_1_1/temp2[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_25_0  ( .A(n1497), .B(n517), .ZN(
        \MC_ARK_ARC_1_1/temp1[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_24_5  ( .A(\MC_ARK_ARC_1_1/temp5[42] ), .B(
        \MC_ARK_ARC_1_1/temp6[42] ), .ZN(\RI1[2][42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_24_5  ( .A(\MC_ARK_ARC_1_1/temp3[42] ), .B(
        \MC_ARK_ARC_1_1/temp4[42] ), .ZN(\MC_ARK_ARC_1_1/temp6[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_24_5  ( .A(\MC_ARK_ARC_1_1/temp1[42] ), .B(
        \MC_ARK_ARC_1_1/temp2[42] ), .ZN(\MC_ARK_ARC_1_1/temp5[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_24_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[78] ), 
        .B(n205), .ZN(\MC_ARK_ARC_1_1/temp4[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_24_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[144] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[108] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_24_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_24_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[36] ), .ZN(\MC_ARK_ARC_1_1/temp1[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_24_4  ( .A(\MC_ARK_ARC_1_1/temp5[43] ), .B(
        \MC_ARK_ARC_1_1/temp6[43] ), .ZN(\RI1[2][43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_24_4  ( .A(\MC_ARK_ARC_1_1/temp3[43] ), .B(
        \MC_ARK_ARC_1_1/temp4[43] ), .ZN(\MC_ARK_ARC_1_1/temp6[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_24_4  ( .A(\MC_ARK_ARC_1_1/temp1[43] ), .B(
        \MC_ARK_ARC_1_1/temp2[43] ), .ZN(\MC_ARK_ARC_1_1/temp5[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_24_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[79] ), 
        .B(n407), .ZN(\MC_ARK_ARC_1_1/temp4[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_24_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_24_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_24_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[37] ), .ZN(\MC_ARK_ARC_1_1/temp1[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_24_3  ( .A(\MC_ARK_ARC_1_1/temp5[44] ), .B(
        \MC_ARK_ARC_1_1/temp6[44] ), .ZN(\RI1[2][44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_24_3  ( .A(\MC_ARK_ARC_1_1/temp3[44] ), .B(
        \MC_ARK_ARC_1_1/temp4[44] ), .ZN(\MC_ARK_ARC_1_1/temp6[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_24_3  ( .A(\MC_ARK_ARC_1_1/temp1[44] ), .B(
        \MC_ARK_ARC_1_1/temp2[44] ), .ZN(\MC_ARK_ARC_1_1/temp5[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_24_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[80] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[33] ), .ZN(\MC_ARK_ARC_1_1/temp4[44] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_24_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[110] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_24_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_24_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[44] ), .ZN(\MC_ARK_ARC_1_1/temp1[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_24_2  ( .A(\MC_ARK_ARC_1_1/temp5[45] ), .B(
        \MC_ARK_ARC_1_1/temp6[45] ), .ZN(\RI1[2][45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_24_2  ( .A(\MC_ARK_ARC_1_1/temp3[45] ), .B(
        \MC_ARK_ARC_1_1/temp4[45] ), .ZN(\MC_ARK_ARC_1_1/temp6[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_24_2  ( .A(\MC_ARK_ARC_1_1/temp2[45] ), .B(
        \MC_ARK_ARC_1_1/temp1[45] ), .ZN(\MC_ARK_ARC_1_1/temp5[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_24_2  ( .A(\RI5[1][81] ), .B(n248), .ZN(
        \MC_ARK_ARC_1_1/temp4[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_24_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[111] ), 
        .B(\RI5[1][147] ), .ZN(\MC_ARK_ARC_1_1/temp3[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_24_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .B(n1486), .ZN(\MC_ARK_ARC_1_1/temp2[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_24_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[39] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[45] ), .ZN(\MC_ARK_ARC_1_1/temp1[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_24_1  ( .A(\MC_ARK_ARC_1_1/temp5[46] ), .B(
        \MC_ARK_ARC_1_1/temp6[46] ), .ZN(\RI1[2][46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_24_1  ( .A(\MC_ARK_ARC_1_1/temp3[46] ), .B(
        \MC_ARK_ARC_1_1/temp4[46] ), .ZN(\MC_ARK_ARC_1_1/temp6[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_24_1  ( .A(\MC_ARK_ARC_1_1/temp2[46] ), .B(
        \MC_ARK_ARC_1_1/temp1[46] ), .ZN(\MC_ARK_ARC_1_1/temp5[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_24_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[82] ), 
        .B(n201), .ZN(\MC_ARK_ARC_1_1/temp4[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_24_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[112] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_24_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[184] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_24_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[46] ), .ZN(\MC_ARK_ARC_1_1/temp1[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_24_0  ( .A(\MC_ARK_ARC_1_1/temp5[47] ), .B(
        \MC_ARK_ARC_1_1/temp6[47] ), .ZN(\RI1[2][47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_24_0  ( .A(\MC_ARK_ARC_1_1/temp3[47] ), .B(
        \MC_ARK_ARC_1_1/temp4[47] ), .ZN(\MC_ARK_ARC_1_1/temp6[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_24_0  ( .A(\MC_ARK_ARC_1_1/temp1[47] ), .B(
        \MC_ARK_ARC_1_1/temp2[47] ), .ZN(\MC_ARK_ARC_1_1/temp5[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_24_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[83] ), 
        .B(n472), .ZN(\MC_ARK_ARC_1_1/temp4[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_24_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[149] ), 
        .B(n807), .ZN(\MC_ARK_ARC_1_1/temp3[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_24_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[185] ), 
        .B(n1643), .ZN(\MC_ARK_ARC_1_1/temp2[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_24_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[47] ), 
        .B(n1498), .ZN(\MC_ARK_ARC_1_1/temp1[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_23_5  ( .A(\MC_ARK_ARC_1_1/temp5[48] ), .B(
        \MC_ARK_ARC_1_1/temp6[48] ), .ZN(\RI1[2][48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_23_5  ( .A(\MC_ARK_ARC_1_1/temp3[48] ), .B(
        \MC_ARK_ARC_1_1/temp4[48] ), .ZN(\MC_ARK_ARC_1_1/temp6[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_23_5  ( .A(\MC_ARK_ARC_1_1/temp1[48] ), .B(
        \MC_ARK_ARC_1_1/temp2[48] ), .ZN(\MC_ARK_ARC_1_1/temp5[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_23_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .B(n490), .ZN(\MC_ARK_ARC_1_1/temp4[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_23_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[114] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_23_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[186] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_23_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_1/temp1[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_23_4  ( .A(\MC_ARK_ARC_1_1/temp5[49] ), .B(
        \MC_ARK_ARC_1_1/temp6[49] ), .ZN(\RI1[2][49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_23_4  ( .A(\MC_ARK_ARC_1_1/temp3[49] ), .B(
        \MC_ARK_ARC_1_1/temp4[49] ), .ZN(\MC_ARK_ARC_1_1/temp6[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_23_4  ( .A(\MC_ARK_ARC_1_1/temp1[49] ), .B(
        \MC_ARK_ARC_1_1/temp2[49] ), .ZN(\MC_ARK_ARC_1_1/temp5[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_23_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[85] ), 
        .B(n408), .ZN(\MC_ARK_ARC_1_1/temp4[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_23_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_23_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[187] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_23_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[43] ), .ZN(\MC_ARK_ARC_1_1/temp1[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_23_3  ( .A(\MC_ARK_ARC_1_1/temp5[50] ), .B(
        \MC_ARK_ARC_1_1/temp6[50] ), .ZN(\RI1[2][50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_23_3  ( .A(\MC_ARK_ARC_1_1/temp3[50] ), .B(
        \MC_ARK_ARC_1_1/temp4[50] ), .ZN(\MC_ARK_ARC_1_1/temp6[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_23_3  ( .A(\MC_ARK_ARC_1_1/temp2[50] ), .B(
        \MC_ARK_ARC_1_1/temp1[50] ), .ZN(\MC_ARK_ARC_1_1/temp5[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_23_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[86] ), 
        .B(n198), .ZN(\MC_ARK_ARC_1_1/temp4[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_23_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_23_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_1/temp2[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_23_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[44] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[50] ), .ZN(\MC_ARK_ARC_1_1/temp1[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_23_2  ( .A(\MC_ARK_ARC_1_1/temp3[51] ), .B(
        \MC_ARK_ARC_1_1/temp4[51] ), .ZN(\MC_ARK_ARC_1_1/temp6[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_23_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[87] ), 
        .B(n384), .ZN(\MC_ARK_ARC_1_1/temp4[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_23_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .B(\RI5[1][117] ), .ZN(\MC_ARK_ARC_1_1/temp3[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_23_2  ( .A(n1935), .B(
        \MC_ARK_ARC_1_1/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_1/temp2[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_23_2  ( .A(\RI5[1][51] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[45] ), .ZN(\MC_ARK_ARC_1_1/temp1[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_23_1  ( .A(\MC_ARK_ARC_1_1/temp6[52] ), .B(
        \MC_ARK_ARC_1_1/temp5[52] ), .ZN(\RI1[2][52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_23_1  ( .A(\MC_ARK_ARC_1_1/temp3[52] ), .B(
        \MC_ARK_ARC_1_1/temp4[52] ), .ZN(\MC_ARK_ARC_1_1/temp6[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_23_1  ( .A(\MC_ARK_ARC_1_1/temp1[52] ), .B(
        \MC_ARK_ARC_1_1/temp2[52] ), .ZN(\MC_ARK_ARC_1_1/temp5[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_23_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[88] ), 
        .B(n287), .ZN(\MC_ARK_ARC_1_1/temp4[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_23_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[118] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_23_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_23_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[46] ), .ZN(\MC_ARK_ARC_1_1/temp1[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_23_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .B(n513), .ZN(\MC_ARK_ARC_1_1/temp4[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_23_0  ( .A(n2153), .B(
        \MC_ARK_ARC_1_1/buf_datainput[119] ), .ZN(\MC_ARK_ARC_1_1/temp3[53] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_23_0  ( .A(n1927), .B(n515), .ZN(
        \MC_ARK_ARC_1_1/temp2[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_23_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[47] ), 
        .B(n838), .ZN(\MC_ARK_ARC_1_1/temp1[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_22_5  ( .A(\MC_ARK_ARC_1_1/temp5[54] ), .B(
        \MC_ARK_ARC_1_1/temp6[54] ), .ZN(\RI1[2][54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_22_5  ( .A(\MC_ARK_ARC_1_1/temp3[54] ), .B(
        \MC_ARK_ARC_1_1/temp4[54] ), .ZN(\MC_ARK_ARC_1_1/temp6[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_22_5  ( .A(\MC_ARK_ARC_1_1/temp1[54] ), .B(
        \MC_ARK_ARC_1_1/temp2[54] ), .ZN(\MC_ARK_ARC_1_1/temp5[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_22_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[90] ), 
        .B(n194), .ZN(\MC_ARK_ARC_1_1/temp4[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_22_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[156] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_22_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_1/temp2[54] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_22_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[48] ), .ZN(\MC_ARK_ARC_1_1/temp1[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_22_4  ( .A(\MC_ARK_ARC_1_1/temp5[55] ), .B(
        \MC_ARK_ARC_1_1/temp6[55] ), .ZN(\RI1[2][55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_22_4  ( .A(\MC_ARK_ARC_1_1/temp3[55] ), .B(
        \MC_ARK_ARC_1_1/temp4[55] ), .ZN(\MC_ARK_ARC_1_1/temp6[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_22_4  ( .A(\MC_ARK_ARC_1_1/temp2[55] ), .B(
        \MC_ARK_ARC_1_1/temp1[55] ), .ZN(\MC_ARK_ARC_1_1/temp5[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_22_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[91] ), 
        .B(n399), .ZN(\MC_ARK_ARC_1_1/temp4[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_22_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[157] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_22_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[1] ), .ZN(\MC_ARK_ARC_1_1/temp2[55] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_22_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[49] ), .ZN(\MC_ARK_ARC_1_1/temp1[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_22_3  ( .A(\MC_ARK_ARC_1_1/temp5[56] ), .B(
        \MC_ARK_ARC_1_1/temp6[56] ), .ZN(\RI1[2][56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_22_3  ( .A(\MC_ARK_ARC_1_1/temp4[56] ), .B(
        \MC_ARK_ARC_1_1/temp3[56] ), .ZN(\MC_ARK_ARC_1_1/temp6[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_22_3  ( .A(\MC_ARK_ARC_1_1/temp1[56] ), .B(
        \MC_ARK_ARC_1_1/temp2[56] ), .ZN(\MC_ARK_ARC_1_1/temp5[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_22_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[92] ), 
        .B(n424), .ZN(\MC_ARK_ARC_1_1/temp4[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_22_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[158] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_22_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_1/temp2[56] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_22_3  ( .A(\RI5[1][56] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[50] ), .ZN(\MC_ARK_ARC_1_1/temp1[56] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_22_2  ( .A(\MC_ARK_ARC_1_1/temp5[57] ), .B(
        \MC_ARK_ARC_1_1/temp6[57] ), .ZN(\RI1[2][57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_22_2  ( .A(\MC_ARK_ARC_1_1/temp3[57] ), .B(
        \MC_ARK_ARC_1_1/temp4[57] ), .ZN(\MC_ARK_ARC_1_1/temp6[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_22_2  ( .A(\MC_ARK_ARC_1_1/temp2[57] ), .B(
        \MC_ARK_ARC_1_1/temp1[57] ), .ZN(\MC_ARK_ARC_1_1/temp5[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_22_2  ( .A(\RI5[1][93] ), .B(n238), .ZN(
        \MC_ARK_ARC_1_1/temp4[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_22_2  ( .A(\RI5[1][123] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[159] ), .ZN(\MC_ARK_ARC_1_1/temp3[57] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_22_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[3] ), .ZN(\MC_ARK_ARC_1_1/temp2[57] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_22_2  ( .A(\RI5[1][51] ), .B(\RI5[1][57] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_22_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .B(n372), .ZN(\MC_ARK_ARC_1_1/temp4[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_22_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_22_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[28] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_1/temp2[58] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_22_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[52] ), .ZN(\MC_ARK_ARC_1_1/temp1[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_22_0  ( .A(\MC_ARK_ARC_1_1/temp3[59] ), .B(
        \MC_ARK_ARC_1_1/temp4[59] ), .ZN(\MC_ARK_ARC_1_1/temp6[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_22_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .B(n326), .ZN(\MC_ARK_ARC_1_1/temp4[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_22_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[161] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[125] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_22_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .B(n1640), .ZN(\MC_ARK_ARC_1_1/temp2[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_21_5  ( .A(\MC_ARK_ARC_1_1/temp5[60] ), .B(
        \MC_ARK_ARC_1_1/temp6[60] ), .ZN(\RI1[2][60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_21_5  ( .A(\MC_ARK_ARC_1_1/temp3[60] ), .B(
        \MC_ARK_ARC_1_1/temp4[60] ), .ZN(\MC_ARK_ARC_1_1/temp6[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_21_5  ( .A(\MC_ARK_ARC_1_1/temp1[60] ), .B(
        \MC_ARK_ARC_1_1/temp2[60] ), .ZN(\MC_ARK_ARC_1_1/temp5[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_21_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[96] ), 
        .B(n280), .ZN(\MC_ARK_ARC_1_1/temp4[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_21_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[162] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[126] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_21_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_1/temp2[60] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_21_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[60] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[54] ), .ZN(\MC_ARK_ARC_1_1/temp1[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_21_4  ( .A(\MC_ARK_ARC_1_1/temp5[61] ), .B(
        \MC_ARK_ARC_1_1/temp6[61] ), .ZN(\RI1[2][61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_21_4  ( .A(\MC_ARK_ARC_1_1/temp3[61] ), .B(
        \MC_ARK_ARC_1_1/temp4[61] ), .ZN(\MC_ARK_ARC_1_1/temp6[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_21_4  ( .A(\MC_ARK_ARC_1_1/temp1[61] ), .B(
        \MC_ARK_ARC_1_1/temp2[61] ), .ZN(\MC_ARK_ARC_1_1/temp5[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_21_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[97] ), 
        .B(n234), .ZN(\MC_ARK_ARC_1_1/temp4[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_21_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[127] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_21_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_1/temp2[61] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_21_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[55] ), .ZN(\MC_ARK_ARC_1_1/temp1[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_21_3  ( .A(\MC_ARK_ARC_1_1/temp5[62] ), .B(
        \MC_ARK_ARC_1_1/temp6[62] ), .ZN(\RI1[2][62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_21_3  ( .A(\MC_ARK_ARC_1_1/temp3[62] ), .B(
        \MC_ARK_ARC_1_1/temp4[62] ), .ZN(\MC_ARK_ARC_1_1/temp6[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_21_3  ( .A(\MC_ARK_ARC_1_1/temp2[62] ), .B(
        \MC_ARK_ARC_1_1/temp1[62] ), .ZN(\MC_ARK_ARC_1_1/temp5[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_21_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[98] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[62] ), .ZN(\MC_ARK_ARC_1_1/temp4[62] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_21_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[128] ), 
        .B(n1625), .ZN(\MC_ARK_ARC_1_1/temp3[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_21_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_1/temp2[62] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_21_3  ( .A(\RI5[1][56] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[62] ), .ZN(\MC_ARK_ARC_1_1/temp1[62] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_21_2  ( .A(\MC_ARK_ARC_1_1/temp3[63] ), .B(
        \MC_ARK_ARC_1_1/temp4[63] ), .ZN(\MC_ARK_ARC_1_1/temp6[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_21_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .B(n322), .ZN(\MC_ARK_ARC_1_1/temp4[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_21_2  ( .A(\RI5[1][129] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[165] ), .ZN(\MC_ARK_ARC_1_1/temp3[63] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_21_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[33] ), 
        .B(\RI5[1][9] ), .ZN(\MC_ARK_ARC_1_1/temp2[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_21_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .B(\RI5[1][57] ), .ZN(\MC_ARK_ARC_1_1/temp1[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_21_1  ( .A(\MC_ARK_ARC_1_1/temp5[64] ), .B(
        \MC_ARK_ARC_1_1/temp6[64] ), .ZN(\RI1[2][64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_21_1  ( .A(\MC_ARK_ARC_1_1/temp3[64] ), .B(
        \MC_ARK_ARC_1_1/temp4[64] ), .ZN(\MC_ARK_ARC_1_1/temp6[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_21_1  ( .A(\MC_ARK_ARC_1_1/temp2[64] ), .B(
        \MC_ARK_ARC_1_1/temp1[64] ), .ZN(\MC_ARK_ARC_1_1/temp5[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_21_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .B(n276), .ZN(\MC_ARK_ARC_1_1/temp4[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_21_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[130] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_21_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_1/temp2[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_21_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[64] ), .ZN(\MC_ARK_ARC_1_1/temp1[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_21_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[101] ), 
        .B(n230), .ZN(\MC_ARK_ARC_1_1/temp4[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_21_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[167] ), 
        .B(n1656), .ZN(\MC_ARK_ARC_1_1/temp3[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_21_0  ( .A(n2104), .B(n517), .ZN(
        \MC_ARK_ARC_1_1/temp2[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_21_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[65] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[59] ), .ZN(\MC_ARK_ARC_1_1/temp1[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_20_5  ( .A(\MC_ARK_ARC_1_1/temp5[66] ), .B(
        \MC_ARK_ARC_1_1/temp6[66] ), .ZN(\RI1[2][66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_20_5  ( .A(\MC_ARK_ARC_1_1/temp3[66] ), .B(
        \MC_ARK_ARC_1_1/temp4[66] ), .ZN(\MC_ARK_ARC_1_1/temp6[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_20_5  ( .A(\MC_ARK_ARC_1_1/temp1[66] ), .B(
        \MC_ARK_ARC_1_1/temp2[66] ), .ZN(\MC_ARK_ARC_1_1/temp5[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_20_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[102] ), 
        .B(n365), .ZN(\MC_ARK_ARC_1_1/temp4[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_20_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .B(\RI5[1][132] ), .ZN(\MC_ARK_ARC_1_1/temp3[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_20_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_1/temp2[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_20_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[60] ), .ZN(\MC_ARK_ARC_1_1/temp1[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_20_4  ( .A(\MC_ARK_ARC_1_1/temp5[67] ), .B(
        \MC_ARK_ARC_1_1/temp6[67] ), .ZN(\RI1[2][67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_20_4  ( .A(\MC_ARK_ARC_1_1/temp3[67] ), .B(
        \MC_ARK_ARC_1_1/temp4[67] ), .ZN(\MC_ARK_ARC_1_1/temp6[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_20_4  ( .A(\MC_ARK_ARC_1_1/temp1[67] ), .B(
        \MC_ARK_ARC_1_1/temp2[67] ), .ZN(\MC_ARK_ARC_1_1/temp5[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_20_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .B(n394), .ZN(\MC_ARK_ARC_1_1/temp4[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_20_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[169] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[133] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_20_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[37] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[13] ), .ZN(\MC_ARK_ARC_1_1/temp2[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_20_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[61] ), .ZN(\MC_ARK_ARC_1_1/temp1[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_20_3  ( .A(\MC_ARK_ARC_1_1/temp5[68] ), .B(
        \MC_ARK_ARC_1_1/temp6[68] ), .ZN(\RI1[2][68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_20_3  ( .A(\MC_ARK_ARC_1_1/temp3[68] ), .B(
        \MC_ARK_ARC_1_1/temp4[68] ), .ZN(\MC_ARK_ARC_1_1/temp6[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_20_3  ( .A(\MC_ARK_ARC_1_1/temp2[68] ), .B(
        \MC_ARK_ARC_1_1/temp1[68] ), .ZN(\MC_ARK_ARC_1_1/temp5[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_20_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[104] ), 
        .B(n272), .ZN(\MC_ARK_ARC_1_1/temp4[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_20_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[170] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_20_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_1/temp2[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_20_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_1/temp1[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_20_2  ( .A(\MC_ARK_ARC_1_1/temp5[69] ), .B(
        \MC_ARK_ARC_1_1/temp6[69] ), .ZN(\RI1[2][69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_20_2  ( .A(\MC_ARK_ARC_1_1/temp4[69] ), .B(
        \MC_ARK_ARC_1_1/temp3[69] ), .ZN(\MC_ARK_ARC_1_1/temp6[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_20_2  ( .A(\MC_ARK_ARC_1_1/temp2[69] ), .B(
        \MC_ARK_ARC_1_1/temp1[69] ), .ZN(\MC_ARK_ARC_1_1/temp5[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_20_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[105] ), 
        .B(n226), .ZN(\MC_ARK_ARC_1_1/temp4[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_20_2  ( .A(\RI5[1][135] ), .B(n1954), .ZN(
        \MC_ARK_ARC_1_1/temp3[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_20_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[39] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[15] ), .ZN(\MC_ARK_ARC_1_1/temp2[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_20_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[69] ), .ZN(\MC_ARK_ARC_1_1/temp1[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_20_1  ( .A(\MC_ARK_ARC_1_1/temp5[70] ), .B(
        \MC_ARK_ARC_1_1/temp6[70] ), .ZN(\RI1[2][70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_20_1  ( .A(\MC_ARK_ARC_1_1/temp3[70] ), .B(
        \MC_ARK_ARC_1_1/temp4[70] ), .ZN(\MC_ARK_ARC_1_1/temp6[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_20_1  ( .A(\MC_ARK_ARC_1_1/temp2[70] ), .B(
        \MC_ARK_ARC_1_1/temp1[70] ), .ZN(\MC_ARK_ARC_1_1/temp5[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_20_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[106] ), 
        .B(n361), .ZN(\MC_ARK_ARC_1_1/temp4[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_20_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_20_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[40] ), .ZN(\MC_ARK_ARC_1_1/temp2[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_20_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_1/temp1[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_20_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[107] ), 
        .B(n505), .ZN(\MC_ARK_ARC_1_1/temp4[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_20_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[137] ), 
        .B(n1937), .ZN(\MC_ARK_ARC_1_1/temp3[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_20_0  ( .A(n1498), .B(
        \MC_ARK_ARC_1_1/buf_datainput[17] ), .ZN(\MC_ARK_ARC_1_1/temp2[71] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_20_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[65] ), 
        .B(n1505), .ZN(\MC_ARK_ARC_1_1/temp1[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_19_5  ( .A(\MC_ARK_ARC_1_1/temp3[72] ), .B(
        \MC_ARK_ARC_1_1/temp4[72] ), .ZN(\MC_ARK_ARC_1_1/temp6[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_19_5  ( .A(\MC_ARK_ARC_1_1/temp1[72] ), .B(
        \MC_ARK_ARC_1_1/temp2[72] ), .ZN(\MC_ARK_ARC_1_1/temp5[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_19_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[108] ), 
        .B(n268), .ZN(\MC_ARK_ARC_1_1/temp4[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_19_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[174] ), 
        .B(\RI5[1][138] ), .ZN(\MC_ARK_ARC_1_1/temp3[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_19_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[18] ), .ZN(\MC_ARK_ARC_1_1/temp2[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_19_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[66] ), .ZN(\MC_ARK_ARC_1_1/temp1[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_19_4  ( .A(\MC_ARK_ARC_1_1/temp5[73] ), .B(
        \MC_ARK_ARC_1_1/temp6[73] ), .ZN(\RI1[2][73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_19_4  ( .A(\MC_ARK_ARC_1_1/temp3[73] ), .B(
        \MC_ARK_ARC_1_1/temp4[73] ), .ZN(\MC_ARK_ARC_1_1/temp6[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_19_4  ( .A(\MC_ARK_ARC_1_1/temp1[73] ), .B(
        \MC_ARK_ARC_1_1/temp2[73] ), .ZN(\MC_ARK_ARC_1_1/temp5[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_19_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[109] ), 
        .B(n222), .ZN(\MC_ARK_ARC_1_1/temp4[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_19_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[139] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_19_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[19] ), .ZN(\MC_ARK_ARC_1_1/temp2[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_19_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[67] ), .ZN(\MC_ARK_ARC_1_1/temp1[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_19_3  ( .A(\MC_ARK_ARC_1_1/temp5[74] ), .B(
        \MC_ARK_ARC_1_1/temp6[74] ), .ZN(\RI1[2][74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_19_3  ( .A(\MC_ARK_ARC_1_1/temp3[74] ), .B(
        \MC_ARK_ARC_1_1/temp4[74] ), .ZN(\MC_ARK_ARC_1_1/temp6[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_19_3  ( .A(\MC_ARK_ARC_1_1/temp2[74] ), .B(
        \MC_ARK_ARC_1_1/temp1[74] ), .ZN(\MC_ARK_ARC_1_1/temp5[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_19_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[74] ), .ZN(\MC_ARK_ARC_1_1/temp4[74] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_19_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_19_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[44] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_1/temp2[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_19_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_1/temp1[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_19_2  ( .A(\MC_ARK_ARC_1_1/temp5[75] ), .B(
        \MC_ARK_ARC_1_1/temp6[75] ), .ZN(\RI1[2][75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_19_2  ( .A(\MC_ARK_ARC_1_1/temp3[75] ), .B(
        \MC_ARK_ARC_1_1/temp4[75] ), .ZN(\MC_ARK_ARC_1_1/temp6[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_19_2  ( .A(\MC_ARK_ARC_1_1/temp1[75] ), .B(
        \MC_ARK_ARC_1_1/temp2[75] ), .ZN(\MC_ARK_ARC_1_1/temp5[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_19_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[111] ), 
        .B(n443), .ZN(\MC_ARK_ARC_1_1/temp4[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_19_2  ( .A(\RI5[1][141] ), .B(\RI5[1][177] ), 
        .ZN(\MC_ARK_ARC_1_1/temp3[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_19_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[45] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_1/temp2[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_19_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[69] ), 
        .B(\RI5[1][75] ), .ZN(\MC_ARK_ARC_1_1/temp1[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_19_1  ( .A(\MC_ARK_ARC_1_1/temp5[76] ), .B(
        \MC_ARK_ARC_1_1/temp6[76] ), .ZN(\RI1[2][76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_19_1  ( .A(\MC_ARK_ARC_1_1/temp3[76] ), .B(
        \MC_ARK_ARC_1_1/temp4[76] ), .ZN(\MC_ARK_ARC_1_1/temp6[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_19_1  ( .A(\MC_ARK_ARC_1_1/temp2[76] ), .B(
        \MC_ARK_ARC_1_1/temp1[76] ), .ZN(\MC_ARK_ARC_1_1/temp5[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_19_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[112] ), 
        .B(n264), .ZN(\MC_ARK_ARC_1_1/temp4[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_19_1  ( .A(n1953), .B(
        \MC_ARK_ARC_1_1/buf_datainput[142] ), .ZN(\MC_ARK_ARC_1_1/temp3[76] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_19_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[46] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[22] ), .ZN(\MC_ARK_ARC_1_1/temp2[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_19_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[76] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_1/temp1[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_19_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[179] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[143] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_19_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[47] ), 
        .B(n1925), .ZN(\MC_ARK_ARC_1_1/temp2[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_19_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[77] ), 
        .B(n1505), .ZN(\MC_ARK_ARC_1_1/temp1[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_18_5  ( .A(\MC_ARK_ARC_1_1/temp5[78] ), .B(
        \MC_ARK_ARC_1_1/temp6[78] ), .ZN(\RI1[2][78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_18_5  ( .A(\MC_ARK_ARC_1_1/temp3[78] ), .B(
        \MC_ARK_ARC_1_1/temp4[78] ), .ZN(\MC_ARK_ARC_1_1/temp6[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_18_5  ( .A(\MC_ARK_ARC_1_1/temp1[78] ), .B(
        \MC_ARK_ARC_1_1/temp2[78] ), .ZN(\MC_ARK_ARC_1_1/temp5[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_18_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[114] ), 
        .B(n447), .ZN(\MC_ARK_ARC_1_1/temp4[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_18_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[180] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[144] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_18_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[24] ), .ZN(\MC_ARK_ARC_1_1/temp2[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_18_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[72] ), .ZN(\MC_ARK_ARC_1_1/temp1[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_18_4  ( .A(\MC_ARK_ARC_1_1/temp5[79] ), .B(
        \MC_ARK_ARC_1_1/temp6[79] ), .ZN(\RI1[2][79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_18_4  ( .A(\MC_ARK_ARC_1_1/temp3[79] ), .B(
        \MC_ARK_ARC_1_1/temp4[79] ), .ZN(\MC_ARK_ARC_1_1/temp6[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_18_4  ( .A(\MC_ARK_ARC_1_1/temp1[79] ), .B(
        \MC_ARK_ARC_1_1/temp2[79] ), .ZN(\MC_ARK_ARC_1_1/temp5[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_18_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[115] ), 
        .B(n397), .ZN(\MC_ARK_ARC_1_1/temp4[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_18_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[145] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_18_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[25] ), .ZN(\MC_ARK_ARC_1_1/temp2[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_18_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[73] ), .ZN(\MC_ARK_ARC_1_1/temp1[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_18_3  ( .A(\MC_ARK_ARC_1_1/temp5[80] ), .B(
        \MC_ARK_ARC_1_1/temp6[80] ), .ZN(\RI1[2][80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_18_3  ( .A(\MC_ARK_ARC_1_1/temp3[80] ), .B(
        \MC_ARK_ARC_1_1/temp4[80] ), .ZN(\MC_ARK_ARC_1_1/temp6[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_18_3  ( .A(\MC_ARK_ARC_1_1/temp2[80] ), .B(
        \MC_ARK_ARC_1_1/temp1[80] ), .ZN(\MC_ARK_ARC_1_1/temp5[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_18_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[116] ), 
        .B(Key[120]), .ZN(\MC_ARK_ARC_1_1/temp4[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_18_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_18_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[50] ), .ZN(\MC_ARK_ARC_1_1/temp2[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_18_3  ( .A(n1646), .B(
        \MC_ARK_ARC_1_1/buf_datainput[74] ), .ZN(\MC_ARK_ARC_1_1/temp1[80] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_18_2  ( .A(\MC_ARK_ARC_1_1/temp5[81] ), .B(
        \MC_ARK_ARC_1_1/temp6[81] ), .ZN(\RI1[2][81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_18_2  ( .A(\MC_ARK_ARC_1_1/temp4[81] ), .B(
        \MC_ARK_ARC_1_1/temp3[81] ), .ZN(\MC_ARK_ARC_1_1/temp6[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_18_2  ( .A(\MC_ARK_ARC_1_1/temp2[81] ), .B(
        \MC_ARK_ARC_1_1/temp1[81] ), .ZN(\MC_ARK_ARC_1_1/temp5[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_18_2  ( .A(\RI5[1][117] ), .B(n433), .ZN(
        \MC_ARK_ARC_1_1/temp4[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_18_2  ( .A(n1958), .B(\RI5[1][147] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_18_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[27] ), 
        .B(\RI5[1][51] ), .ZN(\MC_ARK_ARC_1_1/temp2[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_18_2  ( .A(\RI5[1][75] ), .B(\RI5[1][81] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_18_1  ( .A(\MC_ARK_ARC_1_1/temp5[82] ), .B(
        \MC_ARK_ARC_1_1/temp6[82] ), .ZN(\RI1[2][82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_18_1  ( .A(\MC_ARK_ARC_1_1/temp3[82] ), .B(
        \MC_ARK_ARC_1_1/temp4[82] ), .ZN(\MC_ARK_ARC_1_1/temp6[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_18_1  ( .A(\MC_ARK_ARC_1_1/temp2[82] ), .B(
        \MC_ARK_ARC_1_1/temp1[82] ), .ZN(\MC_ARK_ARC_1_1/temp5[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_18_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[118] ), 
        .B(n466), .ZN(\MC_ARK_ARC_1_1/temp4[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_18_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[184] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[148] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_18_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[28] ), .ZN(\MC_ARK_ARC_1_1/temp2[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_18_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[76] ), .ZN(\MC_ARK_ARC_1_1/temp1[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_18_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[119] ), 
        .B(n502), .ZN(\MC_ARK_ARC_1_1/temp4[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_18_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[185] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[149] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_18_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .B(n837), .ZN(\MC_ARK_ARC_1_1/temp2[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_18_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[77] ), 
        .B(n813), .ZN(\MC_ARK_ARC_1_1/temp1[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_17_5  ( .A(\MC_ARK_ARC_1_1/temp5[84] ), .B(
        \MC_ARK_ARC_1_1/temp6[84] ), .ZN(\RI1[2][84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_17_5  ( .A(\MC_ARK_ARC_1_1/temp3[84] ), .B(
        \MC_ARK_ARC_1_1/temp4[84] ), .ZN(\MC_ARK_ARC_1_1/temp6[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_17_5  ( .A(\MC_ARK_ARC_1_1/temp1[84] ), .B(
        \MC_ARK_ARC_1_1/temp2[84] ), .ZN(\MC_ARK_ARC_1_1/temp5[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_17_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[120] ), 
        .B(n256), .ZN(\MC_ARK_ARC_1_1/temp4[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_17_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[150] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_17_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[30] ), .ZN(\MC_ARK_ARC_1_1/temp2[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_17_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[78] ), .ZN(\MC_ARK_ARC_1_1/temp1[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_17_4  ( .A(\MC_ARK_ARC_1_1/temp5[85] ), .B(
        \MC_ARK_ARC_1_1/temp6[85] ), .ZN(\RI1[2][85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_17_4  ( .A(\MC_ARK_ARC_1_1/temp3[85] ), .B(
        \MC_ARK_ARC_1_1/temp4[85] ), .ZN(\MC_ARK_ARC_1_1/temp6[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_17_4  ( .A(\MC_ARK_ARC_1_1/temp1[85] ), .B(
        \MC_ARK_ARC_1_1/temp2[85] ), .ZN(\MC_ARK_ARC_1_1/temp5[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_17_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[121] ), 
        .B(n405), .ZN(\MC_ARK_ARC_1_1/temp4[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_17_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[151] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_17_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[31] ), .ZN(\MC_ARK_ARC_1_1/temp2[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_17_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[79] ), .ZN(\MC_ARK_ARC_1_1/temp1[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_17_3  ( .A(\MC_ARK_ARC_1_1/temp5[86] ), .B(
        \MC_ARK_ARC_1_1/temp6[86] ), .ZN(\RI1[2][86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_17_3  ( .A(\MC_ARK_ARC_1_1/temp3[86] ), .B(
        \MC_ARK_ARC_1_1/temp4[86] ), .ZN(\MC_ARK_ARC_1_1/temp6[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_17_3  ( .A(\MC_ARK_ARC_1_1/temp1[86] ), .B(
        \MC_ARK_ARC_1_1/temp2[86] ), .ZN(\MC_ARK_ARC_1_1/temp5[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_17_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[122] ), 
        .B(n345), .ZN(\MC_ARK_ARC_1_1/temp4[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_17_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_17_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[32] ), 
        .B(\RI5[1][56] ), .ZN(\MC_ARK_ARC_1_1/temp2[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_17_3  ( .A(n1645), .B(
        \MC_ARK_ARC_1_1/buf_datainput[86] ), .ZN(\MC_ARK_ARC_1_1/temp1[86] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_17_2  ( .A(\MC_ARK_ARC_1_1/temp5[87] ), .B(
        \MC_ARK_ARC_1_1/temp6[87] ), .ZN(\RI1[2][87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_17_2  ( .A(\MC_ARK_ARC_1_1/temp3[87] ), .B(
        \MC_ARK_ARC_1_1/temp4[87] ), .ZN(\MC_ARK_ARC_1_1/temp6[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_17_2  ( .A(\MC_ARK_ARC_1_1/temp1[87] ), .B(
        \MC_ARK_ARC_1_1/temp2[87] ), .ZN(\MC_ARK_ARC_1_1/temp5[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_17_2  ( .A(\RI5[1][123] ), .B(n299), .ZN(
        \MC_ARK_ARC_1_1/temp4[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_17_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .B(n1934), .ZN(\MC_ARK_ARC_1_1/temp3[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_17_2  ( .A(\RI5[1][57] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_1/temp2[87] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_17_2  ( .A(\RI5[1][81] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[87] ), .ZN(\MC_ARK_ARC_1_1/temp1[87] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_17_1  ( .A(\MC_ARK_ARC_1_1/temp5[88] ), .B(
        \MC_ARK_ARC_1_1/temp6[88] ), .ZN(\RI1[2][88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_17_1  ( .A(\MC_ARK_ARC_1_1/temp3[88] ), .B(
        \MC_ARK_ARC_1_1/temp4[88] ), .ZN(\MC_ARK_ARC_1_1/temp6[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_17_1  ( .A(\MC_ARK_ARC_1_1/temp1[88] ), .B(
        \MC_ARK_ARC_1_1/temp2[88] ), .ZN(\MC_ARK_ARC_1_1/temp5[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_17_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[124] ), 
        .B(n442), .ZN(\MC_ARK_ARC_1_1/temp4[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_17_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[190] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_17_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[34] ), .ZN(\MC_ARK_ARC_1_1/temp2[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_17_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_1/temp1[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_17_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[125] ), 
        .B(n484), .ZN(\MC_ARK_ARC_1_1/temp4[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_17_0  ( .A(n2152), .B(n514), .ZN(
        \MC_ARK_ARC_1_1/temp3[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_17_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[59] ), 
        .B(n517), .ZN(\MC_ARK_ARC_1_1/temp2[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_17_0  ( .A(n813), .B(
        \MC_ARK_ARC_1_1/buf_datainput[89] ), .ZN(\MC_ARK_ARC_1_1/temp1[89] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_16_5  ( .A(\MC_ARK_ARC_1_1/temp5[90] ), .B(
        \MC_ARK_ARC_1_1/temp6[90] ), .ZN(\RI1[2][90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_16_5  ( .A(\MC_ARK_ARC_1_1/temp3[90] ), .B(
        \MC_ARK_ARC_1_1/temp4[90] ), .ZN(\MC_ARK_ARC_1_1/temp6[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_16_5  ( .A(\MC_ARK_ARC_1_1/temp1[90] ), .B(
        \MC_ARK_ARC_1_1/temp2[90] ), .ZN(\MC_ARK_ARC_1_1/temp5[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_16_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[126] ), 
        .B(n464), .ZN(\MC_ARK_ARC_1_1/temp4[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_16_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[156] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_16_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[60] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[36] ), .ZN(\MC_ARK_ARC_1_1/temp2[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_16_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[84] ), .ZN(\MC_ARK_ARC_1_1/temp1[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_16_4  ( .A(\MC_ARK_ARC_1_1/temp5[91] ), .B(
        \MC_ARK_ARC_1_1/temp6[91] ), .ZN(\RI1[2][91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_16_4  ( .A(\MC_ARK_ARC_1_1/temp4[91] ), .B(
        \MC_ARK_ARC_1_1/temp3[91] ), .ZN(\MC_ARK_ARC_1_1/temp6[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_16_4  ( .A(\MC_ARK_ARC_1_1/temp2[91] ), .B(
        \MC_ARK_ARC_1_1/temp1[91] ), .ZN(\MC_ARK_ARC_1_1/temp5[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_16_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[127] ), 
        .B(n296), .ZN(\MC_ARK_ARC_1_1/temp4[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_16_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[157] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_16_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[37] ), .ZN(\MC_ARK_ARC_1_1/temp2[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_16_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[85] ), .ZN(\MC_ARK_ARC_1_1/temp1[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_16_3  ( .A(\MC_ARK_ARC_1_1/temp5[92] ), .B(
        \MC_ARK_ARC_1_1/temp6[92] ), .ZN(\RI1[2][92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_16_3  ( .A(\MC_ARK_ARC_1_1/temp3[92] ), .B(
        \MC_ARK_ARC_1_1/temp4[92] ), .ZN(\MC_ARK_ARC_1_1/temp6[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_16_3  ( .A(\MC_ARK_ARC_1_1/temp1[92] ), .B(
        \MC_ARK_ARC_1_1/temp2[92] ), .ZN(\MC_ARK_ARC_1_1/temp5[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_16_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[128] ), 
        .B(n249), .ZN(\MC_ARK_ARC_1_1/temp4[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_16_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[158] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_1/temp3[92] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_16_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_1/temp2[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_16_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[92] ), .ZN(\MC_ARK_ARC_1_1/temp1[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_16_2  ( .A(\MC_ARK_ARC_1_1/temp5[93] ), .B(
        \MC_ARK_ARC_1_1/temp6[93] ), .ZN(\RI1[2][93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_16_2  ( .A(\MC_ARK_ARC_1_1/temp3[93] ), .B(
        \MC_ARK_ARC_1_1/temp4[93] ), .ZN(\MC_ARK_ARC_1_1/temp6[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_16_2  ( .A(\MC_ARK_ARC_1_1/temp1[93] ), .B(
        \MC_ARK_ARC_1_1/temp2[93] ), .ZN(\MC_ARK_ARC_1_1/temp5[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_16_2  ( .A(\RI5[1][129] ), .B(n202), .ZN(
        \MC_ARK_ARC_1_1/temp4[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_16_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[159] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[3] ), .ZN(\MC_ARK_ARC_1_1/temp3[93] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_16_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[39] ), .ZN(\MC_ARK_ARC_1_1/temp2[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_16_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[87] ), 
        .B(\RI5[1][93] ), .ZN(\MC_ARK_ARC_1_1/temp1[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_16_1  ( .A(\MC_ARK_ARC_1_1/temp2[94] ), .B(
        \MC_ARK_ARC_1_1/temp1[94] ), .ZN(\MC_ARK_ARC_1_1/temp5[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_16_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[130] ), 
        .B(n480), .ZN(\MC_ARK_ARC_1_1/temp4[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_16_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_16_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[64] ), .ZN(\MC_ARK_ARC_1_1/temp2[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_16_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_1/temp1[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_16_0  ( .A(\MC_ARK_ARC_1_1/temp5[95] ), .B(
        \MC_ARK_ARC_1_1/temp6[95] ), .ZN(\RI1[2][95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_16_0  ( .A(\MC_ARK_ARC_1_1/temp3[95] ), .B(
        \MC_ARK_ARC_1_1/temp4[95] ), .ZN(\MC_ARK_ARC_1_1/temp6[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_16_0  ( .A(\MC_ARK_ARC_1_1/temp1[95] ), .B(
        \MC_ARK_ARC_1_1/temp2[95] ), .ZN(\MC_ARK_ARC_1_1/temp5[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_16_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[131] ), 
        .B(n450), .ZN(\MC_ARK_ARC_1_1/temp4[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_16_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[161] ), 
        .B(n1640), .ZN(\MC_ARK_ARC_1_1/temp3[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_16_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[65] ), 
        .B(n1497), .ZN(\MC_ARK_ARC_1_1/temp2[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_16_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[95] ), .ZN(\MC_ARK_ARC_1_1/temp1[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_15_5  ( .A(\MC_ARK_ARC_1_1/temp5[96] ), .B(
        \MC_ARK_ARC_1_1/temp6[96] ), .ZN(\RI1[2][96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_15_5  ( .A(\MC_ARK_ARC_1_1/temp4[96] ), .B(
        \MC_ARK_ARC_1_1/temp3[96] ), .ZN(\MC_ARK_ARC_1_1/temp6[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_15_5  ( .A(\MC_ARK_ARC_1_1/temp1[96] ), .B(
        \MC_ARK_ARC_1_1/temp2[96] ), .ZN(\MC_ARK_ARC_1_1/temp5[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_15_5  ( .A(\RI5[1][132] ), .B(n376), .ZN(
        \MC_ARK_ARC_1_1/temp4[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_15_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_15_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_1/temp2[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_15_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[90] ), .ZN(\MC_ARK_ARC_1_1/temp1[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_15_4  ( .A(\MC_ARK_ARC_1_1/temp5[97] ), .B(
        \MC_ARK_ARC_1_1/temp6[97] ), .ZN(\RI1[2][97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_15_4  ( .A(\MC_ARK_ARC_1_1/temp3[97] ), .B(
        \MC_ARK_ARC_1_1/temp4[97] ), .ZN(\MC_ARK_ARC_1_1/temp6[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_15_4  ( .A(\MC_ARK_ARC_1_1/temp1[97] ), .B(
        \MC_ARK_ARC_1_1/temp2[97] ), .ZN(\MC_ARK_ARC_1_1/temp5[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_15_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[133] ), 
        .B(n199), .ZN(\MC_ARK_ARC_1_1/temp4[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_15_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[7] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[163] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_15_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[43] ), .ZN(\MC_ARK_ARC_1_1/temp2[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_15_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[97] ), .ZN(\MC_ARK_ARC_1_1/temp1[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_15_3  ( .A(\MC_ARK_ARC_1_1/temp5[98] ), .B(
        \MC_ARK_ARC_1_1/temp6[98] ), .ZN(\RI1[2][98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_15_3  ( .A(\MC_ARK_ARC_1_1/temp4[98] ), .B(
        \MC_ARK_ARC_1_1/temp3[98] ), .ZN(\MC_ARK_ARC_1_1/temp6[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_15_3  ( .A(\MC_ARK_ARC_1_1/temp2[98] ), .B(
        \MC_ARK_ARC_1_1/temp1[98] ), .ZN(\MC_ARK_ARC_1_1/temp5[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_15_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[134] ), 
        .B(n335), .ZN(\MC_ARK_ARC_1_1/temp4[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_15_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[8] ), 
        .B(n1625), .ZN(\MC_ARK_ARC_1_1/temp3[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_15_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[68] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[44] ), .ZN(\MC_ARK_ARC_1_1/temp2[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_15_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[98] ), .ZN(\MC_ARK_ARC_1_1/temp1[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_15_2  ( .A(\MC_ARK_ARC_1_1/temp5[99] ), .B(
        \MC_ARK_ARC_1_1/temp6[99] ), .ZN(\RI1[2][99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_15_2  ( .A(\MC_ARK_ARC_1_1/temp3[99] ), .B(
        \MC_ARK_ARC_1_1/temp4[99] ), .ZN(\MC_ARK_ARC_1_1/temp6[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_15_2  ( .A(\MC_ARK_ARC_1_1/temp2[99] ), .B(
        \MC_ARK_ARC_1_1/temp1[99] ), .ZN(\MC_ARK_ARC_1_1/temp5[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_15_2  ( .A(\RI5[1][135] ), .B(n423), .ZN(
        \MC_ARK_ARC_1_1/temp4[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_15_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[165] ), 
        .B(\RI5[1][9] ), .ZN(\MC_ARK_ARC_1_1/temp3[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_15_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[45] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[69] ), .ZN(\MC_ARK_ARC_1_1/temp2[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_15_2  ( .A(\RI5[1][93] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[99] ), .ZN(\MC_ARK_ARC_1_1/temp1[99] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_15_1  ( .A(\MC_ARK_ARC_1_1/temp5[100] ), .B(
        \MC_ARK_ARC_1_1/temp6[100] ), .ZN(\RI1[2][100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_15_1  ( .A(\MC_ARK_ARC_1_1/temp3[100] ), .B(
        \MC_ARK_ARC_1_1/temp4[100] ), .ZN(\MC_ARK_ARC_1_1/temp6[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_15_1  ( .A(\MC_ARK_ARC_1_1/temp2[100] ), .B(
        \MC_ARK_ARC_1_1/temp1[100] ), .ZN(\MC_ARK_ARC_1_1/temp5[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_15_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[136] ), 
        .B(n487), .ZN(\MC_ARK_ARC_1_1/temp4[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_15_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_15_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[46] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_15_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[94] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_15_0  ( .A(\MC_ARK_ARC_1_1/temp5[101] ), .B(
        \MC_ARK_ARC_1_1/temp6[101] ), .ZN(\RI1[2][101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_15_0  ( .A(\MC_ARK_ARC_1_1/temp3[101] ), .B(
        \MC_ARK_ARC_1_1/temp4[101] ), .ZN(\MC_ARK_ARC_1_1/temp6[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_15_0  ( .A(\MC_ARK_ARC_1_1/temp1[101] ), .B(
        \MC_ARK_ARC_1_1/temp2[101] ), .ZN(\MC_ARK_ARC_1_1/temp5[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_15_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[137] ), 
        .B(n195), .ZN(\MC_ARK_ARC_1_1/temp4[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_15_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[167] ), 
        .B(n2105), .ZN(\MC_ARK_ARC_1_1/temp3[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_15_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[47] ), 
        .B(n1952), .ZN(\MC_ARK_ARC_1_1/temp2[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_15_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .B(n2124), .ZN(\MC_ARK_ARC_1_1/temp1[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_14_5  ( .A(\MC_ARK_ARC_1_1/temp5[102] ), .B(
        \MC_ARK_ARC_1_1/temp6[102] ), .ZN(\RI1[2][102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_14_5  ( .A(\MC_ARK_ARC_1_1/temp4[102] ), .B(
        \MC_ARK_ARC_1_1/temp3[102] ), .ZN(\MC_ARK_ARC_1_1/temp6[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_14_5  ( .A(\MC_ARK_ARC_1_1/temp1[102] ), .B(
        \MC_ARK_ARC_1_1/temp2[102] ), .ZN(\MC_ARK_ARC_1_1/temp5[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_14_5  ( .A(\RI5[1][138] ), .B(n331), .ZN(
        \MC_ARK_ARC_1_1/temp4[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_14_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_14_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[48] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_14_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[96] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_14_4  ( .A(\MC_ARK_ARC_1_1/temp5[103] ), .B(
        \MC_ARK_ARC_1_1/temp6[103] ), .ZN(\RI1[2][103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_14_4  ( .A(\MC_ARK_ARC_1_1/temp3[103] ), .B(
        \MC_ARK_ARC_1_1/temp4[103] ), .ZN(\MC_ARK_ARC_1_1/temp6[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_14_4  ( .A(\MC_ARK_ARC_1_1/temp1[103] ), .B(
        \MC_ARK_ARC_1_1/temp2[103] ), .ZN(\MC_ARK_ARC_1_1/temp5[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_14_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .B(n284), .ZN(\MC_ARK_ARC_1_1/temp4[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_14_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[169] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_14_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[49] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_14_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[97] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_14_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[140] ), 
        .B(n239), .ZN(\MC_ARK_ARC_1_1/temp4[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_14_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[170] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_14_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[74] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_14_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[98] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_14_2  ( .A(\MC_ARK_ARC_1_1/temp2[105] ), .B(
        \MC_ARK_ARC_1_1/temp1[105] ), .ZN(\MC_ARK_ARC_1_1/temp5[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_14_2  ( .A(\RI5[1][141] ), .B(
        \MC_ARK_ARC_1_1/buf_keyinput[105] ), .ZN(\MC_ARK_ARC_1_1/temp4[105] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_14_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .B(n1954), .ZN(\MC_ARK_ARC_1_1/temp3[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_14_2  ( .A(\RI5[1][51] ), .B(\RI5[1][75] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_14_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[99] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_14_1  ( .A(\MC_ARK_ARC_1_1/temp5[106] ), .B(
        \MC_ARK_ARC_1_1/temp6[106] ), .ZN(\RI1[2][106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_14_1  ( .A(\MC_ARK_ARC_1_1/temp3[106] ), .B(
        \MC_ARK_ARC_1_1/temp4[106] ), .ZN(\MC_ARK_ARC_1_1/temp6[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_14_1  ( .A(\MC_ARK_ARC_1_1/temp1[106] ), .B(
        \MC_ARK_ARC_1_1/temp2[106] ), .ZN(\MC_ARK_ARC_1_1/temp5[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_14_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[106] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_14_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_14_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[76] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_14_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_14_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[143] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[107] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_14_0  ( .A(n1936), .B(n1642), .ZN(
        \MC_ARK_ARC_1_1/temp3[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_14_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[77] ), 
        .B(n837), .ZN(\MC_ARK_ARC_1_1/temp2[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_14_0  ( .A(n2125), .B(n852), .ZN(
        \MC_ARK_ARC_1_1/temp1[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_13_5  ( .A(\MC_ARK_ARC_1_1/temp5[108] ), .B(
        \MC_ARK_ARC_1_1/temp6[108] ), .ZN(\RI1[2][108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_13_5  ( .A(\MC_ARK_ARC_1_1/temp3[108] ), .B(
        \MC_ARK_ARC_1_1/temp4[108] ), .ZN(\MC_ARK_ARC_1_1/temp6[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_13_5  ( .A(\MC_ARK_ARC_1_1/temp1[108] ), .B(
        \MC_ARK_ARC_1_1/temp2[108] ), .ZN(\MC_ARK_ARC_1_1/temp5[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_13_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[144] ), 
        .B(n491), .ZN(\MC_ARK_ARC_1_1/temp4[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_13_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[174] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_13_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[54] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_13_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[108] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[102] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_13_4  ( .A(\MC_ARK_ARC_1_1/temp5[109] ), .B(
        \MC_ARK_ARC_1_1/temp6[109] ), .ZN(\RI1[2][109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_13_4  ( .A(\MC_ARK_ARC_1_1/temp3[109] ), .B(
        \MC_ARK_ARC_1_1/temp4[109] ), .ZN(\MC_ARK_ARC_1_1/temp6[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_13_4  ( .A(\MC_ARK_ARC_1_1/temp1[109] ), .B(
        \MC_ARK_ARC_1_1/temp2[109] ), .ZN(\MC_ARK_ARC_1_1/temp5[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_13_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[145] ), 
        .B(n369), .ZN(\MC_ARK_ARC_1_1/temp4[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_13_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_13_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[55] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_13_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_13_3  ( .A(\MC_ARK_ARC_1_1/temp2[110] ), .B(
        \MC_ARK_ARC_1_1/temp1[110] ), .ZN(\MC_ARK_ARC_1_1/temp5[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_13_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[166] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_13_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_13_3  ( .A(n1645), .B(\RI5[1][56] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_13_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_13_2  ( .A(\MC_ARK_ARC_1_1/temp5[111] ), .B(
        \MC_ARK_ARC_1_1/temp6[111] ), .ZN(\RI1[2][111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_13_2  ( .A(\MC_ARK_ARC_1_1/temp3[111] ), .B(
        \MC_ARK_ARC_1_1/temp4[111] ), .ZN(\MC_ARK_ARC_1_1/temp6[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_13_2  ( .A(\MC_ARK_ARC_1_1/temp2[111] ), .B(
        \MC_ARK_ARC_1_1/temp1[111] ), .ZN(\MC_ARK_ARC_1_1/temp5[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_13_2  ( .A(\RI5[1][147] ), .B(n378), .ZN(
        \MC_ARK_ARC_1_1/temp4[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_13_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[21] ), 
        .B(\RI5[1][177] ), .ZN(\MC_ARK_ARC_1_1/temp3[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_13_2  ( .A(\RI5[1][57] ), .B(\RI5[1][81] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_13_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[111] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[105] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_13_1  ( .A(\MC_ARK_ARC_1_1/temp6[112] ), .B(
        \MC_ARK_ARC_1_1/temp5[112] ), .ZN(\RI1[2][112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_13_1  ( .A(\MC_ARK_ARC_1_1/temp3[112] ), .B(
        \MC_ARK_ARC_1_1/temp4[112] ), .ZN(\MC_ARK_ARC_1_1/temp6[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_13_1  ( .A(\MC_ARK_ARC_1_1/temp2[112] ), .B(
        \MC_ARK_ARC_1_1/temp1[112] ), .ZN(\MC_ARK_ARC_1_1/temp5[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_13_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[148] ), 
        .B(n485), .ZN(\MC_ARK_ARC_1_1/temp4[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_13_1  ( .A(n1953), .B(
        \MC_ARK_ARC_1_1/buf_datainput[22] ), .ZN(\MC_ARK_ARC_1_1/temp3[112] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_13_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[82] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_13_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[112] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_13_0  ( .A(\MC_ARK_ARC_1_1/temp6[113] ), .B(
        \MC_ARK_ARC_1_1/temp5[113] ), .ZN(\RI1[2][113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_13_0  ( .A(\MC_ARK_ARC_1_1/temp3[113] ), .B(
        \MC_ARK_ARC_1_1/temp4[113] ), .ZN(\MC_ARK_ARC_1_1/temp6[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_13_0  ( .A(\MC_ARK_ARC_1_1/temp2[113] ), .B(
        \MC_ARK_ARC_1_1/temp1[113] ), .ZN(\MC_ARK_ARC_1_1/temp5[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_13_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[149] ), 
        .B(n503), .ZN(\MC_ARK_ARC_1_1/temp4[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_13_0  ( .A(n1926), .B(
        \MC_ARK_ARC_1_1/buf_datainput[179] ), .ZN(\MC_ARK_ARC_1_1/temp3[113] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_13_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[59] ), 
        .B(n813), .ZN(\MC_ARK_ARC_1_1/temp2[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_13_0  ( .A(n852), .B(n807), .ZN(
        \MC_ARK_ARC_1_1/temp1[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_12_5  ( .A(\MC_ARK_ARC_1_1/temp5[114] ), .B(
        \MC_ARK_ARC_1_1/temp6[114] ), .ZN(\RI1[2][114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_12_5  ( .A(\MC_ARK_ARC_1_1/temp3[114] ), .B(
        \MC_ARK_ARC_1_1/temp4[114] ), .ZN(\MC_ARK_ARC_1_1/temp6[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_12_5  ( .A(\MC_ARK_ARC_1_1/temp1[114] ), .B(
        \MC_ARK_ARC_1_1/temp2[114] ), .ZN(\MC_ARK_ARC_1_1/temp5[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_12_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .B(n482), .ZN(\MC_ARK_ARC_1_1/temp4[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_12_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_12_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[60] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_12_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[108] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_12_4  ( .A(\MC_ARK_ARC_1_1/temp5[115] ), .B(
        \MC_ARK_ARC_1_1/temp6[115] ), .ZN(\RI1[2][115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_12_4  ( .A(\MC_ARK_ARC_1_1/temp3[115] ), .B(
        \MC_ARK_ARC_1_1/temp4[115] ), .ZN(\MC_ARK_ARC_1_1/temp6[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_12_4  ( .A(\MC_ARK_ARC_1_1/temp1[115] ), .B(
        \MC_ARK_ARC_1_1/temp2[115] ), .ZN(\MC_ARK_ARC_1_1/temp5[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_12_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .B(n273), .ZN(\MC_ARK_ARC_1_1/temp4[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_12_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_12_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[61] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_12_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_12_3  ( .A(\MC_ARK_ARC_1_1/temp5[116] ), .B(
        \MC_ARK_ARC_1_1/temp6[116] ), .ZN(\RI1[2][116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_12_3  ( .A(\MC_ARK_ARC_1_1/temp3[116] ), .B(
        \MC_ARK_ARC_1_1/temp4[116] ), .ZN(\MC_ARK_ARC_1_1/temp6[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_12_3  ( .A(\MC_ARK_ARC_1_1/temp2[116] ), .B(
        \MC_ARK_ARC_1_1/temp1[116] ), .ZN(\MC_ARK_ARC_1_1/temp5[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_12_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[152] ), 
        .B(n377), .ZN(\MC_ARK_ARC_1_1/temp4[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_12_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[26] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_12_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[62] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_12_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[116] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_12_2  ( .A(\MC_ARK_ARC_1_1/temp5[117] ), .B(
        \MC_ARK_ARC_1_1/temp6[117] ), .ZN(\RI1[2][117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_12_2  ( .A(\MC_ARK_ARC_1_1/temp3[117] ), .B(
        \MC_ARK_ARC_1_1/temp4[117] ), .ZN(\MC_ARK_ARC_1_1/temp6[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_12_2  ( .A(\MC_ARK_ARC_1_1/temp1[117] ), .B(
        \MC_ARK_ARC_1_1/temp2[117] ), .ZN(\MC_ARK_ARC_1_1/temp5[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_12_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .B(n362), .ZN(\MC_ARK_ARC_1_1/temp4[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_12_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[27] ), 
        .B(n1958), .ZN(\MC_ARK_ARC_1_1/temp3[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_12_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[87] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_12_2  ( .A(\RI5[1][117] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[111] ), .ZN(\MC_ARK_ARC_1_1/temp1[117] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_12_1  ( .A(\MC_ARK_ARC_1_1/temp5[118] ), .B(
        \MC_ARK_ARC_1_1/temp6[118] ), .ZN(\RI1[2][118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_12_1  ( .A(\MC_ARK_ARC_1_1/temp3[118] ), .B(
        \MC_ARK_ARC_1_1/temp4[118] ), .ZN(\MC_ARK_ARC_1_1/temp6[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_12_1  ( .A(\MC_ARK_ARC_1_1/temp1[118] ), .B(
        \MC_ARK_ARC_1_1/temp2[118] ), .ZN(\MC_ARK_ARC_1_1/temp5[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_12_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[154] ), 
        .B(n500), .ZN(\MC_ARK_ARC_1_1/temp4[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_12_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[184] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[28] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_12_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[88] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_12_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[118] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[112] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_12_0  ( .A(\MC_ARK_ARC_1_1/temp3[119] ), .B(
        \MC_ARK_ARC_1_1/temp4[119] ), .ZN(\MC_ARK_ARC_1_1/temp6[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_12_0  ( .A(\MC_ARK_ARC_1_1/temp2[119] ), .B(
        \MC_ARK_ARC_1_1/temp1[119] ), .ZN(\MC_ARK_ARC_1_1/temp5[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_12_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[155] ), 
        .B(n509), .ZN(\MC_ARK_ARC_1_1/temp4[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_12_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[185] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[29] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_12_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[65] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_12_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[119] ), 
        .B(n808), .ZN(\MC_ARK_ARC_1_1/temp1[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_11_5  ( .A(\MC_ARK_ARC_1_1/temp3[120] ), .B(
        \MC_ARK_ARC_1_1/temp4[120] ), .ZN(\MC_ARK_ARC_1_1/temp6[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_11_5  ( .A(\MC_ARK_ARC_1_1/temp1[120] ), .B(
        \MC_ARK_ARC_1_1/temp2[120] ), .ZN(\MC_ARK_ARC_1_1/temp5[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_11_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[156] ), 
        .B(n223), .ZN(\MC_ARK_ARC_1_1/temp4[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_11_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[186] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_11_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[66] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_11_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[114] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_11_4  ( .A(\MC_ARK_ARC_1_1/temp5[121] ), .B(
        \MC_ARK_ARC_1_1/temp6[121] ), .ZN(\RI1[2][121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_11_4  ( .A(\MC_ARK_ARC_1_1/temp3[121] ), .B(
        \MC_ARK_ARC_1_1/temp4[121] ), .ZN(\MC_ARK_ARC_1_1/temp6[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_11_4  ( .A(\MC_ARK_ARC_1_1/temp1[121] ), .B(
        \MC_ARK_ARC_1_1/temp2[121] ), .ZN(\MC_ARK_ARC_1_1/temp5[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_11_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[157] ), 
        .B(n393), .ZN(\MC_ARK_ARC_1_1/temp4[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_11_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[187] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_11_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[67] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_11_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_11_3  ( .A(\MC_ARK_ARC_1_1/temp5[122] ), .B(
        \MC_ARK_ARC_1_1/temp6[122] ), .ZN(\RI1[2][122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_11_3  ( .A(\MC_ARK_ARC_1_1/temp3[122] ), .B(
        \MC_ARK_ARC_1_1/temp4[122] ), .ZN(\MC_ARK_ARC_1_1/temp6[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_11_3  ( .A(\MC_ARK_ARC_1_1/temp2[122] ), .B(
        \MC_ARK_ARC_1_1/temp1[122] ), .ZN(\MC_ARK_ARC_1_1/temp5[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_11_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[158] ), 
        .B(n312), .ZN(\MC_ARK_ARC_1_1/temp4[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_11_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[32] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_11_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[68] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_11_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[122] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_11_2  ( .A(\MC_ARK_ARC_1_1/temp5[123] ), .B(
        \MC_ARK_ARC_1_1/temp6[123] ), .ZN(\RI1[2][123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_11_2  ( .A(\MC_ARK_ARC_1_1/temp3[123] ), .B(
        \MC_ARK_ARC_1_1/temp4[123] ), .ZN(\MC_ARK_ARC_1_1/temp6[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_11_2  ( .A(\MC_ARK_ARC_1_1/temp2[123] ), .B(
        \MC_ARK_ARC_1_1/temp1[123] ), .ZN(\MC_ARK_ARC_1_1/temp5[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_11_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[159] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[123] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_11_2  ( .A(n1935), .B(
        \MC_ARK_ARC_1_1/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_1/temp3[123] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_11_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[69] ), 
        .B(\RI5[1][93] ), .ZN(\MC_ARK_ARC_1_1/temp2[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_11_2  ( .A(\RI5[1][117] ), .B(\RI5[1][123] ), 
        .ZN(\MC_ARK_ARC_1_1/temp1[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_11_1  ( .A(\MC_ARK_ARC_1_1/temp5[124] ), .B(
        \MC_ARK_ARC_1_1/temp6[124] ), .ZN(\RI1[2][124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_11_1  ( .A(\MC_ARK_ARC_1_1/temp3[124] ), .B(
        \MC_ARK_ARC_1_1/temp4[124] ), .ZN(\MC_ARK_ARC_1_1/temp6[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_11_1  ( .A(\MC_ARK_ARC_1_1/temp1[124] ), .B(
        \MC_ARK_ARC_1_1/temp2[124] ), .ZN(\MC_ARK_ARC_1_1/temp5[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_11_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .B(n441), .ZN(\MC_ARK_ARC_1_1/temp4[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_11_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_11_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[70] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_11_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[118] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_11_0  ( .A(\MC_ARK_ARC_1_1/temp4[125] ), .B(
        \MC_ARK_ARC_1_1/temp3[125] ), .ZN(\MC_ARK_ARC_1_1/temp6[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_11_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[161] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[125] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_11_0  ( .A(n519), .B(n514), .ZN(
        \MC_ARK_ARC_1_1/temp3[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_11_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .B(n1952), .ZN(\MC_ARK_ARC_1_1/temp2[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_11_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[119] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[125] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_10_5  ( .A(\MC_ARK_ARC_1_1/temp5[126] ), .B(
        \MC_ARK_ARC_1_1/temp6[126] ), .ZN(\RI1[2][126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_10_5  ( .A(\MC_ARK_ARC_1_1/temp3[126] ), .B(
        \MC_ARK_ARC_1_1/temp4[126] ), .ZN(\MC_ARK_ARC_1_1/temp6[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_10_5  ( .A(\MC_ARK_ARC_1_1/temp1[126] ), .B(
        \MC_ARK_ARC_1_1/temp2[126] ), .ZN(\MC_ARK_ARC_1_1/temp5[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_10_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[162] ), 
        .B(n308), .ZN(\MC_ARK_ARC_1_1/temp4[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_10_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_1/temp3[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_10_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[72] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_10_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_10_4  ( .A(\MC_ARK_ARC_1_1/temp5[127] ), .B(
        \MC_ARK_ARC_1_1/temp6[127] ), .ZN(\RI1[2][127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_10_4  ( .A(\MC_ARK_ARC_1_1/temp3[127] ), .B(
        \MC_ARK_ARC_1_1/temp4[127] ), .ZN(\MC_ARK_ARC_1_1/temp6[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_10_4  ( .A(\MC_ARK_ARC_1_1/temp1[127] ), .B(
        \MC_ARK_ARC_1_1/temp2[127] ), .ZN(\MC_ARK_ARC_1_1/temp5[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_10_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .B(n402), .ZN(\MC_ARK_ARC_1_1/temp4[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_10_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[37] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[1] ), .ZN(\MC_ARK_ARC_1_1/temp3[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_10_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[73] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_10_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_10_3  ( .A(\MC_ARK_ARC_1_1/temp4[128] ), .B(
        \MC_ARK_ARC_1_1/temp3[128] ), .ZN(\MC_ARK_ARC_1_1/temp6[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_10_3  ( .A(n1624), .B(n215), .ZN(
        \MC_ARK_ARC_1_1/temp4[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_10_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_1/temp3[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_10_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[98] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_10_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[122] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_10_2  ( .A(\MC_ARK_ARC_1_1/temp5[129] ), .B(
        \MC_ARK_ARC_1_1/temp6[129] ), .ZN(\RI1[2][129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_10_2  ( .A(\MC_ARK_ARC_1_1/temp3[129] ), .B(
        \MC_ARK_ARC_1_1/temp4[129] ), .ZN(\MC_ARK_ARC_1_1/temp6[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_10_2  ( .A(\MC_ARK_ARC_1_1/temp1[129] ), .B(
        \MC_ARK_ARC_1_1/temp2[129] ), .ZN(\MC_ARK_ARC_1_1/temp5[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_10_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[165] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[129] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_10_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[39] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[3] ), .ZN(\MC_ARK_ARC_1_1/temp3[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_10_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .B(\RI5[1][75] ), .ZN(\MC_ARK_ARC_1_1/temp2[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_10_2  ( .A(\RI5[1][123] ), .B(\RI5[1][129] ), 
        .ZN(\MC_ARK_ARC_1_1/temp1[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_10_1  ( .A(\MC_ARK_ARC_1_1/temp5[130] ), .B(
        \MC_ARK_ARC_1_1/temp6[130] ), .ZN(\RI1[2][130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_10_1  ( .A(\MC_ARK_ARC_1_1/temp3[130] ), .B(
        \MC_ARK_ARC_1_1/temp4[130] ), .ZN(\MC_ARK_ARC_1_1/temp6[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_10_1  ( .A(\MC_ARK_ARC_1_1/temp1[130] ), .B(
        \MC_ARK_ARC_1_1/temp2[130] ), .ZN(\MC_ARK_ARC_1_1/temp5[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_10_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[166] ), 
        .B(n497), .ZN(\MC_ARK_ARC_1_1/temp4[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_10_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_1/temp3[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_10_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[76] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_10_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[130] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_10_0  ( .A(\MC_ARK_ARC_1_1/temp5[131] ), .B(
        \MC_ARK_ARC_1_1/temp6[131] ), .ZN(\RI1[2][131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_10_0  ( .A(\MC_ARK_ARC_1_1/temp4[131] ), .B(
        \MC_ARK_ARC_1_1/temp3[131] ), .ZN(\MC_ARK_ARC_1_1/temp6[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_10_0  ( .A(\MC_ARK_ARC_1_1/temp1[131] ), .B(
        \MC_ARK_ARC_1_1/temp2[131] ), .ZN(\MC_ARK_ARC_1_1/temp5[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_10_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[167] ), 
        .B(n257), .ZN(\MC_ARK_ARC_1_1/temp4[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_10_0  ( .A(n1498), .B(
        \MC_ARK_ARC_1_1/buf_datainput[5] ), .ZN(\MC_ARK_ARC_1_1/temp3[131] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_10_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[77] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[101] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_10_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[125] ), 
        .B(n1655), .ZN(\MC_ARK_ARC_1_1/temp1[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_9_5  ( .A(\MC_ARK_ARC_1_1/temp5[132] ), .B(
        \MC_ARK_ARC_1_1/temp6[132] ), .ZN(\RI1[2][132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_9_5  ( .A(\MC_ARK_ARC_1_1/temp3[132] ), .B(
        \MC_ARK_ARC_1_1/temp4[132] ), .ZN(\MC_ARK_ARC_1_1/temp6[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_9_5  ( .A(\MC_ARK_ARC_1_1/temp1[132] ), .B(
        \MC_ARK_ARC_1_1/temp2[132] ), .ZN(\MC_ARK_ARC_1_1/temp5[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_9_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .B(n470), .ZN(\MC_ARK_ARC_1_1/temp4[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_9_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_1/temp3[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_9_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[78] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_9_5  ( .A(\RI5[1][132] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[126] ), .ZN(\MC_ARK_ARC_1_1/temp1[132] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_9_4  ( .A(\MC_ARK_ARC_1_1/temp5[133] ), .B(
        \MC_ARK_ARC_1_1/temp6[133] ), .ZN(\RI1[2][133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_9_4  ( .A(\MC_ARK_ARC_1_1/temp3[133] ), .B(
        \MC_ARK_ARC_1_1/temp4[133] ), .ZN(\MC_ARK_ARC_1_1/temp6[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_9_4  ( .A(\MC_ARK_ARC_1_1/temp1[133] ), .B(
        \MC_ARK_ARC_1_1/temp2[133] ), .ZN(\MC_ARK_ARC_1_1/temp5[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_9_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[169] ), 
        .B(n403), .ZN(\MC_ARK_ARC_1_1/temp4[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_9_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_1/temp3[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_9_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[79] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_9_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[133] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[127] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_9_3  ( .A(\MC_ARK_ARC_1_1/temp1[134] ), .B(
        \MC_ARK_ARC_1_1/temp2[134] ), .ZN(\MC_ARK_ARC_1_1/temp5[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_9_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[170] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[134] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_9_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[44] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_1/temp3[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_9_3  ( .A(n1646), .B(
        \MC_ARK_ARC_1_1/buf_datainput[104] ), .ZN(\MC_ARK_ARC_1_1/temp2[134] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_9_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[134] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_9_2  ( .A(\MC_ARK_ARC_1_1/temp5[135] ), .B(
        \MC_ARK_ARC_1_1/temp6[135] ), .ZN(\RI1[2][135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_9_2  ( .A(\MC_ARK_ARC_1_1/temp3[135] ), .B(
        \MC_ARK_ARC_1_1/temp4[135] ), .ZN(\MC_ARK_ARC_1_1/temp6[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_9_2  ( .A(\MC_ARK_ARC_1_1/temp1[135] ), .B(
        \MC_ARK_ARC_1_1/temp2[135] ), .ZN(\MC_ARK_ARC_1_1/temp5[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_9_2  ( .A(n1954), .B(n253), .ZN(
        \MC_ARK_ARC_1_1/temp4[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_9_2  ( .A(\RI5[1][9] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[45] ), .ZN(\MC_ARK_ARC_1_1/temp3[135] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_9_2  ( .A(\RI5[1][81] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[105] ), .ZN(\MC_ARK_ARC_1_1/temp2[135] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_9_2  ( .A(\RI5[1][129] ), .B(\RI5[1][135] ), 
        .ZN(\MC_ARK_ARC_1_1/temp1[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_9_1  ( .A(\MC_ARK_ARC_1_1/temp5[136] ), .B(
        \MC_ARK_ARC_1_1/temp6[136] ), .ZN(\RI1[2][136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_9_1  ( .A(\MC_ARK_ARC_1_1/temp3[136] ), .B(
        \MC_ARK_ARC_1_1/temp4[136] ), .ZN(\MC_ARK_ARC_1_1/temp6[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_9_1  ( .A(\MC_ARK_ARC_1_1/temp2[136] ), .B(
        \MC_ARK_ARC_1_1/temp1[136] ), .ZN(\MC_ARK_ARC_1_1/temp5[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_9_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[172] ), 
        .B(n421), .ZN(\MC_ARK_ARC_1_1/temp4[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_9_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[46] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[10] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_9_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[106] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_9_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_9_0  ( .A(\MC_ARK_ARC_1_1/temp6[137] ), .B(
        \MC_ARK_ARC_1_1/temp5[137] ), .ZN(\RI1[2][137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_9_0  ( .A(\MC_ARK_ARC_1_1/temp3[137] ), .B(
        \MC_ARK_ARC_1_1/temp4[137] ), .ZN(\MC_ARK_ARC_1_1/temp6[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_9_0  ( .A(\MC_ARK_ARC_1_1/temp1[137] ), .B(
        \MC_ARK_ARC_1_1/temp2[137] ), .ZN(\MC_ARK_ARC_1_1/temp5[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_9_0  ( .A(n1937), .B(n504), .ZN(
        \MC_ARK_ARC_1_1/temp4[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_9_0  ( .A(n2104), .B(
        \MC_ARK_ARC_1_1/buf_datainput[47] ), .ZN(\MC_ARK_ARC_1_1/temp3[137] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_9_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[83] ), 
        .B(n853), .ZN(\MC_ARK_ARC_1_1/temp2[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_9_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[137] ), 
        .B(n1655), .ZN(\MC_ARK_ARC_1_1/temp1[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_8_5  ( .A(\MC_ARK_ARC_1_1/temp5[138] ), .B(
        \MC_ARK_ARC_1_1/temp6[138] ), .ZN(\RI1[2][138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_8_5  ( .A(\MC_ARK_ARC_1_1/temp3[138] ), .B(
        \MC_ARK_ARC_1_1/temp4[138] ), .ZN(\MC_ARK_ARC_1_1/temp6[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_8_5  ( .A(\MC_ARK_ARC_1_1/temp1[138] ), .B(
        \MC_ARK_ARC_1_1/temp2[138] ), .ZN(\MC_ARK_ARC_1_1/temp5[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_8_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[174] ), 
        .B(n297), .ZN(\MC_ARK_ARC_1_1/temp4[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_8_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[12] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_8_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[108] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[84] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_8_5  ( .A(\RI5[1][138] ), .B(\RI5[1][132] ), 
        .ZN(\MC_ARK_ARC_1_1/temp1[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_8_4  ( .A(\MC_ARK_ARC_1_1/temp5[139] ), .B(
        \MC_ARK_ARC_1_1/temp6[139] ), .ZN(\RI1[2][139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_8_4  ( .A(\MC_ARK_ARC_1_1/temp3[139] ), .B(
        \MC_ARK_ARC_1_1/temp4[139] ), .ZN(\MC_ARK_ARC_1_1/temp6[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_8_4  ( .A(\MC_ARK_ARC_1_1/temp1[139] ), .B(
        \MC_ARK_ARC_1_1/temp2[139] ), .ZN(\MC_ARK_ARC_1_1/temp5[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_8_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[175] ), 
        .B(n250), .ZN(\MC_ARK_ARC_1_1/temp4[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_8_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[13] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_8_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[85] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_8_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[133] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_8_3  ( .A(\MC_ARK_ARC_1_1/temp5[140] ), .B(
        \MC_ARK_ARC_1_1/temp6[140] ), .ZN(\RI1[2][140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_8_3  ( .A(\MC_ARK_ARC_1_1/temp3[140] ), .B(
        \MC_ARK_ARC_1_1/temp4[140] ), .ZN(\MC_ARK_ARC_1_1/temp6[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_8_3  ( .A(\MC_ARK_ARC_1_1/temp2[140] ), .B(
        \MC_ARK_ARC_1_1/temp1[140] ), .ZN(\MC_ARK_ARC_1_1/temp5[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_8_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[129] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_8_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[50] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_8_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[110] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_8_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[140] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_8_2  ( .A(\MC_ARK_ARC_1_1/temp5[141] ), .B(
        \MC_ARK_ARC_1_1/temp6[141] ), .ZN(\RI1[2][141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_8_2  ( .A(\MC_ARK_ARC_1_1/temp3[141] ), .B(
        \MC_ARK_ARC_1_1/temp4[141] ), .ZN(\MC_ARK_ARC_1_1/temp6[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_8_2  ( .A(\MC_ARK_ARC_1_1/temp1[141] ), .B(
        \MC_ARK_ARC_1_1/temp2[141] ), .ZN(\MC_ARK_ARC_1_1/temp5[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_8_2  ( .A(\RI5[1][177] ), .B(n339), .ZN(
        \MC_ARK_ARC_1_1/temp4[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_8_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .B(\RI5[1][51] ), .ZN(\MC_ARK_ARC_1_1/temp3[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_8_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[111] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[87] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_8_2  ( .A(\RI5[1][141] ), .B(\RI5[1][135] ), 
        .ZN(\MC_ARK_ARC_1_1/temp1[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_8_1  ( .A(\MC_ARK_ARC_1_1/temp5[142] ), .B(
        \MC_ARK_ARC_1_1/temp6[142] ), .ZN(\RI1[2][142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_8_1  ( .A(\MC_ARK_ARC_1_1/temp4[142] ), .B(
        \MC_ARK_ARC_1_1/temp3[142] ), .ZN(\MC_ARK_ARC_1_1/temp6[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_8_1  ( .A(\MC_ARK_ARC_1_1/temp2[142] ), .B(
        \MC_ARK_ARC_1_1/temp1[142] ), .ZN(\MC_ARK_ARC_1_1/temp5[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_8_1  ( .A(n1953), .B(n293), .ZN(
        \MC_ARK_ARC_1_1/temp4[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_8_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[52] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_8_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[88] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_8_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[136] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_8_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[179] ), 
        .B(n510), .ZN(\MC_ARK_ARC_1_1/temp4[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_8_0  ( .A(n1643), .B(n837), .ZN(
        \MC_ARK_ARC_1_1/temp3[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_8_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .B(n808), .ZN(\MC_ARK_ARC_1_1/temp2[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_8_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[143] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_7_5  ( .A(\MC_ARK_ARC_1_1/temp5[144] ), .B(
        \MC_ARK_ARC_1_1/temp6[144] ), .ZN(\RI1[2][144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_7_5  ( .A(\MC_ARK_ARC_1_1/temp3[144] ), .B(
        \MC_ARK_ARC_1_1/temp4[144] ), .ZN(\MC_ARK_ARC_1_1/temp6[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_7_5  ( .A(\MC_ARK_ARC_1_1/temp1[144] ), .B(
        \MC_ARK_ARC_1_1/temp2[144] ), .ZN(\MC_ARK_ARC_1_1/temp5[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_7_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[180] ), 
        .B(n474), .ZN(\MC_ARK_ARC_1_1/temp4[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_7_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[18] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_7_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[90] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_7_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[144] ), 
        .B(\RI5[1][138] ), .ZN(\MC_ARK_ARC_1_1/temp1[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_7_4  ( .A(\MC_ARK_ARC_1_1/temp5[145] ), .B(
        \MC_ARK_ARC_1_1/temp6[145] ), .ZN(\RI1[2][145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_7_4  ( .A(\MC_ARK_ARC_1_1/temp3[145] ), .B(
        \MC_ARK_ARC_1_1/temp4[145] ), .ZN(\MC_ARK_ARC_1_1/temp6[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_7_4  ( .A(\MC_ARK_ARC_1_1/temp1[145] ), .B(
        \MC_ARK_ARC_1_1/temp2[145] ), .ZN(\MC_ARK_ARC_1_1/temp5[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_7_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[181] ), 
        .B(n336), .ZN(\MC_ARK_ARC_1_1/temp4[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_7_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[19] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_7_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[91] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_7_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[139] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_7_3  ( .A(\MC_ARK_ARC_1_1/temp5[146] ), .B(
        \MC_ARK_ARC_1_1/temp6[146] ), .ZN(\RI1[2][146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_7_3  ( .A(\MC_ARK_ARC_1_1/temp3[146] ), .B(
        \MC_ARK_ARC_1_1/temp4[146] ), .ZN(\MC_ARK_ARC_1_1/temp6[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_7_3  ( .A(\MC_ARK_ARC_1_1/temp2[146] ), .B(
        \MC_ARK_ARC_1_1/temp1[146] ), .ZN(\MC_ARK_ARC_1_1/temp5[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_7_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[182] ), 
        .B(n289), .ZN(\MC_ARK_ARC_1_1/temp4[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_7_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[20] ), 
        .B(\RI5[1][56] ), .ZN(\MC_ARK_ARC_1_1/temp3[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_7_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[92] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_7_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[146] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_7_2  ( .A(\MC_ARK_ARC_1_1/temp5[147] ), .B(
        \MC_ARK_ARC_1_1/temp6[147] ), .ZN(\RI1[2][147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_7_2  ( .A(\MC_ARK_ARC_1_1/temp3[147] ), .B(
        \MC_ARK_ARC_1_1/temp4[147] ), .ZN(\MC_ARK_ARC_1_1/temp6[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_7_2  ( .A(\MC_ARK_ARC_1_1/temp2[147] ), .B(
        \MC_ARK_ARC_1_1/temp1[147] ), .ZN(\MC_ARK_ARC_1_1/temp5[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_7_2  ( .A(n1958), .B(n243), .ZN(
        \MC_ARK_ARC_1_1/temp4[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_7_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[21] ), 
        .B(\RI5[1][57] ), .ZN(\MC_ARK_ARC_1_1/temp3[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_7_2  ( .A(\RI5[1][117] ), .B(\RI5[1][93] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_7_2  ( .A(\RI5[1][147] ), .B(\RI5[1][141] ), 
        .ZN(\MC_ARK_ARC_1_1/temp1[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_7_1  ( .A(\MC_ARK_ARC_1_1/temp5[148] ), .B(
        \MC_ARK_ARC_1_1/temp6[148] ), .ZN(\RI1[2][148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_7_1  ( .A(\MC_ARK_ARC_1_1/temp3[148] ), .B(
        \MC_ARK_ARC_1_1/temp4[148] ), .ZN(\MC_ARK_ARC_1_1/temp6[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_7_1  ( .A(\MC_ARK_ARC_1_1/temp2[148] ), .B(
        \MC_ARK_ARC_1_1/temp1[148] ), .ZN(\MC_ARK_ARC_1_1/temp5[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_7_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[184] ), 
        .B(n498), .ZN(\MC_ARK_ARC_1_1/temp4[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_7_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[22] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_7_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[118] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[94] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_7_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[142] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_7_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[185] ), 
        .B(n453), .ZN(\MC_ARK_ARC_1_1/temp4[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_7_0  ( .A(n1925), .B(
        \MC_ARK_ARC_1_1/buf_datainput[59] ), .ZN(\MC_ARK_ARC_1_1/temp3[149] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_7_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[119] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_7_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[149] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[143] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_6_5  ( .A(\MC_ARK_ARC_1_1/temp5[150] ), .B(
        \MC_ARK_ARC_1_1/temp6[150] ), .ZN(\RI1[2][150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_6_5  ( .A(\MC_ARK_ARC_1_1/temp3[150] ), .B(
        \MC_ARK_ARC_1_1/temp4[150] ), .ZN(\MC_ARK_ARC_1_1/temp6[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_6_5  ( .A(\MC_ARK_ARC_1_1/temp1[150] ), .B(
        \MC_ARK_ARC_1_1/temp2[150] ), .ZN(\MC_ARK_ARC_1_1/temp5[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_6_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[186] ), 
        .B(n285), .ZN(\MC_ARK_ARC_1_1/temp4[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_6_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[60] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[24] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_6_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[96] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_6_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[144] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_6_4  ( .A(\MC_ARK_ARC_1_1/temp5[151] ), .B(
        \MC_ARK_ARC_1_1/temp6[151] ), .ZN(\RI1[2][151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_6_4  ( .A(\MC_ARK_ARC_1_1/temp3[151] ), .B(
        \MC_ARK_ARC_1_1/temp4[151] ), .ZN(\MC_ARK_ARC_1_1/temp6[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_6_4  ( .A(\MC_ARK_ARC_1_1/temp2[151] ), .B(
        \MC_ARK_ARC_1_1/temp1[151] ), .ZN(\MC_ARK_ARC_1_1/temp5[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_6_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .B(n395), .ZN(\MC_ARK_ARC_1_1/temp4[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_6_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[25] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_6_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[97] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_6_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[145] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_6_3  ( .A(\MC_ARK_ARC_1_1/temp6[152] ), .B(
        \MC_ARK_ARC_1_1/temp5[152] ), .ZN(\RI1[2][152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_6_3  ( .A(\MC_ARK_ARC_1_1/temp4[152] ), .B(
        \MC_ARK_ARC_1_1/temp3[152] ), .ZN(\MC_ARK_ARC_1_1/temp6[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_6_3  ( .A(\MC_ARK_ARC_1_1/temp2[152] ), .B(
        \MC_ARK_ARC_1_1/temp1[152] ), .ZN(\MC_ARK_ARC_1_1/temp5[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_6_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[152] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_6_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[26] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_6_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[98] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[122] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_6_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_6_2  ( .A(\MC_ARK_ARC_1_1/temp5[153] ), .B(
        \MC_ARK_ARC_1_1/temp6[153] ), .ZN(\RI1[2][153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_6_2  ( .A(\MC_ARK_ARC_1_1/temp3[153] ), .B(
        \MC_ARK_ARC_1_1/temp4[153] ), .ZN(\MC_ARK_ARC_1_1/temp6[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_6_2  ( .A(\MC_ARK_ARC_1_1/temp2[153] ), .B(
        \MC_ARK_ARC_1_1/temp1[153] ), .ZN(\MC_ARK_ARC_1_1/temp5[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_6_2  ( .A(n1934), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[76] ), .ZN(\MC_ARK_ARC_1_1/temp4[153] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_6_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[63] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_6_2  ( .A(\RI5[1][123] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[99] ), .ZN(\MC_ARK_ARC_1_1/temp2[153] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_6_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .B(\RI5[1][147] ), .ZN(\MC_ARK_ARC_1_1/temp1[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_6_1  ( .A(\MC_ARK_ARC_1_1/temp5[154] ), .B(
        \MC_ARK_ARC_1_1/temp6[154] ), .ZN(\RI1[2][154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_6_1  ( .A(\MC_ARK_ARC_1_1/temp3[154] ), .B(
        \MC_ARK_ARC_1_1/temp4[154] ), .ZN(\MC_ARK_ARC_1_1/temp6[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_6_1  ( .A(\MC_ARK_ARC_1_1/temp1[154] ), .B(
        \MC_ARK_ARC_1_1/temp2[154] ), .ZN(\MC_ARK_ARC_1_1/temp5[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_6_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[190] ), 
        .B(n282), .ZN(\MC_ARK_ARC_1_1/temp4[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_6_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[28] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_6_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_6_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_6_0  ( .A(n514), .B(n236), .ZN(
        \MC_ARK_ARC_1_1/temp4[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_6_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[65] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_6_0  ( .A(n2124), .B(
        \MC_ARK_ARC_1_1/buf_datainput[125] ), .ZN(\MC_ARK_ARC_1_1/temp2[155] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_6_0  ( .A(n2152), .B(
        \MC_ARK_ARC_1_1/buf_datainput[149] ), .ZN(\MC_ARK_ARC_1_1/temp1[155] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_5_5  ( .A(\MC_ARK_ARC_1_1/temp5[156] ), .B(
        \MC_ARK_ARC_1_1/temp6[156] ), .ZN(\RI1[2][156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_5_5  ( .A(\MC_ARK_ARC_1_1/temp3[156] ), .B(
        \MC_ARK_ARC_1_1/temp4[156] ), .ZN(\MC_ARK_ARC_1_1/temp6[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_5_5  ( .A(\MC_ARK_ARC_1_1/temp1[156] ), .B(
        \MC_ARK_ARC_1_1/temp2[156] ), .ZN(\MC_ARK_ARC_1_1/temp5[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_5_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .B(n432), .ZN(\MC_ARK_ARC_1_1/temp4[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_5_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[30] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_5_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[102] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_5_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[156] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[150] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_5_4  ( .A(\MC_ARK_ARC_1_1/temp5[157] ), .B(
        \MC_ARK_ARC_1_1/temp6[157] ), .ZN(\RI1[2][157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_5_4  ( .A(\MC_ARK_ARC_1_1/temp3[157] ), .B(
        \MC_ARK_ARC_1_1/temp4[157] ), .ZN(\MC_ARK_ARC_1_1/temp6[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_5_4  ( .A(\MC_ARK_ARC_1_1/temp1[157] ), .B(
        \MC_ARK_ARC_1_1/temp2[157] ), .ZN(\MC_ARK_ARC_1_1/temp5[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_5_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .B(n324), .ZN(\MC_ARK_ARC_1_1/temp4[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_5_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[31] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_5_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_5_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[157] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[151] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_5_3  ( .A(\MC_ARK_ARC_1_1/temp3[158] ), .B(
        \MC_ARK_ARC_1_1/temp4[158] ), .ZN(\MC_ARK_ARC_1_1/temp6[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_5_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[2] ), 
        .B(n278), .ZN(\MC_ARK_ARC_1_1/temp4[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_5_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[68] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_5_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_5_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[158] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_5_2  ( .A(\MC_ARK_ARC_1_1/temp2[159] ), .B(
        \MC_ARK_ARC_1_1/temp1[159] ), .ZN(\MC_ARK_ARC_1_1/temp5[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_5_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[3] ), 
        .B(n232), .ZN(\MC_ARK_ARC_1_1/temp4[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_5_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[69] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_5_2  ( .A(\RI5[1][129] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[105] ), .ZN(\MC_ARK_ARC_1_1/temp2[159] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_5_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[159] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_5_1  ( .A(\MC_ARK_ARC_1_1/temp5[160] ), .B(
        \MC_ARK_ARC_1_1/temp6[160] ), .ZN(\RI1[2][160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_5_1  ( .A(\MC_ARK_ARC_1_1/temp3[160] ), .B(
        \MC_ARK_ARC_1_1/temp4[160] ), .ZN(\MC_ARK_ARC_1_1/temp6[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_5_1  ( .A(\MC_ARK_ARC_1_1/temp1[160] ), .B(
        \MC_ARK_ARC_1_1/temp2[160] ), .ZN(\MC_ARK_ARC_1_1/temp5[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_5_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .B(n499), .ZN(\MC_ARK_ARC_1_1/temp4[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_5_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[34] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_5_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[130] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[106] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_5_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_5_0  ( .A(\MC_ARK_ARC_1_1/temp5[161] ), .B(
        \MC_ARK_ARC_1_1/temp6[161] ), .ZN(\RI1[2][161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_5_0  ( .A(\MC_ARK_ARC_1_1/temp3[161] ), .B(
        \MC_ARK_ARC_1_1/temp4[161] ), .ZN(\MC_ARK_ARC_1_1/temp6[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_5_0  ( .A(\MC_ARK_ARC_1_1/temp1[161] ), .B(
        \MC_ARK_ARC_1_1/temp2[161] ), .ZN(\MC_ARK_ARC_1_1/temp5[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_5_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[5] ), 
        .B(n444), .ZN(\MC_ARK_ARC_1_1/temp4[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_5_0  ( .A(n1505), .B(n519), .ZN(
        \MC_ARK_ARC_1_1/temp3[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_5_0  ( .A(n1655), .B(n853), .ZN(
        \MC_ARK_ARC_1_1/temp2[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_5_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[161] ), 
        .B(n2152), .ZN(\MC_ARK_ARC_1_1/temp1[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_4_5  ( .A(\MC_ARK_ARC_1_1/temp5[162] ), .B(
        \MC_ARK_ARC_1_1/temp6[162] ), .ZN(\RI1[2][162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_4_5  ( .A(\MC_ARK_ARC_1_1/temp3[162] ), .B(
        \MC_ARK_ARC_1_1/temp4[162] ), .ZN(\MC_ARK_ARC_1_1/temp6[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_4_5  ( .A(\MC_ARK_ARC_1_1/temp1[162] ), .B(
        \MC_ARK_ARC_1_1/temp2[162] ), .ZN(\MC_ARK_ARC_1_1/temp5[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_4_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[6] ), 
        .B(n446), .ZN(\MC_ARK_ARC_1_1/temp4[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_4_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[36] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_4_5  ( .A(\RI5[1][132] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[108] ), .ZN(\MC_ARK_ARC_1_1/temp2[162] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_4_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[162] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[156] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_4_4  ( .A(\MC_ARK_ARC_1_1/temp5[163] ), .B(
        \MC_ARK_ARC_1_1/temp6[163] ), .ZN(\RI1[2][163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_4_4  ( .A(\MC_ARK_ARC_1_1/temp3[163] ), .B(
        \MC_ARK_ARC_1_1/temp4[163] ), .ZN(\MC_ARK_ARC_1_1/temp6[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_4_4  ( .A(\MC_ARK_ARC_1_1/temp1[163] ), .B(
        \MC_ARK_ARC_1_1/temp2[163] ), .ZN(\MC_ARK_ARC_1_1/temp5[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_4_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[7] ), 
        .B(n228), .ZN(\MC_ARK_ARC_1_1/temp4[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_4_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[37] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_4_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[133] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_4_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[157] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_4_3  ( .A(\MC_ARK_ARC_1_1/temp6[164] ), .B(
        \MC_ARK_ARC_1_1/temp5[164] ), .ZN(\RI1[2][164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_4_3  ( .A(\MC_ARK_ARC_1_1/temp3[164] ), .B(
        \MC_ARK_ARC_1_1/temp4[164] ), .ZN(\MC_ARK_ARC_1_1/temp6[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_4_3  ( .A(\MC_ARK_ARC_1_1/temp2[164] ), .B(
        \MC_ARK_ARC_1_1/temp1[164] ), .ZN(\MC_ARK_ARC_1_1/temp5[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_4_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[8] ), 
        .B(n363), .ZN(\MC_ARK_ARC_1_1/temp4[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_4_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[38] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_4_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[110] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_4_3  ( .A(n1624), .B(
        \MC_ARK_ARC_1_1/buf_datainput[158] ), .ZN(\MC_ARK_ARC_1_1/temp1[164] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_4_2  ( .A(\MC_ARK_ARC_1_1/temp5[165] ), .B(
        \MC_ARK_ARC_1_1/temp6[165] ), .ZN(\RI1[2][165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_4_2  ( .A(\MC_ARK_ARC_1_1/temp3[165] ), .B(
        \MC_ARK_ARC_1_1/temp4[165] ), .ZN(\MC_ARK_ARC_1_1/temp6[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_4_2  ( .A(\MC_ARK_ARC_1_1/temp1[165] ), .B(
        \MC_ARK_ARC_1_1/temp2[165] ), .ZN(\MC_ARK_ARC_1_1/temp5[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_4_2  ( .A(\RI5[1][9] ), .B(
        \MC_ARK_ARC_1_1/buf_keyinput[165] ), .ZN(\MC_ARK_ARC_1_1/temp4[165] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_4_2  ( .A(\RI5[1][75] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[39] ), .ZN(\MC_ARK_ARC_1_1/temp3[165] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_4_2  ( .A(\RI5[1][135] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[111] ), .ZN(\MC_ARK_ARC_1_1/temp2[165] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_4_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[165] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[159] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_4_1  ( .A(\MC_ARK_ARC_1_1/temp5[166] ), .B(
        \MC_ARK_ARC_1_1/temp6[166] ), .ZN(\RI1[2][166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_4_1  ( .A(\MC_ARK_ARC_1_1/temp3[166] ), .B(
        \MC_ARK_ARC_1_1/temp4[166] ), .ZN(\MC_ARK_ARC_1_1/temp6[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_4_1  ( .A(\MC_ARK_ARC_1_1/temp1[166] ), .B(
        \MC_ARK_ARC_1_1/temp2[166] ), .ZN(\MC_ARK_ARC_1_1/temp5[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_4_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[10] ), 
        .B(n501), .ZN(\MC_ARK_ARC_1_1/temp4[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_4_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[76] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[40] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_4_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[112] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_4_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_4_0  ( .A(\MC_ARK_ARC_1_1/temp3[167] ), .B(
        \MC_ARK_ARC_1_1/temp4[167] ), .ZN(\MC_ARK_ARC_1_1/temp6[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_4_0  ( .A(\MC_ARK_ARC_1_1/temp1[167] ), .B(
        \MC_ARK_ARC_1_1/temp2[167] ), .ZN(\MC_ARK_ARC_1_1/temp5[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_4_0  ( .A(n2105), .B(n224), .ZN(
        \MC_ARK_ARC_1_1/temp4[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_4_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[77] ), 
        .B(n1498), .ZN(\MC_ARK_ARC_1_1/temp3[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_4_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[137] ), 
        .B(n807), .ZN(\MC_ARK_ARC_1_1/temp2[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_4_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[161] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[167] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_3_5  ( .A(\MC_ARK_ARC_1_1/temp5[168] ), .B(
        \MC_ARK_ARC_1_1/temp6[168] ), .ZN(\RI1[2][168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_3_5  ( .A(\MC_ARK_ARC_1_1/temp3[168] ), .B(
        \MC_ARK_ARC_1_1/temp4[168] ), .ZN(\MC_ARK_ARC_1_1/temp6[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_3_5  ( .A(\MC_ARK_ARC_1_1/temp1[168] ), .B(
        \MC_ARK_ARC_1_1/temp2[168] ), .ZN(\MC_ARK_ARC_1_1/temp5[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_3_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[12] ), 
        .B(n452), .ZN(\MC_ARK_ARC_1_1/temp4[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_3_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[42] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_3_5  ( .A(\RI5[1][138] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[114] ), .ZN(\MC_ARK_ARC_1_1/temp2[168] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_3_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_3_4  ( .A(\MC_ARK_ARC_1_1/temp5[169] ), .B(
        \MC_ARK_ARC_1_1/temp6[169] ), .ZN(\RI1[2][169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_3_4  ( .A(\MC_ARK_ARC_1_1/temp3[169] ), .B(
        \MC_ARK_ARC_1_1/temp4[169] ), .ZN(\MC_ARK_ARC_1_1/temp6[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_3_4  ( .A(\MC_ARK_ARC_1_1/temp1[169] ), .B(
        \MC_ARK_ARC_1_1/temp2[169] ), .ZN(\MC_ARK_ARC_1_1/temp5[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_3_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[13] ), 
        .B(n313), .ZN(\MC_ARK_ARC_1_1/temp4[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_3_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[43] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_3_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_3_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[169] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[163] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_3_3  ( .A(\MC_ARK_ARC_1_1/temp5[170] ), .B(
        \MC_ARK_ARC_1_1/temp6[170] ), .ZN(\RI1[2][170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_3_3  ( .A(\MC_ARK_ARC_1_1/temp3[170] ), .B(
        \MC_ARK_ARC_1_1/temp4[170] ), .ZN(\MC_ARK_ARC_1_1/temp6[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_3_3  ( .A(\MC_ARK_ARC_1_1/temp2[170] ), .B(
        \MC_ARK_ARC_1_1/temp1[170] ), .ZN(\MC_ARK_ARC_1_1/temp5[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_3_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[170] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_3_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[44] ), 
        .B(n1645), .ZN(\MC_ARK_ARC_1_1/temp3[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_3_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[116] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_3_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[170] ), 
        .B(n1625), .ZN(\MC_ARK_ARC_1_1/temp1[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_3_2  ( .A(\MC_ARK_ARC_1_1/temp5[171] ), .B(
        \MC_ARK_ARC_1_1/temp6[171] ), .ZN(\RI1[2][171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_3_2  ( .A(\MC_ARK_ARC_1_1/temp3[171] ), .B(
        \MC_ARK_ARC_1_1/temp4[171] ), .ZN(\MC_ARK_ARC_1_1/temp6[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_3_2  ( .A(\MC_ARK_ARC_1_1/temp2[171] ), .B(
        \MC_ARK_ARC_1_1/temp1[171] ), .ZN(\MC_ARK_ARC_1_1/temp5[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_3_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .B(n220), .ZN(\MC_ARK_ARC_1_1/temp4[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_3_2  ( .A(\RI5[1][81] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[45] ), .ZN(\MC_ARK_ARC_1_1/temp3[171] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_3_2  ( .A(\RI5[1][141] ), .B(\RI5[1][117] ), 
        .ZN(\MC_ARK_ARC_1_1/temp2[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_3_2  ( .A(n1954), .B(
        \MC_ARK_ARC_1_1/buf_datainput[165] ), .ZN(\MC_ARK_ARC_1_1/temp1[171] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_3_1  ( .A(\MC_ARK_ARC_1_1/temp5[172] ), .B(
        \MC_ARK_ARC_1_1/temp6[172] ), .ZN(\RI1[2][172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_3_1  ( .A(\MC_ARK_ARC_1_1/temp3[172] ), .B(
        \MC_ARK_ARC_1_1/temp4[172] ), .ZN(\MC_ARK_ARC_1_1/temp6[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_3_1  ( .A(\MC_ARK_ARC_1_1/temp2[172] ), .B(
        \MC_ARK_ARC_1_1/temp1[172] ), .ZN(\MC_ARK_ARC_1_1/temp5[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_3_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[16] ), 
        .B(n355), .ZN(\MC_ARK_ARC_1_1/temp4[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_3_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[46] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_3_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[118] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_3_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_3_0  ( .A(\MC_ARK_ARC_1_1/temp5[173] ), .B(
        \MC_ARK_ARC_1_1/temp6[173] ), .ZN(\RI1[2][173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_3_0  ( .A(\MC_ARK_ARC_1_1/temp3[173] ), .B(
        \MC_ARK_ARC_1_1/temp4[173] ), .ZN(\MC_ARK_ARC_1_1/temp6[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_3_0  ( .A(\MC_ARK_ARC_1_1/temp2[173] ), .B(
        \MC_ARK_ARC_1_1/temp1[173] ), .ZN(\MC_ARK_ARC_1_1/temp5[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_3_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[17] ), 
        .B(n309), .ZN(\MC_ARK_ARC_1_1/temp4[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_3_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[47] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[83] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_3_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[119] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[143] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_3_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[167] ), 
        .B(n1936), .ZN(\MC_ARK_ARC_1_1/temp1[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_2_5  ( .A(\MC_ARK_ARC_1_1/temp5[174] ), .B(
        \MC_ARK_ARC_1_1/temp6[174] ), .ZN(\RI1[2][174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_2_5  ( .A(\MC_ARK_ARC_1_1/temp3[174] ), .B(
        \MC_ARK_ARC_1_1/temp4[174] ), .ZN(\MC_ARK_ARC_1_1/temp6[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_2_5  ( .A(\MC_ARK_ARC_1_1/temp1[174] ), .B(
        \MC_ARK_ARC_1_1/temp2[174] ), .ZN(\MC_ARK_ARC_1_1/temp5[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_2_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[18] ), 
        .B(n262), .ZN(\MC_ARK_ARC_1_1/temp4[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_2_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[48] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_2_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[144] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_2_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[174] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_2_4  ( .A(\MC_ARK_ARC_1_1/temp5[175] ), .B(
        \MC_ARK_ARC_1_1/temp6[175] ), .ZN(\RI1[2][175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_2_4  ( .A(\MC_ARK_ARC_1_1/temp3[175] ), .B(
        \MC_ARK_ARC_1_1/temp4[175] ), .ZN(\MC_ARK_ARC_1_1/temp6[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_2_4  ( .A(\MC_ARK_ARC_1_1/temp1[175] ), .B(
        \MC_ARK_ARC_1_1/temp2[175] ), .ZN(\MC_ARK_ARC_1_1/temp5[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_2_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[19] ), 
        .B(n216), .ZN(\MC_ARK_ARC_1_1/temp4[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_2_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[49] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_2_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_2_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[169] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_2_3  ( .A(\MC_ARK_ARC_1_1/temp5[176] ), .B(
        \MC_ARK_ARC_1_1/temp6[176] ), .ZN(\RI1[2][176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_2_3  ( .A(\MC_ARK_ARC_1_1/temp4[176] ), .B(
        \MC_ARK_ARC_1_1/temp3[176] ), .ZN(\MC_ARK_ARC_1_1/temp6[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_2_3  ( .A(\MC_ARK_ARC_1_1/temp2[176] ), .B(
        \MC_ARK_ARC_1_1/temp1[176] ), .ZN(\MC_ARK_ARC_1_1/temp5[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_2_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[176] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_2_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[86] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_2_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[146] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_2_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[170] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_2_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[21] ), 
        .B(n305), .ZN(\MC_ARK_ARC_1_1/temp4[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_2_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[87] ), 
        .B(\RI5[1][51] ), .ZN(\MC_ARK_ARC_1_1/temp3[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_2_2  ( .A(\RI5[1][123] ), .B(\RI5[1][147] ), 
        .ZN(\MC_ARK_ARC_1_1/temp2[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_2_2  ( .A(\RI5[1][177] ), .B(n1954), .ZN(
        \MC_ARK_ARC_1_1/temp1[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_2_1  ( .A(\MC_ARK_ARC_1_1/temp6[178] ), .B(
        \MC_ARK_ARC_1_1/temp5[178] ), .ZN(\RI1[2][178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_2_1  ( .A(\MC_ARK_ARC_1_1/temp3[178] ), .B(
        \MC_ARK_ARC_1_1/temp4[178] ), .ZN(\MC_ARK_ARC_1_1/temp6[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_2_1  ( .A(\MC_ARK_ARC_1_1/temp2[178] ), .B(
        \MC_ARK_ARC_1_1/temp1[178] ), .ZN(\MC_ARK_ARC_1_1/temp5[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_2_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .B(n258), .ZN(\MC_ARK_ARC_1_1/temp4[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_2_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[52] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_2_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_2_1  ( .A(n1953), .B(
        \MC_ARK_ARC_1_1/buf_datainput[172] ), .ZN(\MC_ARK_ARC_1_1/temp1[178] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_2_0  ( .A(n1926), .B(n212), .ZN(
        \MC_ARK_ARC_1_1/temp4[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_2_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .B(n838), .ZN(\MC_ARK_ARC_1_1/temp3[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_2_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[149] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[125] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_2_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[179] ), 
        .B(n1937), .ZN(\MC_ARK_ARC_1_1/temp1[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_1_5  ( .A(\MC_ARK_ARC_1_1/temp5[180] ), .B(
        \MC_ARK_ARC_1_1/temp6[180] ), .ZN(\RI1[2][180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_1_5  ( .A(\MC_ARK_ARC_1_1/temp3[180] ), .B(
        \MC_ARK_ARC_1_1/temp4[180] ), .ZN(\MC_ARK_ARC_1_1/temp6[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_1_5  ( .A(\MC_ARK_ARC_1_1/temp1[180] ), .B(
        \MC_ARK_ARC_1_1/temp2[180] ), .ZN(\MC_ARK_ARC_1_1/temp5[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_1_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[24] ), 
        .B(n448), .ZN(\MC_ARK_ARC_1_1/temp4[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_1_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[54] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_1_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[126] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_1_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[180] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[174] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_1_4  ( .A(\MC_ARK_ARC_1_1/temp5[181] ), .B(
        \MC_ARK_ARC_1_1/temp6[181] ), .ZN(\RI1[2][181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_1_4  ( .A(\MC_ARK_ARC_1_1/temp3[181] ), .B(
        \MC_ARK_ARC_1_1/temp4[181] ), .ZN(\MC_ARK_ARC_1_1/temp6[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_1_4  ( .A(\MC_ARK_ARC_1_1/temp1[181] ), .B(
        \MC_ARK_ARC_1_1/temp2[181] ), .ZN(\MC_ARK_ARC_1_1/temp5[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_1_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[25] ), 
        .B(n301), .ZN(\MC_ARK_ARC_1_1/temp4[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_1_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[55] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_1_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[127] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_1_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_1_3  ( .A(\MC_ARK_ARC_1_1/temp6[182] ), .B(
        \MC_ARK_ARC_1_1/temp5[182] ), .ZN(\RI1[2][182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_1_3  ( .A(\MC_ARK_ARC_1_1/temp3[182] ), .B(
        \MC_ARK_ARC_1_1/temp4[182] ), .ZN(\MC_ARK_ARC_1_1/temp6[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_1_3  ( .A(\MC_ARK_ARC_1_1/temp1[182] ), .B(
        \MC_ARK_ARC_1_1/temp2[182] ), .ZN(\MC_ARK_ARC_1_1/temp5[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_1_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[26] ), 
        .B(n383), .ZN(\MC_ARK_ARC_1_1/temp4[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_1_3  ( .A(\RI5[1][56] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[92] ), .ZN(\MC_ARK_ARC_1_1/temp3[182] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_1_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_1_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_1_2  ( .A(\MC_ARK_ARC_1_1/temp5[183] ), .B(
        \MC_ARK_ARC_1_1/temp6[183] ), .ZN(\RI1[2][183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_1_2  ( .A(\MC_ARK_ARC_1_1/temp3[183] ), .B(
        \MC_ARK_ARC_1_1/temp4[183] ), .ZN(\MC_ARK_ARC_1_1/temp6[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_1_2  ( .A(\MC_ARK_ARC_1_1/temp2[183] ), .B(
        \MC_ARK_ARC_1_1/temp1[183] ), .ZN(\MC_ARK_ARC_1_1/temp5[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_1_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[183] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_1_2  ( .A(\RI5[1][57] ), .B(\RI5[1][93] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_1_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .B(\RI5[1][129] ), .ZN(\MC_ARK_ARC_1_1/temp2[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_1_2  ( .A(\RI5[1][177] ), .B(n1958), .ZN(
        \MC_ARK_ARC_1_1/temp1[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_1_1  ( .A(\MC_ARK_ARC_1_1/temp5[184] ), .B(
        \MC_ARK_ARC_1_1/temp6[184] ), .ZN(\RI1[2][184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_1_1  ( .A(\MC_ARK_ARC_1_1/temp3[184] ), .B(
        \MC_ARK_ARC_1_1/temp4[184] ), .ZN(\MC_ARK_ARC_1_1/temp6[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_1_1  ( .A(\MC_ARK_ARC_1_1/temp1[184] ), .B(
        \MC_ARK_ARC_1_1/temp2[184] ), .ZN(\MC_ARK_ARC_1_1/temp5[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_1_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[28] ), 
        .B(n460), .ZN(\MC_ARK_ARC_1_1/temp4[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_1_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[58] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_1_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_1_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[184] ), 
        .B(n1953), .ZN(\MC_ARK_ARC_1_1/temp1[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_1_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .B(n488), .ZN(\MC_ARK_ARC_1_1/temp4[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_1_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[59] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_1_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[155] ), 
        .B(n1656), .ZN(\MC_ARK_ARC_1_1/temp2[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_1_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[179] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[185] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_0_5  ( .A(\MC_ARK_ARC_1_1/temp3[186] ), .B(
        \MC_ARK_ARC_1_1/temp4[186] ), .ZN(\MC_ARK_ARC_1_1/temp6[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_0_5  ( .A(\MC_ARK_ARC_1_1/temp1[186] ), .B(
        \MC_ARK_ARC_1_1/temp2[186] ), .ZN(\MC_ARK_ARC_1_1/temp5[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_0_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[30] ), 
        .B(n471), .ZN(\MC_ARK_ARC_1_1/temp4[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_0_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[60] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_0_5  ( .A(\RI5[1][132] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[156] ), .ZN(\MC_ARK_ARC_1_1/temp2[186] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_0_5  ( .A(\MC_ARK_ARC_1_1/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_0_4  ( .A(\MC_ARK_ARC_1_1/temp5[187] ), .B(
        \MC_ARK_ARC_1_1/temp6[187] ), .ZN(\RI1[2][187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_0_4  ( .A(\MC_ARK_ARC_1_1/temp3[187] ), .B(
        \MC_ARK_ARC_1_1/temp4[187] ), .ZN(\MC_ARK_ARC_1_1/temp6[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_0_4  ( .A(\MC_ARK_ARC_1_1/temp1[187] ), .B(
        \MC_ARK_ARC_1_1/temp2[187] ), .ZN(\MC_ARK_ARC_1_1/temp5[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_0_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .B(n204), .ZN(\MC_ARK_ARC_1_1/temp4[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_0_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[61] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_0_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[157] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[133] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_0_4  ( .A(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_0_3  ( .A(\MC_ARK_ARC_1_1/temp2[188] ), .B(
        \MC_ARK_ARC_1_1/temp1[188] ), .ZN(\MC_ARK_ARC_1_1/temp5[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_0_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[32] ), 
        .B(Key[36]), .ZN(\MC_ARK_ARC_1_1/temp4[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_0_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[98] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[62] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_0_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[158] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[134] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_0_3  ( .A(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_0_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[189] ), .ZN(
        \MC_ARK_ARC_1_1/temp4[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_0_2  ( .A(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[63] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_0_2  ( .A(\RI5[1][135] ), .B(
        \MC_ARK_ARC_1_1/buf_datainput[159] ), .ZN(\MC_ARK_ARC_1_1/temp2[189] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_0_2  ( .A(n1486), .B(n1935), .ZN(
        \MC_ARK_ARC_1_1/temp1[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X7_0_1  ( .A(\MC_ARK_ARC_1_1/temp5[190] ), .B(
        \MC_ARK_ARC_1_1/temp6[190] ), .ZN(\RI1[2][190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X6_0_1  ( .A(\MC_ARK_ARC_1_1/temp3[190] ), .B(
        \MC_ARK_ARC_1_1/temp4[190] ), .ZN(\MC_ARK_ARC_1_1/temp6[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X5_0_1  ( .A(\MC_ARK_ARC_1_1/temp2[190] ), .B(
        \MC_ARK_ARC_1_1/temp1[190] ), .ZN(\MC_ARK_ARC_1_1/temp5[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_0_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .B(n451), .ZN(\MC_ARK_ARC_1_1/temp4[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_0_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_1/temp3[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_0_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[136] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_0_1  ( .A(\MC_ARK_ARC_1_1/buf_datainput[190] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[184] ), .ZN(
        \MC_ARK_ARC_1_1/temp1[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X4_0_0  ( .A(n519), .B(n508), .ZN(
        \MC_ARK_ARC_1_1/temp4[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X3_0_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[65] ), 
        .B(n2124), .ZN(\MC_ARK_ARC_1_1/temp3[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X2_0_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_1/buf_datainput[161] ), .ZN(
        \MC_ARK_ARC_1_1/temp2[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_1/X1_0_0  ( .A(\MC_ARK_ARC_1_1/buf_datainput[185] ), 
        .B(n515), .ZN(\MC_ARK_ARC_1_1/temp1[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_31_5  ( .A(\MC_ARK_ARC_1_2/temp5[0] ), .B(
        \MC_ARK_ARC_1_2/temp6[0] ), .ZN(\RI1[3][0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_31_5  ( .A(\MC_ARK_ARC_1_2/temp3[0] ), .B(
        \MC_ARK_ARC_1_2/temp4[0] ), .ZN(\MC_ARK_ARC_1_2/temp6[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_31_5  ( .A(\MC_ARK_ARC_1_2/temp1[0] ), .B(
        \MC_ARK_ARC_1_2/temp2[0] ), .ZN(\MC_ARK_ARC_1_2/temp5[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_31_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[36] ), 
        .B(n286), .ZN(\MC_ARK_ARC_1_2/temp4[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_31_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[66] ), .ZN(\MC_ARK_ARC_1_2/temp3[0] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_31_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[138] ), .ZN(\MC_ARK_ARC_1_2/temp2[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_31_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[186] ), .ZN(\MC_ARK_ARC_1_2/temp1[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_31_4  ( .A(\MC_ARK_ARC_1_2/temp5[1] ), .B(
        \MC_ARK_ARC_1_2/temp6[1] ), .ZN(\RI1[3][1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_31_4  ( .A(\MC_ARK_ARC_1_2/temp3[1] ), .B(
        \MC_ARK_ARC_1_2/temp4[1] ), .ZN(\MC_ARK_ARC_1_2/temp6[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_31_4  ( .A(\MC_ARK_ARC_1_2/temp1[1] ), .B(
        \MC_ARK_ARC_1_2/temp2[1] ), .ZN(\MC_ARK_ARC_1_2/temp5[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_31_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[37] ), 
        .B(n325), .ZN(\MC_ARK_ARC_1_2/temp4[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_31_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[67] ), .ZN(\MC_ARK_ARC_1_2/temp3[1] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_31_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[163] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[139] ), .ZN(\MC_ARK_ARC_1_2/temp2[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_31_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[1] ), 
        .B(\RI5[2][187] ), .ZN(\MC_ARK_ARC_1_2/temp1[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_31_3  ( .A(\MC_ARK_ARC_1_2/temp6[2] ), .B(
        \MC_ARK_ARC_1_2/temp5[2] ), .ZN(\RI1[3][2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_31_3  ( .A(\MC_ARK_ARC_1_2/temp3[2] ), .B(
        \MC_ARK_ARC_1_2/temp4[2] ), .ZN(\MC_ARK_ARC_1_2/temp6[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_31_3  ( .A(\MC_ARK_ARC_1_2/temp1[2] ), .B(
        \MC_ARK_ARC_1_2/temp2[2] ), .ZN(\MC_ARK_ARC_1_2/temp5[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_31_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .B(n398), .ZN(\MC_ARK_ARC_1_2/temp4[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_31_3  ( .A(n2123), .B(
        \MC_ARK_ARC_1_2/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_2/temp3[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_31_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[164] ), .ZN(\MC_ARK_ARC_1_2/temp2[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_31_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[188] ), 
        .B(\RI5[2][2] ), .ZN(\MC_ARK_ARC_1_2/temp1[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_31_2  ( .A(\MC_ARK_ARC_1_2/temp5[3] ), .B(
        \MC_ARK_ARC_1_2/temp6[3] ), .ZN(\RI1[3][3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_31_2  ( .A(\MC_ARK_ARC_1_2/temp3[3] ), .B(
        \MC_ARK_ARC_1_2/temp4[3] ), .ZN(\MC_ARK_ARC_1_2/temp6[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_31_2  ( .A(\MC_ARK_ARC_1_2/temp1[3] ), .B(
        \MC_ARK_ARC_1_2/temp2[3] ), .ZN(\MC_ARK_ARC_1_2/temp5[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_31_2  ( .A(\RI5[2][39] ), .B(n221), .ZN(
        \MC_ARK_ARC_1_2/temp4[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_31_2  ( .A(\RI5[2][69] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[105] ), .ZN(\MC_ARK_ARC_1_2/temp3[3] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_31_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[165] ), 
        .B(n1951), .ZN(\MC_ARK_ARC_1_2/temp2[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_31_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[189] ), 
        .B(\RI5[2][3] ), .ZN(\MC_ARK_ARC_1_2/temp1[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_31_1  ( .A(\MC_ARK_ARC_1_2/temp5[4] ), .B(
        \MC_ARK_ARC_1_2/temp6[4] ), .ZN(\RI1[3][4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_31_1  ( .A(\MC_ARK_ARC_1_2/temp3[4] ), .B(
        \MC_ARK_ARC_1_2/temp4[4] ), .ZN(\MC_ARK_ARC_1_2/temp6[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_31_1  ( .A(\MC_ARK_ARC_1_2/temp1[4] ), .B(
        \MC_ARK_ARC_1_2/temp2[4] ), .ZN(\MC_ARK_ARC_1_2/temp5[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_31_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .B(n259), .ZN(\MC_ARK_ARC_1_2/temp4[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_31_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_2/temp3[4] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_31_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[166] ), .ZN(\MC_ARK_ARC_1_2/temp2[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_31_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[190] ), .ZN(\MC_ARK_ARC_1_2/temp1[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_31_0  ( .A(\MC_ARK_ARC_1_2/temp5[5] ), .B(
        \MC_ARK_ARC_1_2/temp6[5] ), .ZN(\RI1[3][5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_31_0  ( .A(\MC_ARK_ARC_1_2/temp3[5] ), .B(
        \MC_ARK_ARC_1_2/temp4[5] ), .ZN(\MC_ARK_ARC_1_2/temp6[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_31_0  ( .A(\MC_ARK_ARC_1_2/temp2[5] ), .B(
        \MC_ARK_ARC_1_2/temp1[5] ), .ZN(\MC_ARK_ARC_1_2/temp5[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_31_0  ( .A(n1502), .B(
        \MC_ARK_ARC_1_2/buf_datainput[107] ), .ZN(\MC_ARK_ARC_1_2/temp3[5] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_31_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .B(n1628), .ZN(\MC_ARK_ARC_1_2/temp2[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_31_0  ( .A(n1634), .B(n829), .ZN(
        \MC_ARK_ARC_1_2/temp1[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_30_5  ( .A(\MC_ARK_ARC_1_2/temp5[6] ), .B(
        \MC_ARK_ARC_1_2/temp6[6] ), .ZN(\RI1[3][6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_30_5  ( .A(\MC_ARK_ARC_1_2/temp3[6] ), .B(
        \MC_ARK_ARC_1_2/temp4[6] ), .ZN(\MC_ARK_ARC_1_2/temp6[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_30_5  ( .A(\MC_ARK_ARC_1_2/temp1[6] ), .B(
        \MC_ARK_ARC_1_2/temp2[6] ), .ZN(\MC_ARK_ARC_1_2/temp5[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_30_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[42] ), 
        .B(n472), .ZN(\MC_ARK_ARC_1_2/temp4[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_30_5  ( .A(\RI5[2][108] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[72] ), .ZN(\MC_ARK_ARC_1_2/temp3[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_30_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[144] ), .ZN(\MC_ARK_ARC_1_2/temp2[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_30_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_2/temp1[6] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_30_4  ( .A(\MC_ARK_ARC_1_2/temp5[7] ), .B(
        \MC_ARK_ARC_1_2/temp6[7] ), .ZN(\RI1[3][7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_30_4  ( .A(\MC_ARK_ARC_1_2/temp3[7] ), .B(
        \MC_ARK_ARC_1_2/temp4[7] ), .ZN(\MC_ARK_ARC_1_2/temp6[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_30_4  ( .A(\MC_ARK_ARC_1_2/temp1[7] ), .B(
        \MC_ARK_ARC_1_2/temp2[7] ), .ZN(\MC_ARK_ARC_1_2/temp5[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_30_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[43] ), 
        .B(n430), .ZN(\MC_ARK_ARC_1_2/temp4[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_30_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[73] ), .ZN(\MC_ARK_ARC_1_2/temp3[7] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_30_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[169] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[145] ), .ZN(\MC_ARK_ARC_1_2/temp2[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_30_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[1] ), .ZN(\MC_ARK_ARC_1_2/temp1[7] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_30_3  ( .A(\MC_ARK_ARC_1_2/temp5[8] ), .B(
        \MC_ARK_ARC_1_2/temp6[8] ), .ZN(\RI1[3][8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_30_3  ( .A(\MC_ARK_ARC_1_2/temp3[8] ), .B(
        \MC_ARK_ARC_1_2/temp4[8] ), .ZN(\MC_ARK_ARC_1_2/temp6[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_30_3  ( .A(\MC_ARK_ARC_1_2/temp2[8] ), .B(
        \MC_ARK_ARC_1_2/temp1[8] ), .ZN(\MC_ARK_ARC_1_2/temp5[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_30_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[44] ), 
        .B(n234), .ZN(\MC_ARK_ARC_1_2/temp4[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_30_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[74] ), .ZN(\MC_ARK_ARC_1_2/temp3[8] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_30_3  ( .A(n2144), .B(
        \MC_ARK_ARC_1_2/buf_datainput[146] ), .ZN(\MC_ARK_ARC_1_2/temp2[8] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_30_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[8] ), 
        .B(\RI5[2][2] ), .ZN(\MC_ARK_ARC_1_2/temp1[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_30_2  ( .A(\MC_ARK_ARC_1_2/temp5[9] ), .B(
        \MC_ARK_ARC_1_2/temp6[9] ), .ZN(\RI1[3][9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_30_2  ( .A(\MC_ARK_ARC_1_2/temp4[9] ), .B(
        \MC_ARK_ARC_1_2/temp3[9] ), .ZN(\MC_ARK_ARC_1_2/temp6[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_30_2  ( .A(\MC_ARK_ARC_1_2/temp1[9] ), .B(
        \MC_ARK_ARC_1_2/temp2[9] ), .ZN(\MC_ARK_ARC_1_2/temp5[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_30_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .B(n272), .ZN(\MC_ARK_ARC_1_2/temp4[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_30_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[75] ), 
        .B(n1950), .ZN(\MC_ARK_ARC_1_2/temp3[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_30_2  ( .A(n2140), .B(\RI5[2][171] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_30_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[9] ), 
        .B(\RI5[2][3] ), .ZN(\MC_ARK_ARC_1_2/temp1[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_30_1  ( .A(\MC_ARK_ARC_1_2/temp5[10] ), .B(
        \MC_ARK_ARC_1_2/temp6[10] ), .ZN(\RI1[3][10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_30_1  ( .A(\MC_ARK_ARC_1_2/temp3[10] ), .B(
        \MC_ARK_ARC_1_2/temp4[10] ), .ZN(\MC_ARK_ARC_1_2/temp6[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_30_1  ( .A(\MC_ARK_ARC_1_2/temp2[10] ), .B(
        \MC_ARK_ARC_1_2/temp1[10] ), .ZN(\MC_ARK_ARC_1_2/temp5[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_30_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[46] ), 
        .B(n443), .ZN(\MC_ARK_ARC_1_2/temp4[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_30_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[76] ), .ZN(\MC_ARK_ARC_1_2/temp3[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_30_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[148] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_30_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_2/temp1[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_30_0  ( .A(\MC_ARK_ARC_1_2/temp3[11] ), .B(
        \MC_ARK_ARC_1_2/temp4[11] ), .ZN(\MC_ARK_ARC_1_2/temp6[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_30_0  ( .A(\MC_ARK_ARC_1_2/temp1[11] ), .B(
        \MC_ARK_ARC_1_2/temp2[11] ), .ZN(\MC_ARK_ARC_1_2/temp5[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_30_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .B(n349), .ZN(\MC_ARK_ARC_1_2/temp4[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_30_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[77] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[113] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_30_0  ( .A(n827), .B(n816), .ZN(
        \MC_ARK_ARC_1_2/temp2[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_30_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[11] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[5] ), .ZN(\MC_ARK_ARC_1_2/temp1[11] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_29_5  ( .A(\MC_ARK_ARC_1_2/temp5[12] ), .B(
        \MC_ARK_ARC_1_2/temp6[12] ), .ZN(\RI1[3][12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_29_5  ( .A(\MC_ARK_ARC_1_2/temp3[12] ), .B(
        \MC_ARK_ARC_1_2/temp4[12] ), .ZN(\MC_ARK_ARC_1_2/temp6[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_29_5  ( .A(\MC_ARK_ARC_1_2/temp1[12] ), .B(
        \MC_ARK_ARC_1_2/temp2[12] ), .ZN(\MC_ARK_ARC_1_2/temp5[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_29_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[48] ), 
        .B(n206), .ZN(\MC_ARK_ARC_1_2/temp4[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_29_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[78] ), .ZN(\MC_ARK_ARC_1_2/temp3[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_29_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[174] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[150] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_29_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_2/temp1[12] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_29_4  ( .A(\MC_ARK_ARC_1_2/temp5[13] ), .B(
        \MC_ARK_ARC_1_2/temp6[13] ), .ZN(\RI1[3][13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_29_4  ( .A(\MC_ARK_ARC_1_2/temp3[13] ), .B(
        \MC_ARK_ARC_1_2/temp4[13] ), .ZN(\MC_ARK_ARC_1_2/temp6[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_29_4  ( .A(\MC_ARK_ARC_1_2/temp1[13] ), .B(
        \MC_ARK_ARC_1_2/temp2[13] ), .ZN(\MC_ARK_ARC_1_2/temp5[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_29_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .B(n245), .ZN(\MC_ARK_ARC_1_2/temp4[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_29_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[79] ), .ZN(\MC_ARK_ARC_1_2/temp3[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_29_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[151] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_29_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_2/temp1[13] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_29_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[50] ), 
        .B(n284), .ZN(\MC_ARK_ARC_1_2/temp4[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_29_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[80] ), .ZN(\MC_ARK_ARC_1_2/temp3[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_29_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_29_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_2/temp1[14] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_29_2  ( .A(\MC_ARK_ARC_1_2/temp3[15] ), .B(
        \MC_ARK_ARC_1_2/temp4[15] ), .ZN(\MC_ARK_ARC_1_2/temp6[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_29_2  ( .A(\RI5[2][51] ), .B(n323), .ZN(
        \MC_ARK_ARC_1_2/temp4[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_29_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[81] ), 
        .B(\RI5[2][117] ), .ZN(\MC_ARK_ARC_1_2/temp3[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_29_2  ( .A(\RI5[2][177] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[153] ), .ZN(\MC_ARK_ARC_1_2/temp2[15] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_29_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[9] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[15] ), .ZN(\MC_ARK_ARC_1_2/temp1[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_29_1  ( .A(\MC_ARK_ARC_1_2/temp5[16] ), .B(
        \MC_ARK_ARC_1_2/temp6[16] ), .ZN(\RI1[3][16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_29_1  ( .A(\MC_ARK_ARC_1_2/temp3[16] ), .B(
        \MC_ARK_ARC_1_2/temp4[16] ), .ZN(\MC_ARK_ARC_1_2/temp6[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_29_1  ( .A(\MC_ARK_ARC_1_2/temp2[16] ), .B(
        \MC_ARK_ARC_1_2/temp1[16] ), .ZN(\MC_ARK_ARC_1_2/temp5[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_29_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .B(n362), .ZN(\MC_ARK_ARC_1_2/temp4[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_29_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .B(n1957), .ZN(\MC_ARK_ARC_1_2/temp3[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_29_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[178] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_29_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_2/temp1[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_29_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[83] ), 
        .B(n812), .ZN(\MC_ARK_ARC_1_2/temp3[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_29_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[11] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[17] ), .ZN(\MC_ARK_ARC_1_2/temp1[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_28_5  ( .A(\MC_ARK_ARC_1_2/temp5[18] ), .B(
        \MC_ARK_ARC_1_2/temp6[18] ), .ZN(\RI1[3][18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_28_5  ( .A(\MC_ARK_ARC_1_2/temp3[18] ), .B(
        \MC_ARK_ARC_1_2/temp4[18] ), .ZN(\MC_ARK_ARC_1_2/temp6[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_28_5  ( .A(\MC_ARK_ARC_1_2/temp1[18] ), .B(
        \MC_ARK_ARC_1_2/temp2[18] ), .ZN(\MC_ARK_ARC_1_2/temp5[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_28_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[54] ), 
        .B(n492), .ZN(\MC_ARK_ARC_1_2/temp4[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_28_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[84] ), .ZN(\MC_ARK_ARC_1_2/temp3[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_28_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[180] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[156] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_28_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_2/temp1[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_28_4  ( .A(\MC_ARK_ARC_1_2/temp5[19] ), .B(
        \MC_ARK_ARC_1_2/temp6[19] ), .ZN(\RI1[3][19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_28_4  ( .A(\MC_ARK_ARC_1_2/temp3[19] ), .B(
        \MC_ARK_ARC_1_2/temp4[19] ), .ZN(\MC_ARK_ARC_1_2/temp6[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_28_4  ( .A(\MC_ARK_ARC_1_2/temp1[19] ), .B(
        \MC_ARK_ARC_1_2/temp2[19] ), .ZN(\MC_ARK_ARC_1_2/temp5[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_28_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[55] ), 
        .B(n297), .ZN(\MC_ARK_ARC_1_2/temp4[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_28_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[85] ), .ZN(\MC_ARK_ARC_1_2/temp3[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_28_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[157] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_28_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[13] ), .ZN(\MC_ARK_ARC_1_2/temp1[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_28_3  ( .A(\MC_ARK_ARC_1_2/temp1[20] ), .B(
        \MC_ARK_ARC_1_2/temp2[20] ), .ZN(\MC_ARK_ARC_1_2/temp5[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_28_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .B(n336), .ZN(\MC_ARK_ARC_1_2/temp4[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_28_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[122] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_28_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[158] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_28_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_2/temp1[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_28_2  ( .A(\MC_ARK_ARC_1_2/temp5[21] ), .B(
        \MC_ARK_ARC_1_2/temp6[21] ), .ZN(\RI1[3][21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_28_2  ( .A(\MC_ARK_ARC_1_2/temp3[21] ), .B(
        \MC_ARK_ARC_1_2/temp4[21] ), .ZN(\MC_ARK_ARC_1_2/temp6[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_28_2  ( .A(\MC_ARK_ARC_1_2/temp2[21] ), .B(
        \MC_ARK_ARC_1_2/temp1[21] ), .ZN(\MC_ARK_ARC_1_2/temp5[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_28_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[57] ), 
        .B(n374), .ZN(\MC_ARK_ARC_1_2/temp4[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_28_2  ( .A(\RI5[2][123] ), .B(\RI5[2][87] ), 
        .ZN(\MC_ARK_ARC_1_2/temp3[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_28_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[183] ), 
        .B(\RI5[2][159] ), .ZN(\MC_ARK_ARC_1_2/temp2[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_28_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[15] ), 
        .B(\RI5[2][21] ), .ZN(\MC_ARK_ARC_1_2/temp1[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_28_1  ( .A(\MC_ARK_ARC_1_2/temp6[22] ), .B(
        \MC_ARK_ARC_1_2/temp5[22] ), .ZN(\RI1[3][22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_28_1  ( .A(\MC_ARK_ARC_1_2/temp4[22] ), .B(
        \MC_ARK_ARC_1_2/temp3[22] ), .ZN(\MC_ARK_ARC_1_2/temp6[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_28_1  ( .A(\MC_ARK_ARC_1_2/temp2[22] ), .B(
        \MC_ARK_ARC_1_2/temp1[22] ), .ZN(\MC_ARK_ARC_1_2/temp5[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_28_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[58] ), 
        .B(n232), .ZN(\MC_ARK_ARC_1_2/temp4[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_28_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_2/temp3[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_28_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[184] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_28_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_2/temp1[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_28_0  ( .A(n792), .B(n501), .ZN(
        \MC_ARK_ARC_1_2/temp4[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_28_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .B(n1956), .ZN(\MC_ARK_ARC_1_2/temp3[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_28_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[161] ), 
        .B(n823), .ZN(\MC_ARK_ARC_1_2/temp2[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_28_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[17] ), 
        .B(n800), .ZN(\MC_ARK_ARC_1_2/temp1[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_27_5  ( .A(\MC_ARK_ARC_1_2/temp5[24] ), .B(
        \MC_ARK_ARC_1_2/temp6[24] ), .ZN(\RI1[3][24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_27_5  ( .A(\MC_ARK_ARC_1_2/temp3[24] ), .B(
        \MC_ARK_ARC_1_2/temp4[24] ), .ZN(\MC_ARK_ARC_1_2/temp6[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_27_5  ( .A(\MC_ARK_ARC_1_2/temp1[24] ), .B(
        \MC_ARK_ARC_1_2/temp2[24] ), .ZN(\MC_ARK_ARC_1_2/temp5[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_27_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[60] ), 
        .B(n309), .ZN(\MC_ARK_ARC_1_2/temp4[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_27_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[90] ), .ZN(\MC_ARK_ARC_1_2/temp3[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_27_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_27_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[18] ), .ZN(\MC_ARK_ARC_1_2/temp1[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_27_4  ( .A(\MC_ARK_ARC_1_2/temp5[25] ), .B(
        \MC_ARK_ARC_1_2/temp6[25] ), .ZN(\RI1[3][25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_27_4  ( .A(\MC_ARK_ARC_1_2/temp3[25] ), .B(
        \MC_ARK_ARC_1_2/temp4[25] ), .ZN(\MC_ARK_ARC_1_2/temp6[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_27_4  ( .A(\MC_ARK_ARC_1_2/temp1[25] ), .B(
        \MC_ARK_ARC_1_2/temp2[25] ), .ZN(\MC_ARK_ARC_1_2/temp5[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_27_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .B(n448), .ZN(\MC_ARK_ARC_1_2/temp4[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_27_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_2/temp3[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_27_4  ( .A(\RI5[2][187] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[163] ), .ZN(\MC_ARK_ARC_1_2/temp2[25] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_27_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[19] ), .ZN(\MC_ARK_ARC_1_2/temp1[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_27_3  ( .A(\MC_ARK_ARC_1_2/temp6[26] ), .B(
        \MC_ARK_ARC_1_2/temp5[26] ), .ZN(\RI1[3][26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_27_3  ( .A(\MC_ARK_ARC_1_2/temp3[26] ), .B(
        \MC_ARK_ARC_1_2/temp4[26] ), .ZN(\MC_ARK_ARC_1_2/temp6[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_27_3  ( .A(\MC_ARK_ARC_1_2/temp2[26] ), .B(
        \MC_ARK_ARC_1_2/temp1[26] ), .ZN(\MC_ARK_ARC_1_2/temp5[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_27_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[62] ), 
        .B(n401), .ZN(\MC_ARK_ARC_1_2/temp4[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_27_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_27_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[188] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_27_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_2/temp1[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_27_2  ( .A(\MC_ARK_ARC_1_2/temp5[27] ), .B(
        \MC_ARK_ARC_1_2/temp6[27] ), .ZN(\RI1[3][27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_27_2  ( .A(\MC_ARK_ARC_1_2/temp4[27] ), .B(
        \MC_ARK_ARC_1_2/temp3[27] ), .ZN(\MC_ARK_ARC_1_2/temp6[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_27_2  ( .A(\MC_ARK_ARC_1_2/temp1[27] ), .B(
        \MC_ARK_ARC_1_2/temp2[27] ), .ZN(\MC_ARK_ARC_1_2/temp5[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_27_2  ( .A(n2101), .B(n244), .ZN(
        \MC_ARK_ARC_1_2/temp4[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_27_2  ( .A(\RI5[2][93] ), .B(n815), .ZN(
        \MC_ARK_ARC_1_2/temp3[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_27_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[165] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[189] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_27_2  ( .A(\RI5[2][21] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[27] ), .ZN(\MC_ARK_ARC_1_2/temp1[27] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_27_1  ( .A(\MC_ARK_ARC_1_2/temp5[28] ), .B(
        \MC_ARK_ARC_1_2/temp6[28] ), .ZN(\RI1[3][28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_27_1  ( .A(\MC_ARK_ARC_1_2/temp3[28] ), .B(
        \MC_ARK_ARC_1_2/temp4[28] ), .ZN(\MC_ARK_ARC_1_2/temp6[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_27_1  ( .A(\MC_ARK_ARC_1_2/temp1[28] ), .B(
        \MC_ARK_ARC_1_2/temp2[28] ), .ZN(\MC_ARK_ARC_1_2/temp5[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_27_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[64] ), 
        .B(n457), .ZN(\MC_ARK_ARC_1_2/temp4[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_27_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_27_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[190] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_27_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .B(n2142), .ZN(\MC_ARK_ARC_1_2/temp1[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_27_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .B(n437), .ZN(\MC_ARK_ARC_1_2/temp4[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_27_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[131] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_27_0  ( .A(n1629), .B(n830), .ZN(
        \MC_ARK_ARC_1_2/temp2[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_27_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[23] ), .ZN(\MC_ARK_ARC_1_2/temp1[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_26_5  ( .A(\MC_ARK_ARC_1_2/temp5[30] ), .B(
        \MC_ARK_ARC_1_2/temp6[30] ), .ZN(\RI1[3][30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_26_5  ( .A(\MC_ARK_ARC_1_2/temp3[30] ), .B(
        \MC_ARK_ARC_1_2/temp4[30] ), .ZN(\MC_ARK_ARC_1_2/temp6[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_26_5  ( .A(\MC_ARK_ARC_1_2/temp1[30] ), .B(
        \MC_ARK_ARC_1_2/temp2[30] ), .ZN(\MC_ARK_ARC_1_2/temp5[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_26_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[66] ), 
        .B(n506), .ZN(\MC_ARK_ARC_1_2/temp4[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_26_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[132] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[96] ), .ZN(\MC_ARK_ARC_1_2/temp3[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_26_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_26_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[24] ), .ZN(\MC_ARK_ARC_1_2/temp1[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_26_4  ( .A(\MC_ARK_ARC_1_2/temp5[31] ), .B(
        \MC_ARK_ARC_1_2/temp6[31] ), .ZN(\RI1[3][31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_26_4  ( .A(\MC_ARK_ARC_1_2/temp3[31] ), .B(
        \MC_ARK_ARC_1_2/temp4[31] ), .ZN(\MC_ARK_ARC_1_2/temp6[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_26_4  ( .A(\MC_ARK_ARC_1_2/temp1[31] ), .B(
        \MC_ARK_ARC_1_2/temp2[31] ), .ZN(\MC_ARK_ARC_1_2/temp5[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_26_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[67] ), 
        .B(n217), .ZN(\MC_ARK_ARC_1_2/temp4[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_26_4  ( .A(\RI5[2][133] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[97] ), .ZN(\MC_ARK_ARC_1_2/temp3[31] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_26_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[1] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[169] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_26_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[25] ), .ZN(\MC_ARK_ARC_1_2/temp1[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_26_3  ( .A(\MC_ARK_ARC_1_2/temp5[32] ), .B(
        \MC_ARK_ARC_1_2/temp6[32] ), .ZN(\RI1[3][32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_26_3  ( .A(\MC_ARK_ARC_1_2/temp3[32] ), .B(
        \MC_ARK_ARC_1_2/temp4[32] ), .ZN(\MC_ARK_ARC_1_2/temp6[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_26_3  ( .A(\MC_ARK_ARC_1_2/temp2[32] ), .B(
        \MC_ARK_ARC_1_2/temp1[32] ), .ZN(\MC_ARK_ARC_1_2/temp5[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_26_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .B(n255), .ZN(\MC_ARK_ARC_1_2/temp4[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_26_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[98] ), .ZN(\MC_ARK_ARC_1_2/temp3[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_26_3  ( .A(n2144), .B(\RI5[2][2] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_26_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[26] ), 
        .B(n1511), .ZN(\MC_ARK_ARC_1_2/temp1[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_26_2  ( .A(\MC_ARK_ARC_1_2/temp6[33] ), .B(
        \MC_ARK_ARC_1_2/temp5[33] ), .ZN(\RI1[3][33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_26_2  ( .A(\MC_ARK_ARC_1_2/temp3[33] ), .B(
        \MC_ARK_ARC_1_2/temp4[33] ), .ZN(\MC_ARK_ARC_1_2/temp6[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_26_2  ( .A(\MC_ARK_ARC_1_2/temp1[33] ), .B(
        \MC_ARK_ARC_1_2/temp2[33] ), .ZN(\MC_ARK_ARC_1_2/temp5[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_26_2  ( .A(\RI5[2][69] ), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[33] ), .ZN(\MC_ARK_ARC_1_2/temp4[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_26_2  ( .A(n2098), .B(\RI5[2][99] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_26_2  ( .A(\RI5[2][3] ), .B(\RI5[2][171] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_26_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[27] ), .ZN(\MC_ARK_ARC_1_2/temp1[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_26_1  ( .A(\MC_ARK_ARC_1_2/temp5[34] ), .B(
        \MC_ARK_ARC_1_2/temp6[34] ), .ZN(\RI1[3][34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_26_1  ( .A(\MC_ARK_ARC_1_2/temp3[34] ), .B(
        \MC_ARK_ARC_1_2/temp4[34] ), .ZN(\MC_ARK_ARC_1_2/temp6[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_26_1  ( .A(\MC_ARK_ARC_1_2/temp2[34] ), .B(
        \MC_ARK_ARC_1_2/temp1[34] ), .ZN(\MC_ARK_ARC_1_2/temp5[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_26_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .B(n384), .ZN(\MC_ARK_ARC_1_2/temp4[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_26_1  ( .A(n1933), .B(
        \MC_ARK_ARC_1_2/buf_datainput[100] ), .ZN(\MC_ARK_ARC_1_2/temp3[34] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_26_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_2/temp2[34] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_26_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .B(n2142), .ZN(\MC_ARK_ARC_1_2/temp1[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_26_0  ( .A(\MC_ARK_ARC_1_2/temp3[35] ), .B(
        \MC_ARK_ARC_1_2/temp4[35] ), .ZN(\MC_ARK_ARC_1_2/temp6[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_26_0  ( .A(\MC_ARK_ARC_1_2/temp1[35] ), .B(
        \MC_ARK_ARC_1_2/temp2[35] ), .ZN(\MC_ARK_ARC_1_2/temp5[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_26_0  ( .A(n1502), .B(n372), .ZN(
        \MC_ARK_ARC_1_2/temp4[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_26_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[101] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_26_0  ( .A(n1634), .B(n827), .ZN(
        \MC_ARK_ARC_1_2/temp2[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_26_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[35] ), .ZN(\MC_ARK_ARC_1_2/temp1[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_25_5  ( .A(\MC_ARK_ARC_1_2/temp5[36] ), .B(
        \MC_ARK_ARC_1_2/temp6[36] ), .ZN(\RI1[3][36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_25_5  ( .A(\MC_ARK_ARC_1_2/temp3[36] ), .B(
        \MC_ARK_ARC_1_2/temp4[36] ), .ZN(\MC_ARK_ARC_1_2/temp6[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_25_5  ( .A(\MC_ARK_ARC_1_2/temp1[36] ), .B(
        \MC_ARK_ARC_1_2/temp2[36] ), .ZN(\MC_ARK_ARC_1_2/temp5[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_25_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[72] ), 
        .B(n230), .ZN(\MC_ARK_ARC_1_2/temp4[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_25_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[138] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[102] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_25_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[174] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_25_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[30] ), .ZN(\MC_ARK_ARC_1_2/temp1[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_25_4  ( .A(\MC_ARK_ARC_1_2/temp5[37] ), .B(
        \MC_ARK_ARC_1_2/temp6[37] ), .ZN(\RI1[3][37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_25_4  ( .A(\MC_ARK_ARC_1_2/temp3[37] ), .B(
        \MC_ARK_ARC_1_2/temp4[37] ), .ZN(\MC_ARK_ARC_1_2/temp6[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_25_4  ( .A(\MC_ARK_ARC_1_2/temp1[37] ), .B(
        \MC_ARK_ARC_1_2/temp2[37] ), .ZN(\MC_ARK_ARC_1_2/temp5[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_25_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[73] ), 
        .B(n435), .ZN(\MC_ARK_ARC_1_2/temp4[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_25_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_25_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_25_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[37] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[31] ), .ZN(\MC_ARK_ARC_1_2/temp1[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_25_3  ( .A(\MC_ARK_ARC_1_2/temp5[38] ), .B(
        \MC_ARK_ARC_1_2/temp6[38] ), .ZN(\RI1[3][38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_25_3  ( .A(\MC_ARK_ARC_1_2/temp3[38] ), .B(
        \MC_ARK_ARC_1_2/temp4[38] ), .ZN(\MC_ARK_ARC_1_2/temp6[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_25_3  ( .A(\MC_ARK_ARC_1_2/temp2[38] ), .B(
        \MC_ARK_ARC_1_2/temp1[38] ), .ZN(\MC_ARK_ARC_1_2/temp5[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_25_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .B(n307), .ZN(\MC_ARK_ARC_1_2/temp4[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_25_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[140] ), 
        .B(n2123), .ZN(\MC_ARK_ARC_1_2/temp3[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_25_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[8] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_25_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .B(n1511), .ZN(\MC_ARK_ARC_1_2/temp1[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_25_2  ( .A(\MC_ARK_ARC_1_2/temp2[39] ), .B(
        \MC_ARK_ARC_1_2/temp1[39] ), .ZN(\MC_ARK_ARC_1_2/temp5[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_25_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[75] ), 
        .B(n345), .ZN(\MC_ARK_ARC_1_2/temp4[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_25_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .B(n1951), .ZN(\MC_ARK_ARC_1_2/temp3[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_25_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[9] ), 
        .B(\RI5[2][177] ), .ZN(\MC_ARK_ARC_1_2/temp2[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_25_2  ( .A(\RI5[2][39] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_2/temp1[39] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_25_1  ( .A(\MC_ARK_ARC_1_2/temp6[40] ), .B(
        \MC_ARK_ARC_1_2/temp5[40] ), .ZN(\RI1[3][40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_25_1  ( .A(\MC_ARK_ARC_1_2/temp3[40] ), .B(
        \MC_ARK_ARC_1_2/temp4[40] ), .ZN(\MC_ARK_ARC_1_2/temp6[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_25_1  ( .A(\MC_ARK_ARC_1_2/temp2[40] ), .B(
        \MC_ARK_ARC_1_2/temp1[40] ), .ZN(\MC_ARK_ARC_1_2/temp5[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_25_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[76] ), 
        .B(n202), .ZN(\MC_ARK_ARC_1_2/temp4[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_25_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[142] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_25_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[178] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_25_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[34] ), .ZN(\MC_ARK_ARC_1_2/temp1[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_25_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[77] ), 
        .B(n487), .ZN(\MC_ARK_ARC_1_2/temp4[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_25_0  ( .A(n1665), .B(
        \MC_ARK_ARC_1_2/buf_datainput[143] ), .ZN(\MC_ARK_ARC_1_2/temp3[41] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_25_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[11] ), 
        .B(n802), .ZN(\MC_ARK_ARC_1_2/temp2[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_25_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[41] ), .ZN(\MC_ARK_ARC_1_2/temp1[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_24_5  ( .A(\MC_ARK_ARC_1_2/temp6[42] ), .B(
        \MC_ARK_ARC_1_2/temp5[42] ), .ZN(\RI1[3][42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_24_5  ( .A(\MC_ARK_ARC_1_2/temp3[42] ), .B(
        \MC_ARK_ARC_1_2/temp4[42] ), .ZN(\MC_ARK_ARC_1_2/temp6[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_24_5  ( .A(\MC_ARK_ARC_1_2/temp1[42] ), .B(
        \MC_ARK_ARC_1_2/temp2[42] ), .ZN(\MC_ARK_ARC_1_2/temp5[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_24_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[78] ), 
        .B(n281), .ZN(\MC_ARK_ARC_1_2/temp4[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_24_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[144] ), 
        .B(\RI5[2][108] ), .ZN(\MC_ARK_ARC_1_2/temp3[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_24_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_24_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[36] ), .ZN(\MC_ARK_ARC_1_2/temp1[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_24_4  ( .A(\MC_ARK_ARC_1_2/temp5[43] ), .B(
        \MC_ARK_ARC_1_2/temp6[43] ), .ZN(\RI1[3][43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_24_4  ( .A(\MC_ARK_ARC_1_2/temp3[43] ), .B(
        \MC_ARK_ARC_1_2/temp4[43] ), .ZN(\MC_ARK_ARC_1_2/temp6[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_24_4  ( .A(\MC_ARK_ARC_1_2/temp2[43] ), .B(
        \MC_ARK_ARC_1_2/temp1[43] ), .ZN(\MC_ARK_ARC_1_2/temp5[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_24_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[79] ), 
        .B(n482), .ZN(\MC_ARK_ARC_1_2/temp4[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_24_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_24_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_24_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[37] ), .ZN(\MC_ARK_ARC_1_2/temp1[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_24_3  ( .A(\MC_ARK_ARC_1_2/temp3[44] ), .B(
        \MC_ARK_ARC_1_2/temp4[44] ), .ZN(\MC_ARK_ARC_1_2/temp6[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_24_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[80] ), 
        .B(n358), .ZN(\MC_ARK_ARC_1_2/temp4[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_24_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[110] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_24_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_24_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[44] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_2/temp1[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_24_2  ( .A(\MC_ARK_ARC_1_2/temp5[45] ), .B(
        \MC_ARK_ARC_1_2/temp6[45] ), .ZN(\RI1[3][45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_24_2  ( .A(\MC_ARK_ARC_1_2/temp4[45] ), .B(
        \MC_ARK_ARC_1_2/temp3[45] ), .ZN(\MC_ARK_ARC_1_2/temp6[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_24_2  ( .A(\MC_ARK_ARC_1_2/temp1[45] ), .B(
        \MC_ARK_ARC_1_2/temp2[45] ), .ZN(\MC_ARK_ARC_1_2/temp5[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_24_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[81] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[45] ), .ZN(\MC_ARK_ARC_1_2/temp4[45] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_24_2  ( .A(n2139), .B(n1950), .ZN(
        \MC_ARK_ARC_1_2/temp3[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_24_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[15] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[183] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_24_2  ( .A(\RI5[2][39] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[45] ), .ZN(\MC_ARK_ARC_1_2/temp1[45] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_24_1  ( .A(\MC_ARK_ARC_1_2/temp5[46] ), .B(
        \MC_ARK_ARC_1_2/temp6[46] ), .ZN(\RI1[3][46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_24_1  ( .A(\MC_ARK_ARC_1_2/temp3[46] ), .B(
        \MC_ARK_ARC_1_2/temp4[46] ), .ZN(\MC_ARK_ARC_1_2/temp6[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_24_1  ( .A(\MC_ARK_ARC_1_2/temp2[46] ), .B(
        \MC_ARK_ARC_1_2/temp1[46] ), .ZN(\MC_ARK_ARC_1_2/temp5[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_24_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .B(n253), .ZN(\MC_ARK_ARC_1_2/temp4[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_24_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[148] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_24_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[184] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_2/temp2[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_24_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[46] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[40] ), .ZN(\MC_ARK_ARC_1_2/temp1[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_24_0  ( .A(\MC_ARK_ARC_1_2/temp3[47] ), .B(
        \MC_ARK_ARC_1_2/temp4[47] ), .ZN(\MC_ARK_ARC_1_2/temp6[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_24_0  ( .A(\MC_ARK_ARC_1_2/temp1[47] ), .B(
        \MC_ARK_ARC_1_2/temp2[47] ), .ZN(\MC_ARK_ARC_1_2/temp5[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_24_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[83] ), 
        .B(n293), .ZN(\MC_ARK_ARC_1_2/temp4[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_24_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[113] ), 
        .B(n817), .ZN(\MC_ARK_ARC_1_2/temp3[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_24_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[17] ), 
        .B(n822), .ZN(\MC_ARK_ARC_1_2/temp2[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_24_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .B(n846), .ZN(\MC_ARK_ARC_1_2/temp1[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_23_5  ( .A(\MC_ARK_ARC_1_2/temp5[48] ), .B(
        \MC_ARK_ARC_1_2/temp6[48] ), .ZN(\RI1[3][48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_23_5  ( .A(\MC_ARK_ARC_1_2/temp3[48] ), .B(
        \MC_ARK_ARC_1_2/temp4[48] ), .ZN(\MC_ARK_ARC_1_2/temp6[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_23_5  ( .A(\MC_ARK_ARC_1_2/temp1[48] ), .B(
        \MC_ARK_ARC_1_2/temp2[48] ), .ZN(\MC_ARK_ARC_1_2/temp5[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_23_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .B(n453), .ZN(\MC_ARK_ARC_1_2/temp4[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_23_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[150] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[114] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_23_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[186] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_23_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_2/temp1[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_23_4  ( .A(\MC_ARK_ARC_1_2/temp5[49] ), .B(
        \MC_ARK_ARC_1_2/temp6[49] ), .ZN(\RI1[3][49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_23_4  ( .A(\MC_ARK_ARC_1_2/temp3[49] ), .B(
        \MC_ARK_ARC_1_2/temp4[49] ), .ZN(\MC_ARK_ARC_1_2/temp6[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_23_4  ( .A(\MC_ARK_ARC_1_2/temp1[49] ), .B(
        \MC_ARK_ARC_1_2/temp2[49] ), .ZN(\MC_ARK_ARC_1_2/temp5[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_23_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[85] ), 
        .B(n370), .ZN(\MC_ARK_ARC_1_2/temp4[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_23_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_23_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[19] ), 
        .B(\RI5[2][187] ), .ZN(\MC_ARK_ARC_1_2/temp2[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_23_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[43] ), .ZN(\MC_ARK_ARC_1_2/temp1[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_23_3  ( .A(\MC_ARK_ARC_1_2/temp1[50] ), .B(
        \MC_ARK_ARC_1_2/temp2[50] ), .ZN(\MC_ARK_ARC_1_2/temp5[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_23_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[86] ), 
        .B(n228), .ZN(\MC_ARK_ARC_1_2/temp4[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_23_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_23_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[188] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_23_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[44] ), .ZN(\MC_ARK_ARC_1_2/temp1[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_23_2  ( .A(\MC_ARK_ARC_1_2/temp5[51] ), .B(
        \MC_ARK_ARC_1_2/temp6[51] ), .ZN(\RI1[3][51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_23_2  ( .A(\MC_ARK_ARC_1_2/temp3[51] ), .B(
        \MC_ARK_ARC_1_2/temp4[51] ), .ZN(\MC_ARK_ARC_1_2/temp6[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_23_2  ( .A(\MC_ARK_ARC_1_2/temp1[51] ), .B(
        \MC_ARK_ARC_1_2/temp2[51] ), .ZN(\MC_ARK_ARC_1_2/temp5[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_23_2  ( .A(\RI5[2][87] ), .B(
        \MC_ARK_ARC_1_1/buf_keyinput[170] ), .ZN(\MC_ARK_ARC_1_2/temp4[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_23_2  ( .A(\RI5[2][117] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[153] ), .ZN(\MC_ARK_ARC_1_2/temp3[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_23_2  ( .A(\RI5[2][21] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[189] ), .ZN(\MC_ARK_ARC_1_2/temp2[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_23_2  ( .A(\RI5[2][51] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[45] ), .ZN(\MC_ARK_ARC_1_2/temp1[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_23_1  ( .A(\MC_ARK_ARC_1_2/temp6[52] ), .B(
        \MC_ARK_ARC_1_2/temp5[52] ), .ZN(\RI1[3][52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_23_1  ( .A(\MC_ARK_ARC_1_2/temp3[52] ), .B(
        \MC_ARK_ARC_1_2/temp4[52] ), .ZN(\MC_ARK_ARC_1_2/temp6[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_23_1  ( .A(\MC_ARK_ARC_1_2/temp1[52] ), .B(
        \MC_ARK_ARC_1_2/temp2[52] ), .ZN(\MC_ARK_ARC_1_2/temp5[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_23_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[88] ), 
        .B(n305), .ZN(\MC_ARK_ARC_1_2/temp4[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_23_1  ( .A(n1957), .B(
        \MC_ARK_ARC_1_2/buf_datainput[154] ), .ZN(\MC_ARK_ARC_1_2/temp3[52] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_23_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[190] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[22] ), .ZN(\MC_ARK_ARC_1_2/temp2[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_23_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[46] ), .ZN(\MC_ARK_ARC_1_2/temp1[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_23_0  ( .A(\MC_ARK_ARC_1_2/temp3[53] ), .B(
        \MC_ARK_ARC_1_2/temp4[53] ), .ZN(\MC_ARK_ARC_1_2/temp6[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_23_0  ( .A(\MC_ARK_ARC_1_2/temp1[53] ), .B(
        \MC_ARK_ARC_1_2/temp2[53] ), .ZN(\MC_ARK_ARC_1_2/temp5[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_23_0  ( .A(n1501), .B(n460), .ZN(
        \MC_ARK_ARC_1_2/temp4[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_23_0  ( .A(n812), .B(n824), .ZN(
        \MC_ARK_ARC_1_2/temp3[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_23_0  ( .A(n800), .B(n830), .ZN(
        \MC_ARK_ARC_1_2/temp2[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_23_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .B(n782), .ZN(\MC_ARK_ARC_1_2/temp1[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_22_5  ( .A(\MC_ARK_ARC_1_2/temp5[54] ), .B(
        \MC_ARK_ARC_1_2/temp6[54] ), .ZN(\RI1[3][54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_22_5  ( .A(\MC_ARK_ARC_1_2/temp3[54] ), .B(
        \MC_ARK_ARC_1_2/temp4[54] ), .ZN(\MC_ARK_ARC_1_2/temp6[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_22_5  ( .A(\MC_ARK_ARC_1_2/temp1[54] ), .B(
        \MC_ARK_ARC_1_2/temp2[54] ), .ZN(\MC_ARK_ARC_1_2/temp5[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_22_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[90] ), 
        .B(n508), .ZN(\MC_ARK_ARC_1_2/temp4[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_22_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_22_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_2/temp2[54] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_22_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[48] ), .ZN(\MC_ARK_ARC_1_2/temp1[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_22_4  ( .A(\MC_ARK_ARC_1_2/temp5[55] ), .B(
        \MC_ARK_ARC_1_2/temp6[55] ), .ZN(\RI1[3][55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_22_4  ( .A(\MC_ARK_ARC_1_2/temp3[55] ), .B(
        \MC_ARK_ARC_1_2/temp4[55] ), .ZN(\MC_ARK_ARC_1_2/temp6[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_22_4  ( .A(\MC_ARK_ARC_1_2/temp1[55] ), .B(
        \MC_ARK_ARC_1_2/temp2[55] ), .ZN(\MC_ARK_ARC_1_2/temp5[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_22_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[91] ), 
        .B(n461), .ZN(\MC_ARK_ARC_1_2/temp4[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_22_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[157] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_22_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[1] ), .ZN(\MC_ARK_ARC_1_2/temp2[55] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_22_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[49] ), .ZN(\MC_ARK_ARC_1_2/temp1[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_22_3  ( .A(\MC_ARK_ARC_1_2/temp1[56] ), .B(
        \MC_ARK_ARC_1_2/temp2[56] ), .ZN(\MC_ARK_ARC_1_2/temp5[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_22_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[92] ), 
        .B(n494), .ZN(\MC_ARK_ARC_1_2/temp4[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_22_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[158] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_22_3  ( .A(\RI5[2][2] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_2/temp2[56] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_22_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[56] ), .ZN(\MC_ARK_ARC_1_2/temp1[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_22_2  ( .A(\MC_ARK_ARC_1_2/temp5[57] ), .B(
        \MC_ARK_ARC_1_2/temp6[57] ), .ZN(\RI1[3][57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_22_2  ( .A(\MC_ARK_ARC_1_2/temp3[57] ), .B(
        \MC_ARK_ARC_1_2/temp4[57] ), .ZN(\MC_ARK_ARC_1_2/temp6[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_22_2  ( .A(\MC_ARK_ARC_1_2/temp2[57] ), .B(
        \MC_ARK_ARC_1_2/temp1[57] ), .ZN(\MC_ARK_ARC_1_2/temp5[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_22_2  ( .A(\RI5[2][93] ), .B(n318), .ZN(
        \MC_ARK_ARC_1_2/temp4[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_22_2  ( .A(\RI5[2][123] ), .B(\RI5[2][159] ), 
        .ZN(\MC_ARK_ARC_1_2/temp3[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_22_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[27] ), 
        .B(\RI5[2][3] ), .ZN(\MC_ARK_ARC_1_2/temp2[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_22_2  ( .A(\RI5[2][51] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[57] ), .ZN(\MC_ARK_ARC_1_2/temp1[57] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_22_1  ( .A(\MC_ARK_ARC_1_2/temp5[58] ), .B(
        \MC_ARK_ARC_1_2/temp6[58] ), .ZN(\RI1[3][58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_22_1  ( .A(\MC_ARK_ARC_1_2/temp3[58] ), .B(
        \MC_ARK_ARC_1_2/temp4[58] ), .ZN(\MC_ARK_ARC_1_2/temp6[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_22_1  ( .A(\MC_ARK_ARC_1_2/temp1[58] ), .B(
        \MC_ARK_ARC_1_2/temp2[58] ), .ZN(\MC_ARK_ARC_1_2/temp5[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_22_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[27] ), .ZN(\MC_ARK_ARC_1_2/temp4[58] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_22_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_22_1  ( .A(n2142), .B(
        \MC_ARK_ARC_1_2/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_2/temp2[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_22_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[58] ), .ZN(\MC_ARK_ARC_1_2/temp1[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_22_0  ( .A(\MC_ARK_ARC_1_2/temp2[59] ), .B(
        \MC_ARK_ARC_1_2/temp1[59] ), .ZN(\MC_ARK_ARC_1_2/temp5[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_22_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .B(n481), .ZN(\MC_ARK_ARC_1_2/temp4[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_22_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .B(n1636), .ZN(\MC_ARK_ARC_1_2/temp3[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_22_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .B(n1633), .ZN(\MC_ARK_ARC_1_2/temp2[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_22_0  ( .A(n781), .B(n793), .ZN(
        \MC_ARK_ARC_1_2/temp1[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_21_5  ( .A(\MC_ARK_ARC_1_2/temp5[60] ), .B(
        \MC_ARK_ARC_1_2/temp6[60] ), .ZN(\RI1[3][60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_21_5  ( .A(\MC_ARK_ARC_1_2/temp3[60] ), .B(
        \MC_ARK_ARC_1_2/temp4[60] ), .ZN(\MC_ARK_ARC_1_2/temp6[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_21_5  ( .A(\MC_ARK_ARC_1_2/temp1[60] ), .B(
        \MC_ARK_ARC_1_2/temp2[60] ), .ZN(\MC_ARK_ARC_1_2/temp5[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_21_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[96] ), 
        .B(n251), .ZN(\MC_ARK_ARC_1_2/temp4[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_21_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[126] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_21_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_2/temp2[60] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_21_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[60] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[54] ), .ZN(\MC_ARK_ARC_1_2/temp1[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_21_4  ( .A(\MC_ARK_ARC_1_2/temp5[61] ), .B(
        \MC_ARK_ARC_1_2/temp6[61] ), .ZN(\RI1[3][61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_21_4  ( .A(\MC_ARK_ARC_1_2/temp3[61] ), .B(
        \MC_ARK_ARC_1_2/temp4[61] ), .ZN(\MC_ARK_ARC_1_2/temp6[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_21_4  ( .A(\MC_ARK_ARC_1_2/temp2[61] ), .B(
        \MC_ARK_ARC_1_2/temp1[61] ), .ZN(\MC_ARK_ARC_1_2/temp5[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_21_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[97] ), 
        .B(n490), .ZN(\MC_ARK_ARC_1_2/temp4[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_21_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[163] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[127] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_21_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[31] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_2/temp2[61] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_21_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[55] ), .ZN(\MC_ARK_ARC_1_2/temp1[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_21_3  ( .A(\MC_ARK_ARC_1_2/temp1[62] ), .B(
        \MC_ARK_ARC_1_2/temp2[62] ), .ZN(\MC_ARK_ARC_1_2/temp5[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_21_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[98] ), 
        .B(n399), .ZN(\MC_ARK_ARC_1_2/temp4[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_21_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[164] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_21_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[8] ), 
        .B(n1511), .ZN(\MC_ARK_ARC_1_2/temp2[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_21_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[56] ), .ZN(\MC_ARK_ARC_1_2/temp1[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_21_2  ( .A(\MC_ARK_ARC_1_2/temp1[63] ), .B(
        \MC_ARK_ARC_1_2/temp2[63] ), .ZN(\MC_ARK_ARC_1_2/temp5[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_21_2  ( .A(\RI5[2][99] ), .B(n368), .ZN(
        \MC_ARK_ARC_1_2/temp4[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_21_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[165] ), 
        .B(n815), .ZN(\MC_ARK_ARC_1_2/temp3[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_21_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_2/temp2[63] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_21_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[57] ), 
        .B(n2101), .ZN(\MC_ARK_ARC_1_2/temp1[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_21_1  ( .A(\MC_ARK_ARC_1_2/temp5[64] ), .B(
        \MC_ARK_ARC_1_2/temp6[64] ), .ZN(\RI1[3][64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_21_1  ( .A(\MC_ARK_ARC_1_2/temp3[64] ), .B(
        \MC_ARK_ARC_1_2/temp4[64] ), .ZN(\MC_ARK_ARC_1_2/temp6[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_21_1  ( .A(\MC_ARK_ARC_1_2/temp2[64] ), .B(
        \MC_ARK_ARC_1_2/temp1[64] ), .ZN(\MC_ARK_ARC_1_2/temp5[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_21_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[100] ), 
        .B(n226), .ZN(\MC_ARK_ARC_1_2/temp4[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_21_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_21_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_2/temp2[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_21_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[58] ), .ZN(\MC_ARK_ARC_1_2/temp1[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_21_0  ( .A(\MC_ARK_ARC_1_2/temp3[65] ), .B(
        \MC_ARK_ARC_1_2/temp4[65] ), .ZN(\MC_ARK_ARC_1_2/temp6[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_21_0  ( .A(\MC_ARK_ARC_1_2/temp2[65] ), .B(
        \MC_ARK_ARC_1_2/temp1[65] ), .ZN(\MC_ARK_ARC_1_2/temp5[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_21_0  ( .A(n2126), .B(n264), .ZN(
        \MC_ARK_ARC_1_2/temp4[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_21_0  ( .A(n1628), .B(
        \MC_ARK_ARC_1_2/buf_datainput[131] ), .ZN(\MC_ARK_ARC_1_2/temp3[65] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_21_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[11] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[35] ), .ZN(\MC_ARK_ARC_1_2/temp2[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_21_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .B(n792), .ZN(\MC_ARK_ARC_1_2/temp1[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_20_5  ( .A(\MC_ARK_ARC_1_2/temp5[66] ), .B(
        \MC_ARK_ARC_1_2/temp6[66] ), .ZN(\RI1[3][66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_20_5  ( .A(\MC_ARK_ARC_1_2/temp3[66] ), .B(
        \MC_ARK_ARC_1_2/temp4[66] ), .ZN(\MC_ARK_ARC_1_2/temp6[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_20_5  ( .A(\MC_ARK_ARC_1_2/temp1[66] ), .B(
        \MC_ARK_ARC_1_2/temp2[66] ), .ZN(\MC_ARK_ARC_1_2/temp5[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_20_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[102] ), 
        .B(n303), .ZN(\MC_ARK_ARC_1_2/temp4[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_20_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[132] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_20_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_2/temp2[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_20_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[60] ), .ZN(\MC_ARK_ARC_1_2/temp1[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_20_4  ( .A(\MC_ARK_ARC_1_2/temp5[67] ), .B(
        \MC_ARK_ARC_1_2/temp6[67] ), .ZN(\RI1[3][67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_20_4  ( .A(\MC_ARK_ARC_1_2/temp3[67] ), .B(
        \MC_ARK_ARC_1_2/temp4[67] ), .ZN(\MC_ARK_ARC_1_2/temp6[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_20_4  ( .A(\MC_ARK_ARC_1_2/temp1[67] ), .B(
        \MC_ARK_ARC_1_2/temp2[67] ), .ZN(\MC_ARK_ARC_1_2/temp5[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_20_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[103] ), 
        .B(n464), .ZN(\MC_ARK_ARC_1_2/temp4[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_20_4  ( .A(\RI5[2][133] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[169] ), .ZN(\MC_ARK_ARC_1_2/temp3[67] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_20_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[37] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[13] ), .ZN(\MC_ARK_ARC_1_2/temp2[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_20_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[61] ), .ZN(\MC_ARK_ARC_1_2/temp1[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_20_3  ( .A(\MC_ARK_ARC_1_2/temp5[68] ), .B(
        \MC_ARK_ARC_1_2/temp6[68] ), .ZN(\RI1[3][68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_20_3  ( .A(\MC_ARK_ARC_1_2/temp3[68] ), .B(
        \MC_ARK_ARC_1_2/temp4[68] ), .ZN(\MC_ARK_ARC_1_2/temp6[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_20_3  ( .A(\MC_ARK_ARC_1_2/temp2[68] ), .B(
        \MC_ARK_ARC_1_2/temp1[68] ), .ZN(\MC_ARK_ARC_1_2/temp5[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_20_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[104] ), 
        .B(n199), .ZN(\MC_ARK_ARC_1_2/temp4[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_20_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[134] ), 
        .B(\RI5[2][170] ), .ZN(\MC_ARK_ARC_1_2/temp3[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_20_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .B(\RI5[2][14] ), .ZN(\MC_ARK_ARC_1_2/temp2[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_20_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .B(\RI5[2][62] ), .ZN(\MC_ARK_ARC_1_2/temp1[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_20_2  ( .A(\MC_ARK_ARC_1_2/temp2[69] ), .B(
        \MC_ARK_ARC_1_2/temp1[69] ), .ZN(\MC_ARK_ARC_1_2/temp5[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_20_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[69] ), .ZN(\MC_ARK_ARC_1_2/temp4[69] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_20_2  ( .A(\RI5[2][171] ), .B(\RI5[2][135] ), 
        .ZN(\MC_ARK_ARC_1_2/temp3[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_20_2  ( .A(\RI5[2][39] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[15] ), .ZN(\MC_ARK_ARC_1_2/temp2[69] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_20_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .B(\RI5[2][69] ), .ZN(\MC_ARK_ARC_1_2/temp1[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_20_1  ( .A(\MC_ARK_ARC_1_2/temp5[70] ), .B(
        \MC_ARK_ARC_1_2/temp6[70] ), .ZN(\RI1[3][70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_20_1  ( .A(\MC_ARK_ARC_1_2/temp3[70] ), .B(
        \MC_ARK_ARC_1_2/temp4[70] ), .ZN(\MC_ARK_ARC_1_2/temp6[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_20_1  ( .A(\MC_ARK_ARC_1_2/temp1[70] ), .B(
        \MC_ARK_ARC_1_2/temp2[70] ), .ZN(\MC_ARK_ARC_1_2/temp5[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_20_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .B(n378), .ZN(\MC_ARK_ARC_1_2/temp4[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_20_1  ( .A(n1933), .B(\RI5[2][172] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_20_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_2/temp2[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_20_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[64] ), .ZN(\MC_ARK_ARC_1_2/temp1[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_20_0  ( .A(\MC_ARK_ARC_1_2/temp2[71] ), .B(
        \MC_ARK_ARC_1_2/temp1[71] ), .ZN(\MC_ARK_ARC_1_2/temp5[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_20_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[107] ), 
        .B(n500), .ZN(\MC_ARK_ARC_1_2/temp4[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_20_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[173] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_20_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[17] ), 
        .B(n846), .ZN(\MC_ARK_ARC_1_2/temp2[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_20_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .B(n1503), .ZN(\MC_ARK_ARC_1_2/temp1[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_19_5  ( .A(\MC_ARK_ARC_1_2/temp5[72] ), .B(
        \MC_ARK_ARC_1_2/temp6[72] ), .ZN(\RI1[3][72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_19_5  ( .A(\MC_ARK_ARC_1_2/temp3[72] ), .B(
        \MC_ARK_ARC_1_2/temp4[72] ), .ZN(\MC_ARK_ARC_1_2/temp6[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_19_5  ( .A(\MC_ARK_ARC_1_2/temp1[72] ), .B(
        \MC_ARK_ARC_1_2/temp2[72] ), .ZN(\MC_ARK_ARC_1_2/temp5[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_19_5  ( .A(\RI5[2][108] ), .B(n354), .ZN(
        \MC_ARK_ARC_1_2/temp4[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_19_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[174] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[138] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_19_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[18] ), .ZN(\MC_ARK_ARC_1_2/temp2[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_19_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[66] ), .ZN(\MC_ARK_ARC_1_2/temp1[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_19_4  ( .A(\MC_ARK_ARC_1_2/temp5[73] ), .B(
        \MC_ARK_ARC_1_2/temp6[73] ), .ZN(\RI1[3][73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_19_4  ( .A(\MC_ARK_ARC_1_2/temp3[73] ), .B(
        \MC_ARK_ARC_1_2/temp4[73] ), .ZN(\MC_ARK_ARC_1_2/temp6[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_19_4  ( .A(\MC_ARK_ARC_1_2/temp1[73] ), .B(
        \MC_ARK_ARC_1_2/temp2[73] ), .ZN(\MC_ARK_ARC_1_2/temp5[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_19_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[109] ), 
        .B(n470), .ZN(\MC_ARK_ARC_1_2/temp4[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_19_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[139] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_19_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[19] ), .ZN(\MC_ARK_ARC_1_2/temp2[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_19_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[67] ), .ZN(\MC_ARK_ARC_1_2/temp1[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_19_3  ( .A(\MC_ARK_ARC_1_2/temp5[74] ), .B(
        \MC_ARK_ARC_1_2/temp6[74] ), .ZN(\RI1[3][74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_19_3  ( .A(\MC_ARK_ARC_1_2/temp3[74] ), .B(
        \MC_ARK_ARC_1_2/temp4[74] ), .ZN(\MC_ARK_ARC_1_2/temp6[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_19_3  ( .A(\MC_ARK_ARC_1_2/temp1[74] ), .B(
        \MC_ARK_ARC_1_2/temp2[74] ), .ZN(\MC_ARK_ARC_1_2/temp5[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_19_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[110] ), 
        .B(n391), .ZN(\MC_ARK_ARC_1_2/temp4[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_19_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_19_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[44] ), .ZN(\MC_ARK_ARC_1_2/temp2[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_19_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[74] ), .ZN(\MC_ARK_ARC_1_2/temp1[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_19_2  ( .A(\MC_ARK_ARC_1_2/temp1[75] ), .B(
        \MC_ARK_ARC_1_2/temp2[75] ), .ZN(\MC_ARK_ARC_1_2/temp5[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_19_2  ( .A(n1950), .B(n289), .ZN(
        \MC_ARK_ARC_1_2/temp4[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_19_2  ( .A(\RI5[2][177] ), .B(n1951), .ZN(
        \MC_ARK_ARC_1_2/temp3[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_19_2  ( .A(\RI5[2][21] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[45] ), .ZN(\MC_ARK_ARC_1_2/temp2[75] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_19_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[75] ), 
        .B(\RI5[2][69] ), .ZN(\MC_ARK_ARC_1_2/temp1[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_19_1  ( .A(\MC_ARK_ARC_1_2/temp5[76] ), .B(
        \MC_ARK_ARC_1_2/temp6[76] ), .ZN(\RI1[3][76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_19_1  ( .A(\MC_ARK_ARC_1_2/temp3[76] ), .B(
        \MC_ARK_ARC_1_2/temp4[76] ), .ZN(\MC_ARK_ARC_1_2/temp6[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_19_1  ( .A(\MC_ARK_ARC_1_2/temp2[76] ), .B(
        \MC_ARK_ARC_1_2/temp1[76] ), .ZN(\MC_ARK_ARC_1_2/temp5[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_19_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[76] ), .ZN(\MC_ARK_ARC_1_2/temp4[76] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_19_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[178] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_19_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[46] ), .ZN(\MC_ARK_ARC_1_2/temp2[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_19_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[76] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_2/temp1[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_19_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[113] ), 
        .B(n499), .ZN(\MC_ARK_ARC_1_2/temp4[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_19_0  ( .A(n803), .B(
        \MC_ARK_ARC_1_2/buf_datainput[143] ), .ZN(\MC_ARK_ARC_1_2/temp3[77] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_19_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .B(n800), .ZN(\MC_ARK_ARC_1_2/temp2[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_19_0  ( .A(n1503), .B(
        \MC_ARK_ARC_1_2/buf_datainput[77] ), .ZN(\MC_ARK_ARC_1_2/temp1[77] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_18_5  ( .A(\MC_ARK_ARC_1_2/temp5[78] ), .B(
        \MC_ARK_ARC_1_2/temp6[78] ), .ZN(\RI1[3][78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_18_5  ( .A(\MC_ARK_ARC_1_2/temp3[78] ), .B(
        \MC_ARK_ARC_1_2/temp4[78] ), .ZN(\MC_ARK_ARC_1_2/temp6[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_18_5  ( .A(\MC_ARK_ARC_1_2/temp2[78] ), .B(
        \MC_ARK_ARC_1_2/temp1[78] ), .ZN(\MC_ARK_ARC_1_2/temp5[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_18_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[114] ), 
        .B(n511), .ZN(\MC_ARK_ARC_1_2/temp4[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_18_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[180] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[144] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_18_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[24] ), .ZN(\MC_ARK_ARC_1_2/temp2[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_18_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[72] ), .ZN(\MC_ARK_ARC_1_2/temp1[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_18_4  ( .A(\MC_ARK_ARC_1_2/temp5[79] ), .B(
        \MC_ARK_ARC_1_2/temp6[79] ), .ZN(\RI1[3][79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_18_4  ( .A(\MC_ARK_ARC_1_2/temp3[79] ), .B(
        \MC_ARK_ARC_1_2/temp4[79] ), .ZN(\MC_ARK_ARC_1_2/temp6[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_18_4  ( .A(\MC_ARK_ARC_1_2/temp1[79] ), .B(
        \MC_ARK_ARC_1_2/temp2[79] ), .ZN(\MC_ARK_ARC_1_2/temp5[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_18_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .B(n439), .ZN(\MC_ARK_ARC_1_2/temp4[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_18_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[145] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_18_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[25] ), .ZN(\MC_ARK_ARC_1_2/temp2[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_18_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[73] ), .ZN(\MC_ARK_ARC_1_2/temp1[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_18_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[116] ), 
        .B(n301), .ZN(\MC_ARK_ARC_1_2/temp4[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_18_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_18_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_2/temp2[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_18_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[80] ), .ZN(\MC_ARK_ARC_1_2/temp1[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_18_2  ( .A(\MC_ARK_ARC_1_2/temp3[81] ), .B(
        \MC_ARK_ARC_1_2/temp4[81] ), .ZN(\MC_ARK_ARC_1_2/temp6[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_18_2  ( .A(\RI5[2][117] ), .B(n340), .ZN(
        \MC_ARK_ARC_1_2/temp4[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_18_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[183] ), 
        .B(n2139), .ZN(\MC_ARK_ARC_1_2/temp3[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_18_2  ( .A(\RI5[2][51] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[27] ), .ZN(\MC_ARK_ARC_1_2/temp2[81] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_18_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[75] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[81] ), .ZN(\MC_ARK_ARC_1_2/temp1[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_18_1  ( .A(\MC_ARK_ARC_1_2/temp6[82] ), .B(
        \MC_ARK_ARC_1_2/temp5[82] ), .ZN(\RI1[3][82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_18_1  ( .A(\MC_ARK_ARC_1_2/temp3[82] ), .B(
        \MC_ARK_ARC_1_2/temp4[82] ), .ZN(\MC_ARK_ARC_1_2/temp6[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_18_1  ( .A(\MC_ARK_ARC_1_2/temp2[82] ), .B(
        \MC_ARK_ARC_1_2/temp1[82] ), .ZN(\MC_ARK_ARC_1_2/temp5[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_18_1  ( .A(n1957), .B(n197), .ZN(
        \MC_ARK_ARC_1_2/temp4[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_18_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[184] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_18_1  ( .A(n2142), .B(
        \MC_ARK_ARC_1_2/buf_datainput[52] ), .ZN(\MC_ARK_ARC_1_2/temp2[82] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_18_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[76] ), .ZN(\MC_ARK_ARC_1_2/temp1[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_18_0  ( .A(\MC_ARK_ARC_1_2/temp5[83] ), .B(
        \MC_ARK_ARC_1_2/temp6[83] ), .ZN(\RI1[3][83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_18_0  ( .A(\MC_ARK_ARC_1_2/temp3[83] ), .B(
        \MC_ARK_ARC_1_2/temp4[83] ), .ZN(\MC_ARK_ARC_1_2/temp6[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_18_0  ( .A(\MC_ARK_ARC_1_2/temp1[83] ), .B(
        \MC_ARK_ARC_1_2/temp2[83] ), .ZN(\MC_ARK_ARC_1_2/temp5[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_18_0  ( .A(n811), .B(n476), .ZN(
        \MC_ARK_ARC_1_2/temp4[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_18_0  ( .A(n822), .B(n817), .ZN(
        \MC_ARK_ARC_1_2/temp3[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_18_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[53] ), .ZN(\MC_ARK_ARC_1_2/temp2[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_18_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[77] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[83] ), .ZN(\MC_ARK_ARC_1_2/temp1[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_17_5  ( .A(\MC_ARK_ARC_1_2/temp5[84] ), .B(
        \MC_ARK_ARC_1_2/temp6[84] ), .ZN(\RI1[3][84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_17_5  ( .A(\MC_ARK_ARC_1_2/temp3[84] ), .B(
        \MC_ARK_ARC_1_2/temp4[84] ), .ZN(\MC_ARK_ARC_1_2/temp6[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_17_5  ( .A(\MC_ARK_ARC_1_2/temp1[84] ), .B(
        \MC_ARK_ARC_1_2/temp2[84] ), .ZN(\MC_ARK_ARC_1_2/temp5[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_17_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[120] ), 
        .B(n495), .ZN(\MC_ARK_ARC_1_2/temp4[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_17_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[150] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_17_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[30] ), .ZN(\MC_ARK_ARC_1_2/temp2[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_17_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[78] ), .ZN(\MC_ARK_ARC_1_2/temp1[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_17_4  ( .A(\MC_ARK_ARC_1_2/temp5[85] ), .B(
        \MC_ARK_ARC_1_2/temp6[85] ), .ZN(\RI1[3][85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_17_4  ( .A(\MC_ARK_ARC_1_2/temp3[85] ), .B(
        \MC_ARK_ARC_1_2/temp4[85] ), .ZN(\MC_ARK_ARC_1_2/temp6[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_17_4  ( .A(\MC_ARK_ARC_1_2/temp1[85] ), .B(
        \MC_ARK_ARC_1_2/temp2[85] ), .ZN(\MC_ARK_ARC_1_2/temp5[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_17_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .B(n455), .ZN(\MC_ARK_ARC_1_2/temp4[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_17_4  ( .A(\RI5[2][187] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[151] ), .ZN(\MC_ARK_ARC_1_2/temp3[85] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_17_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[31] ), .ZN(\MC_ARK_ARC_1_2/temp2[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_17_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[79] ), .ZN(\MC_ARK_ARC_1_2/temp1[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_17_3  ( .A(\MC_ARK_ARC_1_2/temp5[86] ), .B(
        \MC_ARK_ARC_1_2/temp6[86] ), .ZN(\RI1[3][86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_17_3  ( .A(\MC_ARK_ARC_1_2/temp3[86] ), .B(
        \MC_ARK_ARC_1_2/temp4[86] ), .ZN(\MC_ARK_ARC_1_2/temp6[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_17_3  ( .A(\MC_ARK_ARC_1_2/temp1[86] ), .B(
        \MC_ARK_ARC_1_2/temp2[86] ), .ZN(\MC_ARK_ARC_1_2/temp5[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_17_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[122] ), 
        .B(n352), .ZN(\MC_ARK_ARC_1_2/temp4[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_17_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[188] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_17_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .B(n1511), .ZN(\MC_ARK_ARC_1_2/temp2[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_17_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[80] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[86] ), .ZN(\MC_ARK_ARC_1_2/temp1[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_17_2  ( .A(\MC_ARK_ARC_1_2/temp5[87] ), .B(
        \MC_ARK_ARC_1_2/temp6[87] ), .ZN(\RI1[3][87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_17_2  ( .A(\MC_ARK_ARC_1_2/temp3[87] ), .B(
        \MC_ARK_ARC_1_2/temp4[87] ), .ZN(\MC_ARK_ARC_1_2/temp6[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_17_2  ( .A(\MC_ARK_ARC_1_2/temp1[87] ), .B(
        \MC_ARK_ARC_1_2/temp2[87] ), .ZN(\MC_ARK_ARC_1_2/temp5[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_17_2  ( .A(\RI5[2][123] ), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[87] ), .ZN(\MC_ARK_ARC_1_2/temp4[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_17_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[189] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[153] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_17_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[57] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_2/temp2[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_17_2  ( .A(\RI5[2][87] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[81] ), .ZN(\MC_ARK_ARC_1_2/temp1[87] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_17_1  ( .A(\MC_ARK_ARC_1_2/temp5[88] ), .B(
        \MC_ARK_ARC_1_2/temp6[88] ), .ZN(\RI1[3][88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_17_1  ( .A(\MC_ARK_ARC_1_2/temp3[88] ), .B(
        \MC_ARK_ARC_1_2/temp4[88] ), .ZN(\MC_ARK_ARC_1_2/temp6[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_17_1  ( .A(\MC_ARK_ARC_1_2/temp2[88] ), .B(
        \MC_ARK_ARC_1_2/temp1[88] ), .ZN(\MC_ARK_ARC_1_2/temp5[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_17_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .B(n248), .ZN(\MC_ARK_ARC_1_2/temp4[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_17_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[190] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_17_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[58] ), .ZN(\MC_ARK_ARC_1_2/temp2[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_17_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_2/temp1[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_17_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .B(n422), .ZN(\MC_ARK_ARC_1_2/temp4[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_17_0  ( .A(n824), .B(
        \MC_ARK_ARC_1_2/buf_datainput[191] ), .ZN(\MC_ARK_ARC_1_2/temp3[89] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_17_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .B(n793), .ZN(\MC_ARK_ARC_1_2/temp2[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_17_0  ( .A(n1501), .B(
        \MC_ARK_ARC_1_2/buf_datainput[83] ), .ZN(\MC_ARK_ARC_1_2/temp1[89] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_16_5  ( .A(\MC_ARK_ARC_1_2/temp5[90] ), .B(
        \MC_ARK_ARC_1_2/temp6[90] ), .ZN(\RI1[3][90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_16_5  ( .A(\MC_ARK_ARC_1_2/temp3[90] ), .B(
        \MC_ARK_ARC_1_2/temp4[90] ), .ZN(\MC_ARK_ARC_1_2/temp6[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_16_5  ( .A(\MC_ARK_ARC_1_2/temp1[90] ), .B(
        \MC_ARK_ARC_1_2/temp2[90] ), .ZN(\MC_ARK_ARC_1_2/temp5[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_16_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[126] ), 
        .B(n326), .ZN(\MC_ARK_ARC_1_2/temp4[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_16_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[156] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_16_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[60] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[36] ), .ZN(\MC_ARK_ARC_1_2/temp2[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_16_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[84] ), .ZN(\MC_ARK_ARC_1_2/temp1[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_16_4  ( .A(\MC_ARK_ARC_1_2/temp5[91] ), .B(
        \MC_ARK_ARC_1_2/temp6[91] ), .ZN(\RI1[3][91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_16_4  ( .A(\MC_ARK_ARC_1_2/temp4[91] ), .B(
        \MC_ARK_ARC_1_2/temp3[91] ), .ZN(\MC_ARK_ARC_1_2/temp6[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_16_4  ( .A(\MC_ARK_ARC_1_2/temp1[91] ), .B(
        \MC_ARK_ARC_1_2/temp2[91] ), .ZN(\MC_ARK_ARC_1_2/temp5[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_16_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[127] ), 
        .B(n456), .ZN(\MC_ARK_ARC_1_2/temp4[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_16_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[1] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[157] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_16_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[37] ), .ZN(\MC_ARK_ARC_1_2/temp2[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_16_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[85] ), .ZN(\MC_ARK_ARC_1_2/temp1[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_16_3  ( .A(\MC_ARK_ARC_1_2/temp2[92] ), .B(
        \MC_ARK_ARC_1_2/temp1[92] ), .ZN(\MC_ARK_ARC_1_2/temp5[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_16_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[128] ), 
        .B(n222), .ZN(\MC_ARK_ARC_1_2/temp4[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_16_3  ( .A(\RI5[2][2] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[158] ), .ZN(\MC_ARK_ARC_1_2/temp3[92] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_16_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_2/temp2[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_16_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[86] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[92] ), .ZN(\MC_ARK_ARC_1_2/temp1[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_16_2  ( .A(\MC_ARK_ARC_1_2/temp5[93] ), .B(
        \MC_ARK_ARC_1_2/temp6[93] ), .ZN(\RI1[3][93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_16_2  ( .A(\MC_ARK_ARC_1_2/temp3[93] ), .B(
        \MC_ARK_ARC_1_2/temp4[93] ), .ZN(\MC_ARK_ARC_1_2/temp6[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_16_2  ( .A(\MC_ARK_ARC_1_2/temp2[93] ), .B(
        \MC_ARK_ARC_1_2/temp1[93] ), .ZN(\MC_ARK_ARC_1_2/temp5[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_16_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[129] ), 
        .B(n260), .ZN(\MC_ARK_ARC_1_2/temp4[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_16_2  ( .A(\RI5[2][3] ), .B(\RI5[2][159] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_16_2  ( .A(\RI5[2][39] ), .B(n2101), .ZN(
        \MC_ARK_ARC_1_2/temp2[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_16_2  ( .A(\RI5[2][87] ), .B(\RI5[2][93] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_16_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[130] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[94] ), .ZN(\MC_ARK_ARC_1_2/temp4[94] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_16_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_16_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[40] ), .ZN(\MC_ARK_ARC_1_2/temp2[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_16_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_2/temp1[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_16_0  ( .A(\MC_ARK_ARC_1_2/temp3[95] ), .B(
        \MC_ARK_ARC_1_2/temp4[95] ), .ZN(\MC_ARK_ARC_1_2/temp6[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_16_0  ( .A(\MC_ARK_ARC_1_2/temp1[95] ), .B(
        \MC_ARK_ARC_1_2/temp2[95] ), .ZN(\MC_ARK_ARC_1_2/temp5[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_16_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .B(n338), .ZN(\MC_ARK_ARC_1_2/temp4[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_16_0  ( .A(n1633), .B(n1635), .ZN(
        \MC_ARK_ARC_1_2/temp3[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_16_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .B(n846), .ZN(\MC_ARK_ARC_1_2/temp2[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_16_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .B(n1956), .ZN(\MC_ARK_ARC_1_2/temp1[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_15_5  ( .A(\MC_ARK_ARC_1_2/temp6[96] ), .B(
        \MC_ARK_ARC_1_2/temp5[96] ), .ZN(\RI1[3][96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_15_5  ( .A(\MC_ARK_ARC_1_2/temp3[96] ), .B(
        \MC_ARK_ARC_1_2/temp4[96] ), .ZN(\MC_ARK_ARC_1_2/temp6[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_15_5  ( .A(\MC_ARK_ARC_1_2/temp1[96] ), .B(
        \MC_ARK_ARC_1_2/temp2[96] ), .ZN(\MC_ARK_ARC_1_2/temp5[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_15_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[132] ), 
        .B(n195), .ZN(\MC_ARK_ARC_1_2/temp4[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_15_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[6] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_15_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_2/temp2[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_15_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[90] ), .ZN(\MC_ARK_ARC_1_2/temp1[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_15_4  ( .A(\MC_ARK_ARC_1_2/temp6[97] ), .B(
        \MC_ARK_ARC_1_2/temp5[97] ), .ZN(\RI1[3][97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_15_4  ( .A(\MC_ARK_ARC_1_2/temp3[97] ), .B(
        \MC_ARK_ARC_1_2/temp4[97] ), .ZN(\MC_ARK_ARC_1_2/temp6[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_15_4  ( .A(\MC_ARK_ARC_1_2/temp1[97] ), .B(
        \MC_ARK_ARC_1_2/temp2[97] ), .ZN(\MC_ARK_ARC_1_2/temp5[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_15_4  ( .A(\RI5[2][133] ), .B(n491), .ZN(
        \MC_ARK_ARC_1_2/temp4[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_15_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[163] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_15_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[43] ), .ZN(\MC_ARK_ARC_1_2/temp2[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_15_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_2/temp1[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_15_3  ( .A(\MC_ARK_ARC_1_2/temp5[98] ), .B(
        \MC_ARK_ARC_1_2/temp6[98] ), .ZN(\RI1[3][98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_15_3  ( .A(\MC_ARK_ARC_1_2/temp3[98] ), .B(
        \MC_ARK_ARC_1_2/temp4[98] ), .ZN(\MC_ARK_ARC_1_2/temp6[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_15_3  ( .A(\MC_ARK_ARC_1_2/temp2[98] ), .B(
        \MC_ARK_ARC_1_2/temp1[98] ), .ZN(\MC_ARK_ARC_1_2/temp5[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_15_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[134] ), 
        .B(n273), .ZN(\MC_ARK_ARC_1_2/temp4[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_15_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[8] ), .ZN(\MC_ARK_ARC_1_2/temp3[98] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_15_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[44] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_2/temp2[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_15_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[98] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[92] ), .ZN(\MC_ARK_ARC_1_2/temp1[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_15_2  ( .A(\MC_ARK_ARC_1_2/temp5[99] ), .B(
        \MC_ARK_ARC_1_2/temp6[99] ), .ZN(\RI1[3][99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_15_2  ( .A(\MC_ARK_ARC_1_2/temp3[99] ), .B(
        \MC_ARK_ARC_1_2/temp4[99] ), .ZN(\MC_ARK_ARC_1_2/temp6[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_15_2  ( .A(\MC_ARK_ARC_1_2/temp2[99] ), .B(
        \MC_ARK_ARC_1_2/temp1[99] ), .ZN(\MC_ARK_ARC_1_2/temp5[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_15_2  ( .A(\RI5[2][135] ), .B(n428), .ZN(
        \MC_ARK_ARC_1_2/temp4[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_15_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[165] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_2/temp3[99] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_15_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .B(\RI5[2][69] ), .ZN(\MC_ARK_ARC_1_2/temp2[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_15_2  ( .A(\RI5[2][93] ), .B(\RI5[2][99] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_15_1  ( .A(\MC_ARK_ARC_1_2/temp6[100] ), .B(
        \MC_ARK_ARC_1_2/temp5[100] ), .ZN(\RI1[3][100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_15_1  ( .A(\MC_ARK_ARC_1_2/temp3[100] ), .B(
        \MC_ARK_ARC_1_2/temp4[100] ), .ZN(\MC_ARK_ARC_1_2/temp6[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_15_1  ( .A(\MC_ARK_ARC_1_2/temp2[100] ), .B(
        \MC_ARK_ARC_1_2/temp1[100] ), .ZN(\MC_ARK_ARC_1_2/temp5[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_15_1  ( .A(n1933), .B(n350), .ZN(
        \MC_ARK_ARC_1_2/temp4[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_15_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_15_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[46] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_15_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[94] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_15_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[137] ), 
        .B(n207), .ZN(\MC_ARK_ARC_1_2/temp4[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_15_0  ( .A(n1628), .B(
        \MC_ARK_ARC_1_2/buf_datainput[11] ), .ZN(\MC_ARK_ARC_1_2/temp3[101] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_15_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .B(n1502), .ZN(\MC_ARK_ARC_1_2/temp2[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_15_0  ( .A(n2126), .B(
        \MC_ARK_ARC_1_2/buf_datainput[95] ), .ZN(\MC_ARK_ARC_1_2/temp1[101] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_14_5  ( .A(\MC_ARK_ARC_1_2/temp5[102] ), .B(
        \MC_ARK_ARC_1_2/temp6[102] ), .ZN(\RI1[3][102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_14_5  ( .A(\MC_ARK_ARC_1_2/temp3[102] ), .B(
        \MC_ARK_ARC_1_2/temp4[102] ), .ZN(\MC_ARK_ARC_1_2/temp6[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_14_5  ( .A(\MC_ARK_ARC_1_2/temp1[102] ), .B(
        \MC_ARK_ARC_1_2/temp2[102] ), .ZN(\MC_ARK_ARC_1_2/temp5[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_14_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[138] ), 
        .B(n510), .ZN(\MC_ARK_ARC_1_2/temp4[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_14_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[12] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_14_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[48] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_14_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[96] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_14_4  ( .A(\MC_ARK_ARC_1_2/temp5[103] ), .B(
        \MC_ARK_ARC_1_2/temp6[103] ), .ZN(\RI1[3][103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_14_4  ( .A(\MC_ARK_ARC_1_2/temp3[103] ), .B(
        \MC_ARK_ARC_1_2/temp4[103] ), .ZN(\MC_ARK_ARC_1_2/temp6[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_14_4  ( .A(\MC_ARK_ARC_1_2/temp1[103] ), .B(
        \MC_ARK_ARC_1_2/temp2[103] ), .ZN(\MC_ARK_ARC_1_2/temp5[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_14_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[139] ), 
        .B(n285), .ZN(\MC_ARK_ARC_1_2/temp4[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_14_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[13] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[169] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_14_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[49] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_14_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[97] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_14_3  ( .A(\MC_ARK_ARC_1_2/temp6[104] ), .B(
        \MC_ARK_ARC_1_2/temp5[104] ), .ZN(\RI1[3][104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_14_3  ( .A(\MC_ARK_ARC_1_2/temp3[104] ), .B(
        \MC_ARK_ARC_1_2/temp4[104] ), .ZN(\MC_ARK_ARC_1_2/temp6[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_14_3  ( .A(\MC_ARK_ARC_1_2/temp1[104] ), .B(
        \MC_ARK_ARC_1_2/temp2[104] ), .ZN(\MC_ARK_ARC_1_2/temp5[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_14_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[140] ), 
        .B(n324), .ZN(\MC_ARK_ARC_1_2/temp4[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_14_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[14] ), 
        .B(n2144), .ZN(\MC_ARK_ARC_1_2/temp3[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_14_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[74] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_14_3  ( .A(n2122), .B(
        \MC_ARK_ARC_1_2/buf_datainput[98] ), .ZN(\MC_ARK_ARC_1_2/temp1[104] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_14_2  ( .A(\MC_ARK_ARC_1_2/temp5[105] ), .B(
        \MC_ARK_ARC_1_2/temp6[105] ), .ZN(\RI1[3][105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_14_2  ( .A(\MC_ARK_ARC_1_2/temp3[105] ), .B(
        \MC_ARK_ARC_1_2/temp4[105] ), .ZN(\MC_ARK_ARC_1_2/temp6[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_14_2  ( .A(\MC_ARK_ARC_1_2/temp1[105] ), .B(
        \MC_ARK_ARC_1_2/temp2[105] ), .ZN(\MC_ARK_ARC_1_2/temp5[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_14_2  ( .A(n1951), .B(n427), .ZN(
        \MC_ARK_ARC_1_2/temp4[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_14_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[15] ), 
        .B(\RI5[2][171] ), .ZN(\MC_ARK_ARC_1_2/temp3[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_14_2  ( .A(\RI5[2][51] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[75] ), .ZN(\MC_ARK_ARC_1_2/temp2[105] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_14_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .B(\RI5[2][99] ), .ZN(\MC_ARK_ARC_1_2/temp1[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_14_1  ( .A(\MC_ARK_ARC_1_2/temp6[106] ), .B(
        \MC_ARK_ARC_1_2/temp5[106] ), .ZN(\RI1[3][106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_14_1  ( .A(\MC_ARK_ARC_1_2/temp3[106] ), .B(
        \MC_ARK_ARC_1_2/temp4[106] ), .ZN(\MC_ARK_ARC_1_2/temp6[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_14_1  ( .A(\MC_ARK_ARC_1_2/temp1[106] ), .B(
        \MC_ARK_ARC_1_2/temp2[106] ), .ZN(\MC_ARK_ARC_1_2/temp5[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_14_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[142] ), 
        .B(n220), .ZN(\MC_ARK_ARC_1_2/temp4[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_14_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[16] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_14_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[76] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_14_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_14_0  ( .A(\MC_ARK_ARC_1_2/temp3[107] ), .B(
        \MC_ARK_ARC_1_2/temp4[107] ), .ZN(\MC_ARK_ARC_1_2/temp6[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_14_0  ( .A(\MC_ARK_ARC_1_2/temp1[107] ), .B(
        \MC_ARK_ARC_1_2/temp2[107] ), .ZN(\MC_ARK_ARC_1_2/temp5[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_14_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[107] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_14_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[17] ), 
        .B(n827), .ZN(\MC_ARK_ARC_1_2/temp3[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_14_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[77] ), 
        .B(n781), .ZN(\MC_ARK_ARC_1_2/temp2[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_14_0  ( .A(n1666), .B(n2127), .ZN(
        \MC_ARK_ARC_1_2/temp1[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_13_5  ( .A(\MC_ARK_ARC_1_2/temp5[108] ), .B(
        \MC_ARK_ARC_1_2/temp6[108] ), .ZN(\RI1[3][108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_13_5  ( .A(\MC_ARK_ARC_1_2/temp3[108] ), .B(
        \MC_ARK_ARC_1_2/temp4[108] ), .ZN(\MC_ARK_ARC_1_2/temp6[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_13_5  ( .A(\MC_ARK_ARC_1_2/temp1[108] ), .B(
        \MC_ARK_ARC_1_2/temp2[108] ), .ZN(\MC_ARK_ARC_1_2/temp5[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_13_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[144] ), 
        .B(n298), .ZN(\MC_ARK_ARC_1_2/temp4[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_13_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[18] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[174] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_13_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[54] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_13_5  ( .A(\RI5[2][108] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[102] ), .ZN(\MC_ARK_ARC_1_2/temp1[108] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_13_4  ( .A(\MC_ARK_ARC_1_2/temp5[109] ), .B(
        \MC_ARK_ARC_1_2/temp6[109] ), .ZN(\RI1[3][109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_13_4  ( .A(\MC_ARK_ARC_1_2/temp3[109] ), .B(
        \MC_ARK_ARC_1_2/temp4[109] ), .ZN(\MC_ARK_ARC_1_2/temp6[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_13_4  ( .A(\MC_ARK_ARC_1_2/temp1[109] ), .B(
        \MC_ARK_ARC_1_2/temp2[109] ), .ZN(\MC_ARK_ARC_1_2/temp5[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_13_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[145] ), 
        .B(n469), .ZN(\MC_ARK_ARC_1_2/temp4[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_13_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[19] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_13_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[55] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_13_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_13_3  ( .A(\MC_ARK_ARC_1_2/temp6[110] ), .B(
        \MC_ARK_ARC_1_2/temp5[110] ), .ZN(\RI1[3][110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_13_3  ( .A(\MC_ARK_ARC_1_2/temp3[110] ), .B(
        \MC_ARK_ARC_1_2/temp4[110] ), .ZN(\MC_ARK_ARC_1_2/temp6[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_13_3  ( .A(\MC_ARK_ARC_1_2/temp2[110] ), .B(
        \MC_ARK_ARC_1_2/temp1[110] ), .ZN(\MC_ARK_ARC_1_2/temp5[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_13_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .B(n193), .ZN(\MC_ARK_ARC_1_2/temp4[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_13_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[20] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_13_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[80] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[56] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_13_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[110] ), 
        .B(n2123), .ZN(\MC_ARK_ARC_1_2/temp1[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_13_2  ( .A(\MC_ARK_ARC_1_2/temp6[111] ), .B(
        \MC_ARK_ARC_1_2/temp5[111] ), .ZN(\RI1[3][111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_13_2  ( .A(\MC_ARK_ARC_1_2/temp3[111] ), .B(
        \MC_ARK_ARC_1_2/temp4[111] ), .ZN(\MC_ARK_ARC_1_2/temp6[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_13_2  ( .A(\MC_ARK_ARC_1_2/temp2[111] ), .B(
        \MC_ARK_ARC_1_2/temp1[111] ), .ZN(\MC_ARK_ARC_1_2/temp5[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_13_2  ( .A(n2140), .B(n233), .ZN(
        \MC_ARK_ARC_1_2/temp4[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_13_2  ( .A(\RI5[2][21] ), .B(\RI5[2][177] ), 
        .ZN(\MC_ARK_ARC_1_2/temp3[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_13_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[81] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[57] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_13_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .B(n1950), .ZN(\MC_ARK_ARC_1_2/temp1[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_13_1  ( .A(\MC_ARK_ARC_1_2/temp5[112] ), .B(
        \MC_ARK_ARC_1_2/temp6[112] ), .ZN(\RI1[3][112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_13_1  ( .A(\MC_ARK_ARC_1_2/temp3[112] ), .B(
        \MC_ARK_ARC_1_2/temp4[112] ), .ZN(\MC_ARK_ARC_1_2/temp6[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_13_1  ( .A(\MC_ARK_ARC_1_2/temp2[112] ), .B(
        \MC_ARK_ARC_1_2/temp1[112] ), .ZN(\MC_ARK_ARC_1_2/temp5[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_13_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[112] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_13_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[178] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[22] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_13_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[58] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_13_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[112] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_13_0  ( .A(\MC_ARK_ARC_1_2/temp5[113] ), .B(
        \MC_ARK_ARC_1_2/temp6[113] ), .ZN(\RI1[3][113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_13_0  ( .A(\MC_ARK_ARC_1_2/temp3[113] ), .B(
        \MC_ARK_ARC_1_2/temp4[113] ), .ZN(\MC_ARK_ARC_1_2/temp6[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_13_0  ( .A(\MC_ARK_ARC_1_2/temp1[113] ), .B(
        \MC_ARK_ARC_1_2/temp2[113] ), .ZN(\MC_ARK_ARC_1_2/temp5[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_13_0  ( .A(n816), .B(n486), .ZN(
        \MC_ARK_ARC_1_2/temp4[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_13_0  ( .A(n803), .B(
        \MC_ARK_ARC_1_2/buf_datainput[23] ), .ZN(\MC_ARK_ARC_1_2/temp3[113] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_13_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[83] ), 
        .B(n792), .ZN(\MC_ARK_ARC_1_2/temp2[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_13_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[113] ), 
        .B(n1666), .ZN(\MC_ARK_ARC_1_2/temp1[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_12_5  ( .A(\MC_ARK_ARC_1_2/temp5[114] ), .B(
        \MC_ARK_ARC_1_2/temp6[114] ), .ZN(\RI1[3][114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_12_5  ( .A(\MC_ARK_ARC_1_2/temp3[114] ), .B(
        \MC_ARK_ARC_1_2/temp4[114] ), .ZN(\MC_ARK_ARC_1_2/temp6[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_12_5  ( .A(\MC_ARK_ARC_1_2/temp1[114] ), .B(
        \MC_ARK_ARC_1_2/temp2[114] ), .ZN(\MC_ARK_ARC_1_2/temp5[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_12_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[150] ), 
        .B(n348), .ZN(\MC_ARK_ARC_1_2/temp4[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_12_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_12_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[60] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_12_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[114] ), 
        .B(\RI5[2][108] ), .ZN(\MC_ARK_ARC_1_2/temp1[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_12_4  ( .A(\MC_ARK_ARC_1_2/temp6[115] ), .B(
        \MC_ARK_ARC_1_2/temp5[115] ), .ZN(\RI1[3][115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_12_4  ( .A(\MC_ARK_ARC_1_2/temp3[115] ), .B(
        \MC_ARK_ARC_1_2/temp4[115] ), .ZN(\MC_ARK_ARC_1_2/temp6[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_12_4  ( .A(\MC_ARK_ARC_1_2/temp1[115] ), .B(
        \MC_ARK_ARC_1_2/temp2[115] ), .ZN(\MC_ARK_ARC_1_2/temp5[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_12_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .B(n436), .ZN(\MC_ARK_ARC_1_2/temp4[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_12_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[25] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[181] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_12_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[61] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_12_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[109] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_12_3  ( .A(\MC_ARK_ARC_1_2/temp5[116] ), .B(
        \MC_ARK_ARC_1_2/temp6[116] ), .ZN(\RI1[3][116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_12_3  ( .A(\MC_ARK_ARC_1_2/temp3[116] ), .B(
        \MC_ARK_ARC_1_2/temp4[116] ), .ZN(\MC_ARK_ARC_1_2/temp6[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_12_3  ( .A(\MC_ARK_ARC_1_2/temp2[116] ), .B(
        \MC_ARK_ARC_1_2/temp1[116] ), .ZN(\MC_ARK_ARC_1_2/temp5[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_12_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[152] ), 
        .B(n408), .ZN(\MC_ARK_ARC_1_2/temp4[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_12_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[26] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_12_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[86] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_12_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[116] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_12_2  ( .A(\MC_ARK_ARC_1_2/temp5[117] ), .B(
        \MC_ARK_ARC_1_2/temp6[117] ), .ZN(\RI1[3][117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_12_2  ( .A(\MC_ARK_ARC_1_2/temp3[117] ), .B(
        \MC_ARK_ARC_1_2/temp4[117] ), .ZN(\MC_ARK_ARC_1_2/temp6[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_12_2  ( .A(\MC_ARK_ARC_1_2/temp1[117] ), .B(
        \MC_ARK_ARC_1_2/temp2[117] ), .ZN(\MC_ARK_ARC_1_2/temp5[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_12_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[153] ), 
        .B(n424), .ZN(\MC_ARK_ARC_1_2/temp4[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_12_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[27] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[183] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_12_2  ( .A(\RI5[2][87] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[63] ), .ZN(\MC_ARK_ARC_1_2/temp2[117] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_12_2  ( .A(n1950), .B(\RI5[2][117] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_12_1  ( .A(\MC_ARK_ARC_1_2/temp6[118] ), .B(
        \MC_ARK_ARC_1_2/temp5[118] ), .ZN(\RI1[3][118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_12_1  ( .A(\MC_ARK_ARC_1_2/temp3[118] ), .B(
        \MC_ARK_ARC_1_2/temp4[118] ), .ZN(\MC_ARK_ARC_1_2/temp6[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_12_1  ( .A(\MC_ARK_ARC_1_2/temp1[118] ), .B(
        \MC_ARK_ARC_1_2/temp2[118] ), .ZN(\MC_ARK_ARC_1_2/temp5[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_12_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[118] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_12_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[184] ), 
        .B(n2142), .ZN(\MC_ARK_ARC_1_2/temp3[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_12_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[64] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_12_1  ( .A(n1957), .B(
        \MC_ARK_ARC_1_2/buf_datainput[112] ), .ZN(\MC_ARK_ARC_1_2/temp1[118] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_12_0  ( .A(\MC_ARK_ARC_1_2/temp5[119] ), .B(
        \MC_ARK_ARC_1_2/temp6[119] ), .ZN(\RI1[3][119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_12_0  ( .A(\MC_ARK_ARC_1_2/temp3[119] ), .B(
        \MC_ARK_ARC_1_2/temp4[119] ), .ZN(\MC_ARK_ARC_1_2/temp6[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_12_0  ( .A(\MC_ARK_ARC_1_2/temp2[119] ), .B(
        \MC_ARK_ARC_1_2/temp1[119] ), .ZN(\MC_ARK_ARC_1_2/temp5[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_12_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[155] ), 
        .B(n361), .ZN(\MC_ARK_ARC_1_2/temp4[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_12_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[185] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_12_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .B(n1956), .ZN(\MC_ARK_ARC_1_2/temp2[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_12_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[113] ), 
        .B(n811), .ZN(\MC_ARK_ARC_1_2/temp1[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_11_5  ( .A(\MC_ARK_ARC_1_2/temp5[120] ), .B(
        \MC_ARK_ARC_1_2/temp6[120] ), .ZN(\RI1[3][120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_11_5  ( .A(\MC_ARK_ARC_1_2/temp3[120] ), .B(
        \MC_ARK_ARC_1_2/temp4[120] ), .ZN(\MC_ARK_ARC_1_2/temp6[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_11_5  ( .A(\MC_ARK_ARC_1_2/temp1[120] ), .B(
        \MC_ARK_ARC_1_2/temp2[120] ), .ZN(\MC_ARK_ARC_1_2/temp5[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_11_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .B(n218), .ZN(\MC_ARK_ARC_1_2/temp4[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_11_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[30] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[186] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_11_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[66] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_11_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[114] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_11_4  ( .A(\MC_ARK_ARC_1_2/temp5[121] ), .B(
        \MC_ARK_ARC_1_2/temp6[121] ), .ZN(\RI1[3][121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_11_4  ( .A(\MC_ARK_ARC_1_2/temp3[121] ), .B(
        \MC_ARK_ARC_1_2/temp4[121] ), .ZN(\MC_ARK_ARC_1_2/temp6[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_11_4  ( .A(\MC_ARK_ARC_1_2/temp1[121] ), .B(
        \MC_ARK_ARC_1_2/temp2[121] ), .ZN(\MC_ARK_ARC_1_2/temp5[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_11_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[157] ), 
        .B(n256), .ZN(\MC_ARK_ARC_1_2/temp4[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_11_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[31] ), 
        .B(\RI5[2][187] ), .ZN(\MC_ARK_ARC_1_2/temp3[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_11_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[67] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_11_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_11_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[158] ), 
        .B(n296), .ZN(\MC_ARK_ARC_1_2/temp4[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_11_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[188] ), 
        .B(n1511), .ZN(\MC_ARK_ARC_1_2/temp3[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_11_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[92] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_11_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[122] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_11_2  ( .A(\RI5[2][159] ), .B(n335), .ZN(
        \MC_ARK_ARC_1_2/temp4[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_11_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[189] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_11_2  ( .A(\RI5[2][69] ), .B(\RI5[2][93] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_11_2  ( .A(\RI5[2][123] ), .B(\RI5[2][117] ), 
        .ZN(\MC_ARK_ARC_1_2/temp1[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_11_1  ( .A(\MC_ARK_ARC_1_2/temp6[124] ), .B(
        \MC_ARK_ARC_1_2/temp5[124] ), .ZN(\RI1[3][124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_11_1  ( .A(\MC_ARK_ARC_1_2/temp3[124] ), .B(
        \MC_ARK_ARC_1_2/temp4[124] ), .ZN(\MC_ARK_ARC_1_2/temp6[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_11_1  ( .A(\MC_ARK_ARC_1_2/temp1[124] ), .B(
        \MC_ARK_ARC_1_2/temp2[124] ), .ZN(\MC_ARK_ARC_1_2/temp5[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_11_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[160] ), 
        .B(n373), .ZN(\MC_ARK_ARC_1_2/temp4[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_11_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_11_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[70] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_11_1  ( .A(n1957), .B(
        \MC_ARK_ARC_1_2/buf_datainput[124] ), .ZN(\MC_ARK_ARC_1_2/temp1[124] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_11_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[161] ), 
        .B(n231), .ZN(\MC_ARK_ARC_1_2/temp4[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_11_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .B(n829), .ZN(\MC_ARK_ARC_1_2/temp3[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_11_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .B(n1502), .ZN(\MC_ARK_ARC_1_2/temp2[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_11_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .B(n811), .ZN(\MC_ARK_ARC_1_2/temp1[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_10_5  ( .A(\MC_ARK_ARC_1_2/temp5[126] ), .B(
        \MC_ARK_ARC_1_2/temp6[126] ), .ZN(\RI1[3][126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_10_5  ( .A(\MC_ARK_ARC_1_2/temp3[126] ), .B(
        \MC_ARK_ARC_1_2/temp4[126] ), .ZN(\MC_ARK_ARC_1_2/temp6[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_10_5  ( .A(\MC_ARK_ARC_1_2/temp2[126] ), .B(
        \MC_ARK_ARC_1_2/temp1[126] ), .ZN(\MC_ARK_ARC_1_2/temp5[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_10_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .B(n509), .ZN(\MC_ARK_ARC_1_2/temp4[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_10_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[36] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[0] ), .ZN(\MC_ARK_ARC_1_2/temp3[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_10_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[72] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_10_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_10_4  ( .A(\MC_ARK_ARC_1_2/temp5[127] ), .B(
        \MC_ARK_ARC_1_2/temp6[127] ), .ZN(\RI1[3][127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_10_4  ( .A(\MC_ARK_ARC_1_2/temp3[127] ), .B(
        \MC_ARK_ARC_1_2/temp4[127] ), .ZN(\MC_ARK_ARC_1_2/temp6[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_10_4  ( .A(\MC_ARK_ARC_1_2/temp1[127] ), .B(
        \MC_ARK_ARC_1_2/temp2[127] ), .ZN(\MC_ARK_ARC_1_2/temp5[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_10_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[163] ), 
        .B(n459), .ZN(\MC_ARK_ARC_1_2/temp4[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_10_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[37] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[1] ), .ZN(\MC_ARK_ARC_1_2/temp3[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_10_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[73] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_10_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_10_3  ( .A(\MC_ARK_ARC_1_2/temp5[128] ), .B(
        \MC_ARK_ARC_1_2/temp6[128] ), .ZN(\RI1[3][128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_10_3  ( .A(\MC_ARK_ARC_1_2/temp3[128] ), .B(
        \MC_ARK_ARC_1_2/temp4[128] ), .ZN(\MC_ARK_ARC_1_2/temp6[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_10_3  ( .A(\MC_ARK_ARC_1_2/temp1[128] ), .B(
        \MC_ARK_ARC_1_2/temp2[128] ), .ZN(\MC_ARK_ARC_1_2/temp5[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_10_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .B(n346), .ZN(\MC_ARK_ARC_1_2/temp4[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_10_3  ( .A(\RI5[2][2] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[38] ), .ZN(\MC_ARK_ARC_1_2/temp3[128] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_10_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[98] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_10_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_10_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[165] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[129] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_10_2  ( .A(\RI5[2][39] ), .B(\RI5[2][3] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_10_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[75] ), 
        .B(\RI5[2][99] ), .ZN(\MC_ARK_ARC_1_2/temp2[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_10_2  ( .A(\RI5[2][123] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[129] ), .ZN(\MC_ARK_ARC_1_2/temp1[129] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_10_1  ( .A(\MC_ARK_ARC_1_2/temp6[130] ), .B(
        \MC_ARK_ARC_1_2/temp5[130] ), .ZN(\RI1[3][130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_10_1  ( .A(\MC_ARK_ARC_1_2/temp3[130] ), .B(
        \MC_ARK_ARC_1_2/temp4[130] ), .ZN(\MC_ARK_ARC_1_2/temp6[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_10_1  ( .A(\MC_ARK_ARC_1_2/temp1[130] ), .B(
        \MC_ARK_ARC_1_2/temp2[130] ), .ZN(\MC_ARK_ARC_1_2/temp5[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_10_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[166] ), 
        .B(n243), .ZN(\MC_ARK_ARC_1_2/temp4[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_10_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_2/temp3[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_10_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[76] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_10_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_10_0  ( .A(\MC_ARK_ARC_1_2/temp1[131] ), .B(
        \MC_ARK_ARC_1_2/temp2[131] ), .ZN(\MC_ARK_ARC_1_2/temp5[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_10_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[167] ), 
        .B(n282), .ZN(\MC_ARK_ARC_1_2/temp4[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_10_0  ( .A(n1633), .B(
        \MC_ARK_ARC_1_2/buf_datainput[41] ), .ZN(\MC_ARK_ARC_1_2/temp3[131] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_10_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[77] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[101] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_10_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[125] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_9_5  ( .A(\MC_ARK_ARC_1_2/temp5[132] ), .B(
        \MC_ARK_ARC_1_2/temp6[132] ), .ZN(\RI1[3][132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_9_5  ( .A(\MC_ARK_ARC_1_2/temp3[132] ), .B(
        \MC_ARK_ARC_1_2/temp4[132] ), .ZN(\MC_ARK_ARC_1_2/temp6[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_9_5  ( .A(\MC_ARK_ARC_1_2/temp1[132] ), .B(
        \MC_ARK_ARC_1_2/temp2[132] ), .ZN(\MC_ARK_ARC_1_2/temp5[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_9_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[168] ), 
        .B(n320), .ZN(\MC_ARK_ARC_1_2/temp4[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_9_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[42] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[6] ), .ZN(\MC_ARK_ARC_1_2/temp3[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_9_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[102] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[78] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_9_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[132] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[126] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_9_4  ( .A(\MC_ARK_ARC_1_2/temp5[133] ), .B(
        \MC_ARK_ARC_1_2/temp6[133] ), .ZN(\RI1[3][133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_9_4  ( .A(\MC_ARK_ARC_1_2/temp3[133] ), .B(
        \MC_ARK_ARC_1_2/temp4[133] ), .ZN(\MC_ARK_ARC_1_2/temp6[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_9_4  ( .A(\MC_ARK_ARC_1_2/temp1[133] ), .B(
        \MC_ARK_ARC_1_2/temp2[133] ), .ZN(\MC_ARK_ARC_1_2/temp5[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_9_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[169] ), 
        .B(n452), .ZN(\MC_ARK_ARC_1_2/temp4[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_9_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[43] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[7] ), .ZN(\MC_ARK_ARC_1_2/temp3[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_9_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[103] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[79] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_9_4  ( .A(\RI5[2][133] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[127] ), .ZN(\MC_ARK_ARC_1_2/temp1[133] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_9_3  ( .A(\MC_ARK_ARC_1_2/temp5[134] ), .B(
        \MC_ARK_ARC_1_2/temp6[134] ), .ZN(\RI1[3][134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_9_3  ( .A(\MC_ARK_ARC_1_2/temp3[134] ), .B(
        \MC_ARK_ARC_1_2/temp4[134] ), .ZN(\MC_ARK_ARC_1_2/temp6[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_9_3  ( .A(\MC_ARK_ARC_1_2/temp2[134] ), .B(
        \MC_ARK_ARC_1_2/temp1[134] ), .ZN(\MC_ARK_ARC_1_2/temp5[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_9_3  ( .A(n2144), .B(n216), .ZN(
        \MC_ARK_ARC_1_2/temp4[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_9_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[8] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[44] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_9_3  ( .A(n2122), .B(
        \MC_ARK_ARC_1_2/buf_datainput[80] ), .ZN(\MC_ARK_ARC_1_2/temp2[134] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_9_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_9_2  ( .A(\MC_ARK_ARC_1_2/temp5[135] ), .B(
        \MC_ARK_ARC_1_2/temp6[135] ), .ZN(\RI1[3][135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_9_2  ( .A(\MC_ARK_ARC_1_2/temp4[135] ), .B(
        \MC_ARK_ARC_1_2/temp3[135] ), .ZN(\MC_ARK_ARC_1_2/temp6[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_9_2  ( .A(\MC_ARK_ARC_1_2/temp2[135] ), .B(
        \MC_ARK_ARC_1_2/temp1[135] ), .ZN(\MC_ARK_ARC_1_2/temp5[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_9_2  ( .A(\RI5[2][171] ), .B(n254), .ZN(
        \MC_ARK_ARC_1_2/temp4[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_9_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[9] ), .ZN(\MC_ARK_ARC_1_2/temp3[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_9_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[81] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_9_2  ( .A(n2098), .B(n815), .ZN(
        \MC_ARK_ARC_1_2/temp1[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_9_1  ( .A(\MC_ARK_ARC_1_2/temp6[136] ), .B(
        \MC_ARK_ARC_1_2/temp5[136] ), .ZN(\RI1[3][136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_9_1  ( .A(\MC_ARK_ARC_1_2/temp3[136] ), .B(
        \MC_ARK_ARC_1_2/temp4[136] ), .ZN(\MC_ARK_ARC_1_2/temp6[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_9_1  ( .A(\MC_ARK_ARC_1_2/temp1[136] ), .B(
        \MC_ARK_ARC_1_2/temp2[136] ), .ZN(\MC_ARK_ARC_1_2/temp5[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_9_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[189] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_9_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[46] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[10] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_9_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[82] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_9_1  ( .A(n1932), .B(
        \MC_ARK_ARC_1_2/buf_datainput[130] ), .ZN(\MC_ARK_ARC_1_2/temp1[136] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_9_0  ( .A(\MC_ARK_ARC_1_2/temp6[137] ), .B(
        \MC_ARK_ARC_1_2/temp5[137] ), .ZN(\RI1[3][137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_9_0  ( .A(\MC_ARK_ARC_1_2/temp3[137] ), .B(
        \MC_ARK_ARC_1_2/temp4[137] ), .ZN(\MC_ARK_ARC_1_2/temp6[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_9_0  ( .A(\MC_ARK_ARC_1_2/temp1[137] ), .B(
        \MC_ARK_ARC_1_2/temp2[137] ), .ZN(\MC_ARK_ARC_1_2/temp5[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_9_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[173] ), 
        .B(n475), .ZN(\MC_ARK_ARC_1_2/temp4[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_9_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[11] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_9_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[83] ), 
        .B(n1665), .ZN(\MC_ARK_ARC_1_2/temp2[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_9_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[137] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_8_5  ( .A(\MC_ARK_ARC_1_2/temp5[138] ), .B(
        \MC_ARK_ARC_1_2/temp6[138] ), .ZN(\RI1[3][138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_8_5  ( .A(\MC_ARK_ARC_1_2/temp3[138] ), .B(
        \MC_ARK_ARC_1_2/temp4[138] ), .ZN(\MC_ARK_ARC_1_2/temp6[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_8_5  ( .A(\MC_ARK_ARC_1_2/temp1[138] ), .B(
        \MC_ARK_ARC_1_2/temp2[138] ), .ZN(\MC_ARK_ARC_1_2/temp5[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_8_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[174] ), 
        .B(n473), .ZN(\MC_ARK_ARC_1_2/temp4[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_8_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[48] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[12] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_8_5  ( .A(\RI5[2][108] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[84] ), .ZN(\MC_ARK_ARC_1_2/temp2[138] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_8_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[138] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[132] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_8_4  ( .A(\MC_ARK_ARC_1_2/temp5[139] ), .B(
        \MC_ARK_ARC_1_2/temp6[139] ), .ZN(\RI1[3][139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_8_4  ( .A(\MC_ARK_ARC_1_2/temp3[139] ), .B(
        \MC_ARK_ARC_1_2/temp4[139] ), .ZN(\MC_ARK_ARC_1_2/temp6[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_8_4  ( .A(\MC_ARK_ARC_1_2/temp1[139] ), .B(
        \MC_ARK_ARC_1_2/temp2[139] ), .ZN(\MC_ARK_ARC_1_2/temp5[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_8_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[175] ), 
        .B(n489), .ZN(\MC_ARK_ARC_1_2/temp4[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_8_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[13] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_8_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[109] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[85] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_8_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[139] ), 
        .B(\RI5[2][133] ), .ZN(\MC_ARK_ARC_1_2/temp1[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_8_3  ( .A(\MC_ARK_ARC_1_2/temp6[140] ), .B(
        \MC_ARK_ARC_1_2/temp5[140] ), .ZN(\RI1[3][140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_8_3  ( .A(\MC_ARK_ARC_1_2/temp3[140] ), .B(
        \MC_ARK_ARC_1_2/temp4[140] ), .ZN(\MC_ARK_ARC_1_2/temp6[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_8_3  ( .A(\MC_ARK_ARC_1_2/temp1[140] ), .B(
        \MC_ARK_ARC_1_2/temp2[140] ), .ZN(\MC_ARK_ARC_1_2/temp5[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_8_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[176] ), 
        .B(n267), .ZN(\MC_ARK_ARC_1_2/temp4[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_8_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[50] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_8_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[86] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_8_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[134] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_8_2  ( .A(\MC_ARK_ARC_1_2/temp6[141] ), .B(
        \MC_ARK_ARC_1_2/temp5[141] ), .ZN(\RI1[3][141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_8_2  ( .A(\MC_ARK_ARC_1_2/temp3[141] ), .B(
        \MC_ARK_ARC_1_2/temp4[141] ), .ZN(\MC_ARK_ARC_1_2/temp6[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_8_2  ( .A(\MC_ARK_ARC_1_2/temp1[141] ), .B(
        \MC_ARK_ARC_1_2/temp2[141] ), .ZN(\MC_ARK_ARC_1_2/temp5[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_8_2  ( .A(\RI5[2][177] ), .B(Key[72]), .ZN(
        \MC_ARK_ARC_1_2/temp4[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_8_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[15] ), 
        .B(\RI5[2][51] ), .ZN(\MC_ARK_ARC_1_2/temp3[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_8_2  ( .A(\RI5[2][87] ), .B(n1950), .ZN(
        \MC_ARK_ARC_1_2/temp2[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_8_2  ( .A(n1951), .B(n2099), .ZN(
        \MC_ARK_ARC_1_2/temp1[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_8_1  ( .A(\MC_ARK_ARC_1_2/temp5[142] ), .B(
        \MC_ARK_ARC_1_2/temp6[142] ), .ZN(\RI1[3][142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_8_1  ( .A(\MC_ARK_ARC_1_2/temp4[142] ), .B(
        \MC_ARK_ARC_1_2/temp3[142] ), .ZN(\MC_ARK_ARC_1_2/temp6[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_8_1  ( .A(\MC_ARK_ARC_1_2/temp1[142] ), .B(
        \MC_ARK_ARC_1_2/temp2[142] ), .ZN(\MC_ARK_ARC_1_2/temp5[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_8_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[178] ), 
        .B(n344), .ZN(\MC_ARK_ARC_1_2/temp4[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_8_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[16] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_8_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[88] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_8_1  ( .A(n1932), .B(
        \MC_ARK_ARC_1_2/buf_datainput[142] ), .ZN(\MC_ARK_ARC_1_2/temp1[142] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_8_0  ( .A(\MC_ARK_ARC_1_2/temp5[143] ), .B(
        \MC_ARK_ARC_1_2/temp6[143] ), .ZN(\RI1[3][143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_8_0  ( .A(\MC_ARK_ARC_1_2/temp3[143] ), .B(
        \MC_ARK_ARC_1_2/temp4[143] ), .ZN(\MC_ARK_ARC_1_2/temp6[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_8_0  ( .A(\MC_ARK_ARC_1_2/temp1[143] ), .B(
        \MC_ARK_ARC_1_2/temp2[143] ), .ZN(\MC_ARK_ARC_1_2/temp5[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_8_0  ( .A(n802), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[143] ), .ZN(\MC_ARK_ARC_1_2/temp4[143] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_8_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[17] ), 
        .B(n782), .ZN(\MC_ARK_ARC_1_2/temp3[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_8_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[113] ), 
        .B(n1956), .ZN(\MC_ARK_ARC_1_2/temp2[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_8_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[143] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_7_5  ( .A(\MC_ARK_ARC_1_2/temp5[144] ), .B(
        \MC_ARK_ARC_1_2/temp6[144] ), .ZN(\RI1[3][144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_7_5  ( .A(\MC_ARK_ARC_1_2/temp3[144] ), .B(
        \MC_ARK_ARC_1_2/temp4[144] ), .ZN(\MC_ARK_ARC_1_2/temp6[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_7_5  ( .A(\MC_ARK_ARC_1_2/temp1[144] ), .B(
        \MC_ARK_ARC_1_2/temp2[144] ), .ZN(\MC_ARK_ARC_1_2/temp5[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_7_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[180] ), 
        .B(n513), .ZN(\MC_ARK_ARC_1_2/temp4[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_7_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[54] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[18] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_7_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[114] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[90] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_7_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[144] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[138] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_7_4  ( .A(\MC_ARK_ARC_1_2/temp5[145] ), .B(
        \MC_ARK_ARC_1_2/temp6[145] ), .ZN(\RI1[3][145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_7_4  ( .A(\MC_ARK_ARC_1_2/temp3[145] ), .B(
        \MC_ARK_ARC_1_2/temp4[145] ), .ZN(\MC_ARK_ARC_1_2/temp6[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_7_4  ( .A(\MC_ARK_ARC_1_2/temp1[145] ), .B(
        \MC_ARK_ARC_1_2/temp2[145] ), .ZN(\MC_ARK_ARC_1_2/temp5[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_7_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[181] ), 
        .B(n463), .ZN(\MC_ARK_ARC_1_2/temp4[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_7_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[55] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[19] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_7_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[91] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_7_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[139] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_7_3  ( .A(\MC_ARK_ARC_1_2/temp5[146] ), .B(
        \MC_ARK_ARC_1_2/temp6[146] ), .ZN(\RI1[3][146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_7_3  ( .A(\MC_ARK_ARC_1_2/temp3[146] ), .B(
        \MC_ARK_ARC_1_2/temp4[146] ), .ZN(\MC_ARK_ARC_1_2/temp6[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_7_3  ( .A(\MC_ARK_ARC_1_2/temp1[146] ), .B(
        \MC_ARK_ARC_1_2/temp2[146] ), .ZN(\MC_ARK_ARC_1_2/temp5[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_7_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[182] ), 
        .B(n319), .ZN(\MC_ARK_ARC_1_2/temp4[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_7_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[56] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_7_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[92] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_7_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[140] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_7_2  ( .A(\MC_ARK_ARC_1_2/temp5[147] ), .B(
        \MC_ARK_ARC_1_2/temp6[147] ), .ZN(\RI1[3][147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_7_2  ( .A(\MC_ARK_ARC_1_2/temp3[147] ), .B(
        \MC_ARK_ARC_1_2/temp4[147] ), .ZN(\MC_ARK_ARC_1_2/temp6[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_7_2  ( .A(\MC_ARK_ARC_1_2/temp1[147] ), .B(
        \MC_ARK_ARC_1_2/temp2[147] ), .ZN(\MC_ARK_ARC_1_2/temp5[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_7_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[183] ), 
        .B(n357), .ZN(\MC_ARK_ARC_1_2/temp4[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_7_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[57] ), 
        .B(\RI5[2][21] ), .ZN(\MC_ARK_ARC_1_2/temp3[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_7_2  ( .A(\RI5[2][117] ), .B(\RI5[2][93] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_7_2  ( .A(n2139), .B(n1951), .ZN(
        \MC_ARK_ARC_1_2/temp1[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_7_1  ( .A(\MC_ARK_ARC_1_2/temp6[148] ), .B(
        \MC_ARK_ARC_1_2/temp5[148] ), .ZN(\RI1[3][148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_7_1  ( .A(\MC_ARK_ARC_1_2/temp3[148] ), .B(
        \MC_ARK_ARC_1_2/temp4[148] ), .ZN(\MC_ARK_ARC_1_2/temp6[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_7_1  ( .A(\MC_ARK_ARC_1_2/temp1[148] ), .B(
        \MC_ARK_ARC_1_2/temp2[148] ), .ZN(\MC_ARK_ARC_1_2/temp5[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_7_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[184] ), 
        .B(n214), .ZN(\MC_ARK_ARC_1_2/temp4[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_7_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[58] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[22] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_7_1  ( .A(n1957), .B(
        \MC_ARK_ARC_1_2/buf_datainput[94] ), .ZN(\MC_ARK_ARC_1_2/temp2[148] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_7_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[142] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_7_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[185] ), 
        .B(n252), .ZN(\MC_ARK_ARC_1_2/temp4[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_7_0  ( .A(n793), .B(n800), .ZN(
        \MC_ARK_ARC_1_2/temp3[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_7_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .B(n812), .ZN(\MC_ARK_ARC_1_2/temp2[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_7_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .B(n816), .ZN(\MC_ARK_ARC_1_2/temp1[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_6_5  ( .A(\MC_ARK_ARC_1_2/temp5[150] ), .B(
        \MC_ARK_ARC_1_2/temp6[150] ), .ZN(\RI1[3][150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_6_5  ( .A(\MC_ARK_ARC_1_2/temp3[150] ), .B(
        \MC_ARK_ARC_1_2/temp4[150] ), .ZN(\MC_ARK_ARC_1_2/temp6[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_6_5  ( .A(\MC_ARK_ARC_1_2/temp1[150] ), .B(
        \MC_ARK_ARC_1_2/temp2[150] ), .ZN(\MC_ARK_ARC_1_2/temp5[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_6_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[186] ), 
        .B(n292), .ZN(\MC_ARK_ARC_1_2/temp4[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_6_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[60] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[24] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_6_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[120] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[96] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_6_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[150] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[144] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_6_4  ( .A(\MC_ARK_ARC_1_2/temp5[151] ), .B(
        \MC_ARK_ARC_1_2/temp6[151] ), .ZN(\RI1[3][151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_6_4  ( .A(\MC_ARK_ARC_1_2/temp3[151] ), .B(
        \MC_ARK_ARC_1_2/temp4[151] ), .ZN(\MC_ARK_ARC_1_2/temp6[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_6_4  ( .A(\MC_ARK_ARC_1_2/temp1[151] ), .B(
        \MC_ARK_ARC_1_2/temp2[151] ), .ZN(\MC_ARK_ARC_1_2/temp5[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_6_4  ( .A(\RI5[2][187] ), .B(n462), .ZN(
        \MC_ARK_ARC_1_2/temp4[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_6_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[25] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_6_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[97] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_6_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[145] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_6_3  ( .A(\MC_ARK_ARC_1_2/temp5[152] ), .B(
        \MC_ARK_ARC_1_2/temp6[152] ), .ZN(\RI1[3][152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_6_3  ( .A(\MC_ARK_ARC_1_2/temp3[152] ), .B(
        \MC_ARK_ARC_1_2/temp4[152] ), .ZN(\MC_ARK_ARC_1_2/temp6[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_6_3  ( .A(\MC_ARK_ARC_1_2/temp2[152] ), .B(
        \MC_ARK_ARC_1_2/temp1[152] ), .ZN(\MC_ARK_ARC_1_2/temp5[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_6_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[188] ), 
        .B(n369), .ZN(\MC_ARK_ARC_1_2/temp4[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_6_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[26] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_6_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[122] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[98] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_6_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[152] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_6_2  ( .A(\MC_ARK_ARC_1_2/temp6[153] ), .B(
        \MC_ARK_ARC_1_2/temp5[153] ), .ZN(\RI1[3][153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_6_2  ( .A(\MC_ARK_ARC_1_2/temp3[153] ), .B(
        \MC_ARK_ARC_1_2/temp4[153] ), .ZN(\MC_ARK_ARC_1_2/temp6[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_6_2  ( .A(\MC_ARK_ARC_1_2/temp2[153] ), .B(
        \MC_ARK_ARC_1_2/temp1[153] ), .ZN(\MC_ARK_ARC_1_2/temp5[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_6_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[189] ), 
        .B(n377), .ZN(\MC_ARK_ARC_1_2/temp4[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_6_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[27] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_6_2  ( .A(\RI5[2][99] ), .B(\RI5[2][123] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_6_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[153] ), 
        .B(\RI5[2][147] ), .ZN(\MC_ARK_ARC_1_2/temp1[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_6_1  ( .A(\MC_ARK_ARC_1_2/temp5[154] ), .B(
        \MC_ARK_ARC_1_2/temp6[154] ), .ZN(\RI1[3][154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_6_1  ( .A(\MC_ARK_ARC_1_2/temp3[154] ), .B(
        \MC_ARK_ARC_1_2/temp4[154] ), .ZN(\MC_ARK_ARC_1_2/temp6[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_6_1  ( .A(\MC_ARK_ARC_1_2/temp1[154] ), .B(
        \MC_ARK_ARC_1_2/temp2[154] ), .ZN(\MC_ARK_ARC_1_2/temp5[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_6_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[190] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[123] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_6_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[64] ), 
        .B(n2142), .ZN(\MC_ARK_ARC_1_2/temp3[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_6_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_6_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_6_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[191] ), 
        .B(n304), .ZN(\MC_ARK_ARC_1_2/temp4[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_6_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[29] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_6_0  ( .A(n2126), .B(
        \MC_ARK_ARC_1_2/buf_datainput[125] ), .ZN(\MC_ARK_ARC_1_2/temp2[155] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_6_0  ( .A(n817), .B(
        \MC_ARK_ARC_1_2/buf_datainput[155] ), .ZN(\MC_ARK_ARC_1_2/temp1[155] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_5_5  ( .A(\MC_ARK_ARC_1_2/temp5[156] ), .B(
        \MC_ARK_ARC_1_2/temp6[156] ), .ZN(\RI1[3][156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_5_5  ( .A(\MC_ARK_ARC_1_2/temp3[156] ), .B(
        \MC_ARK_ARC_1_2/temp4[156] ), .ZN(\MC_ARK_ARC_1_2/temp6[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_5_5  ( .A(\MC_ARK_ARC_1_2/temp1[156] ), .B(
        \MC_ARK_ARC_1_2/temp2[156] ), .ZN(\MC_ARK_ARC_1_2/temp5[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_5_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .B(n504), .ZN(\MC_ARK_ARC_1_2/temp4[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_5_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[66] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[30] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_5_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[126] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[102] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_5_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[150] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_5_4  ( .A(\MC_ARK_ARC_1_2/temp5[157] ), .B(
        \MC_ARK_ARC_1_2/temp6[157] ), .ZN(\RI1[3][157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_5_4  ( .A(\MC_ARK_ARC_1_2/temp3[157] ), .B(
        \MC_ARK_ARC_1_2/temp4[157] ), .ZN(\MC_ARK_ARC_1_2/temp6[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_5_4  ( .A(\MC_ARK_ARC_1_2/temp1[157] ), .B(
        \MC_ARK_ARC_1_2/temp2[157] ), .ZN(\MC_ARK_ARC_1_2/temp5[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_5_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[1] ), 
        .B(n474), .ZN(\MC_ARK_ARC_1_2/temp4[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_5_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[67] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[31] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_5_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[127] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[103] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_5_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[157] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[151] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_5_3  ( .A(\MC_ARK_ARC_1_2/temp5[158] ), .B(
        \MC_ARK_ARC_1_2/temp6[158] ), .ZN(\RI1[3][158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_5_3  ( .A(\MC_ARK_ARC_1_2/temp3[158] ), .B(
        \MC_ARK_ARC_1_2/temp4[158] ), .ZN(\MC_ARK_ARC_1_2/temp6[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_5_3  ( .A(\MC_ARK_ARC_1_2/temp2[158] ), .B(
        \MC_ARK_ARC_1_2/temp1[158] ), .ZN(\MC_ARK_ARC_1_2/temp5[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_5_3  ( .A(\RI5[2][2] ), .B(n240), .ZN(
        \MC_ARK_ARC_1_2/temp4[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_5_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .B(n1511), .ZN(\MC_ARK_ARC_1_2/temp3[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_5_3  ( .A(n2122), .B(
        \MC_ARK_ARC_1_2/buf_datainput[128] ), .ZN(\MC_ARK_ARC_1_2/temp2[158] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_5_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[152] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[158] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_5_2  ( .A(\MC_ARK_ARC_1_2/temp6[159] ), .B(
        \MC_ARK_ARC_1_2/temp5[159] ), .ZN(\RI1[3][159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_5_2  ( .A(\MC_ARK_ARC_1_2/temp3[159] ), .B(
        \MC_ARK_ARC_1_2/temp4[159] ), .ZN(\MC_ARK_ARC_1_2/temp6[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_5_2  ( .A(\MC_ARK_ARC_1_2/temp1[159] ), .B(
        \MC_ARK_ARC_1_2/temp2[159] ), .ZN(\MC_ARK_ARC_1_2/temp5[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_5_2  ( .A(\RI5[2][3] ), .B(n278), .ZN(
        \MC_ARK_ARC_1_2/temp4[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_5_2  ( .A(\RI5[2][69] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[33] ), .ZN(\MC_ARK_ARC_1_2/temp3[159] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_5_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[129] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_5_2  ( .A(\RI5[2][159] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[153] ), .ZN(\MC_ARK_ARC_1_2/temp1[159] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_5_1  ( .A(\MC_ARK_ARC_1_2/temp5[160] ), .B(
        \MC_ARK_ARC_1_2/temp6[160] ), .ZN(\RI1[3][160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_5_1  ( .A(\MC_ARK_ARC_1_2/temp3[160] ), .B(
        \MC_ARK_ARC_1_2/temp4[160] ), .ZN(\MC_ARK_ARC_1_2/temp6[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_5_1  ( .A(\MC_ARK_ARC_1_2/temp1[160] ), .B(
        \MC_ARK_ARC_1_2/temp2[160] ), .ZN(\MC_ARK_ARC_1_2/temp5[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_5_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .B(n317), .ZN(\MC_ARK_ARC_1_2/temp4[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_5_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[70] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_5_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_5_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[160] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_5_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[5] ), 
        .B(n355), .ZN(\MC_ARK_ARC_1_2/temp4[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_5_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .B(n1503), .ZN(\MC_ARK_ARC_1_2/temp3[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_5_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .B(n1665), .ZN(\MC_ARK_ARC_1_2/temp2[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_5_0  ( .A(n1635), .B(
        \MC_ARK_ARC_1_2/buf_datainput[155] ), .ZN(\MC_ARK_ARC_1_2/temp1[161] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_4_5  ( .A(\MC_ARK_ARC_1_2/temp5[162] ), .B(
        \MC_ARK_ARC_1_2/temp6[162] ), .ZN(\RI1[3][162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_4_5  ( .A(\MC_ARK_ARC_1_2/temp3[162] ), .B(
        \MC_ARK_ARC_1_2/temp4[162] ), .ZN(\MC_ARK_ARC_1_2/temp6[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_4_5  ( .A(\MC_ARK_ARC_1_2/temp2[162] ), .B(
        \MC_ARK_ARC_1_2/temp1[162] ), .ZN(\MC_ARK_ARC_1_2/temp5[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_4_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[6] ), 
        .B(n212), .ZN(\MC_ARK_ARC_1_2/temp4[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_4_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[72] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[36] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_4_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[132] ), 
        .B(\RI5[2][108] ), .ZN(\MC_ARK_ARC_1_2/temp2[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_4_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[156] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_4_4  ( .A(\MC_ARK_ARC_1_2/temp5[163] ), .B(
        \MC_ARK_ARC_1_2/temp6[163] ), .ZN(\RI1[3][163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_4_4  ( .A(\MC_ARK_ARC_1_2/temp3[163] ), .B(
        \MC_ARK_ARC_1_2/temp4[163] ), .ZN(\MC_ARK_ARC_1_2/temp6[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_4_4  ( .A(\MC_ARK_ARC_1_2/temp1[163] ), .B(
        \MC_ARK_ARC_1_2/temp2[163] ), .ZN(\MC_ARK_ARC_1_2/temp5[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_4_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .B(n471), .ZN(\MC_ARK_ARC_1_2/temp4[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_4_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[73] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[37] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_4_4  ( .A(\RI5[2][133] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[109] ), .ZN(\MC_ARK_ARC_1_2/temp2[163] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_4_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[163] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[157] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_4_3  ( .A(\MC_ARK_ARC_1_2/temp5[164] ), .B(
        \MC_ARK_ARC_1_2/temp6[164] ), .ZN(\RI1[3][164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_4_3  ( .A(\MC_ARK_ARC_1_2/temp3[164] ), .B(
        \MC_ARK_ARC_1_2/temp4[164] ), .ZN(\MC_ARK_ARC_1_2/temp6[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_4_3  ( .A(\MC_ARK_ARC_1_2/temp1[164] ), .B(
        \MC_ARK_ARC_1_2/temp2[164] ), .ZN(\MC_ARK_ARC_1_2/temp5[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_4_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[8] ), 
        .B(n290), .ZN(\MC_ARK_ARC_1_2/temp4[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_4_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[74] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_4_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[110] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_4_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[158] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_4_2  ( .A(\MC_ARK_ARC_1_2/temp5[165] ), .B(
        \MC_ARK_ARC_1_2/temp6[165] ), .ZN(\RI1[3][165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_4_2  ( .A(\MC_ARK_ARC_1_2/temp3[165] ), .B(
        \MC_ARK_ARC_1_2/temp4[165] ), .ZN(\MC_ARK_ARC_1_2/temp6[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_4_2  ( .A(\MC_ARK_ARC_1_2/temp1[165] ), .B(
        \MC_ARK_ARC_1_2/temp2[165] ), .ZN(\MC_ARK_ARC_1_2/temp5[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_4_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[9] ), 
        .B(n329), .ZN(\MC_ARK_ARC_1_2/temp4[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_4_2  ( .A(\RI5[2][39] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[75] ), .ZN(\MC_ARK_ARC_1_2/temp3[165] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_4_2  ( .A(n2099), .B(n1950), .ZN(
        \MC_ARK_ARC_1_2/temp2[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_4_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[165] ), 
        .B(\RI5[2][159] ), .ZN(\MC_ARK_ARC_1_2/temp1[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_4_1  ( .A(\MC_ARK_ARC_1_2/temp5[166] ), .B(
        \MC_ARK_ARC_1_2/temp6[166] ), .ZN(\RI1[3][166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_4_1  ( .A(\MC_ARK_ARC_1_2/temp3[166] ), .B(
        \MC_ARK_ARC_1_2/temp4[166] ), .ZN(\MC_ARK_ARC_1_2/temp6[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_4_1  ( .A(\MC_ARK_ARC_1_2/temp1[166] ), .B(
        \MC_ARK_ARC_1_2/temp2[166] ), .ZN(\MC_ARK_ARC_1_2/temp5[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_4_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[10] ), 
        .B(n468), .ZN(\MC_ARK_ARC_1_2/temp4[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_4_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[76] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_4_1  ( .A(n1932), .B(
        \MC_ARK_ARC_1_2/buf_datainput[112] ), .ZN(\MC_ARK_ARC_1_2/temp2[166] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_4_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[160] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_4_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[11] ), 
        .B(n225), .ZN(\MC_ARK_ARC_1_2/temp4[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_4_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[77] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[41] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_4_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[113] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[137] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_4_0  ( .A(n1629), .B(n1636), .ZN(
        \MC_ARK_ARC_1_2/temp1[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_3_5  ( .A(\MC_ARK_ARC_1_2/temp5[168] ), .B(
        \MC_ARK_ARC_1_2/temp6[168] ), .ZN(\RI1[3][168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_3_5  ( .A(\MC_ARK_ARC_1_2/temp3[168] ), .B(
        \MC_ARK_ARC_1_2/temp4[168] ), .ZN(\MC_ARK_ARC_1_2/temp6[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_3_5  ( .A(\MC_ARK_ARC_1_2/temp1[168] ), .B(
        \MC_ARK_ARC_1_2/temp2[168] ), .ZN(\MC_ARK_ARC_1_2/temp5[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_3_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[12] ), 
        .B(n263), .ZN(\MC_ARK_ARC_1_2/temp4[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_3_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[78] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[42] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_3_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[138] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[114] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_3_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[168] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[162] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_3_4  ( .A(\MC_ARK_ARC_1_2/temp5[169] ), .B(
        \MC_ARK_ARC_1_2/temp6[169] ), .ZN(\RI1[3][169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_3_4  ( .A(\MC_ARK_ARC_1_2/temp4[169] ), .B(
        \MC_ARK_ARC_1_2/temp3[169] ), .ZN(\MC_ARK_ARC_1_2/temp6[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_3_4  ( .A(\MC_ARK_ARC_1_2/temp1[169] ), .B(
        \MC_ARK_ARC_1_2/temp2[169] ), .ZN(\MC_ARK_ARC_1_2/temp5[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_3_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[13] ), 
        .B(n458), .ZN(\MC_ARK_ARC_1_2/temp4[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_3_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[79] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[43] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_3_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[139] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[115] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_3_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[169] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[163] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_3_3  ( .A(\MC_ARK_ARC_1_2/temp6[170] ), .B(
        \MC_ARK_ARC_1_2/temp5[170] ), .ZN(\RI1[3][170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_3_3  ( .A(\MC_ARK_ARC_1_2/temp4[170] ), .B(
        \MC_ARK_ARC_1_2/temp3[170] ), .ZN(\MC_ARK_ARC_1_2/temp6[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_3_3  ( .A(\MC_ARK_ARC_1_2/temp1[170] ), .B(
        \MC_ARK_ARC_1_2/temp2[170] ), .ZN(\MC_ARK_ARC_1_2/temp5[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_3_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[14] ), 
        .B(n407), .ZN(\MC_ARK_ARC_1_2/temp4[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_3_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[80] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[44] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_3_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[140] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[116] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_3_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .B(n2144), .ZN(\MC_ARK_ARC_1_2/temp1[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_3_2  ( .A(\MC_ARK_ARC_1_2/temp5[171] ), .B(
        \MC_ARK_ARC_1_2/temp6[171] ), .ZN(\RI1[3][171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_3_2  ( .A(\MC_ARK_ARC_1_2/temp3[171] ), .B(
        \MC_ARK_ARC_1_2/temp4[171] ), .ZN(\MC_ARK_ARC_1_2/temp6[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_3_2  ( .A(\MC_ARK_ARC_1_2/temp2[171] ), .B(
        \MC_ARK_ARC_1_2/temp1[171] ), .ZN(\MC_ARK_ARC_1_2/temp5[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_3_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[15] ), 
        .B(n198), .ZN(\MC_ARK_ARC_1_2/temp4[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_3_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[81] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[45] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_3_2  ( .A(n1951), .B(\RI5[2][117] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_3_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[165] ), 
        .B(\RI5[2][171] ), .ZN(\MC_ARK_ARC_1_2/temp1[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_3_1  ( .A(\MC_ARK_ARC_1_2/temp5[172] ), .B(
        \MC_ARK_ARC_1_2/temp6[172] ), .ZN(\RI1[3][172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_3_1  ( .A(\MC_ARK_ARC_1_2/temp3[172] ), .B(
        \MC_ARK_ARC_1_2/temp4[172] ), .ZN(\MC_ARK_ARC_1_2/temp6[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_3_1  ( .A(\MC_ARK_ARC_1_2/temp1[172] ), .B(
        \MC_ARK_ARC_1_2/temp2[172] ), .ZN(\MC_ARK_ARC_1_2/temp5[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_3_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[172] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_3_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[46] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[82] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_3_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[142] ), 
        .B(n1957), .ZN(\MC_ARK_ARC_1_2/temp2[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_3_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_3_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[17] ), 
        .B(n276), .ZN(\MC_ARK_ARC_1_2/temp4[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_3_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[83] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_3_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .B(n811), .ZN(\MC_ARK_ARC_1_2/temp2[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_3_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[167] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[173] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_2_5  ( .A(\MC_ARK_ARC_1_2/temp5[174] ), .B(
        \MC_ARK_ARC_1_2/temp6[174] ), .ZN(\RI1[3][174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_2_5  ( .A(\MC_ARK_ARC_1_2/temp3[174] ), .B(
        \MC_ARK_ARC_1_2/temp4[174] ), .ZN(\MC_ARK_ARC_1_2/temp6[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_2_5  ( .A(\MC_ARK_ARC_1_2/temp1[174] ), .B(
        \MC_ARK_ARC_1_2/temp2[174] ), .ZN(\MC_ARK_ARC_1_2/temp5[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_2_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[18] ), 
        .B(n505), .ZN(\MC_ARK_ARC_1_2/temp4[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_2_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[48] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_2_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[144] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[120] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_2_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[174] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[168] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_2_4  ( .A(\MC_ARK_ARC_1_2/temp2[175] ), .B(
        \MC_ARK_ARC_1_2/temp1[175] ), .ZN(\MC_ARK_ARC_1_2/temp5[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_2_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[19] ), 
        .B(n447), .ZN(\MC_ARK_ARC_1_2/temp4[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_2_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[85] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[49] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_2_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[145] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[121] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_2_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[175] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[169] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_2_3  ( .A(\MC_ARK_ARC_1_2/temp5[176] ), .B(
        \MC_ARK_ARC_1_2/temp6[176] ), .ZN(\RI1[3][176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_2_3  ( .A(\MC_ARK_ARC_1_2/temp3[176] ), .B(
        \MC_ARK_ARC_1_2/temp4[176] ), .ZN(\MC_ARK_ARC_1_2/temp6[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_2_3  ( .A(\MC_ARK_ARC_1_2/temp1[176] ), .B(
        \MC_ARK_ARC_1_2/temp2[176] ), .ZN(\MC_ARK_ARC_1_2/temp5[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_2_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[20] ), 
        .B(n405), .ZN(\MC_ARK_ARC_1_2/temp4[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_2_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[50] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[86] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_2_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[122] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_2_3  ( .A(n2144), .B(
        \MC_ARK_ARC_1_2/buf_datainput[176] ), .ZN(\MC_ARK_ARC_1_2/temp1[176] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_2_2  ( .A(\MC_ARK_ARC_1_2/temp5[177] ), .B(
        \MC_ARK_ARC_1_2/temp6[177] ), .ZN(\RI1[3][177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_2_2  ( .A(\MC_ARK_ARC_1_2/temp3[177] ), .B(
        \MC_ARK_ARC_1_2/temp4[177] ), .ZN(\MC_ARK_ARC_1_2/temp6[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_2_2  ( .A(\MC_ARK_ARC_1_2/temp2[177] ), .B(
        \MC_ARK_ARC_1_2/temp1[177] ), .ZN(\MC_ARK_ARC_1_2/temp5[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_2_2  ( .A(\RI5[2][21] ), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[177] ), .ZN(\MC_ARK_ARC_1_2/temp4[177] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_2_2  ( .A(\RI5[2][51] ), .B(\RI5[2][87] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_2_2  ( .A(\RI5[2][147] ), .B(\RI5[2][123] ), 
        .ZN(\MC_ARK_ARC_1_2/temp2[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_2_2  ( .A(\RI5[2][171] ), .B(\RI5[2][177] ), 
        .ZN(\MC_ARK_ARC_1_2/temp1[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_2_1  ( .A(\MC_ARK_ARC_1_2/temp5[178] ), .B(
        \MC_ARK_ARC_1_2/temp6[178] ), .ZN(\RI1[3][178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_2_1  ( .A(\MC_ARK_ARC_1_2/temp3[178] ), .B(
        \MC_ARK_ARC_1_2/temp4[178] ), .ZN(\MC_ARK_ARC_1_2/temp6[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_2_1  ( .A(\MC_ARK_ARC_1_2/temp1[178] ), .B(
        \MC_ARK_ARC_1_2/temp2[178] ), .ZN(\MC_ARK_ARC_1_2/temp5[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_2_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .B(n288), .ZN(\MC_ARK_ARC_1_2/temp4[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_2_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[52] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_2_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[124] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_2_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[178] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_2_0  ( .A(\MC_ARK_ARC_1_2/temp5[179] ), .B(
        \MC_ARK_ARC_1_2/temp6[179] ), .ZN(\RI1[3][179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_2_0  ( .A(\MC_ARK_ARC_1_2/temp3[179] ), .B(
        \MC_ARK_ARC_1_2/temp4[179] ), .ZN(\MC_ARK_ARC_1_2/temp6[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_2_0  ( .A(\MC_ARK_ARC_1_2/temp2[179] ), .B(
        \MC_ARK_ARC_1_2/temp1[179] ), .ZN(\MC_ARK_ARC_1_2/temp5[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_2_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[23] ), 
        .B(n327), .ZN(\MC_ARK_ARC_1_2/temp4[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_2_0  ( .A(n1501), .B(n781), .ZN(
        \MC_ARK_ARC_1_2/temp3[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_2_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .B(n816), .ZN(\MC_ARK_ARC_1_2/temp2[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_2_0  ( .A(n827), .B(n803), .ZN(
        \MC_ARK_ARC_1_2/temp1[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_1_5  ( .A(\MC_ARK_ARC_1_2/temp5[180] ), .B(
        \MC_ARK_ARC_1_2/temp6[180] ), .ZN(\RI1[3][180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_1_5  ( .A(\MC_ARK_ARC_1_2/temp3[180] ), .B(
        \MC_ARK_ARC_1_2/temp4[180] ), .ZN(\MC_ARK_ARC_1_2/temp6[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_1_5  ( .A(\MC_ARK_ARC_1_2/temp1[180] ), .B(
        \MC_ARK_ARC_1_2/temp2[180] ), .ZN(\MC_ARK_ARC_1_2/temp5[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_1_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .B(n503), .ZN(\MC_ARK_ARC_1_2/temp4[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_1_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[90] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[54] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_1_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[150] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[126] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_1_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[180] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[174] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_1_4  ( .A(\MC_ARK_ARC_1_2/temp5[181] ), .B(
        \MC_ARK_ARC_1_2/temp6[181] ), .ZN(\RI1[3][181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_1_4  ( .A(\MC_ARK_ARC_1_2/temp4[181] ), .B(
        \MC_ARK_ARC_1_2/temp3[181] ), .ZN(\MC_ARK_ARC_1_2/temp6[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_1_4  ( .A(\MC_ARK_ARC_1_2/temp1[181] ), .B(
        \MC_ARK_ARC_1_2/temp2[181] ), .ZN(\MC_ARK_ARC_1_2/temp5[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_1_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[25] ), 
        .B(n223), .ZN(\MC_ARK_ARC_1_2/temp4[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_1_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[91] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[55] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_1_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[127] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_1_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[181] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[175] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_1_3  ( .A(\MC_ARK_ARC_1_2/temp5[182] ), .B(
        \MC_ARK_ARC_1_2/temp6[182] ), .ZN(\RI1[3][182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_1_3  ( .A(\MC_ARK_ARC_1_2/temp3[182] ), .B(
        \MC_ARK_ARC_1_2/temp4[182] ), .ZN(\MC_ARK_ARC_1_2/temp6[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_1_3  ( .A(\MC_ARK_ARC_1_2/temp1[182] ), .B(
        \MC_ARK_ARC_1_2/temp2[182] ), .ZN(\MC_ARK_ARC_1_2/temp5[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_1_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[26] ), 
        .B(n402), .ZN(\MC_ARK_ARC_1_2/temp4[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_1_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[92] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[56] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_1_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[152] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[128] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_1_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[176] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_1_2  ( .A(\MC_ARK_ARC_1_2/temp5[183] ), .B(
        \MC_ARK_ARC_1_2/temp6[183] ), .ZN(\RI1[3][183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_1_2  ( .A(\MC_ARK_ARC_1_2/temp3[183] ), .B(
        \MC_ARK_ARC_1_2/temp4[183] ), .ZN(\MC_ARK_ARC_1_2/temp6[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_1_2  ( .A(\MC_ARK_ARC_1_2/temp1[183] ), .B(
        \MC_ARK_ARC_1_2/temp2[183] ), .ZN(\MC_ARK_ARC_1_2/temp5[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_1_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[27] ), 
        .B(n300), .ZN(\MC_ARK_ARC_1_2/temp4[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_1_2  ( .A(\RI5[2][93] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[57] ), .ZN(\MC_ARK_ARC_1_2/temp3[183] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_1_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[153] ), 
        .B(n815), .ZN(\MC_ARK_ARC_1_2/temp2[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_1_2  ( .A(\RI5[2][177] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[183] ), .ZN(\MC_ARK_ARC_1_2/temp1[183] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_1_1  ( .A(\MC_ARK_ARC_1_2/temp5[184] ), .B(
        \MC_ARK_ARC_1_2/temp6[184] ), .ZN(\RI1[3][184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_1_1  ( .A(\MC_ARK_ARC_1_2/temp3[184] ), .B(
        \MC_ARK_ARC_1_2/temp4[184] ), .ZN(\MC_ARK_ARC_1_2/temp6[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_1_1  ( .A(\MC_ARK_ARC_1_2/temp1[184] ), .B(
        \MC_ARK_ARC_1_2/temp2[184] ), .ZN(\MC_ARK_ARC_1_2/temp5[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_1_1  ( .A(n2142), .B(
        \MC_ARK_ARC_1_2/buf_keyinput[184] ), .ZN(\MC_ARK_ARC_1_2/temp4[184] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_1_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[94] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[58] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_1_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[154] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[130] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_1_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[184] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[178] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_1_0  ( .A(\MC_ARK_ARC_1_2/temp3[185] ), .B(
        \MC_ARK_ARC_1_2/temp4[185] ), .ZN(\MC_ARK_ARC_1_2/temp6[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_1_0  ( .A(\MC_ARK_ARC_1_2/temp2[185] ), .B(
        \MC_ARK_ARC_1_2/temp1[185] ), .ZN(\MC_ARK_ARC_1_2/temp5[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_1_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .B(n498), .ZN(\MC_ARK_ARC_1_2/temp4[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_1_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .B(n792), .ZN(\MC_ARK_ARC_1_2/temp3[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_1_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .B(n824), .ZN(\MC_ARK_ARC_1_2/temp2[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_1_0  ( .A(n802), .B(n823), .ZN(
        \MC_ARK_ARC_1_2/temp1[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_0_5  ( .A(\MC_ARK_ARC_1_2/temp5[186] ), .B(
        \MC_ARK_ARC_1_2/temp6[186] ), .ZN(\RI1[3][186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_0_5  ( .A(\MC_ARK_ARC_1_2/temp3[186] ), .B(
        \MC_ARK_ARC_1_2/temp4[186] ), .ZN(\MC_ARK_ARC_1_2/temp6[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_0_5  ( .A(\MC_ARK_ARC_1_2/temp1[186] ), .B(
        \MC_ARK_ARC_1_2/temp2[186] ), .ZN(\MC_ARK_ARC_1_2/temp5[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_0_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[30] ), 
        .B(n507), .ZN(\MC_ARK_ARC_1_2/temp4[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_0_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[96] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[60] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_0_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[132] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_0_5  ( .A(\MC_ARK_ARC_1_2/buf_datainput[186] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[180] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_0_4  ( .A(\MC_ARK_ARC_1_2/temp5[187] ), .B(
        \MC_ARK_ARC_1_2/temp6[187] ), .ZN(\RI1[3][187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_0_4  ( .A(\MC_ARK_ARC_1_2/temp3[187] ), .B(
        \MC_ARK_ARC_1_2/temp4[187] ), .ZN(\MC_ARK_ARC_1_2/temp6[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_0_4  ( .A(\MC_ARK_ARC_1_2/temp1[187] ), .B(
        \MC_ARK_ARC_1_2/temp2[187] ), .ZN(\MC_ARK_ARC_1_2/temp5[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_0_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[31] ), 
        .B(n446), .ZN(\MC_ARK_ARC_1_2/temp4[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_0_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[97] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[61] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_0_4  ( .A(\MC_ARK_ARC_1_2/buf_datainput[157] ), 
        .B(\RI5[2][133] ), .ZN(\MC_ARK_ARC_1_2/temp2[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_0_4  ( .A(\RI5[2][187] ), .B(
        \MC_ARK_ARC_1_2/buf_datainput[181] ), .ZN(\MC_ARK_ARC_1_2/temp1[187] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_0_3  ( .A(\MC_ARK_ARC_1_2/temp5[188] ), .B(
        \MC_ARK_ARC_1_2/temp6[188] ), .ZN(\RI1[3][188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_0_3  ( .A(\MC_ARK_ARC_1_2/temp3[188] ), .B(
        \MC_ARK_ARC_1_2/temp4[188] ), .ZN(\MC_ARK_ARC_1_2/temp6[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_0_3  ( .A(\MC_ARK_ARC_1_2/temp1[188] ), .B(
        \MC_ARK_ARC_1_2/temp2[188] ), .ZN(\MC_ARK_ARC_1_2/temp5[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_0_3  ( .A(n1511), .B(n404), .ZN(
        \MC_ARK_ARC_1_2/temp4[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_0_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[62] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[98] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_0_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[134] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[158] ), .ZN(
        \MC_ARK_ARC_1_2/temp2[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_0_3  ( .A(\MC_ARK_ARC_1_2/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[188] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_0_2  ( .A(\MC_ARK_ARC_1_2/temp6[189] ), .B(
        \MC_ARK_ARC_1_2/temp5[189] ), .ZN(\RI1[3][189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_0_2  ( .A(\MC_ARK_ARC_1_2/temp3[189] ), .B(
        \MC_ARK_ARC_1_2/temp4[189] ), .ZN(\MC_ARK_ARC_1_2/temp6[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_0_2  ( .A(\MC_ARK_ARC_1_2/temp2[189] ), .B(
        \MC_ARK_ARC_1_2/temp1[189] ), .ZN(\MC_ARK_ARC_1_2/temp5[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_0_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[33] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[176] ), .ZN(
        \MC_ARK_ARC_1_2/temp4[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_0_2  ( .A(\RI5[2][99] ), .B(n2101), .ZN(
        \MC_ARK_ARC_1_2/temp3[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_0_2  ( .A(\RI5[2][159] ), .B(n2098), .ZN(
        \MC_ARK_ARC_1_2/temp2[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_0_2  ( .A(\MC_ARK_ARC_1_2/buf_datainput[189] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[183] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X7_0_1  ( .A(\MC_ARK_ARC_1_2/temp5[190] ), .B(
        \MC_ARK_ARC_1_2/temp6[190] ), .ZN(\RI1[3][190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X6_0_1  ( .A(\MC_ARK_ARC_1_2/temp3[190] ), .B(
        \MC_ARK_ARC_1_2/temp4[190] ), .ZN(\MC_ARK_ARC_1_2/temp6[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X5_0_1  ( .A(\MC_ARK_ARC_1_2/temp1[190] ), .B(
        \MC_ARK_ARC_1_2/temp2[190] ), .ZN(\MC_ARK_ARC_1_2/temp5[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_0_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .B(n208), .ZN(\MC_ARK_ARC_1_2/temp4[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_0_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[64] ), .ZN(
        \MC_ARK_ARC_1_2/temp3[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_0_1  ( .A(n1933), .B(
        \MC_ARK_ARC_1_2/buf_datainput[160] ), .ZN(\MC_ARK_ARC_1_2/temp2[190] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_0_1  ( .A(\MC_ARK_ARC_1_2/buf_datainput[184] ), 
        .B(\MC_ARK_ARC_1_2/buf_datainput[190] ), .ZN(
        \MC_ARK_ARC_1_2/temp1[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X4_0_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .B(n247), .ZN(\MC_ARK_ARC_1_2/temp4[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X3_0_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .B(n2127), .ZN(\MC_ARK_ARC_1_2/temp3[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X2_0_0  ( .A(\MC_ARK_ARC_1_2/buf_datainput[137] ), 
        .B(n1635), .ZN(\MC_ARK_ARC_1_2/temp2[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_2/X1_0_0  ( .A(n822), .B(n829), .ZN(
        \MC_ARK_ARC_1_2/temp1[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_31_5  ( .A(\MC_ARK_ARC_1_3/temp5[0] ), .B(
        \MC_ARK_ARC_1_3/temp6[0] ), .ZN(\RI1[4][0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_31_5  ( .A(\MC_ARK_ARC_1_3/temp3[0] ), .B(
        \MC_ARK_ARC_1_3/temp4[0] ), .ZN(\MC_ARK_ARC_1_3/temp6[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_31_5  ( .A(\MC_ARK_ARC_1_3/temp1[0] ), .B(
        \MC_ARK_ARC_1_3/temp2[0] ), .ZN(\MC_ARK_ARC_1_3/temp5[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_31_5  ( .A(\RI5[3][36] ), .B(n512), .ZN(
        \MC_ARK_ARC_1_3/temp4[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_31_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .B(\RI5[3][66] ), .ZN(\MC_ARK_ARC_1_3/temp3[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_31_5  ( .A(\RI5[3][162] ), .B(n818), .ZN(
        \MC_ARK_ARC_1_3/temp2[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_31_5  ( .A(\RI5[3][0] ), .B(\RI5[3][186] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[0] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_31_4  ( .A(\MC_ARK_ARC_1_3/temp5[1] ), .B(
        \MC_ARK_ARC_1_3/temp6[1] ), .ZN(\RI1[4][1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_31_4  ( .A(\MC_ARK_ARC_1_3/temp3[1] ), .B(
        \MC_ARK_ARC_1_3/temp4[1] ), .ZN(\MC_ARK_ARC_1_3/temp6[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_31_4  ( .A(\MC_ARK_ARC_1_3/temp1[1] ), .B(
        \MC_ARK_ARC_1_3/temp2[1] ), .ZN(\MC_ARK_ARC_1_3/temp5[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_31_4  ( .A(\RI5[3][37] ), .B(n206), .ZN(
        \MC_ARK_ARC_1_3/temp4[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_31_4  ( .A(\RI5[3][103] ), .B(\RI5[3][67] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_31_4  ( .A(\RI5[3][163] ), .B(\RI5[3][139] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_31_4  ( .A(\RI5[3][1] ), .B(\RI5[3][187] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[1] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_31_3  ( .A(\MC_ARK_ARC_1_3/temp5[2] ), .B(
        \MC_ARK_ARC_1_3/temp6[2] ), .ZN(\RI1[4][2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_31_3  ( .A(\MC_ARK_ARC_1_3/temp4[2] ), .B(
        \MC_ARK_ARC_1_3/temp3[2] ), .ZN(\MC_ARK_ARC_1_3/temp6[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_31_3  ( .A(\MC_ARK_ARC_1_3/temp2[2] ), .B(
        \MC_ARK_ARC_1_3/temp1[2] ), .ZN(\MC_ARK_ARC_1_3/temp5[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_31_3  ( .A(\RI5[3][38] ), .B(n297), .ZN(
        \MC_ARK_ARC_1_3/temp4[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_31_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[104] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_3/temp3[2] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_31_3  ( .A(n1627), .B(\RI5[3][140] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_31_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[2] ), 
        .B(\RI5[3][188] ), .ZN(\MC_ARK_ARC_1_3/temp1[2] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_31_2  ( .A(\MC_ARK_ARC_1_3/temp6[3] ), .B(
        \MC_ARK_ARC_1_3/temp5[3] ), .ZN(\RI1[4][3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_31_2  ( .A(\MC_ARK_ARC_1_3/temp3[3] ), .B(
        \MC_ARK_ARC_1_3/temp4[3] ), .ZN(\MC_ARK_ARC_1_3/temp6[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_31_2  ( .A(\MC_ARK_ARC_1_3/temp1[3] ), .B(
        \MC_ARK_ARC_1_3/temp2[3] ), .ZN(\MC_ARK_ARC_1_3/temp5[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_31_2  ( .A(\RI5[3][39] ), .B(n401), .ZN(
        \MC_ARK_ARC_1_3/temp4[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_31_2  ( .A(\RI5[3][105] ), .B(\RI5[3][69] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_31_2  ( .A(\RI5[3][165] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[141] ), .ZN(\MC_ARK_ARC_1_3/temp2[3] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_31_2  ( .A(\RI5[3][3] ), .B(\RI5[3][189] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[3] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_31_1  ( .A(\MC_ARK_ARC_1_3/temp5[4] ), .B(
        \MC_ARK_ARC_1_3/temp6[4] ), .ZN(\RI1[4][4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_31_1  ( .A(\MC_ARK_ARC_1_3/temp3[4] ), .B(
        \MC_ARK_ARC_1_3/temp4[4] ), .ZN(\MC_ARK_ARC_1_3/temp6[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_31_1  ( .A(\MC_ARK_ARC_1_3/temp1[4] ), .B(
        \MC_ARK_ARC_1_3/temp2[4] ), .ZN(\MC_ARK_ARC_1_3/temp5[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_31_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[40] ), 
        .B(n295), .ZN(\MC_ARK_ARC_1_3/temp4[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_31_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[106] ), .ZN(\MC_ARK_ARC_1_3/temp3[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_31_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[166] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[142] ), .ZN(\MC_ARK_ARC_1_3/temp2[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_31_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[4] ), 
        .B(\RI5[3][190] ), .ZN(\MC_ARK_ARC_1_3/temp1[4] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_31_0  ( .A(n2111), .B(
        \MC_ARK_ARC_1_0/buf_keyinput[80] ), .ZN(\MC_ARK_ARC_1_3/temp4[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_31_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .B(n2108), .ZN(\MC_ARK_ARC_1_3/temp3[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_31_0  ( .A(n1661), .B(n1947), .ZN(
        \MC_ARK_ARC_1_3/temp2[5] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_31_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[191] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[5] ), .ZN(\MC_ARK_ARC_1_3/temp1[5] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_30_5  ( .A(\MC_ARK_ARC_1_3/temp5[6] ), .B(
        \MC_ARK_ARC_1_3/temp6[6] ), .ZN(\RI1[4][6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_30_5  ( .A(\MC_ARK_ARC_1_3/temp3[6] ), .B(
        \MC_ARK_ARC_1_3/temp4[6] ), .ZN(\MC_ARK_ARC_1_3/temp6[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_30_5  ( .A(\MC_ARK_ARC_1_3/temp1[6] ), .B(
        \MC_ARK_ARC_1_3/temp2[6] ), .ZN(\MC_ARK_ARC_1_3/temp5[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_30_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[42] ), 
        .B(n438), .ZN(\MC_ARK_ARC_1_3/temp4[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_30_5  ( .A(\RI5[3][108] ), .B(\RI5[3][72] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_30_5  ( .A(\RI5[3][168] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[144] ), .ZN(\MC_ARK_ARC_1_3/temp2[6] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_30_5  ( .A(\RI5[3][6] ), .B(\RI5[3][0] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[6] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_30_4  ( .A(\MC_ARK_ARC_1_3/temp5[7] ), .B(
        \MC_ARK_ARC_1_3/temp6[7] ), .ZN(\RI1[4][7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_30_4  ( .A(\MC_ARK_ARC_1_3/temp3[7] ), .B(
        \MC_ARK_ARC_1_3/temp4[7] ), .ZN(\MC_ARK_ARC_1_3/temp6[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_30_4  ( .A(\MC_ARK_ARC_1_3/temp1[7] ), .B(
        \MC_ARK_ARC_1_3/temp2[7] ), .ZN(\MC_ARK_ARC_1_3/temp5[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_30_4  ( .A(\RI5[3][43] ), .B(n200), .ZN(
        \MC_ARK_ARC_1_3/temp4[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_30_4  ( .A(\RI5[3][109] ), .B(\RI5[3][73] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_30_4  ( .A(\RI5[3][169] ), .B(\RI5[3][145] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_30_4  ( .A(\RI5[3][7] ), .B(\RI5[3][1] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[7] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_30_3  ( .A(\MC_ARK_ARC_1_3/temp5[8] ), .B(
        \MC_ARK_ARC_1_3/temp6[8] ), .ZN(\RI1[4][8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_30_3  ( .A(\MC_ARK_ARC_1_3/temp3[8] ), .B(
        \MC_ARK_ARC_1_3/temp4[8] ), .ZN(\MC_ARK_ARC_1_3/temp6[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_30_3  ( .A(\MC_ARK_ARC_1_3/temp2[8] ), .B(
        \MC_ARK_ARC_1_3/temp1[8] ), .ZN(\MC_ARK_ARC_1_3/temp5[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_30_3  ( .A(\RI5[3][44] ), .B(n490), .ZN(
        \MC_ARK_ARC_1_3/temp4[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_30_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[110] ), .ZN(\MC_ARK_ARC_1_3/temp3[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_30_3  ( .A(\RI5[3][170] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[146] ), .ZN(\MC_ARK_ARC_1_3/temp2[8] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_30_3  ( .A(\RI5[3][8] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_3/temp1[8] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_30_2  ( .A(\MC_ARK_ARC_1_3/temp5[9] ), .B(
        \MC_ARK_ARC_1_3/temp6[9] ), .ZN(\RI1[4][9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_30_2  ( .A(\MC_ARK_ARC_1_3/temp3[9] ), .B(
        \MC_ARK_ARC_1_3/temp4[9] ), .ZN(\MC_ARK_ARC_1_3/temp6[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_30_2  ( .A(\MC_ARK_ARC_1_3/temp1[9] ), .B(
        \MC_ARK_ARC_1_3/temp2[9] ), .ZN(\MC_ARK_ARC_1_3/temp5[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_30_2  ( .A(\RI5[3][45] ), .B(n199), .ZN(
        \MC_ARK_ARC_1_3/temp4[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_30_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[111] ), 
        .B(\RI5[3][75] ), .ZN(\MC_ARK_ARC_1_3/temp3[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_30_2  ( .A(\RI5[3][171] ), .B(\RI5[3][147] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_30_2  ( .A(\RI5[3][9] ), .B(\RI5[3][3] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[9] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_30_1  ( .A(\MC_ARK_ARC_1_3/temp5[10] ), .B(
        \MC_ARK_ARC_1_3/temp6[10] ), .ZN(\RI1[4][10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_30_1  ( .A(\MC_ARK_ARC_1_3/temp3[10] ), .B(
        \MC_ARK_ARC_1_3/temp4[10] ), .ZN(\MC_ARK_ARC_1_3/temp6[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_30_1  ( .A(\MC_ARK_ARC_1_3/temp1[10] ), .B(
        \MC_ARK_ARC_1_3/temp2[10] ), .ZN(\MC_ARK_ARC_1_3/temp5[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_30_1  ( .A(\RI5[3][46] ), .B(n289), .ZN(
        \MC_ARK_ARC_1_3/temp4[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_30_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[76] ), .ZN(\MC_ARK_ARC_1_3/temp3[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_30_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[172] ), 
        .B(n1510), .ZN(\MC_ARK_ARC_1_3/temp2[10] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_30_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_3/temp1[10] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_30_0  ( .A(\MC_ARK_ARC_1_3/temp5[11] ), .B(
        \MC_ARK_ARC_1_3/temp6[11] ), .ZN(\RI1[4][11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_30_0  ( .A(\MC_ARK_ARC_1_3/temp3[11] ), .B(
        \MC_ARK_ARC_1_3/temp4[11] ), .ZN(\MC_ARK_ARC_1_3/temp6[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_30_0  ( .A(\MC_ARK_ARC_1_3/temp1[11] ), .B(
        \MC_ARK_ARC_1_3/temp2[11] ), .ZN(\MC_ARK_ARC_1_3/temp5[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_30_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[77] ), 
        .B(n797), .ZN(\MC_ARK_ARC_1_3/temp3[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_30_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[173] ), 
        .B(n849), .ZN(\MC_ARK_ARC_1_3/temp2[11] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_30_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[11] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[5] ), .ZN(\MC_ARK_ARC_1_3/temp1[11] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_29_5  ( .A(\MC_ARK_ARC_1_3/temp6[12] ), .B(
        \MC_ARK_ARC_1_3/temp5[12] ), .ZN(\RI1[4][12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_29_5  ( .A(\MC_ARK_ARC_1_3/temp3[12] ), .B(
        \MC_ARK_ARC_1_3/temp4[12] ), .ZN(\MC_ARK_ARC_1_3/temp6[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_29_5  ( .A(\MC_ARK_ARC_1_3/temp1[12] ), .B(
        \MC_ARK_ARC_1_3/temp2[12] ), .ZN(\MC_ARK_ARC_1_3/temp5[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_29_5  ( .A(\RI5[3][48] ), .B(n287), .ZN(
        \MC_ARK_ARC_1_3/temp4[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_29_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[114] ), 
        .B(\RI5[3][78] ), .ZN(\MC_ARK_ARC_1_3/temp3[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_29_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .B(\RI5[3][150] ), .ZN(\MC_ARK_ARC_1_3/temp2[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_29_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[12] ), 
        .B(\RI5[3][6] ), .ZN(\MC_ARK_ARC_1_3/temp1[12] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_29_4  ( .A(\MC_ARK_ARC_1_3/temp5[13] ), .B(
        \MC_ARK_ARC_1_3/temp6[13] ), .ZN(\RI1[4][13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_29_4  ( .A(\MC_ARK_ARC_1_3/temp3[13] ), .B(
        \MC_ARK_ARC_1_3/temp4[13] ), .ZN(\MC_ARK_ARC_1_3/temp6[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_29_4  ( .A(\MC_ARK_ARC_1_3/temp1[13] ), .B(
        \MC_ARK_ARC_1_3/temp2[13] ), .ZN(\MC_ARK_ARC_1_3/temp5[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_29_4  ( .A(\RI5[3][49] ), .B(n195), .ZN(
        \MC_ARK_ARC_1_3/temp4[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_29_4  ( .A(\RI5[3][115] ), .B(\RI5[3][79] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_29_4  ( .A(\RI5[3][175] ), .B(\RI5[3][151] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_29_4  ( .A(\RI5[3][13] ), .B(\RI5[3][7] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[13] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_29_3  ( .A(\MC_ARK_ARC_1_3/temp5[14] ), .B(
        \MC_ARK_ARC_1_3/temp6[14] ), .ZN(\RI1[4][14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_29_3  ( .A(\MC_ARK_ARC_1_3/temp3[14] ), .B(
        \MC_ARK_ARC_1_3/temp4[14] ), .ZN(\MC_ARK_ARC_1_3/temp6[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_29_3  ( .A(\MC_ARK_ARC_1_3/temp1[14] ), .B(
        \MC_ARK_ARC_1_3/temp2[14] ), .ZN(\MC_ARK_ARC_1_3/temp5[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_29_3  ( .A(\RI5[3][50] ), .B(n285), .ZN(
        \MC_ARK_ARC_1_3/temp4[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_29_3  ( .A(\RI5[3][80] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[116] ), .ZN(\MC_ARK_ARC_1_3/temp3[14] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_29_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .B(\RI5[3][152] ), .ZN(\MC_ARK_ARC_1_3/temp2[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_29_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .B(\RI5[3][8] ), .ZN(\MC_ARK_ARC_1_3/temp1[14] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_29_2  ( .A(\MC_ARK_ARC_1_3/temp5[15] ), .B(
        \MC_ARK_ARC_1_3/temp6[15] ), .ZN(\RI1[4][15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_29_2  ( .A(\MC_ARK_ARC_1_3/temp3[15] ), .B(
        \MC_ARK_ARC_1_3/temp4[15] ), .ZN(\MC_ARK_ARC_1_3/temp6[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_29_2  ( .A(\MC_ARK_ARC_1_3/temp1[15] ), .B(
        \MC_ARK_ARC_1_3/temp2[15] ), .ZN(\MC_ARK_ARC_1_3/temp5[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_29_2  ( .A(\RI5[3][51] ), .B(n406), .ZN(
        \MC_ARK_ARC_1_3/temp4[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_29_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[117] ), 
        .B(\RI5[3][81] ), .ZN(\MC_ARK_ARC_1_3/temp3[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_29_2  ( .A(\RI5[3][177] ), .B(\RI5[3][153] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_29_2  ( .A(\RI5[3][15] ), .B(\RI5[3][9] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[15] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_29_1  ( .A(\MC_ARK_ARC_1_3/temp3[16] ), .B(
        \MC_ARK_ARC_1_3/temp4[16] ), .ZN(\MC_ARK_ARC_1_3/temp6[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_29_1  ( .A(\MC_ARK_ARC_1_3/temp1[16] ), .B(
        \MC_ARK_ARC_1_3/temp2[16] ), .ZN(\MC_ARK_ARC_1_3/temp5[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_29_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[52] ), 
        .B(n424), .ZN(\MC_ARK_ARC_1_3/temp4[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_29_1  ( .A(\RI5[3][118] ), .B(\RI5[3][82] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_29_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[154] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_29_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_3/temp1[16] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_29_0  ( .A(\MC_ARK_ARC_1_3/temp6[17] ), .B(
        \MC_ARK_ARC_1_3/temp5[17] ), .ZN(\RI1[4][17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_29_0  ( .A(\MC_ARK_ARC_1_3/temp3[17] ), .B(
        \MC_ARK_ARC_1_3/temp4[17] ), .ZN(\MC_ARK_ARC_1_3/temp6[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_29_0  ( .A(\MC_ARK_ARC_1_3/temp2[17] ), .B(
        \MC_ARK_ARC_1_3/temp1[17] ), .ZN(\MC_ARK_ARC_1_3/temp5[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_29_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .B(n373), .ZN(\MC_ARK_ARC_1_3/temp4[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_29_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[83] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[119] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_29_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .B(n2121), .ZN(\MC_ARK_ARC_1_3/temp2[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_29_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[11] ), .ZN(\MC_ARK_ARC_1_3/temp1[17] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_28_5  ( .A(\MC_ARK_ARC_1_3/temp5[18] ), .B(
        \MC_ARK_ARC_1_3/temp6[18] ), .ZN(\RI1[4][18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_28_5  ( .A(\MC_ARK_ARC_1_3/temp3[18] ), .B(
        \MC_ARK_ARC_1_3/temp4[18] ), .ZN(\MC_ARK_ARC_1_3/temp6[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_28_5  ( .A(\MC_ARK_ARC_1_3/temp1[18] ), .B(
        \MC_ARK_ARC_1_3/temp2[18] ), .ZN(\MC_ARK_ARC_1_3/temp5[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_28_5  ( .A(\RI5[3][54] ), .B(n282), .ZN(
        \MC_ARK_ARC_1_3/temp4[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_28_5  ( .A(\RI5[3][120] ), .B(\RI5[3][84] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_28_5  ( .A(\RI5[3][180] ), .B(\RI5[3][156] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[18] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_28_5  ( .A(\RI5[3][18] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_3/temp1[18] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_28_4  ( .A(\MC_ARK_ARC_1_3/temp5[19] ), .B(
        \MC_ARK_ARC_1_3/temp6[19] ), .ZN(\RI1[4][19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_28_4  ( .A(\MC_ARK_ARC_1_3/temp3[19] ), .B(
        \MC_ARK_ARC_1_3/temp4[19] ), .ZN(\MC_ARK_ARC_1_3/temp6[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_28_4  ( .A(\MC_ARK_ARC_1_3/temp1[19] ), .B(
        \MC_ARK_ARC_1_3/temp2[19] ), .ZN(\MC_ARK_ARC_1_3/temp5[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_28_4  ( .A(\RI5[3][55] ), .B(n473), .ZN(
        \MC_ARK_ARC_1_3/temp4[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_28_4  ( .A(\RI5[3][121] ), .B(\RI5[3][85] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_28_4  ( .A(\RI5[3][181] ), .B(\RI5[3][157] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_28_4  ( .A(\RI5[3][19] ), .B(\RI5[3][13] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[19] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_28_3  ( .A(\MC_ARK_ARC_1_3/temp5[20] ), .B(
        \MC_ARK_ARC_1_3/temp6[20] ), .ZN(\RI1[4][20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_28_3  ( .A(\MC_ARK_ARC_1_3/temp3[20] ), .B(
        \MC_ARK_ARC_1_3/temp4[20] ), .ZN(\MC_ARK_ARC_1_3/temp6[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_28_3  ( .A(\MC_ARK_ARC_1_3/temp1[20] ), .B(
        \MC_ARK_ARC_1_3/temp2[20] ), .ZN(\MC_ARK_ARC_1_3/temp5[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_28_3  ( .A(\RI5[3][56] ), .B(n463), .ZN(
        \MC_ARK_ARC_1_3/temp4[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_28_3  ( .A(n1930), .B(\RI5[3][86] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_28_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .B(n1955), .ZN(\MC_ARK_ARC_1_3/temp2[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_28_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_3/temp1[20] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_28_2  ( .A(\MC_ARK_ARC_1_3/temp5[21] ), .B(
        \MC_ARK_ARC_1_3/temp6[21] ), .ZN(\RI1[4][21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_28_2  ( .A(\MC_ARK_ARC_1_3/temp3[21] ), .B(
        \MC_ARK_ARC_1_3/temp4[21] ), .ZN(\MC_ARK_ARC_1_3/temp6[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_28_2  ( .A(\MC_ARK_ARC_1_3/temp1[21] ), .B(
        \MC_ARK_ARC_1_3/temp2[21] ), .ZN(\MC_ARK_ARC_1_3/temp5[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_28_2  ( .A(\RI5[3][57] ), .B(n369), .ZN(
        \MC_ARK_ARC_1_3/temp4[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_28_2  ( .A(\RI5[3][123] ), .B(\RI5[3][87] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_28_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[183] ), 
        .B(\RI5[3][159] ), .ZN(\MC_ARK_ARC_1_3/temp2[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_28_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .B(\RI5[3][15] ), .ZN(\MC_ARK_ARC_1_3/temp1[21] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_28_1  ( .A(\MC_ARK_ARC_1_3/temp5[22] ), .B(
        \MC_ARK_ARC_1_3/temp6[22] ), .ZN(\RI1[4][22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_28_1  ( .A(\MC_ARK_ARC_1_3/temp3[22] ), .B(
        \MC_ARK_ARC_1_3/temp4[22] ), .ZN(\MC_ARK_ARC_1_3/temp6[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_28_1  ( .A(\MC_ARK_ARC_1_3/temp2[22] ), .B(
        \MC_ARK_ARC_1_3/temp1[22] ), .ZN(\MC_ARK_ARC_1_3/temp5[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_28_1  ( .A(\RI5[3][58] ), .B(Key[102]), .ZN(
        \MC_ARK_ARC_1_3/temp4[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_28_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_3/temp3[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_28_1  ( .A(\RI5[3][184] ), .B(\RI5[3][160] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_28_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_3/temp1[22] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_28_0  ( .A(\MC_ARK_ARC_1_3/temp5[23] ), .B(
        \MC_ARK_ARC_1_3/temp6[23] ), .ZN(\RI1[4][23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_28_0  ( .A(\MC_ARK_ARC_1_3/temp3[23] ), .B(
        \MC_ARK_ARC_1_3/temp4[23] ), .ZN(\MC_ARK_ARC_1_3/temp6[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_28_0  ( .A(\MC_ARK_ARC_1_3/temp2[23] ), .B(
        \MC_ARK_ARC_1_3/temp1[23] ), .ZN(\MC_ARK_ARC_1_3/temp5[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_28_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[59] ), 
        .B(n468), .ZN(\MC_ARK_ARC_1_3/temp4[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_28_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[89] ), 
        .B(n521), .ZN(\MC_ARK_ARC_1_3/temp3[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_28_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[161] ), 
        .B(n839), .ZN(\MC_ARK_ARC_1_3/temp2[23] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_28_0  ( .A(n1653), .B(
        \MC_ARK_ARC_1_3/buf_datainput[17] ), .ZN(\MC_ARK_ARC_1_3/temp1[23] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_27_5  ( .A(\MC_ARK_ARC_1_3/temp5[24] ), .B(
        \MC_ARK_ARC_1_3/temp6[24] ), .ZN(\RI1[4][24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_27_5  ( .A(\MC_ARK_ARC_1_3/temp3[24] ), .B(
        \MC_ARK_ARC_1_3/temp4[24] ), .ZN(\MC_ARK_ARC_1_3/temp6[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_27_5  ( .A(\MC_ARK_ARC_1_3/temp1[24] ), .B(
        \MC_ARK_ARC_1_3/temp2[24] ), .ZN(\MC_ARK_ARC_1_3/temp5[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_27_5  ( .A(\RI5[3][60] ), .B(n477), .ZN(
        \MC_ARK_ARC_1_3/temp4[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_27_5  ( .A(n1654), .B(\RI5[3][90] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_27_5  ( .A(\RI5[3][186] ), .B(\RI5[3][162] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_27_5  ( .A(\RI5[3][24] ), .B(\RI5[3][18] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[24] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_27_4  ( .A(\MC_ARK_ARC_1_3/temp5[25] ), .B(
        \MC_ARK_ARC_1_3/temp6[25] ), .ZN(\RI1[4][25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_27_4  ( .A(\MC_ARK_ARC_1_3/temp3[25] ), .B(
        \MC_ARK_ARC_1_3/temp4[25] ), .ZN(\MC_ARK_ARC_1_3/temp6[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_27_4  ( .A(\MC_ARK_ARC_1_3/temp1[25] ), .B(
        \MC_ARK_ARC_1_3/temp2[25] ), .ZN(\MC_ARK_ARC_1_3/temp5[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_27_4  ( .A(\RI5[3][61] ), .B(n366), .ZN(
        \MC_ARK_ARC_1_3/temp4[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_27_4  ( .A(\RI5[3][127] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_3/temp3[25] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_27_4  ( .A(\RI5[3][187] ), .B(\RI5[3][163] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_27_4  ( .A(\RI5[3][25] ), .B(\RI5[3][19] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[25] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_27_3  ( .A(\MC_ARK_ARC_1_3/temp3[26] ), .B(
        \MC_ARK_ARC_1_3/temp4[26] ), .ZN(\MC_ARK_ARC_1_3/temp6[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_27_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[62] ), 
        .B(n446), .ZN(\MC_ARK_ARC_1_3/temp4[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_27_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[128] ), 
        .B(\RI5[3][92] ), .ZN(\MC_ARK_ARC_1_3/temp3[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_27_3  ( .A(\RI5[3][188] ), .B(\RI5[3][164] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_27_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_3/temp1[26] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_27_2  ( .A(\MC_ARK_ARC_1_3/temp5[27] ), .B(
        \MC_ARK_ARC_1_3/temp6[27] ), .ZN(\RI1[4][27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_27_2  ( .A(\MC_ARK_ARC_1_3/temp3[27] ), .B(
        \MC_ARK_ARC_1_3/temp4[27] ), .ZN(\MC_ARK_ARC_1_3/temp6[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_27_2  ( .A(\MC_ARK_ARC_1_3/temp1[27] ), .B(
        \MC_ARK_ARC_1_3/temp2[27] ), .ZN(\MC_ARK_ARC_1_3/temp5[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_27_2  ( .A(\RI5[3][63] ), .B(n364), .ZN(
        \MC_ARK_ARC_1_3/temp4[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_27_2  ( .A(\RI5[3][129] ), .B(\RI5[3][93] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_27_2  ( .A(\RI5[3][189] ), .B(\RI5[3][165] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[27] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_27_2  ( .A(\RI5[3][27] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_3/temp1[27] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_27_1  ( .A(\MC_ARK_ARC_1_3/temp5[28] ), .B(
        \MC_ARK_ARC_1_3/temp6[28] ), .ZN(\RI1[4][28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_27_1  ( .A(\MC_ARK_ARC_1_3/temp3[28] ), .B(
        \MC_ARK_ARC_1_3/temp4[28] ), .ZN(\MC_ARK_ARC_1_3/temp6[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_27_1  ( .A(\MC_ARK_ARC_1_3/temp1[28] ), .B(
        \MC_ARK_ARC_1_3/temp2[28] ), .ZN(\MC_ARK_ARC_1_3/temp5[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_27_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[64] ), 
        .B(Key[108]), .ZN(\MC_ARK_ARC_1_3/temp4[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_27_1  ( .A(n1944), .B(\RI5[3][94] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_27_1  ( .A(\RI5[3][190] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[166] ), .ZN(\MC_ARK_ARC_1_3/temp2[28] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_27_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .B(\RI5[3][28] ), .ZN(\MC_ARK_ARC_1_3/temp1[28] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_27_0  ( .A(\MC_ARK_ARC_1_3/temp3[29] ), .B(
        \MC_ARK_ARC_1_3/temp4[29] ), .ZN(\MC_ARK_ARC_1_3/temp6[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_27_0  ( .A(\MC_ARK_ARC_1_3/temp2[29] ), .B(
        \MC_ARK_ARC_1_3/temp1[29] ), .ZN(\MC_ARK_ARC_1_3/temp5[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_27_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[65] ), 
        .B(n362), .ZN(\MC_ARK_ARC_1_3/temp4[29] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_27_0  ( .A(n2145), .B(
        \MC_ARK_ARC_1_3/buf_datainput[131] ), .ZN(\MC_ARK_ARC_1_3/temp3[29] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_27_0  ( .A(n1948), .B(
        \MC_ARK_ARC_1_3/buf_datainput[191] ), .ZN(\MC_ARK_ARC_1_3/temp2[29] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_27_0  ( .A(n1653), .B(
        \MC_ARK_ARC_1_3/buf_datainput[29] ), .ZN(\MC_ARK_ARC_1_3/temp1[29] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_26_5  ( .A(\MC_ARK_ARC_1_3/temp5[30] ), .B(
        \MC_ARK_ARC_1_3/temp6[30] ), .ZN(\RI1[4][30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_26_5  ( .A(\MC_ARK_ARC_1_3/temp3[30] ), .B(
        \MC_ARK_ARC_1_3/temp4[30] ), .ZN(\MC_ARK_ARC_1_3/temp6[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_26_5  ( .A(\MC_ARK_ARC_1_3/temp1[30] ), .B(
        \MC_ARK_ARC_1_3/temp2[30] ), .ZN(\MC_ARK_ARC_1_3/temp5[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_26_5  ( .A(\RI5[3][66] ), .B(n270), .ZN(
        \MC_ARK_ARC_1_3/temp4[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_26_5  ( .A(\RI5[3][0] ), .B(\RI5[3][168] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_26_5  ( .A(\RI5[3][30] ), .B(\RI5[3][24] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[30] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_26_4  ( .A(\MC_ARK_ARC_1_3/temp5[31] ), .B(
        \MC_ARK_ARC_1_3/temp6[31] ), .ZN(\RI1[4][31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_26_4  ( .A(\MC_ARK_ARC_1_3/temp3[31] ), .B(
        \MC_ARK_ARC_1_3/temp4[31] ), .ZN(\MC_ARK_ARC_1_3/temp6[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_26_4  ( .A(\MC_ARK_ARC_1_3/temp1[31] ), .B(
        \MC_ARK_ARC_1_3/temp2[31] ), .ZN(\MC_ARK_ARC_1_3/temp5[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_26_4  ( .A(\RI5[3][67] ), .B(n506), .ZN(
        \MC_ARK_ARC_1_3/temp4[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_26_4  ( .A(\RI5[3][133] ), .B(\RI5[3][97] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_26_4  ( .A(\RI5[3][1] ), .B(\RI5[3][169] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_26_4  ( .A(\RI5[3][31] ), .B(\RI5[3][25] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[31] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_26_3  ( .A(\MC_ARK_ARC_1_3/temp5[32] ), .B(
        \MC_ARK_ARC_1_3/temp6[32] ), .ZN(\RI1[4][32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_26_3  ( .A(\MC_ARK_ARC_1_3/temp3[32] ), .B(
        \MC_ARK_ARC_1_3/temp4[32] ), .ZN(\MC_ARK_ARC_1_3/temp6[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_26_3  ( .A(\MC_ARK_ARC_1_3/temp1[32] ), .B(
        \MC_ARK_ARC_1_3/temp2[32] ), .ZN(\MC_ARK_ARC_1_3/temp5[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_26_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[68] ), 
        .B(n268), .ZN(\MC_ARK_ARC_1_3/temp4[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_26_3  ( .A(\RI5[3][134] ), .B(\RI5[3][98] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_26_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[2] ), 
        .B(\RI5[3][170] ), .ZN(\MC_ARK_ARC_1_3/temp2[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_26_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[32] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_3/temp1[32] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_26_2  ( .A(\MC_ARK_ARC_1_3/temp5[33] ), .B(
        \MC_ARK_ARC_1_3/temp6[33] ), .ZN(\RI1[4][33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_26_2  ( .A(\MC_ARK_ARC_1_3/temp3[33] ), .B(
        \MC_ARK_ARC_1_3/temp4[33] ), .ZN(\MC_ARK_ARC_1_3/temp6[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_26_2  ( .A(\MC_ARK_ARC_1_3/temp1[33] ), .B(
        \MC_ARK_ARC_1_3/temp2[33] ), .ZN(\MC_ARK_ARC_1_3/temp5[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_26_2  ( .A(\RI5[3][69] ), .B(n393), .ZN(
        \MC_ARK_ARC_1_3/temp4[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_26_2  ( .A(\RI5[3][135] ), .B(\RI5[3][99] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_26_2  ( .A(\RI5[3][3] ), .B(\RI5[3][171] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_26_2  ( .A(\RI5[3][33] ), .B(\RI5[3][27] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[33] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_26_1  ( .A(\MC_ARK_ARC_1_3/temp6[34] ), .B(
        \MC_ARK_ARC_1_3/temp5[34] ), .ZN(\RI1[4][34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_26_1  ( .A(\MC_ARK_ARC_1_3/temp3[34] ), .B(
        \MC_ARK_ARC_1_3/temp4[34] ), .ZN(\MC_ARK_ARC_1_3/temp6[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_26_1  ( .A(\MC_ARK_ARC_1_3/temp1[34] ), .B(
        \MC_ARK_ARC_1_3/temp2[34] ), .ZN(\MC_ARK_ARC_1_3/temp5[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_26_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[70] ), 
        .B(n266), .ZN(\MC_ARK_ARC_1_3/temp4[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_26_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_26_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_26_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[34] ), 
        .B(\RI5[3][28] ), .ZN(\MC_ARK_ARC_1_3/temp1[34] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_26_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .B(n356), .ZN(\MC_ARK_ARC_1_3/temp4[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_26_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[137] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_26_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[173] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[5] ), .ZN(\MC_ARK_ARC_1_3/temp2[35] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_26_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[35] ), .ZN(\MC_ARK_ARC_1_3/temp1[35] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_25_5  ( .A(\MC_ARK_ARC_1_3/temp5[36] ), .B(
        \MC_ARK_ARC_1_3/temp6[36] ), .ZN(\RI1[4][36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_25_5  ( .A(\MC_ARK_ARC_1_3/temp3[36] ), .B(
        \MC_ARK_ARC_1_3/temp4[36] ), .ZN(\MC_ARK_ARC_1_3/temp6[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_25_5  ( .A(\MC_ARK_ARC_1_3/temp1[36] ), .B(
        \MC_ARK_ARC_1_3/temp2[36] ), .ZN(\MC_ARK_ARC_1_3/temp5[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_25_5  ( .A(\RI5[3][72] ), .B(n467), .ZN(
        \MC_ARK_ARC_1_3/temp4[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_25_5  ( .A(\RI5[3][138] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[102] ), .ZN(\MC_ARK_ARC_1_3/temp3[36] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_25_5  ( .A(\RI5[3][6] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[174] ), .ZN(\MC_ARK_ARC_1_3/temp2[36] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_25_5  ( .A(\RI5[3][36] ), .B(\RI5[3][30] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[36] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_25_4  ( .A(\MC_ARK_ARC_1_3/temp3[37] ), .B(
        \MC_ARK_ARC_1_3/temp4[37] ), .ZN(\MC_ARK_ARC_1_3/temp6[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_25_4  ( .A(\RI5[3][73] ), .B(n354), .ZN(
        \MC_ARK_ARC_1_3/temp4[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_25_4  ( .A(\RI5[3][139] ), .B(\RI5[3][103] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_25_4  ( .A(\RI5[3][7] ), .B(\RI5[3][175] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_25_4  ( .A(\RI5[3][37] ), .B(\RI5[3][31] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[37] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_25_3  ( .A(\MC_ARK_ARC_1_3/temp6[38] ), .B(
        \MC_ARK_ARC_1_3/temp5[38] ), .ZN(\RI1[4][38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_25_3  ( .A(\MC_ARK_ARC_1_3/temp3[38] ), .B(
        \MC_ARK_ARC_1_3/temp4[38] ), .ZN(\MC_ARK_ARC_1_3/temp6[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_25_3  ( .A(\MC_ARK_ARC_1_3/temp1[38] ), .B(
        \MC_ARK_ARC_1_3/temp2[38] ), .ZN(\MC_ARK_ARC_1_3/temp5[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_25_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .B(n262), .ZN(\MC_ARK_ARC_1_3/temp4[38] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_25_3  ( .A(\RI5[3][140] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[104] ), .ZN(\MC_ARK_ARC_1_3/temp3[38] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_25_3  ( .A(\RI5[3][8] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[176] ), .ZN(\MC_ARK_ARC_1_3/temp2[38] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_25_3  ( .A(\RI5[3][38] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[32] ), .ZN(\MC_ARK_ARC_1_3/temp1[38] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_25_2  ( .A(\MC_ARK_ARC_1_3/temp5[39] ), .B(
        \MC_ARK_ARC_1_3/temp6[39] ), .ZN(\RI1[4][39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_25_2  ( .A(\MC_ARK_ARC_1_3/temp3[39] ), .B(
        \MC_ARK_ARC_1_3/temp4[39] ), .ZN(\MC_ARK_ARC_1_3/temp6[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_25_2  ( .A(\MC_ARK_ARC_1_3/temp1[39] ), .B(
        \MC_ARK_ARC_1_3/temp2[39] ), .ZN(\MC_ARK_ARC_1_3/temp5[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_25_2  ( .A(\RI5[3][75] ), .B(n352), .ZN(
        \MC_ARK_ARC_1_3/temp4[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_25_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[141] ), 
        .B(\RI5[3][105] ), .ZN(\MC_ARK_ARC_1_3/temp3[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_25_2  ( .A(\RI5[3][9] ), .B(\RI5[3][177] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_25_2  ( .A(\RI5[3][39] ), .B(\RI5[3][33] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[39] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_25_1  ( .A(\MC_ARK_ARC_1_3/temp5[40] ), .B(
        \MC_ARK_ARC_1_3/temp6[40] ), .ZN(\RI1[4][40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_25_1  ( .A(\MC_ARK_ARC_1_3/temp3[40] ), .B(
        \MC_ARK_ARC_1_3/temp4[40] ), .ZN(\MC_ARK_ARC_1_3/temp6[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_25_1  ( .A(\MC_ARK_ARC_1_3/temp2[40] ), .B(
        \MC_ARK_ARC_1_3/temp1[40] ), .ZN(\MC_ARK_ARC_1_3/temp5[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_25_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[76] ), 
        .B(n260), .ZN(\MC_ARK_ARC_1_3/temp4[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_25_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[106] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_25_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[178] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_25_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[34] ), .ZN(\MC_ARK_ARC_1_3/temp1[40] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_25_0  ( .A(\MC_ARK_ARC_1_3/temp5[41] ), .B(
        \MC_ARK_ARC_1_3/temp6[41] ), .ZN(\RI1[4][41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_25_0  ( .A(\MC_ARK_ARC_1_3/temp3[41] ), .B(
        \MC_ARK_ARC_1_3/temp4[41] ), .ZN(\MC_ARK_ARC_1_3/temp6[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_25_0  ( .A(\MC_ARK_ARC_1_3/temp2[41] ), .B(
        \MC_ARK_ARC_1_3/temp1[41] ), .ZN(\MC_ARK_ARC_1_3/temp5[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_25_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[77] ), 
        .B(n350), .ZN(\MC_ARK_ARC_1_3/temp4[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_25_0  ( .A(n1661), .B(n2108), .ZN(
        \MC_ARK_ARC_1_3/temp3[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_25_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[11] ), .ZN(\MC_ARK_ARC_1_3/temp2[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_25_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[35] ), 
        .B(n2111), .ZN(\MC_ARK_ARC_1_3/temp1[41] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_24_5  ( .A(\MC_ARK_ARC_1_3/temp5[42] ), .B(
        \MC_ARK_ARC_1_3/temp6[42] ), .ZN(\RI1[4][42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_24_5  ( .A(\MC_ARK_ARC_1_3/temp3[42] ), .B(
        \MC_ARK_ARC_1_3/temp4[42] ), .ZN(\MC_ARK_ARC_1_3/temp6[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_24_5  ( .A(\MC_ARK_ARC_1_3/temp1[42] ), .B(
        \MC_ARK_ARC_1_3/temp2[42] ), .ZN(\MC_ARK_ARC_1_3/temp5[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_24_5  ( .A(\RI5[3][78] ), .B(n258), .ZN(
        \MC_ARK_ARC_1_3/temp4[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_24_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[12] ), 
        .B(\RI5[3][180] ), .ZN(\MC_ARK_ARC_1_3/temp2[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_24_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[42] ), 
        .B(\RI5[3][36] ), .ZN(\MC_ARK_ARC_1_3/temp1[42] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_24_4  ( .A(\MC_ARK_ARC_1_3/temp3[43] ), .B(
        \MC_ARK_ARC_1_3/temp4[43] ), .ZN(\MC_ARK_ARC_1_3/temp6[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_24_4  ( .A(\RI5[3][79] ), .B(n348), .ZN(
        \MC_ARK_ARC_1_3/temp4[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_24_4  ( .A(\RI5[3][145] ), .B(\RI5[3][109] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_24_4  ( .A(\RI5[3][13] ), .B(\RI5[3][181] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_24_4  ( .A(\RI5[3][43] ), .B(\RI5[3][37] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[43] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_24_3  ( .A(\MC_ARK_ARC_1_3/temp5[44] ), .B(
        \MC_ARK_ARC_1_3/temp6[44] ), .ZN(\RI1[4][44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_24_3  ( .A(\MC_ARK_ARC_1_3/temp3[44] ), .B(
        \MC_ARK_ARC_1_3/temp4[44] ), .ZN(\MC_ARK_ARC_1_3/temp6[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_24_3  ( .A(\MC_ARK_ARC_1_3/temp2[44] ), .B(
        \MC_ARK_ARC_1_3/temp1[44] ), .ZN(\MC_ARK_ARC_1_3/temp5[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_24_3  ( .A(\RI5[3][80] ), .B(
        \MC_ARK_ARC_1_3/buf_keyinput[44] ), .ZN(\MC_ARK_ARC_1_3/temp4[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_24_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[146] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[110] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_24_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_24_3  ( .A(\RI5[3][44] ), .B(\RI5[3][38] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[44] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_24_2  ( .A(\MC_ARK_ARC_1_3/temp5[45] ), .B(
        \MC_ARK_ARC_1_3/temp6[45] ), .ZN(\RI1[4][45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_24_2  ( .A(\MC_ARK_ARC_1_3/temp3[45] ), .B(
        \MC_ARK_ARC_1_3/temp4[45] ), .ZN(\MC_ARK_ARC_1_3/temp6[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_24_2  ( .A(\MC_ARK_ARC_1_3/temp1[45] ), .B(
        \MC_ARK_ARC_1_3/temp2[45] ), .ZN(\MC_ARK_ARC_1_3/temp5[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_24_2  ( .A(\RI5[3][81] ), .B(n346), .ZN(
        \MC_ARK_ARC_1_3/temp4[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_24_2  ( .A(\RI5[3][147] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[111] ), .ZN(\MC_ARK_ARC_1_3/temp3[45] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_24_2  ( .A(\RI5[3][15] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[183] ), .ZN(\MC_ARK_ARC_1_3/temp2[45] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_24_2  ( .A(\RI5[3][45] ), .B(\RI5[3][39] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[45] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_24_1  ( .A(\MC_ARK_ARC_1_3/temp5[46] ), .B(
        \MC_ARK_ARC_1_3/temp6[46] ), .ZN(\RI1[4][46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_24_1  ( .A(\MC_ARK_ARC_1_3/temp3[46] ), .B(
        \MC_ARK_ARC_1_3/temp4[46] ), .ZN(\MC_ARK_ARC_1_3/temp6[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_24_1  ( .A(\MC_ARK_ARC_1_3/temp1[46] ), .B(
        \MC_ARK_ARC_1_3/temp2[46] ), .ZN(\MC_ARK_ARC_1_3/temp5[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_24_1  ( .A(\RI5[3][82] ), .B(n383), .ZN(
        \MC_ARK_ARC_1_3/temp4[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_24_1  ( .A(n1510), .B(
        \MC_ARK_ARC_1_3/buf_datainput[112] ), .ZN(\MC_ARK_ARC_1_3/temp3[46] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_24_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[16] ), 
        .B(\RI5[3][184] ), .ZN(\MC_ARK_ARC_1_3/temp2[46] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_24_1  ( .A(\RI5[3][46] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[40] ), .ZN(\MC_ARK_ARC_1_3/temp1[46] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_24_0  ( .A(\MC_ARK_ARC_1_3/temp5[47] ), .B(
        \MC_ARK_ARC_1_3/temp6[47] ), .ZN(\RI1[4][47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_24_0  ( .A(\MC_ARK_ARC_1_3/temp3[47] ), .B(
        \MC_ARK_ARC_1_3/temp4[47] ), .ZN(\MC_ARK_ARC_1_3/temp6[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_24_0  ( .A(\MC_ARK_ARC_1_3/temp1[47] ), .B(
        \MC_ARK_ARC_1_3/temp2[47] ), .ZN(\MC_ARK_ARC_1_3/temp5[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_24_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[83] ), 
        .B(n344), .ZN(\MC_ARK_ARC_1_3/temp4[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_24_0  ( .A(n849), .B(n796), .ZN(
        \MC_ARK_ARC_1_3/temp3[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_24_0  ( .A(n839), .B(
        \MC_ARK_ARC_1_3/buf_datainput[17] ), .ZN(\MC_ARK_ARC_1_3/temp2[47] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_24_0  ( .A(n2111), .B(n842), .ZN(
        \MC_ARK_ARC_1_3/temp1[47] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_23_5  ( .A(\MC_ARK_ARC_1_3/temp5[48] ), .B(
        \MC_ARK_ARC_1_3/temp6[48] ), .ZN(\RI1[4][48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_23_5  ( .A(\MC_ARK_ARC_1_3/temp3[48] ), .B(
        \MC_ARK_ARC_1_3/temp4[48] ), .ZN(\MC_ARK_ARC_1_3/temp6[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_23_5  ( .A(\MC_ARK_ARC_1_3/temp2[48] ), .B(
        \MC_ARK_ARC_1_3/temp1[48] ), .ZN(\MC_ARK_ARC_1_3/temp5[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_23_5  ( .A(\RI5[3][84] ), .B(n252), .ZN(
        \MC_ARK_ARC_1_3/temp4[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_23_5  ( .A(\RI5[3][150] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[114] ), .ZN(\MC_ARK_ARC_1_3/temp3[48] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_23_5  ( .A(\RI5[3][18] ), .B(\RI5[3][186] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[48] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_23_5  ( .A(\RI5[3][48] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_3/temp1[48] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_23_4  ( .A(\MC_ARK_ARC_1_3/temp5[49] ), .B(
        \MC_ARK_ARC_1_3/temp6[49] ), .ZN(\RI1[4][49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_23_4  ( .A(\MC_ARK_ARC_1_3/temp3[49] ), .B(
        \MC_ARK_ARC_1_3/temp4[49] ), .ZN(\MC_ARK_ARC_1_3/temp6[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_23_4  ( .A(\MC_ARK_ARC_1_3/temp1[49] ), .B(
        \MC_ARK_ARC_1_3/temp2[49] ), .ZN(\MC_ARK_ARC_1_3/temp5[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_23_4  ( .A(\RI5[3][85] ), .B(n504), .ZN(
        \MC_ARK_ARC_1_3/temp4[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_23_4  ( .A(\RI5[3][151] ), .B(\RI5[3][115] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_23_4  ( .A(\RI5[3][19] ), .B(\RI5[3][187] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_23_4  ( .A(\RI5[3][49] ), .B(\RI5[3][43] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[49] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_23_3  ( .A(\MC_ARK_ARC_1_3/temp5[50] ), .B(
        \MC_ARK_ARC_1_3/temp6[50] ), .ZN(\RI1[4][50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_23_3  ( .A(\MC_ARK_ARC_1_3/temp3[50] ), .B(
        \MC_ARK_ARC_1_3/temp4[50] ), .ZN(\MC_ARK_ARC_1_3/temp6[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_23_3  ( .A(\MC_ARK_ARC_1_3/temp1[50] ), .B(
        \MC_ARK_ARC_1_3/temp2[50] ), .ZN(\MC_ARK_ARC_1_3/temp5[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_23_3  ( .A(\RI5[3][86] ), .B(n471), .ZN(
        \MC_ARK_ARC_1_3/temp4[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_23_3  ( .A(\RI5[3][152] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[116] ), .ZN(\MC_ARK_ARC_1_3/temp3[50] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_23_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[20] ), 
        .B(\RI5[3][188] ), .ZN(\MC_ARK_ARC_1_3/temp2[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_23_3  ( .A(n2128), .B(\RI5[3][44] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[50] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_23_2  ( .A(\MC_ARK_ARC_1_3/temp5[51] ), .B(
        \MC_ARK_ARC_1_3/temp6[51] ), .ZN(\RI1[4][51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_23_2  ( .A(\MC_ARK_ARC_1_3/temp3[51] ), .B(
        \MC_ARK_ARC_1_3/temp4[51] ), .ZN(\MC_ARK_ARC_1_3/temp6[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_23_2  ( .A(\MC_ARK_ARC_1_3/temp2[51] ), .B(
        \MC_ARK_ARC_1_3/temp1[51] ), .ZN(\MC_ARK_ARC_1_3/temp5[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_23_2  ( .A(\RI5[3][87] ), .B(n407), .ZN(
        \MC_ARK_ARC_1_3/temp4[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_23_2  ( .A(\RI5[3][153] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[117] ), .ZN(\MC_ARK_ARC_1_3/temp3[51] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_23_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .B(\RI5[3][189] ), .ZN(\MC_ARK_ARC_1_3/temp2[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_23_2  ( .A(\RI5[3][51] ), .B(\RI5[3][45] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[51] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_23_1  ( .A(\MC_ARK_ARC_1_3/temp5[52] ), .B(
        \MC_ARK_ARC_1_3/temp6[52] ), .ZN(\RI1[4][52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_23_1  ( .A(\MC_ARK_ARC_1_3/temp3[52] ), .B(
        \MC_ARK_ARC_1_3/temp4[52] ), .ZN(\MC_ARK_ARC_1_3/temp6[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_23_1  ( .A(\MC_ARK_ARC_1_3/temp1[52] ), .B(
        \MC_ARK_ARC_1_3/temp2[52] ), .ZN(\MC_ARK_ARC_1_3/temp5[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_23_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[177] ), .ZN(\MC_ARK_ARC_1_3/temp4[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_23_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[154] ), 
        .B(\RI5[3][118] ), .ZN(\MC_ARK_ARC_1_3/temp3[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_23_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .B(\RI5[3][190] ), .ZN(\MC_ARK_ARC_1_3/temp2[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_23_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[52] ), 
        .B(\RI5[3][46] ), .ZN(\MC_ARK_ARC_1_3/temp1[52] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_23_0  ( .A(\MC_ARK_ARC_1_3/temp5[53] ), .B(
        \MC_ARK_ARC_1_3/temp6[53] ), .ZN(\RI1[4][53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_23_0  ( .A(\MC_ARK_ARC_1_3/temp3[53] ), .B(
        \MC_ARK_ARC_1_3/temp4[53] ), .ZN(\MC_ARK_ARC_1_3/temp6[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_23_0  ( .A(\MC_ARK_ARC_1_3/temp1[53] ), .B(
        \MC_ARK_ARC_1_3/temp2[53] ), .ZN(\MC_ARK_ARC_1_3/temp5[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_23_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[89] ), 
        .B(n339), .ZN(\MC_ARK_ARC_1_3/temp4[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_23_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .B(n2121), .ZN(\MC_ARK_ARC_1_3/temp3[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_23_0  ( .A(n1653), .B(
        \MC_ARK_ARC_1_3/buf_datainput[191] ), .ZN(\MC_ARK_ARC_1_3/temp2[53] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_23_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .B(n842), .ZN(\MC_ARK_ARC_1_3/temp1[53] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_22_5  ( .A(\MC_ARK_ARC_1_3/temp5[54] ), .B(
        \MC_ARK_ARC_1_3/temp6[54] ), .ZN(\RI1[4][54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_22_5  ( .A(\MC_ARK_ARC_1_3/temp3[54] ), .B(
        \MC_ARK_ARC_1_3/temp4[54] ), .ZN(\MC_ARK_ARC_1_3/temp6[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_22_5  ( .A(\MC_ARK_ARC_1_3/temp1[54] ), .B(
        \MC_ARK_ARC_1_3/temp2[54] ), .ZN(\MC_ARK_ARC_1_3/temp5[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_22_5  ( .A(\RI5[3][90] ), .B(n247), .ZN(
        \MC_ARK_ARC_1_3/temp4[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_22_5  ( .A(\RI5[3][156] ), .B(\RI5[3][120] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_22_5  ( .A(\RI5[3][24] ), .B(\RI5[3][0] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_22_5  ( .A(\RI5[3][54] ), .B(\RI5[3][48] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[54] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_22_4  ( .A(\MC_ARK_ARC_1_3/temp5[55] ), .B(
        \MC_ARK_ARC_1_3/temp6[55] ), .ZN(\RI1[4][55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_22_4  ( .A(\MC_ARK_ARC_1_3/temp3[55] ), .B(
        \MC_ARK_ARC_1_3/temp4[55] ), .ZN(\MC_ARK_ARC_1_3/temp6[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_22_4  ( .A(\MC_ARK_ARC_1_3/temp1[55] ), .B(
        \MC_ARK_ARC_1_3/temp2[55] ), .ZN(\MC_ARK_ARC_1_3/temp5[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_22_4  ( .A(\MC_ARK_ARC_1_3/buf_datainput[91] ), 
        .B(n337), .ZN(\MC_ARK_ARC_1_3/temp4[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_22_4  ( .A(\RI5[3][157] ), .B(\RI5[3][121] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_22_4  ( .A(\RI5[3][25] ), .B(\RI5[3][1] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_22_4  ( .A(\RI5[3][55] ), .B(\RI5[3][49] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[55] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_22_3  ( .A(\MC_ARK_ARC_1_3/temp5[56] ), .B(
        \MC_ARK_ARC_1_3/temp6[56] ), .ZN(\RI1[4][56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_22_3  ( .A(\MC_ARK_ARC_1_3/temp3[56] ), .B(
        \MC_ARK_ARC_1_3/temp4[56] ), .ZN(\MC_ARK_ARC_1_3/temp6[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_22_3  ( .A(\MC_ARK_ARC_1_3/temp1[56] ), .B(
        \MC_ARK_ARC_1_3/temp2[56] ), .ZN(\MC_ARK_ARC_1_3/temp5[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_22_3  ( .A(\RI5[3][92] ), .B(n376), .ZN(
        \MC_ARK_ARC_1_3/temp4[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_22_3  ( .A(n1955), .B(n1930), .ZN(
        \MC_ARK_ARC_1_3/temp3[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_22_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_3/temp2[56] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_22_3  ( .A(\RI5[3][56] ), .B(n2128), .ZN(
        \MC_ARK_ARC_1_3/temp1[56] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_22_2  ( .A(\MC_ARK_ARC_1_3/temp5[57] ), .B(
        \MC_ARK_ARC_1_3/temp6[57] ), .ZN(\RI1[4][57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_22_2  ( .A(\MC_ARK_ARC_1_3/temp3[57] ), .B(
        \MC_ARK_ARC_1_3/temp4[57] ), .ZN(\MC_ARK_ARC_1_3/temp6[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_22_2  ( .A(\MC_ARK_ARC_1_3/temp1[57] ), .B(
        \MC_ARK_ARC_1_3/temp2[57] ), .ZN(\MC_ARK_ARC_1_3/temp5[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_22_2  ( .A(\RI5[3][93] ), .B(n400), .ZN(
        \MC_ARK_ARC_1_3/temp4[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_22_2  ( .A(\RI5[3][159] ), .B(\RI5[3][123] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_22_2  ( .A(\RI5[3][27] ), .B(\RI5[3][3] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_22_2  ( .A(\RI5[3][57] ), .B(\RI5[3][51] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[57] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_22_1  ( .A(\MC_ARK_ARC_1_3/temp5[58] ), .B(
        \MC_ARK_ARC_1_3/temp6[58] ), .ZN(\RI1[4][58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_22_1  ( .A(\MC_ARK_ARC_1_3/temp3[58] ), .B(
        \MC_ARK_ARC_1_3/temp4[58] ), .ZN(\MC_ARK_ARC_1_3/temp6[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_22_1  ( .A(\MC_ARK_ARC_1_3/temp2[58] ), .B(
        \MC_ARK_ARC_1_3/temp1[58] ), .ZN(\MC_ARK_ARC_1_3/temp5[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_22_1  ( .A(\RI5[3][94] ), .B(Key[138]), .ZN(
        \MC_ARK_ARC_1_3/temp4[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_22_1  ( .A(\RI5[3][160] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[124] ), .ZN(\MC_ARK_ARC_1_3/temp3[58] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_22_1  ( .A(\RI5[3][28] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[4] ), .ZN(\MC_ARK_ARC_1_3/temp2[58] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_22_1  ( .A(n2103), .B(
        \MC_ARK_ARC_1_3/buf_datainput[52] ), .ZN(\MC_ARK_ARC_1_3/temp1[58] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_22_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[95] ), 
        .B(n334), .ZN(\MC_ARK_ARC_1_3/temp4[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_22_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[161] ), 
        .B(n520), .ZN(\MC_ARK_ARC_1_3/temp3[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_22_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[5] ), .ZN(\MC_ARK_ARC_1_3/temp2[59] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_22_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[59] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[53] ), .ZN(\MC_ARK_ARC_1_3/temp1[59] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_21_5  ( .A(\MC_ARK_ARC_1_3/temp5[60] ), .B(
        \MC_ARK_ARC_1_3/temp6[60] ), .ZN(\RI1[4][60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_21_5  ( .A(\MC_ARK_ARC_1_3/temp3[60] ), .B(
        \MC_ARK_ARC_1_3/temp4[60] ), .ZN(\MC_ARK_ARC_1_3/temp6[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_21_5  ( .A(\MC_ARK_ARC_1_3/temp1[60] ), .B(
        \MC_ARK_ARC_1_3/temp2[60] ), .ZN(\MC_ARK_ARC_1_3/temp5[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_21_5  ( .A(\RI5[3][96] ), .B(n242), .ZN(
        \MC_ARK_ARC_1_3/temp4[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_21_5  ( .A(\RI5[3][162] ), .B(\RI5[3][126] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_21_5  ( .A(\RI5[3][30] ), .B(\RI5[3][6] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_21_5  ( .A(\RI5[3][60] ), .B(\RI5[3][54] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[60] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_21_4  ( .A(\MC_ARK_ARC_1_3/temp5[61] ), .B(
        \MC_ARK_ARC_1_3/temp6[61] ), .ZN(\RI1[4][61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_21_4  ( .A(\MC_ARK_ARC_1_3/temp3[61] ), .B(
        \MC_ARK_ARC_1_3/temp4[61] ), .ZN(\MC_ARK_ARC_1_3/temp6[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_21_4  ( .A(\MC_ARK_ARC_1_3/temp2[61] ), .B(
        \MC_ARK_ARC_1_3/temp1[61] ), .ZN(\MC_ARK_ARC_1_3/temp5[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_21_4  ( .A(\RI5[3][97] ), .B(n332), .ZN(
        \MC_ARK_ARC_1_3/temp4[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_21_4  ( .A(\RI5[3][163] ), .B(\RI5[3][127] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_21_4  ( .A(\RI5[3][31] ), .B(\RI5[3][7] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_21_4  ( .A(\RI5[3][61] ), .B(\RI5[3][55] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[61] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_21_3  ( .A(\MC_ARK_ARC_1_3/temp5[62] ), .B(
        \MC_ARK_ARC_1_3/temp6[62] ), .ZN(\RI1[4][62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_21_3  ( .A(\MC_ARK_ARC_1_3/temp3[62] ), .B(
        \MC_ARK_ARC_1_3/temp4[62] ), .ZN(\MC_ARK_ARC_1_3/temp6[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_21_3  ( .A(\MC_ARK_ARC_1_3/temp1[62] ), .B(
        \MC_ARK_ARC_1_3/temp2[62] ), .ZN(\MC_ARK_ARC_1_3/temp5[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_21_3  ( .A(\RI5[3][98] ), .B(n461), .ZN(
        \MC_ARK_ARC_1_3/temp4[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_21_3  ( .A(n1626), .B(
        \MC_ARK_ARC_1_3/buf_datainput[128] ), .ZN(\MC_ARK_ARC_1_3/temp3[62] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_21_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[32] ), 
        .B(\RI5[3][8] ), .ZN(\MC_ARK_ARC_1_3/temp2[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_21_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[62] ), 
        .B(\RI5[3][56] ), .ZN(\MC_ARK_ARC_1_3/temp1[62] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_21_2  ( .A(\MC_ARK_ARC_1_3/temp5[63] ), .B(
        \MC_ARK_ARC_1_3/temp6[63] ), .ZN(\RI1[4][63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_21_2  ( .A(\MC_ARK_ARC_1_3/temp3[63] ), .B(
        \MC_ARK_ARC_1_3/temp4[63] ), .ZN(\MC_ARK_ARC_1_3/temp6[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_21_2  ( .A(\MC_ARK_ARC_1_3/temp1[63] ), .B(
        \MC_ARK_ARC_1_3/temp2[63] ), .ZN(\MC_ARK_ARC_1_3/temp5[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_21_2  ( .A(\RI5[3][99] ), .B(n330), .ZN(
        \MC_ARK_ARC_1_3/temp4[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_21_2  ( .A(\RI5[3][165] ), .B(\RI5[3][129] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_21_2  ( .A(\RI5[3][33] ), .B(\RI5[3][9] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_21_2  ( .A(\RI5[3][63] ), .B(\RI5[3][57] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[63] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_21_1  ( .A(\MC_ARK_ARC_1_3/temp3[64] ), .B(
        \MC_ARK_ARC_1_3/temp4[64] ), .ZN(\MC_ARK_ARC_1_3/temp6[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_21_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[166] ), 
        .B(n1943), .ZN(\MC_ARK_ARC_1_3/temp3[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_21_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[34] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_3/temp2[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_21_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[64] ), 
        .B(n2102), .ZN(\MC_ARK_ARC_1_3/temp1[64] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_21_0  ( .A(\MC_ARK_ARC_1_3/temp5[65] ), .B(
        \MC_ARK_ARC_1_3/temp6[65] ), .ZN(\RI1[4][65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_21_0  ( .A(\MC_ARK_ARC_1_3/temp3[65] ), .B(
        \MC_ARK_ARC_1_3/temp4[65] ), .ZN(\MC_ARK_ARC_1_3/temp6[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_21_0  ( .A(\MC_ARK_ARC_1_3/temp2[65] ), .B(
        \MC_ARK_ARC_1_3/temp1[65] ), .ZN(\MC_ARK_ARC_1_3/temp5[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_21_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .B(n328), .ZN(\MC_ARK_ARC_1_3/temp4[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_21_0  ( .A(n1947), .B(
        \MC_ARK_ARC_1_3/buf_datainput[131] ), .ZN(\MC_ARK_ARC_1_3/temp3[65] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_21_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[35] ), 
        .B(n1650), .ZN(\MC_ARK_ARC_1_3/temp2[65] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_21_0  ( .A(n2112), .B(
        \MC_ARK_ARC_1_3/buf_datainput[59] ), .ZN(\MC_ARK_ARC_1_3/temp1[65] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_20_5  ( .A(\MC_ARK_ARC_1_3/temp5[66] ), .B(
        \MC_ARK_ARC_1_3/temp6[66] ), .ZN(\RI1[4][66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_20_5  ( .A(\MC_ARK_ARC_1_3/temp3[66] ), .B(
        \MC_ARK_ARC_1_3/temp4[66] ), .ZN(\MC_ARK_ARC_1_3/temp6[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_20_5  ( .A(\MC_ARK_ARC_1_3/temp1[66] ), .B(
        \MC_ARK_ARC_1_3/temp2[66] ), .ZN(\MC_ARK_ARC_1_3/temp5[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_20_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .B(n237), .ZN(\MC_ARK_ARC_1_3/temp4[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_20_5  ( .A(\RI5[3][168] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[132] ), .ZN(\MC_ARK_ARC_1_3/temp3[66] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_20_5  ( .A(\RI5[3][36] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_3/temp2[66] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_20_5  ( .A(\RI5[3][66] ), .B(\RI5[3][60] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[66] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_20_4  ( .A(\MC_ARK_ARC_1_3/temp5[67] ), .B(
        \MC_ARK_ARC_1_3/temp6[67] ), .ZN(\RI1[4][67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_20_4  ( .A(\MC_ARK_ARC_1_3/temp3[67] ), .B(
        \MC_ARK_ARC_1_3/temp4[67] ), .ZN(\MC_ARK_ARC_1_3/temp6[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_20_4  ( .A(\MC_ARK_ARC_1_3/temp1[67] ), .B(
        \MC_ARK_ARC_1_3/temp2[67] ), .ZN(\MC_ARK_ARC_1_3/temp5[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_20_4  ( .A(\RI5[3][103] ), .B(n496), .ZN(
        \MC_ARK_ARC_1_3/temp4[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_20_4  ( .A(\RI5[3][169] ), .B(\RI5[3][133] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_20_4  ( .A(\RI5[3][37] ), .B(\RI5[3][13] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_20_4  ( .A(\RI5[3][67] ), .B(\RI5[3][61] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[67] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_20_3  ( .A(\MC_ARK_ARC_1_3/temp6[68] ), .B(
        \MC_ARK_ARC_1_3/temp5[68] ), .ZN(\RI1[4][68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_20_3  ( .A(\MC_ARK_ARC_1_3/temp3[68] ), .B(
        \MC_ARK_ARC_1_3/temp4[68] ), .ZN(\MC_ARK_ARC_1_3/temp6[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_20_3  ( .A(\MC_ARK_ARC_1_3/temp1[68] ), .B(
        \MC_ARK_ARC_1_3/temp2[68] ), .ZN(\MC_ARK_ARC_1_3/temp5[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_20_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[104] ), 
        .B(n235), .ZN(\MC_ARK_ARC_1_3/temp4[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_20_3  ( .A(\RI5[3][170] ), .B(\RI5[3][134] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_20_3  ( .A(\RI5[3][38] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[14] ), .ZN(\MC_ARK_ARC_1_3/temp2[68] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_20_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[68] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[62] ), .ZN(\MC_ARK_ARC_1_3/temp1[68] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_20_2  ( .A(\MC_ARK_ARC_1_3/temp5[69] ), .B(
        \MC_ARK_ARC_1_3/temp6[69] ), .ZN(\RI1[4][69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_20_2  ( .A(\MC_ARK_ARC_1_3/temp3[69] ), .B(
        \MC_ARK_ARC_1_3/temp4[69] ), .ZN(\MC_ARK_ARC_1_3/temp6[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_20_2  ( .A(\MC_ARK_ARC_1_3/temp1[69] ), .B(
        \MC_ARK_ARC_1_3/temp2[69] ), .ZN(\MC_ARK_ARC_1_3/temp5[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_20_2  ( .A(\RI5[3][105] ), .B(n324), .ZN(
        \MC_ARK_ARC_1_3/temp4[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_20_2  ( .A(\RI5[3][171] ), .B(\RI5[3][135] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_20_2  ( .A(\RI5[3][39] ), .B(\RI5[3][15] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_20_2  ( .A(\RI5[3][69] ), .B(\RI5[3][63] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[69] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_20_1  ( .A(\MC_ARK_ARC_1_3/temp3[70] ), .B(
        \MC_ARK_ARC_1_3/temp4[70] ), .ZN(\MC_ARK_ARC_1_3/temp6[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_20_1  ( .A(\MC_ARK_ARC_1_3/temp1[70] ), .B(
        \MC_ARK_ARC_1_3/temp2[70] ), .ZN(\MC_ARK_ARC_1_3/temp5[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_20_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[70] ), .ZN(\MC_ARK_ARC_1_3/temp4[70] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_20_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[136] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_20_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[40] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[16] ), .ZN(\MC_ARK_ARC_1_3/temp2[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_20_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[64] ), .ZN(\MC_ARK_ARC_1_3/temp1[70] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_20_0  ( .A(\MC_ARK_ARC_1_3/temp5[71] ), .B(
        \MC_ARK_ARC_1_3/temp6[71] ), .ZN(\RI1[4][71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_20_0  ( .A(\MC_ARK_ARC_1_3/temp3[71] ), .B(
        \MC_ARK_ARC_1_3/temp4[71] ), .ZN(\MC_ARK_ARC_1_3/temp6[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_20_0  ( .A(\MC_ARK_ARC_1_3/temp2[71] ), .B(
        \MC_ARK_ARC_1_3/temp1[71] ), .ZN(\MC_ARK_ARC_1_3/temp5[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_20_0  ( .A(n2109), .B(n322), .ZN(
        \MC_ARK_ARC_1_3/temp4[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_20_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[173] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[137] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_20_0  ( .A(n2111), .B(
        \MC_ARK_ARC_1_3/buf_datainput[17] ), .ZN(\MC_ARK_ARC_1_3/temp2[71] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_20_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .B(n2112), .ZN(\MC_ARK_ARC_1_3/temp1[71] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_19_5  ( .A(\MC_ARK_ARC_1_3/temp3[72] ), .B(
        \MC_ARK_ARC_1_3/temp4[72] ), .ZN(\MC_ARK_ARC_1_3/temp6[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_19_5  ( .A(\RI5[3][108] ), .B(n231), .ZN(
        \MC_ARK_ARC_1_3/temp4[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_19_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .B(\RI5[3][138] ), .ZN(\MC_ARK_ARC_1_3/temp3[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_19_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[42] ), 
        .B(\RI5[3][18] ), .ZN(\MC_ARK_ARC_1_3/temp2[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_19_5  ( .A(\RI5[3][72] ), .B(\RI5[3][66] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[72] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_19_4  ( .A(\MC_ARK_ARC_1_3/temp5[73] ), .B(
        \MC_ARK_ARC_1_3/temp6[73] ), .ZN(\RI1[4][73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_19_4  ( .A(\MC_ARK_ARC_1_3/temp3[73] ), .B(
        \MC_ARK_ARC_1_3/temp4[73] ), .ZN(\MC_ARK_ARC_1_3/temp6[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_19_4  ( .A(\MC_ARK_ARC_1_3/temp1[73] ), .B(
        \MC_ARK_ARC_1_3/temp2[73] ), .ZN(\MC_ARK_ARC_1_3/temp5[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_19_4  ( .A(\RI5[3][109] ), .B(n320), .ZN(
        \MC_ARK_ARC_1_3/temp4[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_19_4  ( .A(\RI5[3][175] ), .B(\RI5[3][139] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_19_4  ( .A(\RI5[3][43] ), .B(\RI5[3][19] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_19_4  ( .A(\RI5[3][73] ), .B(\RI5[3][67] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[73] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_19_3  ( .A(\MC_ARK_ARC_1_3/temp5[74] ), .B(
        \MC_ARK_ARC_1_3/temp6[74] ), .ZN(\RI1[4][74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_19_3  ( .A(\MC_ARK_ARC_1_3/temp3[74] ), .B(
        \MC_ARK_ARC_1_3/temp4[74] ), .ZN(\MC_ARK_ARC_1_3/temp6[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_19_3  ( .A(\MC_ARK_ARC_1_3/temp2[74] ), .B(
        \MC_ARK_ARC_1_3/temp1[74] ), .ZN(\MC_ARK_ARC_1_3/temp5[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_19_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[110] ), 
        .B(n229), .ZN(\MC_ARK_ARC_1_3/temp4[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_19_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .B(\RI5[3][140] ), .ZN(\MC_ARK_ARC_1_3/temp3[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_19_3  ( .A(\RI5[3][44] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_3/temp2[74] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_19_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_3/temp1[74] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_19_2  ( .A(\MC_ARK_ARC_1_3/temp5[75] ), .B(
        \MC_ARK_ARC_1_3/temp6[75] ), .ZN(\RI1[4][75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_19_2  ( .A(\MC_ARK_ARC_1_3/temp4[75] ), .B(
        \MC_ARK_ARC_1_3/temp3[75] ), .ZN(\MC_ARK_ARC_1_3/temp6[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_19_2  ( .A(\MC_ARK_ARC_1_3/temp1[75] ), .B(
        \MC_ARK_ARC_1_3/temp2[75] ), .ZN(\MC_ARK_ARC_1_3/temp5[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_19_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[111] ), 
        .B(n319), .ZN(\MC_ARK_ARC_1_3/temp4[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_19_2  ( .A(\RI5[3][177] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[141] ), .ZN(\MC_ARK_ARC_1_3/temp3[75] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_19_2  ( .A(\RI5[3][45] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_3/temp2[75] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_19_2  ( .A(\RI5[3][75] ), .B(\RI5[3][69] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[75] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_19_1  ( .A(\MC_ARK_ARC_1_3/temp3[76] ), .B(
        \MC_ARK_ARC_1_3/temp4[76] ), .ZN(\MC_ARK_ARC_1_3/temp6[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_19_1  ( .A(\MC_ARK_ARC_1_3/temp2[76] ), .B(
        \MC_ARK_ARC_1_3/temp1[76] ), .ZN(\MC_ARK_ARC_1_3/temp5[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_19_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[112] ), 
        .B(n227), .ZN(\MC_ARK_ARC_1_3/temp4[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_19_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[142] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_19_1  ( .A(\RI5[3][46] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[22] ), .ZN(\MC_ARK_ARC_1_3/temp2[76] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_19_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[76] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_3/temp1[76] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_19_0  ( .A(n797), .B(
        \MC_ARK_ARC_1_1/buf_keyinput[165] ), .ZN(\MC_ARK_ARC_1_3/temp4[77] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_19_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .B(n1661), .ZN(\MC_ARK_ARC_1_3/temp3[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_19_0  ( .A(n1653), .B(
        \MC_ARK_ARC_1_3/buf_datainput[47] ), .ZN(\MC_ARK_ARC_1_3/temp2[77] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_19_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[77] ), .ZN(\MC_ARK_ARC_1_3/temp1[77] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_18_5  ( .A(\MC_ARK_ARC_1_3/temp5[78] ), .B(
        \MC_ARK_ARC_1_3/temp6[78] ), .ZN(\RI1[4][78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_18_5  ( .A(\MC_ARK_ARC_1_3/temp3[78] ), .B(
        \MC_ARK_ARC_1_3/temp4[78] ), .ZN(\MC_ARK_ARC_1_3/temp6[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_18_5  ( .A(\MC_ARK_ARC_1_3/temp2[78] ), .B(
        \MC_ARK_ARC_1_3/temp1[78] ), .ZN(\MC_ARK_ARC_1_3/temp5[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_18_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[114] ), 
        .B(n225), .ZN(\MC_ARK_ARC_1_3/temp4[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_18_5  ( .A(\RI5[3][180] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[144] ), .ZN(\MC_ARK_ARC_1_3/temp3[78] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_18_5  ( .A(\RI5[3][48] ), .B(\RI5[3][24] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_18_5  ( .A(\RI5[3][78] ), .B(\RI5[3][72] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[78] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_18_4  ( .A(\MC_ARK_ARC_1_3/temp3[79] ), .B(
        \MC_ARK_ARC_1_3/temp4[79] ), .ZN(\MC_ARK_ARC_1_3/temp6[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_18_4  ( .A(\RI5[3][115] ), .B(n315), .ZN(
        \MC_ARK_ARC_1_3/temp4[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_18_4  ( .A(\RI5[3][181] ), .B(\RI5[3][145] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_18_4  ( .A(\RI5[3][49] ), .B(\RI5[3][25] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_18_4  ( .A(\RI5[3][79] ), .B(\RI5[3][73] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[79] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_18_3  ( .A(\MC_ARK_ARC_1_3/temp5[80] ), .B(
        \MC_ARK_ARC_1_3/temp6[80] ), .ZN(\RI1[4][80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_18_3  ( .A(\MC_ARK_ARC_1_3/temp3[80] ), .B(
        \MC_ARK_ARC_1_3/temp4[80] ), .ZN(\MC_ARK_ARC_1_3/temp6[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_18_3  ( .A(\MC_ARK_ARC_1_3/temp1[80] ), .B(
        \MC_ARK_ARC_1_3/temp2[80] ), .ZN(\MC_ARK_ARC_1_3/temp5[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_18_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[116] ), 
        .B(Key[160]), .ZN(\MC_ARK_ARC_1_3/temp4[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_18_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[146] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_18_3  ( .A(n2129), .B(
        \MC_ARK_ARC_1_3/buf_datainput[26] ), .ZN(\MC_ARK_ARC_1_3/temp2[80] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_18_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .B(\RI5[3][80] ), .ZN(\MC_ARK_ARC_1_3/temp1[80] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_18_2  ( .A(\MC_ARK_ARC_1_3/temp5[81] ), .B(
        \MC_ARK_ARC_1_3/temp6[81] ), .ZN(\RI1[4][81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_18_2  ( .A(\MC_ARK_ARC_1_3/temp3[81] ), .B(
        \MC_ARK_ARC_1_3/temp4[81] ), .ZN(\MC_ARK_ARC_1_3/temp6[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_18_2  ( .A(\MC_ARK_ARC_1_3/temp1[81] ), .B(
        \MC_ARK_ARC_1_3/temp2[81] ), .ZN(\MC_ARK_ARC_1_3/temp5[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_18_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[117] ), 
        .B(n313), .ZN(\MC_ARK_ARC_1_3/temp4[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_18_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[183] ), 
        .B(\RI5[3][147] ), .ZN(\MC_ARK_ARC_1_3/temp3[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_18_2  ( .A(\RI5[3][51] ), .B(\RI5[3][27] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_18_2  ( .A(n1658), .B(\RI5[3][75] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[81] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_18_1  ( .A(\MC_ARK_ARC_1_3/temp3[82] ), .B(
        \MC_ARK_ARC_1_3/temp4[82] ), .ZN(\MC_ARK_ARC_1_3/temp6[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_18_1  ( .A(\RI5[3][118] ), .B(
        \MC_ARK_ARC_1_0/buf_keyinput[187] ), .ZN(\MC_ARK_ARC_1_3/temp4[82] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_18_1  ( .A(\RI5[3][184] ), .B(n1510), .ZN(
        \MC_ARK_ARC_1_3/temp3[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_18_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[52] ), 
        .B(\RI5[3][28] ), .ZN(\MC_ARK_ARC_1_3/temp2[82] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_18_1  ( .A(\RI5[3][82] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[76] ), .ZN(\MC_ARK_ARC_1_3/temp1[82] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_18_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .B(n311), .ZN(\MC_ARK_ARC_1_3/temp4[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_18_0  ( .A(n850), .B(
        \MC_ARK_ARC_1_3/buf_datainput[185] ), .ZN(\MC_ARK_ARC_1_3/temp3[83] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_18_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[29] ), .ZN(\MC_ARK_ARC_1_3/temp2[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_18_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[83] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[77] ), .ZN(\MC_ARK_ARC_1_3/temp1[83] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_17_5  ( .A(\MC_ARK_ARC_1_3/temp5[84] ), .B(
        \MC_ARK_ARC_1_3/temp6[84] ), .ZN(\RI1[4][84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_17_5  ( .A(\MC_ARK_ARC_1_3/temp3[84] ), .B(
        \MC_ARK_ARC_1_3/temp4[84] ), .ZN(\MC_ARK_ARC_1_3/temp6[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_17_5  ( .A(\MC_ARK_ARC_1_3/temp1[84] ), .B(
        \MC_ARK_ARC_1_3/temp2[84] ), .ZN(\MC_ARK_ARC_1_3/temp5[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_17_5  ( .A(\RI5[3][120] ), .B(n219), .ZN(
        \MC_ARK_ARC_1_3/temp4[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_17_5  ( .A(\RI5[3][186] ), .B(\RI5[3][150] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_17_5  ( .A(\RI5[3][54] ), .B(\RI5[3][30] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_17_5  ( .A(n2130), .B(\RI5[3][78] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[84] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_17_4  ( .A(\MC_ARK_ARC_1_3/temp5[85] ), .B(
        \MC_ARK_ARC_1_3/temp6[85] ), .ZN(\RI1[4][85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_17_4  ( .A(\MC_ARK_ARC_1_3/temp3[85] ), .B(
        \MC_ARK_ARC_1_3/temp4[85] ), .ZN(\MC_ARK_ARC_1_3/temp6[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_17_4  ( .A(\MC_ARK_ARC_1_3/temp1[85] ), .B(
        \MC_ARK_ARC_1_3/temp2[85] ), .ZN(\MC_ARK_ARC_1_3/temp5[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_17_4  ( .A(\RI5[3][121] ), .B(n449), .ZN(
        \MC_ARK_ARC_1_3/temp4[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_17_4  ( .A(\RI5[3][187] ), .B(\RI5[3][151] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_17_4  ( .A(\RI5[3][55] ), .B(\RI5[3][31] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_17_4  ( .A(\RI5[3][85] ), .B(\RI5[3][79] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[85] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_17_3  ( .A(\MC_ARK_ARC_1_3/temp3[86] ), .B(
        \MC_ARK_ARC_1_3/temp4[86] ), .ZN(\MC_ARK_ARC_1_3/temp6[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_17_3  ( .A(n1929), .B(n431), .ZN(
        \MC_ARK_ARC_1_3/temp4[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_17_3  ( .A(\RI5[3][188] ), .B(\RI5[3][152] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_17_3  ( .A(\RI5[3][56] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[32] ), .ZN(\MC_ARK_ARC_1_3/temp2[86] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_17_3  ( .A(\RI5[3][86] ), .B(\RI5[3][80] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[86] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_17_2  ( .A(\MC_ARK_ARC_1_3/temp5[87] ), .B(
        \MC_ARK_ARC_1_3/temp6[87] ), .ZN(\RI1[4][87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_17_2  ( .A(\MC_ARK_ARC_1_3/temp3[87] ), .B(
        \MC_ARK_ARC_1_3/temp4[87] ), .ZN(\MC_ARK_ARC_1_3/temp6[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_17_2  ( .A(\MC_ARK_ARC_1_3/temp1[87] ), .B(
        \MC_ARK_ARC_1_3/temp2[87] ), .ZN(\MC_ARK_ARC_1_3/temp5[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_17_2  ( .A(\RI5[3][123] ), .B(n397), .ZN(
        \MC_ARK_ARC_1_3/temp4[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_17_2  ( .A(\RI5[3][189] ), .B(\RI5[3][153] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_17_2  ( .A(\RI5[3][57] ), .B(\RI5[3][33] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_17_2  ( .A(\RI5[3][87] ), .B(n1658), .ZN(
        \MC_ARK_ARC_1_3/temp1[87] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_17_1  ( .A(\MC_ARK_ARC_1_3/temp3[88] ), .B(
        \MC_ARK_ARC_1_3/temp4[88] ), .ZN(\MC_ARK_ARC_1_3/temp6[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_17_1  ( .A(\MC_ARK_ARC_1_3/temp2[88] ), .B(
        \MC_ARK_ARC_1_3/temp1[88] ), .ZN(\MC_ARK_ARC_1_3/temp5[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_17_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_2/buf_keyinput[45] ), .ZN(\MC_ARK_ARC_1_3/temp4[88] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_17_1  ( .A(\RI5[3][190] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[154] ), .ZN(\MC_ARK_ARC_1_3/temp3[88] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_17_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[34] ), 
        .B(n2103), .ZN(\MC_ARK_ARC_1_3/temp2[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_17_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[88] ), 
        .B(\RI5[3][82] ), .ZN(\MC_ARK_ARC_1_3/temp1[88] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_17_0  ( .A(\MC_ARK_ARC_1_3/temp5[89] ), .B(
        \MC_ARK_ARC_1_3/temp6[89] ), .ZN(\RI1[4][89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_17_0  ( .A(\MC_ARK_ARC_1_3/temp3[89] ), .B(
        \MC_ARK_ARC_1_3/temp4[89] ), .ZN(\MC_ARK_ARC_1_3/temp6[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_17_0  ( .A(\MC_ARK_ARC_1_3/temp2[89] ), .B(
        \MC_ARK_ARC_1_3/temp1[89] ), .ZN(\MC_ARK_ARC_1_3/temp5[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_17_0  ( .A(n521), .B(
        \MC_ARK_ARC_1_3/buf_keyinput[89] ), .ZN(\MC_ARK_ARC_1_3/temp4[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_17_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[191] ), 
        .B(n2120), .ZN(\MC_ARK_ARC_1_3/temp3[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_17_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[35] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[59] ), .ZN(\MC_ARK_ARC_1_3/temp2[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_17_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[83] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[89] ), .ZN(\MC_ARK_ARC_1_3/temp1[89] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_16_5  ( .A(\MC_ARK_ARC_1_3/temp5[90] ), .B(
        \MC_ARK_ARC_1_3/temp6[90] ), .ZN(\RI1[4][90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_16_5  ( .A(\MC_ARK_ARC_1_3/temp3[90] ), .B(
        \MC_ARK_ARC_1_3/temp4[90] ), .ZN(\MC_ARK_ARC_1_3/temp6[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_16_5  ( .A(\MC_ARK_ARC_1_3/temp1[90] ), .B(
        \MC_ARK_ARC_1_3/temp2[90] ), .ZN(\MC_ARK_ARC_1_3/temp5[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_16_5  ( .A(\RI5[3][126] ), .B(n481), .ZN(
        \MC_ARK_ARC_1_3/temp4[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_16_5  ( .A(\RI5[3][0] ), .B(\RI5[3][156] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_16_5  ( .A(\RI5[3][60] ), .B(\RI5[3][36] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_16_5  ( .A(\RI5[3][90] ), .B(n2130), .ZN(
        \MC_ARK_ARC_1_3/temp1[90] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_16_4  ( .A(\MC_ARK_ARC_1_3/temp5[91] ), .B(
        \MC_ARK_ARC_1_3/temp6[91] ), .ZN(\RI1[4][91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_16_4  ( .A(\MC_ARK_ARC_1_3/temp3[91] ), .B(
        \MC_ARK_ARC_1_3/temp4[91] ), .ZN(\MC_ARK_ARC_1_3/temp6[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_16_4  ( .A(\MC_ARK_ARC_1_3/temp1[91] ), .B(
        \MC_ARK_ARC_1_3/temp2[91] ), .ZN(\MC_ARK_ARC_1_3/temp5[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_16_4  ( .A(\RI5[3][127] ), .B(n502), .ZN(
        \MC_ARK_ARC_1_3/temp4[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_16_4  ( .A(\RI5[3][1] ), .B(\RI5[3][157] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_16_4  ( .A(\RI5[3][61] ), .B(\RI5[3][37] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_16_4  ( .A(\MC_ARK_ARC_1_3/buf_datainput[91] ), 
        .B(\RI5[3][85] ), .ZN(\MC_ARK_ARC_1_3/temp1[91] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_16_3  ( .A(\MC_ARK_ARC_1_3/temp1[92] ), .B(
        \MC_ARK_ARC_1_3/temp2[92] ), .ZN(\MC_ARK_ARC_1_3/temp5[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_16_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[128] ), 
        .B(n211), .ZN(\MC_ARK_ARC_1_3/temp4[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_16_3  ( .A(n2119), .B(
        \MC_ARK_ARC_1_3/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_3/temp3[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_16_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[62] ), 
        .B(\RI5[3][38] ), .ZN(\MC_ARK_ARC_1_3/temp2[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_16_3  ( .A(\RI5[3][92] ), .B(\RI5[3][86] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[92] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_16_2  ( .A(\MC_ARK_ARC_1_3/temp5[93] ), .B(
        \MC_ARK_ARC_1_3/temp6[93] ), .ZN(\RI1[4][93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_16_2  ( .A(\MC_ARK_ARC_1_3/temp3[93] ), .B(
        \MC_ARK_ARC_1_3/temp4[93] ), .ZN(\MC_ARK_ARC_1_3/temp6[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_16_2  ( .A(\MC_ARK_ARC_1_3/temp1[93] ), .B(
        \MC_ARK_ARC_1_3/temp2[93] ), .ZN(\MC_ARK_ARC_1_3/temp5[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_16_2  ( .A(\RI5[3][129] ), .B(n387), .ZN(
        \MC_ARK_ARC_1_3/temp4[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_16_2  ( .A(\RI5[3][3] ), .B(\RI5[3][159] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_16_2  ( .A(\RI5[3][63] ), .B(\RI5[3][39] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_16_2  ( .A(\RI5[3][93] ), .B(\RI5[3][87] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[93] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_16_1  ( .A(\MC_ARK_ARC_1_3/temp3[94] ), .B(
        \MC_ARK_ARC_1_3/temp4[94] ), .ZN(\MC_ARK_ARC_1_3/temp6[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_16_1  ( .A(n1942), .B(n209), .ZN(
        \MC_ARK_ARC_1_3/temp4[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_16_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[4] ), 
        .B(\RI5[3][160] ), .ZN(\MC_ARK_ARC_1_3/temp3[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_16_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[64] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[40] ), .ZN(\MC_ARK_ARC_1_3/temp2[94] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_16_1  ( .A(\RI5[3][94] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[88] ), .ZN(\MC_ARK_ARC_1_3/temp1[94] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_16_0  ( .A(\MC_ARK_ARC_1_3/temp5[95] ), .B(
        \MC_ARK_ARC_1_3/temp6[95] ), .ZN(\RI1[4][95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_16_0  ( .A(\MC_ARK_ARC_1_3/temp4[95] ), .B(
        \MC_ARK_ARC_1_3/temp3[95] ), .ZN(\MC_ARK_ARC_1_3/temp6[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_16_0  ( .A(\MC_ARK_ARC_1_3/temp1[95] ), .B(
        \MC_ARK_ARC_1_3/temp2[95] ), .ZN(\MC_ARK_ARC_1_3/temp5[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_16_0  ( .A(n801), .B(n299), .ZN(
        \MC_ARK_ARC_1_3/temp4[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_16_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[161] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[5] ), .ZN(\MC_ARK_ARC_1_3/temp3[95] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_16_0  ( .A(n2111), .B(n2112), .ZN(
        \MC_ARK_ARC_1_3/temp2[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_16_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[89] ), 
        .B(n2145), .ZN(\MC_ARK_ARC_1_3/temp1[95] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_15_5  ( .A(\MC_ARK_ARC_1_3/temp5[96] ), .B(
        \MC_ARK_ARC_1_3/temp6[96] ), .ZN(\RI1[4][96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_15_5  ( .A(\MC_ARK_ARC_1_3/temp3[96] ), .B(
        \MC_ARK_ARC_1_3/temp4[96] ), .ZN(\MC_ARK_ARC_1_3/temp6[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_15_5  ( .A(\MC_ARK_ARC_1_3/temp1[96] ), .B(
        \MC_ARK_ARC_1_3/temp2[96] ), .ZN(\MC_ARK_ARC_1_3/temp5[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_15_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[132] ), 
        .B(n207), .ZN(\MC_ARK_ARC_1_3/temp4[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_15_5  ( .A(\RI5[3][6] ), .B(\RI5[3][162] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_15_5  ( .A(\RI5[3][66] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_3/temp2[96] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_15_5  ( .A(\RI5[3][96] ), .B(\RI5[3][90] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[96] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_15_4  ( .A(\MC_ARK_ARC_1_3/temp5[97] ), .B(
        \MC_ARK_ARC_1_3/temp6[97] ), .ZN(\RI1[4][97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_15_4  ( .A(\MC_ARK_ARC_1_3/temp3[97] ), .B(
        \MC_ARK_ARC_1_3/temp4[97] ), .ZN(\MC_ARK_ARC_1_3/temp6[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_15_4  ( .A(\MC_ARK_ARC_1_3/temp1[97] ), .B(
        \MC_ARK_ARC_1_3/temp2[97] ), .ZN(\MC_ARK_ARC_1_3/temp5[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_15_4  ( .A(\RI5[3][133] ), .B(n298), .ZN(
        \MC_ARK_ARC_1_3/temp4[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_15_4  ( .A(\RI5[3][7] ), .B(\RI5[3][163] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_15_4  ( .A(\RI5[3][67] ), .B(\RI5[3][43] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[97] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_15_4  ( .A(\RI5[3][97] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_3/temp1[97] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_15_3  ( .A(\MC_ARK_ARC_1_3/temp5[98] ), .B(
        \MC_ARK_ARC_1_3/temp6[98] ), .ZN(\RI1[4][98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_15_3  ( .A(\MC_ARK_ARC_1_3/temp3[98] ), .B(
        \MC_ARK_ARC_1_3/temp4[98] ), .ZN(\MC_ARK_ARC_1_3/temp6[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_15_3  ( .A(\MC_ARK_ARC_1_3/temp1[98] ), .B(
        \MC_ARK_ARC_1_3/temp2[98] ), .ZN(\MC_ARK_ARC_1_3/temp5[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_15_3  ( .A(\RI5[3][134] ), .B(n436), .ZN(
        \MC_ARK_ARC_1_3/temp4[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_15_3  ( .A(\RI5[3][8] ), .B(n1626), .ZN(
        \MC_ARK_ARC_1_3/temp3[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_15_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[68] ), 
        .B(\RI5[3][44] ), .ZN(\MC_ARK_ARC_1_3/temp2[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_15_3  ( .A(\RI5[3][98] ), .B(\RI5[3][92] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[98] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_15_2  ( .A(\MC_ARK_ARC_1_3/temp5[99] ), .B(
        \MC_ARK_ARC_1_3/temp6[99] ), .ZN(\RI1[4][99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_15_2  ( .A(\MC_ARK_ARC_1_3/temp3[99] ), .B(
        \MC_ARK_ARC_1_3/temp4[99] ), .ZN(\MC_ARK_ARC_1_3/temp6[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_15_2  ( .A(\MC_ARK_ARC_1_3/temp1[99] ), .B(
        \MC_ARK_ARC_1_3/temp2[99] ), .ZN(\MC_ARK_ARC_1_3/temp5[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_15_2  ( .A(\RI5[3][135] ), .B(n296), .ZN(
        \MC_ARK_ARC_1_3/temp4[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_15_2  ( .A(\RI5[3][9] ), .B(\RI5[3][165] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_15_2  ( .A(\RI5[3][69] ), .B(\RI5[3][45] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_15_2  ( .A(\RI5[3][99] ), .B(\RI5[3][93] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[99] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_15_1  ( .A(\MC_ARK_ARC_1_3/temp5[100] ), .B(
        \MC_ARK_ARC_1_3/temp6[100] ), .ZN(\RI1[4][100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_15_1  ( .A(\MC_ARK_ARC_1_3/temp3[100] ), .B(
        \MC_ARK_ARC_1_3/temp4[100] ), .ZN(\MC_ARK_ARC_1_3/temp6[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_15_1  ( .A(\MC_ARK_ARC_1_3/temp1[100] ), .B(
        \MC_ARK_ARC_1_3/temp2[100] ), .ZN(\MC_ARK_ARC_1_3/temp5[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_15_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[136] ), 
        .B(n203), .ZN(\MC_ARK_ARC_1_3/temp4[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_15_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_15_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[70] ), 
        .B(\RI5[3][46] ), .ZN(\MC_ARK_ARC_1_3/temp2[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_15_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[100] ), 
        .B(\RI5[3][94] ), .ZN(\MC_ARK_ARC_1_3/temp1[100] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_15_0  ( .A(\MC_ARK_ARC_1_3/temp5[101] ), .B(
        \MC_ARK_ARC_1_3/temp6[101] ), .ZN(\RI1[4][101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_15_0  ( .A(\MC_ARK_ARC_1_3/temp3[101] ), .B(
        \MC_ARK_ARC_1_3/temp4[101] ), .ZN(\MC_ARK_ARC_1_3/temp6[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_15_0  ( .A(\MC_ARK_ARC_1_3/temp1[101] ), .B(
        \MC_ARK_ARC_1_3/temp2[101] ), .ZN(\MC_ARK_ARC_1_3/temp5[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_15_0  ( .A(n1946), .B(
        \MC_ARK_ARC_1_3/buf_datainput[11] ), .ZN(\MC_ARK_ARC_1_3/temp3[101] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_15_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .B(n842), .ZN(\MC_ARK_ARC_1_3/temp2[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_15_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[95] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[101] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_14_5  ( .A(\MC_ARK_ARC_1_3/temp5[102] ), .B(
        \MC_ARK_ARC_1_3/temp6[102] ), .ZN(\RI1[4][102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_14_5  ( .A(\MC_ARK_ARC_1_3/temp3[102] ), .B(
        \MC_ARK_ARC_1_3/temp4[102] ), .ZN(\MC_ARK_ARC_1_3/temp6[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_14_5  ( .A(\MC_ARK_ARC_1_3/temp1[102] ), .B(
        \MC_ARK_ARC_1_3/temp2[102] ), .ZN(\MC_ARK_ARC_1_3/temp5[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_14_5  ( .A(\RI5[3][138] ), .B(n201), .ZN(
        \MC_ARK_ARC_1_3/temp4[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_14_5  ( .A(\RI5[3][72] ), .B(\RI5[3][48] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_14_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .B(\RI5[3][96] ), .ZN(\MC_ARK_ARC_1_3/temp1[102] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_14_4  ( .A(\MC_ARK_ARC_1_3/temp5[103] ), .B(
        \MC_ARK_ARC_1_3/temp6[103] ), .ZN(\RI1[4][103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_14_4  ( .A(\MC_ARK_ARC_1_3/temp3[103] ), .B(
        \MC_ARK_ARC_1_3/temp4[103] ), .ZN(\MC_ARK_ARC_1_3/temp6[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_14_4  ( .A(\MC_ARK_ARC_1_3/temp1[103] ), .B(
        \MC_ARK_ARC_1_3/temp2[103] ), .ZN(\MC_ARK_ARC_1_3/temp5[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_14_4  ( .A(\RI5[3][139] ), .B(n292), .ZN(
        \MC_ARK_ARC_1_3/temp4[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_14_4  ( .A(\RI5[3][13] ), .B(\RI5[3][169] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_14_4  ( .A(\RI5[3][73] ), .B(\RI5[3][49] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_14_4  ( .A(\RI5[3][103] ), .B(\RI5[3][97] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[103] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_14_3  ( .A(\MC_ARK_ARC_1_3/temp5[104] ), .B(
        \MC_ARK_ARC_1_3/temp6[104] ), .ZN(\RI1[4][104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_14_3  ( .A(\MC_ARK_ARC_1_3/temp3[104] ), .B(
        \MC_ARK_ARC_1_3/temp4[104] ), .ZN(\MC_ARK_ARC_1_3/temp6[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_14_3  ( .A(\MC_ARK_ARC_1_3/temp1[104] ), .B(
        \MC_ARK_ARC_1_3/temp2[104] ), .ZN(\MC_ARK_ARC_1_3/temp5[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_14_3  ( .A(\RI5[3][140] ), .B(n474), .ZN(
        \MC_ARK_ARC_1_3/temp4[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_14_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .B(\RI5[3][170] ), .ZN(\MC_ARK_ARC_1_3/temp3[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_14_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .B(\RI5[3][50] ), .ZN(\MC_ARK_ARC_1_3/temp2[104] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_14_3  ( .A(\RI5[3][98] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[104] ), .ZN(\MC_ARK_ARC_1_3/temp1[104] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_14_2  ( .A(\MC_ARK_ARC_1_3/temp5[105] ), .B(
        \MC_ARK_ARC_1_3/temp6[105] ), .ZN(\RI1[4][105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_14_2  ( .A(\MC_ARK_ARC_1_3/temp3[105] ), .B(
        \MC_ARK_ARC_1_3/temp4[105] ), .ZN(\MC_ARK_ARC_1_3/temp6[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_14_2  ( .A(\MC_ARK_ARC_1_3/temp1[105] ), .B(
        \MC_ARK_ARC_1_3/temp2[105] ), .ZN(\MC_ARK_ARC_1_3/temp5[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_14_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[141] ), 
        .B(n290), .ZN(\MC_ARK_ARC_1_3/temp4[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_14_2  ( .A(\RI5[3][15] ), .B(\RI5[3][171] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_14_2  ( .A(\RI5[3][75] ), .B(\RI5[3][51] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_14_2  ( .A(\RI5[3][105] ), .B(\RI5[3][99] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[105] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_14_1  ( .A(\MC_ARK_ARC_1_3/temp5[106] ), .B(
        \MC_ARK_ARC_1_3/temp6[106] ), .ZN(\RI1[4][106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_14_1  ( .A(\MC_ARK_ARC_1_3/temp3[106] ), .B(
        \MC_ARK_ARC_1_3/temp4[106] ), .ZN(\MC_ARK_ARC_1_3/temp6[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_14_1  ( .A(\MC_ARK_ARC_1_3/temp1[106] ), .B(
        \MC_ARK_ARC_1_3/temp2[106] ), .ZN(\MC_ARK_ARC_1_3/temp5[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_14_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .B(Key[186]), .ZN(\MC_ARK_ARC_1_3/temp4[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_14_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_14_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[76] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[52] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_14_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[106] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[106] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_14_0  ( .A(\MC_ARK_ARC_1_3/temp5[107] ), .B(
        \MC_ARK_ARC_1_3/temp6[107] ), .ZN(\RI1[4][107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_14_0  ( .A(\MC_ARK_ARC_1_3/temp3[107] ), .B(
        \MC_ARK_ARC_1_3/temp4[107] ), .ZN(\MC_ARK_ARC_1_3/temp6[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_14_0  ( .A(\MC_ARK_ARC_1_3/temp2[107] ), .B(
        \MC_ARK_ARC_1_3/temp1[107] ), .ZN(\MC_ARK_ARC_1_3/temp5[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_14_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[143] ), 
        .B(n423), .ZN(\MC_ARK_ARC_1_3/temp4[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_14_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[173] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[17] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_14_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[77] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_14_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .B(n2109), .ZN(\MC_ARK_ARC_1_3/temp1[107] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_13_5  ( .A(\MC_ARK_ARC_1_3/temp5[108] ), .B(
        \MC_ARK_ARC_1_3/temp6[108] ), .ZN(\RI1[4][108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_13_5  ( .A(\MC_ARK_ARC_1_3/temp3[108] ), .B(
        \MC_ARK_ARC_1_3/temp4[108] ), .ZN(\MC_ARK_ARC_1_3/temp6[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_13_5  ( .A(\MC_ARK_ARC_1_3/temp1[108] ), .B(
        \MC_ARK_ARC_1_3/temp2[108] ), .ZN(\MC_ARK_ARC_1_3/temp5[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_13_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[144] ), 
        .B(n196), .ZN(\MC_ARK_ARC_1_3/temp4[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_13_5  ( .A(\RI5[3][18] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[174] ), .ZN(\MC_ARK_ARC_1_3/temp3[108] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_13_5  ( .A(\RI5[3][78] ), .B(\RI5[3][54] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[108] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_13_5  ( .A(\RI5[3][108] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[102] ), .ZN(\MC_ARK_ARC_1_3/temp1[108] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_13_4  ( .A(\MC_ARK_ARC_1_3/temp5[109] ), .B(
        \MC_ARK_ARC_1_3/temp6[109] ), .ZN(\RI1[4][109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_13_4  ( .A(\MC_ARK_ARC_1_3/temp3[109] ), .B(
        \MC_ARK_ARC_1_3/temp4[109] ), .ZN(\MC_ARK_ARC_1_3/temp6[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_13_4  ( .A(\MC_ARK_ARC_1_3/temp1[109] ), .B(
        \MC_ARK_ARC_1_3/temp2[109] ), .ZN(\MC_ARK_ARC_1_3/temp5[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_13_4  ( .A(\RI5[3][145] ), .B(n286), .ZN(
        \MC_ARK_ARC_1_3/temp4[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_13_4  ( .A(\RI5[3][19] ), .B(\RI5[3][175] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_13_4  ( .A(\RI5[3][79] ), .B(\RI5[3][55] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_13_4  ( .A(\RI5[3][109] ), .B(\RI5[3][103] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[109] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_13_3  ( .A(\MC_ARK_ARC_1_3/temp5[110] ), .B(
        \MC_ARK_ARC_1_3/temp6[110] ), .ZN(\RI1[4][110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_13_3  ( .A(\MC_ARK_ARC_1_3/temp3[110] ), .B(
        \MC_ARK_ARC_1_3/temp4[110] ), .ZN(\MC_ARK_ARC_1_3/temp6[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_13_3  ( .A(\MC_ARK_ARC_1_3/temp1[110] ), .B(
        \MC_ARK_ARC_1_3/temp2[110] ), .ZN(\MC_ARK_ARC_1_3/temp5[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_13_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[146] ), 
        .B(n194), .ZN(\MC_ARK_ARC_1_3/temp4[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_13_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[20] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_13_3  ( .A(\RI5[3][80] ), .B(\RI5[3][56] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_13_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[110] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[110] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_13_2  ( .A(\MC_ARK_ARC_1_3/temp5[111] ), .B(
        \MC_ARK_ARC_1_3/temp6[111] ), .ZN(\RI1[4][111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_13_2  ( .A(\MC_ARK_ARC_1_3/temp3[111] ), .B(
        \MC_ARK_ARC_1_3/temp4[111] ), .ZN(\MC_ARK_ARC_1_3/temp6[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_13_2  ( .A(\MC_ARK_ARC_1_3/temp2[111] ), .B(
        \MC_ARK_ARC_1_3/temp1[111] ), .ZN(\MC_ARK_ARC_1_3/temp5[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_13_2  ( .A(\RI5[3][147] ), .B(n479), .ZN(
        \MC_ARK_ARC_1_3/temp4[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_13_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .B(\RI5[3][177] ), .ZN(\MC_ARK_ARC_1_3/temp3[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_13_2  ( .A(n1658), .B(\RI5[3][57] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_13_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[111] ), 
        .B(\RI5[3][105] ), .ZN(\MC_ARK_ARC_1_3/temp1[111] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_13_1  ( .A(\MC_ARK_ARC_1_3/temp5[112] ), .B(
        \MC_ARK_ARC_1_3/temp6[112] ), .ZN(\RI1[4][112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_13_1  ( .A(\MC_ARK_ARC_1_3/temp3[112] ), .B(
        \MC_ARK_ARC_1_3/temp4[112] ), .ZN(\MC_ARK_ARC_1_3/temp6[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_13_1  ( .A(\MC_ARK_ARC_1_3/temp2[112] ), .B(
        \MC_ARK_ARC_1_3/temp1[112] ), .ZN(\MC_ARK_ARC_1_3/temp5[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_13_1  ( .A(n1510), .B(n374), .ZN(
        \MC_ARK_ARC_1_3/temp4[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_13_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[178] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_13_1  ( .A(\RI5[3][82] ), .B(n2102), .ZN(
        \MC_ARK_ARC_1_3/temp2[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_13_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[106] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[112] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_13_0  ( .A(\MC_ARK_ARC_1_3/temp3[113] ), .B(
        \MC_ARK_ARC_1_3/temp4[113] ), .ZN(\MC_ARK_ARC_1_3/temp6[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_13_0  ( .A(\MC_ARK_ARC_1_3/temp2[113] ), .B(
        \MC_ARK_ARC_1_3/temp1[113] ), .ZN(\MC_ARK_ARC_1_3/temp5[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_13_0  ( .A(n850), .B(n457), .ZN(
        \MC_ARK_ARC_1_3/temp4[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_13_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[23] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_13_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[59] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[83] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_13_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[107] ), 
        .B(n796), .ZN(\MC_ARK_ARC_1_3/temp1[113] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_12_5  ( .A(\MC_ARK_ARC_1_3/temp5[114] ), .B(
        \MC_ARK_ARC_1_3/temp6[114] ), .ZN(\RI1[4][114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_12_5  ( .A(\MC_ARK_ARC_1_3/temp3[114] ), .B(
        \MC_ARK_ARC_1_3/temp4[114] ), .ZN(\MC_ARK_ARC_1_3/temp6[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_12_5  ( .A(\MC_ARK_ARC_1_3/temp2[114] ), .B(
        \MC_ARK_ARC_1_3/temp1[114] ), .ZN(\MC_ARK_ARC_1_3/temp5[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_12_5  ( .A(\RI5[3][150] ), .B(n372), .ZN(
        \MC_ARK_ARC_1_3/temp4[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_12_5  ( .A(\RI5[3][24] ), .B(\RI5[3][180] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_12_5  ( .A(n2130), .B(\RI5[3][60] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_12_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[114] ), 
        .B(\RI5[3][108] ), .ZN(\MC_ARK_ARC_1_3/temp1[114] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_12_4  ( .A(\MC_ARK_ARC_1_3/temp5[115] ), .B(
        \MC_ARK_ARC_1_3/temp6[115] ), .ZN(\RI1[4][115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_12_4  ( .A(\MC_ARK_ARC_1_3/temp3[115] ), .B(
        \MC_ARK_ARC_1_3/temp4[115] ), .ZN(\MC_ARK_ARC_1_3/temp6[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_12_4  ( .A(\MC_ARK_ARC_1_3/temp1[115] ), .B(
        \MC_ARK_ARC_1_3/temp2[115] ), .ZN(\MC_ARK_ARC_1_3/temp5[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_12_4  ( .A(\RI5[3][151] ), .B(n281), .ZN(
        \MC_ARK_ARC_1_3/temp4[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_12_4  ( .A(\RI5[3][25] ), .B(\RI5[3][181] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_12_4  ( .A(\RI5[3][85] ), .B(\RI5[3][61] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_12_4  ( .A(\RI5[3][115] ), .B(\RI5[3][109] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[115] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_12_3  ( .A(\MC_ARK_ARC_1_3/temp5[116] ), .B(
        \MC_ARK_ARC_1_3/temp6[116] ), .ZN(\RI1[4][116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_12_3  ( .A(\MC_ARK_ARC_1_3/temp3[116] ), .B(
        \MC_ARK_ARC_1_3/temp4[116] ), .ZN(\MC_ARK_ARC_1_3/temp6[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_12_3  ( .A(\MC_ARK_ARC_1_3/temp2[116] ), .B(
        \MC_ARK_ARC_1_3/temp1[116] ), .ZN(\MC_ARK_ARC_1_3/temp5[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_12_3  ( .A(\RI5[3][152] ), .B(n370), .ZN(
        \MC_ARK_ARC_1_3/temp4[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_12_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[182] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_12_3  ( .A(\RI5[3][86] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[62] ), .ZN(\MC_ARK_ARC_1_3/temp2[116] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_12_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[116] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[110] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[116] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_12_2  ( .A(\MC_ARK_ARC_1_3/temp5[117] ), .B(
        \MC_ARK_ARC_1_3/temp6[117] ), .ZN(\RI1[4][117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_12_2  ( .A(\MC_ARK_ARC_1_3/temp3[117] ), .B(
        \MC_ARK_ARC_1_3/temp4[117] ), .ZN(\MC_ARK_ARC_1_3/temp6[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_12_2  ( .A(\MC_ARK_ARC_1_3/temp1[117] ), .B(
        \MC_ARK_ARC_1_3/temp2[117] ), .ZN(\MC_ARK_ARC_1_3/temp5[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_12_2  ( .A(\RI5[3][153] ), .B(n279), .ZN(
        \MC_ARK_ARC_1_3/temp4[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_12_2  ( .A(\RI5[3][27] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[183] ), .ZN(\MC_ARK_ARC_1_3/temp3[117] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_12_2  ( .A(\RI5[3][87] ), .B(\RI5[3][63] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_12_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[117] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[111] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[117] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_12_1  ( .A(\MC_ARK_ARC_1_3/temp5[118] ), .B(
        \MC_ARK_ARC_1_3/temp6[118] ), .ZN(\RI1[4][118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_12_1  ( .A(\MC_ARK_ARC_1_3/temp3[118] ), .B(
        \MC_ARK_ARC_1_3/temp4[118] ), .ZN(\MC_ARK_ARC_1_3/temp6[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_12_1  ( .A(\MC_ARK_ARC_1_3/temp1[118] ), .B(
        \MC_ARK_ARC_1_3/temp2[118] ), .ZN(\MC_ARK_ARC_1_3/temp5[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_12_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[154] ), 
        .B(n368), .ZN(\MC_ARK_ARC_1_3/temp4[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_12_1  ( .A(\RI5[3][28] ), .B(\RI5[3][184] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_12_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[64] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[118] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_12_1  ( .A(\RI5[3][118] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[112] ), .ZN(\MC_ARK_ARC_1_3/temp1[118] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_12_0  ( .A(\MC_ARK_ARC_1_3/temp5[119] ), .B(
        \MC_ARK_ARC_1_3/temp6[119] ), .ZN(\RI1[4][119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_12_0  ( .A(\MC_ARK_ARC_1_3/temp3[119] ), .B(
        \MC_ARK_ARC_1_3/temp4[119] ), .ZN(\MC_ARK_ARC_1_3/temp6[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_12_0  ( .A(\MC_ARK_ARC_1_3/temp2[119] ), .B(
        \MC_ARK_ARC_1_3/temp1[119] ), .ZN(\MC_ARK_ARC_1_3/temp5[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_12_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[155] ), 
        .B(n277), .ZN(\MC_ARK_ARC_1_3/temp4[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_12_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[185] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_12_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[89] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[65] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_12_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .B(n797), .ZN(\MC_ARK_ARC_1_3/temp1[119] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_11_5  ( .A(\MC_ARK_ARC_1_3/temp5[120] ), .B(
        \MC_ARK_ARC_1_3/temp6[120] ), .ZN(\RI1[4][120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_11_5  ( .A(\MC_ARK_ARC_1_3/temp3[120] ), .B(
        \MC_ARK_ARC_1_3/temp4[120] ), .ZN(\MC_ARK_ARC_1_3/temp6[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_11_5  ( .A(\MC_ARK_ARC_1_3/temp2[120] ), .B(
        \MC_ARK_ARC_1_3/temp1[120] ), .ZN(\MC_ARK_ARC_1_3/temp5[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_11_5  ( .A(\RI5[3][156] ), .B(n367), .ZN(
        \MC_ARK_ARC_1_3/temp4[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_11_5  ( .A(\RI5[3][30] ), .B(\RI5[3][186] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_11_5  ( .A(\RI5[3][90] ), .B(\RI5[3][66] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[120] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_11_5  ( .A(\RI5[3][120] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[114] ), .ZN(\MC_ARK_ARC_1_3/temp1[120] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_11_4  ( .A(\MC_ARK_ARC_1_3/temp3[121] ), .B(
        \MC_ARK_ARC_1_3/temp4[121] ), .ZN(\MC_ARK_ARC_1_3/temp6[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_11_4  ( .A(\RI5[3][157] ), .B(n275), .ZN(
        \MC_ARK_ARC_1_3/temp4[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_11_4  ( .A(\RI5[3][31] ), .B(\RI5[3][187] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_11_4  ( .A(\MC_ARK_ARC_1_3/buf_datainput[91] ), 
        .B(\RI5[3][67] ), .ZN(\MC_ARK_ARC_1_3/temp2[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_11_4  ( .A(\RI5[3][121] ), .B(\RI5[3][115] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[121] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_11_3  ( .A(\MC_ARK_ARC_1_3/temp5[122] ), .B(
        \MC_ARK_ARC_1_3/temp6[122] ), .ZN(\RI1[4][122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_11_3  ( .A(\MC_ARK_ARC_1_3/temp3[122] ), .B(
        \MC_ARK_ARC_1_3/temp4[122] ), .ZN(\MC_ARK_ARC_1_3/temp6[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_11_3  ( .A(\MC_ARK_ARC_1_3/temp1[122] ), .B(
        \MC_ARK_ARC_1_3/temp2[122] ), .ZN(\MC_ARK_ARC_1_3/temp5[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_11_3  ( .A(n2119), .B(n365), .ZN(
        \MC_ARK_ARC_1_3/temp4[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_11_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[32] ), 
        .B(\RI5[3][188] ), .ZN(\MC_ARK_ARC_1_3/temp3[122] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_11_3  ( .A(\RI5[3][92] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[68] ), .ZN(\MC_ARK_ARC_1_3/temp2[122] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_11_3  ( .A(n1929), .B(
        \MC_ARK_ARC_1_3/buf_datainput[116] ), .ZN(\MC_ARK_ARC_1_3/temp1[122] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_11_2  ( .A(\MC_ARK_ARC_1_3/temp3[123] ), .B(
        \MC_ARK_ARC_1_3/temp4[123] ), .ZN(\MC_ARK_ARC_1_3/temp6[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_11_2  ( .A(\RI5[3][159] ), .B(n273), .ZN(
        \MC_ARK_ARC_1_3/temp4[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_11_2  ( .A(\RI5[3][33] ), .B(\RI5[3][189] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_11_2  ( .A(\RI5[3][93] ), .B(\RI5[3][69] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[123] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_11_2  ( .A(\RI5[3][123] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[117] ), .ZN(\MC_ARK_ARC_1_3/temp1[123] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_11_1  ( .A(\MC_ARK_ARC_1_3/temp3[124] ), .B(
        \MC_ARK_ARC_1_3/temp4[124] ), .ZN(\MC_ARK_ARC_1_3/temp6[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_11_1  ( .A(\MC_ARK_ARC_1_3/temp1[124] ), .B(
        \MC_ARK_ARC_1_3/temp2[124] ), .ZN(\MC_ARK_ARC_1_3/temp5[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_11_1  ( .A(\RI5[3][160] ), .B(n427), .ZN(
        \MC_ARK_ARC_1_3/temp4[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_11_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[34] ), 
        .B(\RI5[3][190] ), .ZN(\MC_ARK_ARC_1_3/temp3[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_11_1  ( .A(\RI5[3][94] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[70] ), .ZN(\MC_ARK_ARC_1_3/temp2[124] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_11_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[124] ), 
        .B(\RI5[3][118] ), .ZN(\MC_ARK_ARC_1_3/temp1[124] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_11_0  ( .A(\MC_ARK_ARC_1_3/temp5[125] ), .B(
        \MC_ARK_ARC_1_3/temp6[125] ), .ZN(\RI1[4][125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_11_0  ( .A(\MC_ARK_ARC_1_3/temp3[125] ), .B(
        \MC_ARK_ARC_1_3/temp4[125] ), .ZN(\MC_ARK_ARC_1_3/temp6[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_11_0  ( .A(\MC_ARK_ARC_1_3/temp1[125] ), .B(
        \MC_ARK_ARC_1_3/temp2[125] ), .ZN(\MC_ARK_ARC_1_3/temp5[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_11_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[161] ), 
        .B(n271), .ZN(\MC_ARK_ARC_1_3/temp4[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_11_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[35] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[191] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_11_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .B(n2145), .ZN(\MC_ARK_ARC_1_3/temp2[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_11_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .B(n521), .ZN(\MC_ARK_ARC_1_3/temp1[125] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_10_5  ( .A(\MC_ARK_ARC_1_3/temp6[126] ), .B(
        \MC_ARK_ARC_1_3/temp5[126] ), .ZN(\RI1[4][126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_10_5  ( .A(\MC_ARK_ARC_1_3/temp3[126] ), .B(
        \MC_ARK_ARC_1_3/temp4[126] ), .ZN(\MC_ARK_ARC_1_3/temp6[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_10_5  ( .A(\MC_ARK_ARC_1_3/temp1[126] ), .B(
        \MC_ARK_ARC_1_3/temp2[126] ), .ZN(\MC_ARK_ARC_1_3/temp5[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_10_5  ( .A(\RI5[3][162] ), .B(n379), .ZN(
        \MC_ARK_ARC_1_3/temp4[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_10_5  ( .A(\RI5[3][36] ), .B(\RI5[3][0] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_10_5  ( .A(\RI5[3][96] ), .B(\RI5[3][72] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_10_5  ( .A(n1654), .B(\RI5[3][120] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[126] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_10_4  ( .A(\MC_ARK_ARC_1_3/temp5[127] ), .B(
        \MC_ARK_ARC_1_3/temp6[127] ), .ZN(\RI1[4][127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_10_4  ( .A(\MC_ARK_ARC_1_3/temp3[127] ), .B(
        \MC_ARK_ARC_1_3/temp4[127] ), .ZN(\MC_ARK_ARC_1_3/temp6[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_10_4  ( .A(\MC_ARK_ARC_1_3/temp1[127] ), .B(
        \MC_ARK_ARC_1_3/temp2[127] ), .ZN(\MC_ARK_ARC_1_3/temp5[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_10_4  ( .A(\RI5[3][163] ), .B(n509), .ZN(
        \MC_ARK_ARC_1_3/temp4[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_10_4  ( .A(\RI5[3][37] ), .B(\RI5[3][1] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_10_4  ( .A(\RI5[3][97] ), .B(\RI5[3][73] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_10_4  ( .A(\RI5[3][127] ), .B(\RI5[3][121] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[127] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_10_3  ( .A(\MC_ARK_ARC_1_3/temp5[128] ), .B(
        \MC_ARK_ARC_1_3/temp6[128] ), .ZN(\RI1[4][128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_10_3  ( .A(\MC_ARK_ARC_1_3/temp3[128] ), .B(
        \MC_ARK_ARC_1_3/temp4[128] ), .ZN(\MC_ARK_ARC_1_3/temp6[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_10_3  ( .A(\MC_ARK_ARC_1_3/temp1[128] ), .B(
        \MC_ARK_ARC_1_3/temp2[128] ), .ZN(\MC_ARK_ARC_1_3/temp5[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_10_3  ( .A(\RI5[3][164] ), .B(n452), .ZN(
        \MC_ARK_ARC_1_3/temp4[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_10_3  ( .A(\RI5[3][38] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[2] ), .ZN(\MC_ARK_ARC_1_3/temp3[128] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_10_3  ( .A(\RI5[3][98] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[74] ), .ZN(\MC_ARK_ARC_1_3/temp2[128] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_10_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[128] ), 
        .B(n1928), .ZN(\MC_ARK_ARC_1_3/temp1[128] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_10_2  ( .A(\MC_ARK_ARC_1_3/temp5[129] ), .B(
        \MC_ARK_ARC_1_3/temp6[129] ), .ZN(\RI1[4][129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_10_2  ( .A(\MC_ARK_ARC_1_3/temp3[129] ), .B(
        \MC_ARK_ARC_1_3/temp4[129] ), .ZN(\MC_ARK_ARC_1_3/temp6[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_10_2  ( .A(\MC_ARK_ARC_1_3/temp2[129] ), .B(
        \MC_ARK_ARC_1_3/temp1[129] ), .ZN(\MC_ARK_ARC_1_3/temp5[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_10_2  ( .A(\RI5[3][165] ), .B(n396), .ZN(
        \MC_ARK_ARC_1_3/temp4[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_10_2  ( .A(\RI5[3][39] ), .B(\RI5[3][3] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_10_2  ( .A(\RI5[3][99] ), .B(\RI5[3][75] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_10_2  ( .A(\RI5[3][129] ), .B(\RI5[3][123] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[129] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_10_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[166] ), 
        .B(n357), .ZN(\MC_ARK_ARC_1_3/temp4[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_10_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[40] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_10_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[76] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[130] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_10_1  ( .A(n1944), .B(
        \MC_ARK_ARC_1_3/buf_datainput[124] ), .ZN(\MC_ARK_ARC_1_3/temp1[130] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_10_0  ( .A(n1948), .B(n265), .ZN(
        \MC_ARK_ARC_1_3/temp4[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_10_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .B(n2111), .ZN(\MC_ARK_ARC_1_3/temp3[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_10_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[77] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_10_0  ( .A(n801), .B(n521), .ZN(
        \MC_ARK_ARC_1_3/temp1[131] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_9_5  ( .A(\MC_ARK_ARC_1_3/temp5[132] ), .B(
        \MC_ARK_ARC_1_3/temp6[132] ), .ZN(\RI1[4][132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_9_5  ( .A(\MC_ARK_ARC_1_3/temp3[132] ), .B(
        \MC_ARK_ARC_1_3/temp4[132] ), .ZN(\MC_ARK_ARC_1_3/temp6[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_9_5  ( .A(\MC_ARK_ARC_1_3/temp2[132] ), .B(
        \MC_ARK_ARC_1_3/temp1[132] ), .ZN(\MC_ARK_ARC_1_3/temp5[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_9_5  ( .A(\RI5[3][168] ), .B(n478), .ZN(
        \MC_ARK_ARC_1_3/temp4[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_9_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[42] ), 
        .B(\RI5[3][6] ), .ZN(\MC_ARK_ARC_1_3/temp3[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_9_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .B(\RI5[3][78] ), .ZN(\MC_ARK_ARC_1_3/temp2[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_9_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[132] ), 
        .B(n1654), .ZN(\MC_ARK_ARC_1_3/temp1[132] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_9_4  ( .A(\MC_ARK_ARC_1_3/temp5[133] ), .B(
        \MC_ARK_ARC_1_3/temp6[133] ), .ZN(\RI1[4][133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_9_4  ( .A(\MC_ARK_ARC_1_3/temp3[133] ), .B(
        \MC_ARK_ARC_1_3/temp4[133] ), .ZN(\MC_ARK_ARC_1_3/temp6[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_9_4  ( .A(\MC_ARK_ARC_1_3/temp1[133] ), .B(
        \MC_ARK_ARC_1_3/temp2[133] ), .ZN(\MC_ARK_ARC_1_3/temp5[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_9_4  ( .A(\RI5[3][169] ), .B(n263), .ZN(
        \MC_ARK_ARC_1_3/temp4[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_9_4  ( .A(\RI5[3][43] ), .B(\RI5[3][7] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_9_4  ( .A(\RI5[3][103] ), .B(\RI5[3][79] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_9_4  ( .A(\RI5[3][133] ), .B(\RI5[3][127] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[133] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_9_3  ( .A(\MC_ARK_ARC_1_3/temp5[134] ), .B(
        \MC_ARK_ARC_1_3/temp6[134] ), .ZN(\RI1[4][134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_9_3  ( .A(\MC_ARK_ARC_1_3/temp3[134] ), .B(
        \MC_ARK_ARC_1_3/temp4[134] ), .ZN(\MC_ARK_ARC_1_3/temp6[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_9_3  ( .A(\MC_ARK_ARC_1_3/temp1[134] ), .B(
        \MC_ARK_ARC_1_3/temp2[134] ), .ZN(\MC_ARK_ARC_1_3/temp5[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_9_3  ( .A(\RI5[3][170] ), .B(n447), .ZN(
        \MC_ARK_ARC_1_3/temp4[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_9_3  ( .A(\RI5[3][44] ), .B(\RI5[3][8] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_9_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[104] ), 
        .B(\RI5[3][80] ), .ZN(\MC_ARK_ARC_1_3/temp2[134] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_9_3  ( .A(\RI5[3][134] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[128] ), .ZN(\MC_ARK_ARC_1_3/temp1[134] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_9_2  ( .A(\MC_ARK_ARC_1_3/temp5[135] ), .B(
        \MC_ARK_ARC_1_3/temp6[135] ), .ZN(\RI1[4][135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_9_2  ( .A(\MC_ARK_ARC_1_3/temp3[135] ), .B(
        \MC_ARK_ARC_1_3/temp4[135] ), .ZN(\MC_ARK_ARC_1_3/temp6[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_9_2  ( .A(\MC_ARK_ARC_1_3/temp2[135] ), .B(
        \MC_ARK_ARC_1_3/temp1[135] ), .ZN(\MC_ARK_ARC_1_3/temp5[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_9_2  ( .A(\RI5[3][171] ), .B(n261), .ZN(
        \MC_ARK_ARC_1_3/temp4[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_9_2  ( .A(\RI5[3][45] ), .B(\RI5[3][9] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_9_2  ( .A(\RI5[3][105] ), .B(\RI5[3][81] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_9_2  ( .A(\RI5[3][135] ), .B(\RI5[3][129] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[135] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_9_1  ( .A(\MC_ARK_ARC_1_3/temp5[136] ), .B(
        \MC_ARK_ARC_1_3/temp6[136] ), .ZN(\RI1[4][136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_9_1  ( .A(\MC_ARK_ARC_1_3/temp3[136] ), .B(
        \MC_ARK_ARC_1_3/temp4[136] ), .ZN(\MC_ARK_ARC_1_3/temp6[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_9_1  ( .A(\MC_ARK_ARC_1_3/temp1[136] ), .B(
        \MC_ARK_ARC_1_3/temp2[136] ), .ZN(\MC_ARK_ARC_1_3/temp5[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_9_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[172] ), 
        .B(n351), .ZN(\MC_ARK_ARC_1_3/temp4[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_9_1  ( .A(\RI5[3][46] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[10] ), .ZN(\MC_ARK_ARC_1_3/temp3[136] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_9_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[106] ), 
        .B(\RI5[3][82] ), .ZN(\MC_ARK_ARC_1_3/temp2[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_9_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[136] ), 
        .B(n1943), .ZN(\MC_ARK_ARC_1_3/temp1[136] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_9_0  ( .A(\MC_ARK_ARC_1_3/temp5[137] ), .B(
        \MC_ARK_ARC_1_3/temp6[137] ), .ZN(\RI1[4][137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_9_0  ( .A(\MC_ARK_ARC_1_3/temp4[137] ), .B(
        \MC_ARK_ARC_1_3/temp3[137] ), .ZN(\MC_ARK_ARC_1_3/temp6[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_9_0  ( .A(\MC_ARK_ARC_1_3/temp2[137] ), .B(
        \MC_ARK_ARC_1_3/temp1[137] ), .ZN(\MC_ARK_ARC_1_3/temp5[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_9_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[173] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[137] ), .ZN(
        \MC_ARK_ARC_1_3/temp4[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_9_0  ( .A(n1650), .B(
        \MC_ARK_ARC_1_3/buf_datainput[47] ), .ZN(\MC_ARK_ARC_1_3/temp3[137] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_9_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[83] ), 
        .B(n2108), .ZN(\MC_ARK_ARC_1_3/temp2[137] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_9_0  ( .A(n784), .B(
        \MC_ARK_ARC_1_3/buf_datainput[131] ), .ZN(\MC_ARK_ARC_1_3/temp1[137] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_8_5  ( .A(\MC_ARK_ARC_1_3/temp5[138] ), .B(
        \MC_ARK_ARC_1_3/temp6[138] ), .ZN(\RI1[4][138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_8_5  ( .A(\MC_ARK_ARC_1_3/temp3[138] ), .B(
        \MC_ARK_ARC_1_3/temp4[138] ), .ZN(\MC_ARK_ARC_1_3/temp6[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_8_5  ( .A(\MC_ARK_ARC_1_3/temp2[138] ), .B(
        \MC_ARK_ARC_1_3/temp1[138] ), .ZN(\MC_ARK_ARC_1_3/temp5[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_8_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .B(n349), .ZN(\MC_ARK_ARC_1_3/temp4[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_8_5  ( .A(\RI5[3][48] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[12] ), .ZN(\MC_ARK_ARC_1_3/temp3[138] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_8_5  ( .A(\RI5[3][108] ), .B(n2130), .ZN(
        \MC_ARK_ARC_1_3/temp2[138] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_8_5  ( .A(n818), .B(
        \MC_ARK_ARC_1_3/buf_datainput[132] ), .ZN(\MC_ARK_ARC_1_3/temp1[138] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_8_4  ( .A(\MC_ARK_ARC_1_3/temp5[139] ), .B(
        \MC_ARK_ARC_1_3/temp6[139] ), .ZN(\RI1[4][139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_8_4  ( .A(\MC_ARK_ARC_1_3/temp3[139] ), .B(
        \MC_ARK_ARC_1_3/temp4[139] ), .ZN(\MC_ARK_ARC_1_3/temp6[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_8_4  ( .A(\MC_ARK_ARC_1_3/temp1[139] ), .B(
        \MC_ARK_ARC_1_3/temp2[139] ), .ZN(\MC_ARK_ARC_1_3/temp5[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_8_4  ( .A(\RI5[3][175] ), .B(n492), .ZN(
        \MC_ARK_ARC_1_3/temp4[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_8_4  ( .A(\RI5[3][49] ), .B(\RI5[3][13] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_8_4  ( .A(\RI5[3][109] ), .B(\RI5[3][85] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_8_4  ( .A(\RI5[3][139] ), .B(\RI5[3][133] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[139] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_8_3  ( .A(\MC_ARK_ARC_1_3/temp5[140] ), .B(
        \MC_ARK_ARC_1_3/temp6[140] ), .ZN(\RI1[4][140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_8_3  ( .A(\MC_ARK_ARC_1_3/temp3[140] ), .B(
        \MC_ARK_ARC_1_3/temp4[140] ), .ZN(\MC_ARK_ARC_1_3/temp6[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_8_3  ( .A(\MC_ARK_ARC_1_3/temp1[140] ), .B(
        \MC_ARK_ARC_1_3/temp2[140] ), .ZN(\MC_ARK_ARC_1_3/temp5[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_8_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .B(n347), .ZN(\MC_ARK_ARC_1_3/temp4[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_8_3  ( .A(n2129), .B(
        \MC_ARK_ARC_1_3/buf_datainput[14] ), .ZN(\MC_ARK_ARC_1_3/temp3[140] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_8_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[110] ), 
        .B(\RI5[3][86] ), .ZN(\MC_ARK_ARC_1_3/temp2[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_8_3  ( .A(\RI5[3][140] ), .B(\RI5[3][134] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[140] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_8_2  ( .A(\MC_ARK_ARC_1_3/temp5[141] ), .B(
        \MC_ARK_ARC_1_3/temp6[141] ), .ZN(\RI1[4][141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_8_2  ( .A(\MC_ARK_ARC_1_3/temp3[141] ), .B(
        \MC_ARK_ARC_1_3/temp4[141] ), .ZN(\MC_ARK_ARC_1_3/temp6[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_8_2  ( .A(\MC_ARK_ARC_1_3/temp1[141] ), .B(
        \MC_ARK_ARC_1_3/temp2[141] ), .ZN(\MC_ARK_ARC_1_3/temp5[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_8_2  ( .A(\RI5[3][177] ), .B(n255), .ZN(
        \MC_ARK_ARC_1_3/temp4[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_8_2  ( .A(\RI5[3][51] ), .B(\RI5[3][15] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_8_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[111] ), 
        .B(\RI5[3][87] ), .ZN(\MC_ARK_ARC_1_3/temp2[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_8_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[141] ), 
        .B(\RI5[3][135] ), .ZN(\MC_ARK_ARC_1_3/temp1[141] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_8_1  ( .A(\MC_ARK_ARC_1_3/temp5[142] ), .B(
        \MC_ARK_ARC_1_3/temp6[142] ), .ZN(\RI1[4][142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_8_1  ( .A(\MC_ARK_ARC_1_3/temp3[142] ), .B(
        \MC_ARK_ARC_1_3/temp4[142] ), .ZN(\MC_ARK_ARC_1_3/temp6[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_8_1  ( .A(\MC_ARK_ARC_1_3/temp1[142] ), .B(
        \MC_ARK_ARC_1_3/temp2[142] ), .ZN(\MC_ARK_ARC_1_3/temp5[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_8_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[142] ), .ZN(
        \MC_ARK_ARC_1_3/temp4[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_8_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[52] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[16] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_8_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[112] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[88] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_8_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[136] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[142] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_8_0  ( .A(\MC_ARK_ARC_1_3/temp6[143] ), .B(
        \MC_ARK_ARC_1_3/temp5[143] ), .ZN(\RI1[4][143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_8_0  ( .A(\MC_ARK_ARC_1_3/temp3[143] ), .B(
        \MC_ARK_ARC_1_3/temp4[143] ), .ZN(\MC_ARK_ARC_1_3/temp6[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_8_0  ( .A(\MC_ARK_ARC_1_3/temp2[143] ), .B(
        \MC_ARK_ARC_1_3/temp1[143] ), .ZN(\MC_ARK_ARC_1_3/temp5[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_8_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .B(n253), .ZN(\MC_ARK_ARC_1_3/temp4[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_8_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[53] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_8_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[89] ), 
        .B(n796), .ZN(\MC_ARK_ARC_1_3/temp2[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_8_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[137] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[143] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[143] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_7_5  ( .A(\MC_ARK_ARC_1_3/temp5[144] ), .B(
        \MC_ARK_ARC_1_3/temp6[144] ), .ZN(\RI1[4][144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_7_5  ( .A(\MC_ARK_ARC_1_3/temp3[144] ), .B(
        \MC_ARK_ARC_1_3/temp4[144] ), .ZN(\MC_ARK_ARC_1_3/temp6[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_7_5  ( .A(\MC_ARK_ARC_1_3/temp2[144] ), .B(
        \MC_ARK_ARC_1_3/temp1[144] ), .ZN(\MC_ARK_ARC_1_3/temp5[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_7_5  ( .A(\RI5[3][180] ), .B(n343), .ZN(
        \MC_ARK_ARC_1_3/temp4[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_7_5  ( .A(\RI5[3][54] ), .B(\RI5[3][18] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_7_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[114] ), 
        .B(\RI5[3][90] ), .ZN(\MC_ARK_ARC_1_3/temp2[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_7_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[144] ), 
        .B(\RI5[3][138] ), .ZN(\MC_ARK_ARC_1_3/temp1[144] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_7_4  ( .A(\MC_ARK_ARC_1_3/temp5[145] ), .B(
        \MC_ARK_ARC_1_3/temp6[145] ), .ZN(\RI1[4][145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_7_4  ( .A(\MC_ARK_ARC_1_3/temp3[145] ), .B(
        \MC_ARK_ARC_1_3/temp4[145] ), .ZN(\MC_ARK_ARC_1_3/temp6[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_7_4  ( .A(\MC_ARK_ARC_1_3/temp1[145] ), .B(
        \MC_ARK_ARC_1_3/temp2[145] ), .ZN(\MC_ARK_ARC_1_3/temp5[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_7_4  ( .A(\RI5[3][181] ), .B(n251), .ZN(
        \MC_ARK_ARC_1_3/temp4[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_7_4  ( .A(\RI5[3][55] ), .B(\RI5[3][19] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_7_4  ( .A(\RI5[3][115] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[91] ), .ZN(\MC_ARK_ARC_1_3/temp2[145] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_7_4  ( .A(\RI5[3][145] ), .B(\RI5[3][139] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[145] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_7_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .B(n341), .ZN(\MC_ARK_ARC_1_3/temp4[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_7_3  ( .A(\RI5[3][56] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[20] ), .ZN(\MC_ARK_ARC_1_3/temp3[146] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_7_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[116] ), 
        .B(\RI5[3][92] ), .ZN(\MC_ARK_ARC_1_3/temp2[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_7_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[146] ), 
        .B(\RI5[3][140] ), .ZN(\MC_ARK_ARC_1_3/temp1[146] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_7_2  ( .A(\MC_ARK_ARC_1_3/temp3[147] ), .B(
        \MC_ARK_ARC_1_3/temp4[147] ), .ZN(\MC_ARK_ARC_1_3/temp6[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_7_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[183] ), 
        .B(n250), .ZN(\MC_ARK_ARC_1_3/temp4[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_7_2  ( .A(\RI5[3][57] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[21] ), .ZN(\MC_ARK_ARC_1_3/temp3[147] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_7_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[117] ), 
        .B(\RI5[3][93] ), .ZN(\MC_ARK_ARC_1_3/temp2[147] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_7_2  ( .A(\RI5[3][147] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[141] ), .ZN(\MC_ARK_ARC_1_3/temp1[147] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_7_1  ( .A(\MC_ARK_ARC_1_3/temp6[148] ), .B(
        \MC_ARK_ARC_1_3/temp5[148] ), .ZN(\RI1[4][148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_7_1  ( .A(\MC_ARK_ARC_1_3/temp3[148] ), .B(
        \MC_ARK_ARC_1_3/temp4[148] ), .ZN(\MC_ARK_ARC_1_3/temp6[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_7_1  ( .A(\MC_ARK_ARC_1_3/temp2[148] ), .B(
        \MC_ARK_ARC_1_3/temp1[148] ), .ZN(\MC_ARK_ARC_1_3/temp5[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_7_1  ( .A(\RI5[3][184] ), .B(n340), .ZN(
        \MC_ARK_ARC_1_3/temp4[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_7_1  ( .A(n2102), .B(
        \MC_ARK_ARC_1_3/buf_datainput[22] ), .ZN(\MC_ARK_ARC_1_3/temp3[148] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_7_1  ( .A(\RI5[3][118] ), .B(\RI5[3][94] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[148] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_7_1  ( .A(n1510), .B(
        \MC_ARK_ARC_1_3/buf_datainput[142] ), .ZN(\MC_ARK_ARC_1_3/temp1[148] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_7_0  ( .A(\MC_ARK_ARC_1_3/temp6[149] ), .B(
        \MC_ARK_ARC_1_3/temp5[149] ), .ZN(\RI1[4][149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_7_0  ( .A(\MC_ARK_ARC_1_3/temp3[149] ), .B(
        \MC_ARK_ARC_1_3/temp4[149] ), .ZN(\MC_ARK_ARC_1_3/temp6[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_7_0  ( .A(\MC_ARK_ARC_1_3/temp2[149] ), .B(
        \MC_ARK_ARC_1_3/temp1[149] ), .ZN(\MC_ARK_ARC_1_3/temp5[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_7_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[185] ), 
        .B(Key[133]), .ZN(\MC_ARK_ARC_1_3/temp4[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_7_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[59] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[23] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_7_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[95] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[149] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_7_0  ( .A(n849), .B(
        \MC_ARK_ARC_1_3/buf_datainput[143] ), .ZN(\MC_ARK_ARC_1_3/temp1[149] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_6_5  ( .A(\MC_ARK_ARC_1_3/temp6[150] ), .B(
        \MC_ARK_ARC_1_3/temp5[150] ), .ZN(\RI1[4][150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_6_5  ( .A(\MC_ARK_ARC_1_3/temp3[150] ), .B(
        \MC_ARK_ARC_1_3/temp4[150] ), .ZN(\MC_ARK_ARC_1_3/temp6[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_6_5  ( .A(\MC_ARK_ARC_1_3/temp2[150] ), .B(
        \MC_ARK_ARC_1_3/temp1[150] ), .ZN(\MC_ARK_ARC_1_3/temp5[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_6_5  ( .A(\RI5[3][186] ), .B(n338), .ZN(
        \MC_ARK_ARC_1_3/temp4[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_6_5  ( .A(\RI5[3][60] ), .B(\RI5[3][24] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_6_5  ( .A(\RI5[3][120] ), .B(\RI5[3][96] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[150] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_6_5  ( .A(\RI5[3][150] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[144] ), .ZN(\MC_ARK_ARC_1_3/temp1[150] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_6_4  ( .A(\MC_ARK_ARC_1_3/temp5[151] ), .B(
        \MC_ARK_ARC_1_3/temp6[151] ), .ZN(\RI1[4][151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_6_4  ( .A(\MC_ARK_ARC_1_3/temp3[151] ), .B(
        \MC_ARK_ARC_1_3/temp4[151] ), .ZN(\MC_ARK_ARC_1_3/temp6[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_6_4  ( .A(\MC_ARK_ARC_1_3/temp1[151] ), .B(
        \MC_ARK_ARC_1_3/temp2[151] ), .ZN(\MC_ARK_ARC_1_3/temp5[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_6_4  ( .A(\RI5[3][187] ), .B(n246), .ZN(
        \MC_ARK_ARC_1_3/temp4[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_6_4  ( .A(\RI5[3][61] ), .B(\RI5[3][25] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_6_4  ( .A(\RI5[3][121] ), .B(\RI5[3][97] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_6_4  ( .A(\RI5[3][151] ), .B(\RI5[3][145] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[151] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_6_3  ( .A(\MC_ARK_ARC_1_3/temp5[152] ), .B(
        \MC_ARK_ARC_1_3/temp6[152] ), .ZN(\RI1[4][152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_6_3  ( .A(\MC_ARK_ARC_1_3/temp3[152] ), .B(
        \MC_ARK_ARC_1_3/temp4[152] ), .ZN(\MC_ARK_ARC_1_3/temp6[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_6_3  ( .A(\MC_ARK_ARC_1_3/temp1[152] ), .B(
        \MC_ARK_ARC_1_3/temp2[152] ), .ZN(\MC_ARK_ARC_1_3/temp5[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_6_3  ( .A(\RI5[3][188] ), .B(n469), .ZN(
        \MC_ARK_ARC_1_3/temp4[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_6_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[26] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[62] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_6_3  ( .A(n1929), .B(\RI5[3][98] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[152] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_6_3  ( .A(\RI5[3][152] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[146] ), .ZN(\MC_ARK_ARC_1_3/temp1[152] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_6_2  ( .A(\MC_ARK_ARC_1_3/temp5[153] ), .B(
        \MC_ARK_ARC_1_3/temp6[153] ), .ZN(\RI1[4][153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_6_2  ( .A(\MC_ARK_ARC_1_3/temp3[153] ), .B(
        \MC_ARK_ARC_1_3/temp4[153] ), .ZN(\MC_ARK_ARC_1_3/temp6[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_6_2  ( .A(\MC_ARK_ARC_1_3/temp1[153] ), .B(
        \MC_ARK_ARC_1_3/temp2[153] ), .ZN(\MC_ARK_ARC_1_3/temp5[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_6_2  ( .A(\RI5[3][189] ), .B(n408), .ZN(
        \MC_ARK_ARC_1_3/temp4[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_6_2  ( .A(\RI5[3][63] ), .B(\RI5[3][27] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_6_2  ( .A(\RI5[3][123] ), .B(\RI5[3][99] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_6_2  ( .A(\RI5[3][147] ), .B(\RI5[3][153] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[153] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_6_1  ( .A(\MC_ARK_ARC_1_3/temp6[154] ), .B(
        \MC_ARK_ARC_1_3/temp5[154] ), .ZN(\RI1[4][154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_6_1  ( .A(\MC_ARK_ARC_1_3/temp3[154] ), .B(
        \MC_ARK_ARC_1_3/temp4[154] ), .ZN(\MC_ARK_ARC_1_3/temp6[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_6_1  ( .A(\MC_ARK_ARC_1_3/temp2[154] ), .B(
        \MC_ARK_ARC_1_3/temp1[154] ), .ZN(\MC_ARK_ARC_1_3/temp5[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_6_1  ( .A(\RI5[3][190] ), .B(
        \MC_ARK_ARC_1_3/buf_keyinput[154] ), .ZN(\MC_ARK_ARC_1_3/temp4[154] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_6_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[64] ), 
        .B(\RI5[3][28] ), .ZN(\MC_ARK_ARC_1_3/temp3[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_6_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[124] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[100] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_6_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[154] ), 
        .B(n1510), .ZN(\MC_ARK_ARC_1_3/temp1[154] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_6_0  ( .A(\MC_ARK_ARC_1_3/temp5[155] ), .B(
        \MC_ARK_ARC_1_3/temp6[155] ), .ZN(\RI1[4][155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_6_0  ( .A(\MC_ARK_ARC_1_3/temp3[155] ), .B(
        \MC_ARK_ARC_1_3/temp4[155] ), .ZN(\MC_ARK_ARC_1_3/temp6[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_6_0  ( .A(\MC_ARK_ARC_1_3/temp2[155] ), .B(
        \MC_ARK_ARC_1_3/temp1[155] ), .ZN(\MC_ARK_ARC_1_3/temp5[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_6_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[191] ), 
        .B(n243), .ZN(\MC_ARK_ARC_1_3/temp4[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_6_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .B(n2112), .ZN(\MC_ARK_ARC_1_3/temp3[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_6_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .B(n521), .ZN(\MC_ARK_ARC_1_3/temp2[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_6_0  ( .A(n850), .B(n2120), .ZN(
        \MC_ARK_ARC_1_3/temp1[155] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_5_5  ( .A(\MC_ARK_ARC_1_3/temp6[156] ), .B(
        \MC_ARK_ARC_1_3/temp5[156] ), .ZN(\RI1[4][156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_5_5  ( .A(\MC_ARK_ARC_1_3/temp3[156] ), .B(
        \MC_ARK_ARC_1_3/temp4[156] ), .ZN(\MC_ARK_ARC_1_3/temp6[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_5_5  ( .A(\MC_ARK_ARC_1_3/temp1[156] ), .B(
        \MC_ARK_ARC_1_3/temp2[156] ), .ZN(\MC_ARK_ARC_1_3/temp5[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_5_5  ( .A(\RI5[3][0] ), .B(n333), .ZN(
        \MC_ARK_ARC_1_3/temp4[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_5_5  ( .A(\RI5[3][66] ), .B(\RI5[3][30] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_5_5  ( .A(n1654), .B(
        \MC_ARK_ARC_1_3/buf_datainput[102] ), .ZN(\MC_ARK_ARC_1_3/temp2[156] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_5_5  ( .A(\RI5[3][156] ), .B(\RI5[3][150] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[156] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_5_4  ( .A(\MC_ARK_ARC_1_3/temp5[157] ), .B(
        \MC_ARK_ARC_1_3/temp6[157] ), .ZN(\RI1[4][157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_5_4  ( .A(\MC_ARK_ARC_1_3/temp3[157] ), .B(
        \MC_ARK_ARC_1_3/temp4[157] ), .ZN(\MC_ARK_ARC_1_3/temp6[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_5_4  ( .A(\MC_ARK_ARC_1_3/temp1[157] ), .B(
        \MC_ARK_ARC_1_3/temp2[157] ), .ZN(\MC_ARK_ARC_1_3/temp5[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_5_4  ( .A(\RI5[3][1] ), .B(n513), .ZN(
        \MC_ARK_ARC_1_3/temp4[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_5_4  ( .A(\RI5[3][67] ), .B(\RI5[3][31] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_5_4  ( .A(\RI5[3][127] ), .B(\RI5[3][103] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_5_4  ( .A(\RI5[3][157] ), .B(\RI5[3][151] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[157] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_5_3  ( .A(\MC_ARK_ARC_1_3/temp5[158] ), .B(
        \MC_ARK_ARC_1_3/temp6[158] ), .ZN(\RI1[4][158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_5_3  ( .A(\MC_ARK_ARC_1_3/temp3[158] ), .B(
        \MC_ARK_ARC_1_3/temp4[158] ), .ZN(\MC_ARK_ARC_1_3/temp6[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_5_3  ( .A(\MC_ARK_ARC_1_3/temp2[158] ), .B(
        \MC_ARK_ARC_1_3/temp1[158] ), .ZN(\MC_ARK_ARC_1_3/temp5[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_5_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[2] ), 
        .B(n462), .ZN(\MC_ARK_ARC_1_3/temp4[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_5_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[68] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[32] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_5_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[128] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[104] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_5_3  ( .A(n1955), .B(\RI5[3][152] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[158] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_5_2  ( .A(\MC_ARK_ARC_1_3/temp5[159] ), .B(
        \MC_ARK_ARC_1_3/temp6[159] ), .ZN(\RI1[4][159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_5_2  ( .A(\MC_ARK_ARC_1_3/temp3[159] ), .B(
        \MC_ARK_ARC_1_3/temp4[159] ), .ZN(\MC_ARK_ARC_1_3/temp6[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_5_2  ( .A(\MC_ARK_ARC_1_3/temp1[159] ), .B(
        \MC_ARK_ARC_1_3/temp2[159] ), .ZN(\MC_ARK_ARC_1_3/temp5[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_5_2  ( .A(\RI5[3][3] ), .B(n240), .ZN(
        \MC_ARK_ARC_1_3/temp4[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_5_2  ( .A(\RI5[3][69] ), .B(\RI5[3][33] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_5_2  ( .A(\RI5[3][129] ), .B(\RI5[3][105] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_5_2  ( .A(\RI5[3][159] ), .B(\RI5[3][153] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[159] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_5_1  ( .A(\MC_ARK_ARC_1_3/temp5[160] ), .B(
        \MC_ARK_ARC_1_3/temp6[160] ), .ZN(\RI1[4][160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_5_1  ( .A(\MC_ARK_ARC_1_3/temp3[160] ), .B(
        \MC_ARK_ARC_1_3/temp4[160] ), .ZN(\MC_ARK_ARC_1_3/temp6[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_5_1  ( .A(\MC_ARK_ARC_1_3/temp2[160] ), .B(
        \MC_ARK_ARC_1_3/temp1[160] ), .ZN(\MC_ARK_ARC_1_3/temp5[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_5_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[4] ), 
        .B(\MC_ARK_ARC_1_1/buf_keyinput[8] ), .ZN(\MC_ARK_ARC_1_3/temp4[160] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_5_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[70] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[34] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[160] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_5_1  ( .A(n1944), .B(
        \MC_ARK_ARC_1_3/buf_datainput[106] ), .ZN(\MC_ARK_ARC_1_3/temp2[160] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_5_1  ( .A(\RI5[3][160] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[154] ), .ZN(\MC_ARK_ARC_1_3/temp1[160] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_5_0  ( .A(\MC_ARK_ARC_1_3/temp5[161] ), .B(
        \MC_ARK_ARC_1_3/temp6[161] ), .ZN(\RI1[4][161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_5_0  ( .A(\MC_ARK_ARC_1_3/temp3[161] ), .B(
        \MC_ARK_ARC_1_3/temp4[161] ), .ZN(\MC_ARK_ARC_1_3/temp6[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_5_0  ( .A(\MC_ARK_ARC_1_3/temp1[161] ), .B(
        \MC_ARK_ARC_1_3/temp2[161] ), .ZN(\MC_ARK_ARC_1_3/temp5[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_5_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .B(n238), .ZN(\MC_ARK_ARC_1_3/temp4[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_5_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[35] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[71] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_5_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[107] ), 
        .B(n801), .ZN(\MC_ARK_ARC_1_3/temp2[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_5_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[155] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[161] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[161] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_4_5  ( .A(\MC_ARK_ARC_1_3/temp5[162] ), .B(
        \MC_ARK_ARC_1_3/temp6[162] ), .ZN(\RI1[4][162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_4_5  ( .A(\MC_ARK_ARC_1_3/temp3[162] ), .B(
        \MC_ARK_ARC_1_3/temp4[162] ), .ZN(\MC_ARK_ARC_1_3/temp6[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_4_5  ( .A(\MC_ARK_ARC_1_3/temp1[162] ), .B(
        \MC_ARK_ARC_1_3/temp2[162] ), .ZN(\MC_ARK_ARC_1_3/temp5[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_4_5  ( .A(\RI5[3][6] ), .B(n327), .ZN(
        \MC_ARK_ARC_1_3/temp4[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_4_5  ( .A(\RI5[3][72] ), .B(\RI5[3][36] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_4_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[132] ), 
        .B(\RI5[3][108] ), .ZN(\MC_ARK_ARC_1_3/temp2[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_4_5  ( .A(\RI5[3][162] ), .B(\RI5[3][156] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[162] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_4_4  ( .A(\MC_ARK_ARC_1_3/temp5[163] ), .B(
        \MC_ARK_ARC_1_3/temp6[163] ), .ZN(\RI1[4][163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_4_4  ( .A(\MC_ARK_ARC_1_3/temp3[163] ), .B(
        \MC_ARK_ARC_1_3/temp4[163] ), .ZN(\MC_ARK_ARC_1_3/temp6[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_4_4  ( .A(\MC_ARK_ARC_1_3/temp1[163] ), .B(
        \MC_ARK_ARC_1_3/temp2[163] ), .ZN(\MC_ARK_ARC_1_3/temp5[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_4_4  ( .A(\RI5[3][7] ), .B(n507), .ZN(
        \MC_ARK_ARC_1_3/temp4[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_4_4  ( .A(\RI5[3][73] ), .B(\RI5[3][37] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_4_4  ( .A(\RI5[3][133] ), .B(\RI5[3][109] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_4_4  ( .A(\RI5[3][163] ), .B(\RI5[3][157] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[163] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_4_3  ( .A(\MC_ARK_ARC_1_3/temp5[164] ), .B(
        \MC_ARK_ARC_1_3/temp6[164] ), .ZN(\RI1[4][164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_4_3  ( .A(\MC_ARK_ARC_1_3/temp3[164] ), .B(
        \MC_ARK_ARC_1_3/temp4[164] ), .ZN(\MC_ARK_ARC_1_3/temp6[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_4_3  ( .A(\MC_ARK_ARC_1_3/temp2[164] ), .B(
        \MC_ARK_ARC_1_3/temp1[164] ), .ZN(\MC_ARK_ARC_1_3/temp5[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_4_3  ( .A(\RI5[3][8] ), .B(n375), .ZN(
        \MC_ARK_ARC_1_3/temp4[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_4_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .B(\RI5[3][38] ), .ZN(\MC_ARK_ARC_1_3/temp3[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_4_3  ( .A(\RI5[3][134] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[110] ), .ZN(\MC_ARK_ARC_1_3/temp2[164] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_4_3  ( .A(n1626), .B(n1955), .ZN(
        \MC_ARK_ARC_1_3/temp1[164] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_4_2  ( .A(\MC_ARK_ARC_1_3/temp5[165] ), .B(
        \MC_ARK_ARC_1_3/temp6[165] ), .ZN(\RI1[4][165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_4_2  ( .A(\MC_ARK_ARC_1_3/temp3[165] ), .B(
        \MC_ARK_ARC_1_3/temp4[165] ), .ZN(\MC_ARK_ARC_1_3/temp6[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_4_2  ( .A(\MC_ARK_ARC_1_3/temp1[165] ), .B(
        \MC_ARK_ARC_1_3/temp2[165] ), .ZN(\MC_ARK_ARC_1_3/temp5[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_4_2  ( .A(\RI5[3][9] ), .B(n234), .ZN(
        \MC_ARK_ARC_1_3/temp4[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_4_2  ( .A(\RI5[3][75] ), .B(\RI5[3][39] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_4_2  ( .A(\RI5[3][135] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[111] ), .ZN(\MC_ARK_ARC_1_3/temp2[165] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_4_2  ( .A(\RI5[3][165] ), .B(\RI5[3][159] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[165] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_4_1  ( .A(\MC_ARK_ARC_1_3/temp5[166] ), .B(
        \MC_ARK_ARC_1_3/temp6[166] ), .ZN(\RI1[4][166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_4_1  ( .A(\MC_ARK_ARC_1_3/temp3[166] ), .B(
        \MC_ARK_ARC_1_3/temp4[166] ), .ZN(\MC_ARK_ARC_1_3/temp6[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_4_1  ( .A(\MC_ARK_ARC_1_3/temp1[166] ), .B(
        \MC_ARK_ARC_1_3/temp2[166] ), .ZN(\MC_ARK_ARC_1_3/temp5[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_4_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[10] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[166] ), .ZN(
        \MC_ARK_ARC_1_3/temp4[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_4_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[76] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[40] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_4_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[136] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[112] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_4_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[166] ), 
        .B(\RI5[3][160] ), .ZN(\MC_ARK_ARC_1_3/temp1[166] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_4_0  ( .A(n1650), .B(n232), .ZN(
        \MC_ARK_ARC_1_3/temp4[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_4_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[77] ), 
        .B(\RI5[3][41] ), .ZN(\MC_ARK_ARC_1_3/temp3[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_4_0  ( .A(n797), .B(n784), .ZN(
        \MC_ARK_ARC_1_3/temp2[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_4_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[161] ), 
        .B(n1947), .ZN(\MC_ARK_ARC_1_3/temp1[167] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_3_5  ( .A(\MC_ARK_ARC_1_3/temp5[168] ), .B(
        \MC_ARK_ARC_1_3/temp6[168] ), .ZN(\RI1[4][168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_3_5  ( .A(\MC_ARK_ARC_1_3/temp3[168] ), .B(
        \MC_ARK_ARC_1_3/temp4[168] ), .ZN(\MC_ARK_ARC_1_3/temp6[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_3_5  ( .A(\MC_ARK_ARC_1_3/temp1[168] ), .B(
        \MC_ARK_ARC_1_3/temp2[168] ), .ZN(\MC_ARK_ARC_1_3/temp5[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_3_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[12] ), 
        .B(n321), .ZN(\MC_ARK_ARC_1_3/temp4[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_3_5  ( .A(\RI5[3][78] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[42] ), .ZN(\MC_ARK_ARC_1_3/temp3[168] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_3_5  ( .A(n818), .B(
        \MC_ARK_ARC_1_3/buf_datainput[114] ), .ZN(\MC_ARK_ARC_1_3/temp2[168] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_3_5  ( .A(\RI5[3][168] ), .B(\RI5[3][162] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[168] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_3_4  ( .A(\MC_ARK_ARC_1_3/temp5[169] ), .B(
        \MC_ARK_ARC_1_3/temp6[169] ), .ZN(\RI1[4][169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_3_4  ( .A(\MC_ARK_ARC_1_3/temp3[169] ), .B(
        \MC_ARK_ARC_1_3/temp4[169] ), .ZN(\MC_ARK_ARC_1_3/temp6[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_3_4  ( .A(\MC_ARK_ARC_1_3/temp1[169] ), .B(
        \MC_ARK_ARC_1_3/temp2[169] ), .ZN(\MC_ARK_ARC_1_3/temp5[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_3_4  ( .A(\RI5[3][13] ), .B(n230), .ZN(
        \MC_ARK_ARC_1_3/temp4[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_3_4  ( .A(\RI5[3][79] ), .B(\RI5[3][43] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_3_4  ( .A(\RI5[3][139] ), .B(\RI5[3][115] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_3_4  ( .A(\RI5[3][169] ), .B(\RI5[3][163] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[169] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_3_3  ( .A(\MC_ARK_ARC_1_3/temp5[170] ), .B(
        \MC_ARK_ARC_1_3/temp6[170] ), .ZN(\RI1[4][170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_3_3  ( .A(\MC_ARK_ARC_1_3/temp3[170] ), .B(
        \MC_ARK_ARC_1_3/temp4[170] ), .ZN(\MC_ARK_ARC_1_3/temp6[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_3_3  ( .A(\MC_ARK_ARC_1_3/temp1[170] ), .B(
        \MC_ARK_ARC_1_3/temp2[170] ), .ZN(\MC_ARK_ARC_1_3/temp5[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_3_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .B(n482), .ZN(\MC_ARK_ARC_1_3/temp4[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_3_3  ( .A(\RI5[3][80] ), .B(\RI5[3][44] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_3_3  ( .A(\RI5[3][140] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[116] ), .ZN(\MC_ARK_ARC_1_3/temp2[170] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_3_3  ( .A(\RI5[3][170] ), .B(n1627), .ZN(
        \MC_ARK_ARC_1_3/temp1[170] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_3_2  ( .A(\MC_ARK_ARC_1_3/temp6[171] ), .B(
        \MC_ARK_ARC_1_3/temp5[171] ), .ZN(\RI1[4][171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_3_2  ( .A(\MC_ARK_ARC_1_3/temp3[171] ), .B(
        \MC_ARK_ARC_1_3/temp4[171] ), .ZN(\MC_ARK_ARC_1_3/temp6[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_3_2  ( .A(\MC_ARK_ARC_1_3/temp1[171] ), .B(
        \MC_ARK_ARC_1_3/temp2[171] ), .ZN(\MC_ARK_ARC_1_3/temp5[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_3_2  ( .A(\RI5[3][15] ), .B(n228), .ZN(
        \MC_ARK_ARC_1_3/temp4[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_3_2  ( .A(n1658), .B(\RI5[3][45] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_3_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[141] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[117] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_3_2  ( .A(\RI5[3][171] ), .B(\RI5[3][165] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[171] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_3_1  ( .A(\MC_ARK_ARC_1_3/temp5[172] ), .B(
        \MC_ARK_ARC_1_3/temp6[172] ), .ZN(\RI1[4][172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_3_1  ( .A(\MC_ARK_ARC_1_3/temp3[172] ), .B(
        \MC_ARK_ARC_1_3/temp4[172] ), .ZN(\MC_ARK_ARC_1_3/temp6[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_3_1  ( .A(\MC_ARK_ARC_1_3/temp1[172] ), .B(
        \MC_ARK_ARC_1_3/temp2[172] ), .ZN(\MC_ARK_ARC_1_3/temp5[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_3_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[16] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[172] ), .ZN(
        \MC_ARK_ARC_1_3/temp4[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_3_1  ( .A(\RI5[3][82] ), .B(\RI5[3][46] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_3_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .B(\RI5[3][118] ), .ZN(\MC_ARK_ARC_1_3/temp2[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_3_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[172] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[166] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[172] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_3_0  ( .A(\MC_ARK_ARC_1_3/temp5[173] ), .B(
        \MC_ARK_ARC_1_3/temp6[173] ), .ZN(\RI1[4][173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_3_0  ( .A(\MC_ARK_ARC_1_3/temp3[173] ), .B(
        \MC_ARK_ARC_1_3/temp4[173] ), .ZN(\MC_ARK_ARC_1_3/temp6[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_3_0  ( .A(\MC_ARK_ARC_1_3/temp1[173] ), .B(
        \MC_ARK_ARC_1_3/temp2[173] ), .ZN(\MC_ARK_ARC_1_3/temp5[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_3_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .B(\MC_ARK_ARC_1_3/buf_keyinput[173] ), .ZN(
        \MC_ARK_ARC_1_3/temp4[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_3_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[83] ), 
        .B(n842), .ZN(\MC_ARK_ARC_1_3/temp3[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_3_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .B(n1661), .ZN(\MC_ARK_ARC_1_3/temp2[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_3_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[173] ), 
        .B(n1946), .ZN(\MC_ARK_ARC_1_3/temp1[173] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_2_5  ( .A(\MC_ARK_ARC_1_3/temp5[174] ), .B(
        \MC_ARK_ARC_1_3/temp6[174] ), .ZN(\RI1[4][174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_2_5  ( .A(\MC_ARK_ARC_1_3/temp3[174] ), .B(
        \MC_ARK_ARC_1_3/temp4[174] ), .ZN(\MC_ARK_ARC_1_3/temp6[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_2_5  ( .A(\MC_ARK_ARC_1_3/temp1[174] ), .B(
        \MC_ARK_ARC_1_3/temp2[174] ), .ZN(\MC_ARK_ARC_1_3/temp5[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_2_5  ( .A(\RI5[3][18] ), .B(n500), .ZN(
        \MC_ARK_ARC_1_3/temp4[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_2_5  ( .A(\RI5[3][84] ), .B(\RI5[3][48] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_2_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[144] ), 
        .B(\RI5[3][120] ), .ZN(\MC_ARK_ARC_1_3/temp2[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_2_5  ( .A(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .B(\RI5[3][168] ), .ZN(\MC_ARK_ARC_1_3/temp1[174] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_2_4  ( .A(\MC_ARK_ARC_1_3/temp5[175] ), .B(
        \MC_ARK_ARC_1_3/temp6[175] ), .ZN(\RI1[4][175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_2_4  ( .A(\MC_ARK_ARC_1_3/temp3[175] ), .B(
        \MC_ARK_ARC_1_3/temp4[175] ), .ZN(\MC_ARK_ARC_1_3/temp6[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_2_4  ( .A(\MC_ARK_ARC_1_3/temp1[175] ), .B(
        \MC_ARK_ARC_1_3/temp2[175] ), .ZN(\MC_ARK_ARC_1_3/temp5[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_2_4  ( .A(\RI5[3][19] ), .B(n511), .ZN(
        \MC_ARK_ARC_1_3/temp4[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_2_4  ( .A(\RI5[3][85] ), .B(\RI5[3][49] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_2_4  ( .A(\RI5[3][145] ), .B(\RI5[3][121] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_2_4  ( .A(\RI5[3][175] ), .B(\RI5[3][169] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[175] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_2_3  ( .A(\MC_ARK_ARC_1_3/temp5[176] ), .B(
        \MC_ARK_ARC_1_3/temp6[176] ), .ZN(\RI1[4][176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_2_3  ( .A(\MC_ARK_ARC_1_3/temp3[176] ), .B(
        \MC_ARK_ARC_1_3/temp4[176] ), .ZN(\MC_ARK_ARC_1_3/temp6[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_2_3  ( .A(\MC_ARK_ARC_1_3/temp1[176] ), .B(
        \MC_ARK_ARC_1_3/temp2[176] ), .ZN(\MC_ARK_ARC_1_3/temp5[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_2_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[20] ), 
        .B(n314), .ZN(\MC_ARK_ARC_1_3/temp4[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_2_3  ( .A(\RI5[3][86] ), .B(n2129), .ZN(
        \MC_ARK_ARC_1_3/temp3[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_2_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[146] ), 
        .B(n1928), .ZN(\MC_ARK_ARC_1_3/temp2[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_2_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .B(\RI5[3][170] ), .ZN(\MC_ARK_ARC_1_3/temp1[176] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_2_2  ( .A(\MC_ARK_ARC_1_3/temp5[177] ), .B(
        \MC_ARK_ARC_1_3/temp6[177] ), .ZN(\RI1[4][177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_2_2  ( .A(\MC_ARK_ARC_1_3/temp3[177] ), .B(
        \MC_ARK_ARC_1_3/temp4[177] ), .ZN(\MC_ARK_ARC_1_3/temp6[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_2_2  ( .A(\MC_ARK_ARC_1_3/temp1[177] ), .B(
        \MC_ARK_ARC_1_3/temp2[177] ), .ZN(\MC_ARK_ARC_1_3/temp5[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_2_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .B(n392), .ZN(\MC_ARK_ARC_1_3/temp4[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_2_2  ( .A(\RI5[3][87] ), .B(\RI5[3][51] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_2_2  ( .A(\RI5[3][147] ), .B(\RI5[3][123] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_2_2  ( .A(\RI5[3][177] ), .B(\RI5[3][171] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[177] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_2_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .B(n428), .ZN(\MC_ARK_ARC_1_3/temp4[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_2_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[88] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[52] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_2_1  ( .A(n1510), .B(
        \MC_ARK_ARC_1_3/buf_datainput[124] ), .ZN(\MC_ARK_ARC_1_3/temp2[178] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_2_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[172] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[178] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_2_0  ( .A(\MC_ARK_ARC_1_3/temp1[179] ), .B(
        \MC_ARK_ARC_1_3/temp2[179] ), .ZN(\MC_ARK_ARC_1_3/temp5[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_2_0  ( .A(n1653), .B(
        \MC_ARK_ARC_1_3/buf_keyinput[179] ), .ZN(\MC_ARK_ARC_1_3/temp4[179] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_2_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[89] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_2_0  ( .A(n850), .B(n520), .ZN(
        \MC_ARK_ARC_1_3/temp2[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_2_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[173] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[179] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_1_5  ( .A(\MC_ARK_ARC_1_3/temp5[180] ), .B(
        \MC_ARK_ARC_1_3/temp6[180] ), .ZN(\RI1[4][180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_1_5  ( .A(\MC_ARK_ARC_1_3/temp3[180] ), .B(
        \MC_ARK_ARC_1_3/temp4[180] ), .ZN(\MC_ARK_ARC_1_3/temp6[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_1_5  ( .A(\MC_ARK_ARC_1_3/temp1[180] ), .B(
        \MC_ARK_ARC_1_3/temp2[180] ), .ZN(\MC_ARK_ARC_1_3/temp5[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_1_5  ( .A(\RI5[3][24] ), .B(n310), .ZN(
        \MC_ARK_ARC_1_3/temp4[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_1_5  ( .A(\RI5[3][90] ), .B(\RI5[3][54] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_1_5  ( .A(\RI5[3][150] ), .B(\RI5[3][126] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[180] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_1_5  ( .A(\RI5[3][180] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[174] ), .ZN(\MC_ARK_ARC_1_3/temp1[180] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_1_4  ( .A(\MC_ARK_ARC_1_3/temp5[181] ), .B(
        \MC_ARK_ARC_1_3/temp6[181] ), .ZN(\RI1[4][181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_1_4  ( .A(\MC_ARK_ARC_1_3/temp3[181] ), .B(
        \MC_ARK_ARC_1_3/temp4[181] ), .ZN(\MC_ARK_ARC_1_3/temp6[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_1_4  ( .A(\MC_ARK_ARC_1_3/temp1[181] ), .B(
        \MC_ARK_ARC_1_3/temp2[181] ), .ZN(\MC_ARK_ARC_1_3/temp5[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_1_4  ( .A(\RI5[3][25] ), .B(n218), .ZN(
        \MC_ARK_ARC_1_3/temp4[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_1_4  ( .A(\MC_ARK_ARC_1_3/buf_datainput[91] ), 
        .B(\RI5[3][55] ), .ZN(\MC_ARK_ARC_1_3/temp3[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_1_4  ( .A(\RI5[3][151] ), .B(\RI5[3][127] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_1_4  ( .A(\RI5[3][181] ), .B(\RI5[3][175] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[181] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_1_3  ( .A(\MC_ARK_ARC_1_3/temp3[182] ), .B(
        \MC_ARK_ARC_1_3/temp4[182] ), .ZN(\MC_ARK_ARC_1_3/temp6[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_1_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[26] ), 
        .B(n459), .ZN(\MC_ARK_ARC_1_3/temp4[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_1_3  ( .A(\RI5[3][92] ), .B(\RI5[3][56] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_1_3  ( .A(\RI5[3][152] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[128] ), .ZN(\MC_ARK_ARC_1_3/temp2[182] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_1_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[176] ), .ZN(
        \MC_ARK_ARC_1_3/temp1[182] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_1_2  ( .A(\MC_ARK_ARC_1_3/temp5[183] ), .B(
        \MC_ARK_ARC_1_3/temp6[183] ), .ZN(\RI1[4][183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_1_2  ( .A(\MC_ARK_ARC_1_3/temp3[183] ), .B(
        \MC_ARK_ARC_1_3/temp4[183] ), .ZN(\MC_ARK_ARC_1_3/temp6[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_1_2  ( .A(\MC_ARK_ARC_1_3/temp1[183] ), .B(
        \MC_ARK_ARC_1_3/temp2[183] ), .ZN(\MC_ARK_ARC_1_3/temp5[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_1_2  ( .A(\RI5[3][27] ), .B(n385), .ZN(
        \MC_ARK_ARC_1_3/temp4[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_1_2  ( .A(\RI5[3][93] ), .B(\RI5[3][57] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_1_2  ( .A(\RI5[3][153] ), .B(\RI5[3][129] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_1_2  ( .A(\MC_ARK_ARC_1_3/buf_datainput[183] ), 
        .B(\RI5[3][177] ), .ZN(\MC_ARK_ARC_1_3/temp1[183] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_1_1  ( .A(\MC_ARK_ARC_1_3/temp5[184] ), .B(
        \MC_ARK_ARC_1_3/temp6[184] ), .ZN(\RI1[4][184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_1_1  ( .A(\MC_ARK_ARC_1_3/temp3[184] ), .B(
        \MC_ARK_ARC_1_3/temp4[184] ), .ZN(\MC_ARK_ARC_1_3/temp6[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_1_1  ( .A(\MC_ARK_ARC_1_3/temp1[184] ), .B(
        \MC_ARK_ARC_1_3/temp2[184] ), .ZN(\MC_ARK_ARC_1_3/temp5[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_1_1  ( .A(\RI5[3][28] ), .B(n306), .ZN(
        \MC_ARK_ARC_1_3/temp4[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_1_1  ( .A(\RI5[3][94] ), .B(\RI5[3][58] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_1_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[154] ), 
        .B(n1942), .ZN(\MC_ARK_ARC_1_3/temp2[184] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_1_1  ( .A(\RI5[3][184] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[178] ), .ZN(\MC_ARK_ARC_1_3/temp1[184] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_1_0  ( .A(\MC_ARK_ARC_1_3/temp5[185] ), .B(
        \MC_ARK_ARC_1_3/temp6[185] ), .ZN(\RI1[4][185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_1_0  ( .A(\MC_ARK_ARC_1_3/temp3[185] ), .B(
        \MC_ARK_ARC_1_3/temp4[185] ), .ZN(\MC_ARK_ARC_1_3/temp6[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_1_0  ( .A(\MC_ARK_ARC_1_3/temp1[185] ), .B(
        \MC_ARK_ARC_1_3/temp2[185] ), .ZN(\MC_ARK_ARC_1_3/temp5[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_1_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .B(n433), .ZN(\MC_ARK_ARC_1_3/temp4[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_1_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[59] ), 
        .B(n2145), .ZN(\MC_ARK_ARC_1_3/temp3[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_1_0  ( .A(n801), .B(n2121), .ZN(
        \MC_ARK_ARC_1_3/temp2[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_1_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .B(n839), .ZN(\MC_ARK_ARC_1_3/temp1[185] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_0_5  ( .A(\MC_ARK_ARC_1_3/temp6[186] ), .B(
        \MC_ARK_ARC_1_3/temp5[186] ), .ZN(\RI1[4][186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_0_5  ( .A(\MC_ARK_ARC_1_3/temp3[186] ), .B(
        \MC_ARK_ARC_1_3/temp4[186] ), .ZN(\MC_ARK_ARC_1_3/temp6[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_0_5  ( .A(\MC_ARK_ARC_1_3/temp1[186] ), .B(
        \MC_ARK_ARC_1_3/temp2[186] ), .ZN(\MC_ARK_ARC_1_3/temp5[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_0_5  ( .A(\RI5[3][30] ), .B(n497), .ZN(
        \MC_ARK_ARC_1_3/temp4[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_0_5  ( .A(\RI5[3][96] ), .B(\RI5[3][60] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_0_5  ( .A(\RI5[3][156] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[132] ), .ZN(\MC_ARK_ARC_1_3/temp2[186] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_0_5  ( .A(\RI5[3][186] ), .B(\RI5[3][180] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[186] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_0_4  ( .A(\MC_ARK_ARC_1_3/temp5[187] ), .B(
        \MC_ARK_ARC_1_3/temp6[187] ), .ZN(\RI1[4][187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_0_4  ( .A(\MC_ARK_ARC_1_3/temp3[187] ), .B(
        \MC_ARK_ARC_1_3/temp4[187] ), .ZN(\MC_ARK_ARC_1_3/temp6[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_0_4  ( .A(\MC_ARK_ARC_1_3/temp1[187] ), .B(
        \MC_ARK_ARC_1_3/temp2[187] ), .ZN(\MC_ARK_ARC_1_3/temp5[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_0_4  ( .A(\RI5[3][31] ), .B(n483), .ZN(
        \MC_ARK_ARC_1_3/temp4[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_0_4  ( .A(\RI5[3][97] ), .B(\RI5[3][61] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_0_4  ( .A(\RI5[3][157] ), .B(\RI5[3][133] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_0_4  ( .A(\RI5[3][187] ), .B(\RI5[3][181] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[187] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_0_3  ( .A(\MC_ARK_ARC_1_3/temp5[188] ), .B(
        \MC_ARK_ARC_1_3/temp6[188] ), .ZN(\RI1[4][188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_0_3  ( .A(\MC_ARK_ARC_1_3/temp3[188] ), .B(
        \MC_ARK_ARC_1_3/temp4[188] ), .ZN(\MC_ARK_ARC_1_3/temp6[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_0_3  ( .A(\MC_ARK_ARC_1_3/temp1[188] ), .B(
        \MC_ARK_ARC_1_3/temp2[188] ), .ZN(\MC_ARK_ARC_1_3/temp5[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_0_3  ( .A(\MC_ARK_ARC_1_3/buf_datainput[32] ), 
        .B(n302), .ZN(\MC_ARK_ARC_1_3/temp4[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_0_3  ( .A(\RI5[3][98] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[62] ), .ZN(\MC_ARK_ARC_1_3/temp3[188] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_0_3  ( .A(n2119), .B(\RI5[3][134] ), .ZN(
        \MC_ARK_ARC_1_3/temp2[188] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_0_3  ( .A(\RI5[3][188] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[182] ), .ZN(\MC_ARK_ARC_1_3/temp1[188] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_0_2  ( .A(\MC_ARK_ARC_1_3/temp5[189] ), .B(
        \MC_ARK_ARC_1_3/temp6[189] ), .ZN(\RI1[4][189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_0_2  ( .A(\MC_ARK_ARC_1_3/temp3[189] ), .B(
        \MC_ARK_ARC_1_3/temp4[189] ), .ZN(\MC_ARK_ARC_1_3/temp6[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_0_2  ( .A(\MC_ARK_ARC_1_3/temp1[189] ), .B(
        \MC_ARK_ARC_1_3/temp2[189] ), .ZN(\MC_ARK_ARC_1_3/temp5[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_0_2  ( .A(\RI5[3][33] ), .B(n405), .ZN(
        \MC_ARK_ARC_1_3/temp4[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_0_2  ( .A(\RI5[3][99] ), .B(\RI5[3][63] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_0_2  ( .A(\RI5[3][159] ), .B(\RI5[3][135] ), 
        .ZN(\MC_ARK_ARC_1_3/temp2[189] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_0_2  ( .A(\RI5[3][189] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[183] ), .ZN(\MC_ARK_ARC_1_3/temp1[189] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_0_1  ( .A(\MC_ARK_ARC_1_3/temp5[190] ), .B(
        \MC_ARK_ARC_1_3/temp6[190] ), .ZN(\RI1[4][190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_0_1  ( .A(\MC_ARK_ARC_1_3/temp3[190] ), .B(
        \MC_ARK_ARC_1_3/temp4[190] ), .ZN(\MC_ARK_ARC_1_3/temp6[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_0_1  ( .A(\MC_ARK_ARC_1_3/temp1[190] ), .B(
        \MC_ARK_ARC_1_3/temp2[190] ), .ZN(\MC_ARK_ARC_1_3/temp5[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_0_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[34] ), 
        .B(n300), .ZN(\MC_ARK_ARC_1_3/temp4[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_0_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[100] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[64] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_0_1  ( .A(\RI5[3][160] ), .B(
        \MC_ARK_ARC_1_3/buf_datainput[136] ), .ZN(\MC_ARK_ARC_1_3/temp2[190] )
         );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_0_1  ( .A(\RI5[3][190] ), .B(\RI5[3][184] ), 
        .ZN(\MC_ARK_ARC_1_3/temp1[190] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_0_0  ( .A(\MC_ARK_ARC_1_3/temp5[191] ), .B(
        \MC_ARK_ARC_1_3/temp6[191] ), .ZN(\RI1[4][191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X6_0_0  ( .A(\MC_ARK_ARC_1_3/temp3[191] ), .B(
        \MC_ARK_ARC_1_3/temp4[191] ), .ZN(\MC_ARK_ARC_1_3/temp6[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X5_0_0  ( .A(\MC_ARK_ARC_1_3/temp2[191] ), .B(
        \MC_ARK_ARC_1_3/temp1[191] ), .ZN(\MC_ARK_ARC_1_3/temp5[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_0_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[35] ), 
        .B(n208), .ZN(\MC_ARK_ARC_1_3/temp4[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X3_0_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .B(\MC_ARK_ARC_1_3/buf_datainput[65] ), .ZN(
        \MC_ARK_ARC_1_3/temp3[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X2_0_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[161] ), 
        .B(n784), .ZN(\MC_ARK_ARC_1_3/temp2[191] ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X1_0_0  ( .A(\MC_ARK_ARC_1_3/buf_datainput[191] ), 
        .B(n839), .ZN(\MC_ARK_ARC_1_3/temp1[191] ) );
  INV_X1 \SB1_0_0/INV_3  ( .A(n3), .ZN(\SB1_0_0/i0[10] ) );
  INV_X1 \SB1_0_0/INV_2  ( .A(n4), .ZN(\SB1_0_0/i0_0 ) );
  INV_X1 \SB1_0_0/INV_1  ( .A(n5), .ZN(\SB1_0_0/i0[6] ) );
  INV_X1 \SB1_0_1/INV_2  ( .A(n10), .ZN(\SB1_0_1/i0_0 ) );
  INV_X1 \SB1_0_2/INV_4  ( .A(n14), .ZN(\SB1_0_2/i0_4 ) );
  INV_X1 \SB1_0_2/INV_3  ( .A(n15), .ZN(\SB1_0_2/i0[10] ) );
  INV_X1 \SB1_0_2/INV_2  ( .A(n16), .ZN(\SB1_0_2/i0_0 ) );
  INV_X1 \SB1_0_2/INV_1  ( .A(n17), .ZN(\SB1_0_2/i0[6] ) );
  INV_X1 \SB1_0_2/INV_0  ( .A(n18), .ZN(\SB1_0_2/i0[9] ) );
  BUF_X1 \SB1_0_2/BUF_5  ( .A(n13), .Z(\SB1_0_2/i1_5 ) );
  BUF_X1 \SB1_0_2/BUF_1  ( .A(n17), .Z(\SB1_0_2/i1_7 ) );
  INV_X1 \SB1_0_3/INV_4  ( .A(n20), .ZN(\SB1_0_3/i0_4 ) );
  INV_X1 \SB1_0_3/INV_3  ( .A(n21), .ZN(\SB1_0_3/i0[10] ) );
  INV_X1 \SB1_0_3/INV_2  ( .A(n22), .ZN(\SB1_0_3/i0_0 ) );
  INV_X1 \SB1_0_3/INV_1  ( .A(n23), .ZN(\SB1_0_3/i0[6] ) );
  INV_X1 \SB1_0_3/INV_0  ( .A(n24), .ZN(\SB1_0_3/i0[9] ) );
  BUF_X1 \SB1_0_3/BUF_5  ( .A(n19), .Z(\SB1_0_3/i1_5 ) );
  INV_X1 \SB1_0_4/INV_4  ( .A(n26), .ZN(\SB1_0_4/i0_4 ) );
  INV_X1 \SB1_0_4/INV_3  ( .A(n27), .ZN(\SB1_0_4/i0[10] ) );
  INV_X1 \SB1_0_4/INV_2  ( .A(n28), .ZN(\SB1_0_4/i0_0 ) );
  INV_X1 \SB1_0_4/INV_1  ( .A(n29), .ZN(\SB1_0_4/i0[6] ) );
  INV_X1 \SB1_0_4/INV_0  ( .A(n30), .ZN(\SB1_0_4/i0[9] ) );
  BUF_X1 \SB1_0_4/BUF_5  ( .A(n25), .Z(\SB1_0_4/i1_5 ) );
  BUF_X1 \SB1_0_4/BUF_1  ( .A(n29), .Z(\SB1_0_4/i1_7 ) );
  INV_X1 \SB1_0_5/INV_4  ( .A(n32), .ZN(\SB1_0_5/i0_4 ) );
  INV_X1 \SB1_0_5/INV_1  ( .A(n35), .ZN(\SB1_0_5/i0[6] ) );
  BUF_X1 \SB1_0_5/BUF_1  ( .A(n35), .Z(\SB1_0_5/i1_7 ) );
  INV_X1 \SB1_0_6/INV_3  ( .A(n39), .ZN(\SB1_0_6/i0[10] ) );
  INV_X1 \SB1_0_6/INV_2  ( .A(n40), .ZN(\SB1_0_6/i0_0 ) );
  INV_X1 \SB1_0_6/INV_1  ( .A(n41), .ZN(\SB1_0_6/i0[6] ) );
  INV_X1 \SB1_0_7/INV_3  ( .A(n45), .ZN(\SB1_0_7/i0[10] ) );
  INV_X1 \SB1_0_7/INV_2  ( .A(n46), .ZN(\SB1_0_7/i0_0 ) );
  INV_X1 \SB1_0_7/INV_1  ( .A(n47), .ZN(\SB1_0_7/i0[6] ) );
  INV_X1 \SB1_0_7/INV_0  ( .A(n48), .ZN(\SB1_0_7/i0[9] ) );
  INV_X1 \SB1_0_8/INV_3  ( .A(n51), .ZN(\SB1_0_8/i0[10] ) );
  INV_X1 \SB1_0_8/INV_2  ( .A(n52), .ZN(\SB1_0_8/i0_0 ) );
  INV_X1 \SB1_0_8/INV_1  ( .A(n53), .ZN(\SB1_0_8/i0[6] ) );
  INV_X1 \SB1_0_8/INV_0  ( .A(n54), .ZN(\SB1_0_8/i0[9] ) );
  INV_X1 \SB1_0_9/INV_3  ( .A(n57), .ZN(\SB1_0_9/i0[10] ) );
  INV_X1 \SB1_0_9/INV_2  ( .A(n58), .ZN(\SB1_0_9/i0_0 ) );
  INV_X1 \SB1_0_9/INV_1  ( .A(n59), .ZN(\SB1_0_9/i0[6] ) );
  INV_X1 \SB1_0_9/INV_0  ( .A(n60), .ZN(\SB1_0_9/i0[9] ) );
  BUF_X1 \SB1_0_9/BUF_5  ( .A(n55), .Z(\SB1_0_9/i1_5 ) );
  BUF_X1 \SB1_0_9/BUF_1  ( .A(n59), .Z(\SB1_0_9/i1_7 ) );
  INV_X1 \SB1_0_10/INV_3  ( .A(n63), .ZN(\SB1_0_10/i0[10] ) );
  INV_X1 \SB1_0_10/INV_2  ( .A(n64), .ZN(\SB1_0_10/i0_0 ) );
  INV_X1 \SB1_0_10/INV_1  ( .A(n65), .ZN(\SB1_0_10/i0[6] ) );
  INV_X1 \SB1_0_10/INV_0  ( .A(n66), .ZN(\SB1_0_10/i0[9] ) );
  BUF_X1 \SB1_0_10/BUF_5  ( .A(n61), .Z(\SB1_0_10/i1_5 ) );
  BUF_X1 \SB1_0_10/BUF_1  ( .A(n65), .Z(\SB1_0_10/i1_7 ) );
  INV_X1 \SB1_0_11/INV_4  ( .A(n68), .ZN(\SB1_0_11/i0_4 ) );
  INV_X1 \SB1_0_11/INV_3  ( .A(n69), .ZN(\SB1_0_11/i0[10] ) );
  INV_X1 \SB1_0_11/INV_2  ( .A(n70), .ZN(\SB1_0_11/i0_0 ) );
  INV_X1 \SB1_0_11/INV_1  ( .A(n71), .ZN(\SB1_0_11/i0[6] ) );
  INV_X1 \SB1_0_11/INV_0  ( .A(n72), .ZN(\SB1_0_11/i0[9] ) );
  BUF_X1 \SB1_0_11/BUF_5  ( .A(n67), .Z(\SB1_0_11/i1_5 ) );
  BUF_X1 \SB1_0_11/BUF_1  ( .A(n71), .Z(\SB1_0_11/i1_7 ) );
  INV_X1 \SB1_0_12/INV_3  ( .A(n75), .ZN(\SB1_0_12/i0[10] ) );
  INV_X1 \SB1_0_12/INV_1  ( .A(n77), .ZN(\SB1_0_12/i0[6] ) );
  BUF_X1 \SB1_0_12/BUF_1  ( .A(n77), .Z(\SB1_0_12/i1_7 ) );
  INV_X1 \SB1_0_13/INV_3  ( .A(n81), .ZN(\SB1_0_13/i0[10] ) );
  INV_X1 \SB1_0_13/INV_2  ( .A(n82), .ZN(\SB1_0_13/i0_0 ) );
  INV_X1 \SB1_0_14/INV_4  ( .A(n86), .ZN(\SB1_0_14/i0_4 ) );
  INV_X1 \SB1_0_14/INV_3  ( .A(n87), .ZN(\SB1_0_14/i0[10] ) );
  INV_X1 \SB1_0_14/INV_1  ( .A(n89), .ZN(\SB1_0_14/i0[6] ) );
  INV_X1 \SB1_0_14/INV_0  ( .A(n90), .ZN(\SB1_0_14/i0[9] ) );
  INV_X1 \SB1_0_15/INV_4  ( .A(n92), .ZN(\SB1_0_15/i0_4 ) );
  INV_X1 \SB1_0_15/INV_3  ( .A(n93), .ZN(\SB1_0_15/i0[10] ) );
  INV_X1 \SB1_0_15/INV_2  ( .A(n94), .ZN(\SB1_0_15/i0_0 ) );
  INV_X1 \SB1_0_15/INV_1  ( .A(n95), .ZN(\SB1_0_15/i0[6] ) );
  INV_X1 \SB1_0_15/INV_0  ( .A(n96), .ZN(\SB1_0_15/i0[9] ) );
  BUF_X1 \SB1_0_15/BUF_5  ( .A(n91), .Z(\SB1_0_15/i1_5 ) );
  INV_X1 \SB1_0_16/INV_3  ( .A(n99), .ZN(\SB1_0_16/i0[10] ) );
  INV_X1 \SB1_0_16/INV_2  ( .A(n100), .ZN(\SB1_0_16/i0_0 ) );
  INV_X1 \SB1_0_16/INV_1  ( .A(n101), .ZN(\SB1_0_16/i0[6] ) );
  INV_X1 \SB1_0_16/INV_0  ( .A(n102), .ZN(\SB1_0_16/i0[9] ) );
  BUF_X1 \SB1_0_16/BUF_5  ( .A(n97), .Z(\SB1_0_16/i1_5 ) );
  INV_X1 \SB1_0_17/INV_4  ( .A(n104), .ZN(\SB1_0_17/i0_4 ) );
  INV_X1 \SB1_0_17/INV_3  ( .A(n105), .ZN(\SB1_0_17/i0[10] ) );
  INV_X1 \SB1_0_17/INV_2  ( .A(n106), .ZN(\SB1_0_17/i0_0 ) );
  INV_X1 \SB1_0_17/INV_1  ( .A(n107), .ZN(\SB1_0_17/i0[6] ) );
  INV_X1 \SB1_0_17/INV_0  ( .A(n108), .ZN(\SB1_0_17/i0[9] ) );
  BUF_X1 \SB1_0_17/BUF_5  ( .A(n103), .Z(\SB1_0_17/i1_5 ) );
  INV_X1 \SB1_0_18/INV_3  ( .A(n111), .ZN(\SB1_0_18/i0[10] ) );
  INV_X1 \SB1_0_18/INV_2  ( .A(n112), .ZN(\SB1_0_18/i0_0 ) );
  INV_X1 \SB1_0_18/INV_1  ( .A(n113), .ZN(\SB1_0_18/i0[6] ) );
  INV_X1 \SB1_0_18/INV_0  ( .A(n114), .ZN(\SB1_0_18/i0[9] ) );
  BUF_X1 \SB1_0_18/BUF_5  ( .A(n109), .Z(\SB1_0_18/i1_5 ) );
  INV_X1 \SB1_0_19/INV_3  ( .A(n117), .ZN(\SB1_0_19/i0[10] ) );
  INV_X1 \SB1_0_19/INV_2  ( .A(n118), .ZN(\SB1_0_19/i0_0 ) );
  INV_X1 \SB1_0_19/INV_1  ( .A(n119), .ZN(\SB1_0_19/i0[6] ) );
  INV_X1 \SB1_0_19/INV_0  ( .A(n120), .ZN(\SB1_0_19/i0[9] ) );
  BUF_X1 \SB1_0_19/BUF_5  ( .A(n115), .Z(\SB1_0_19/i1_5 ) );
  BUF_X1 \SB1_0_19/BUF_1  ( .A(n119), .Z(\SB1_0_19/i1_7 ) );
  INV_X1 \SB1_0_20/INV_4  ( .A(n122), .ZN(\SB1_0_20/i0_4 ) );
  INV_X1 \SB1_0_20/INV_3  ( .A(n123), .ZN(\SB1_0_20/i0[10] ) );
  INV_X1 \SB1_0_20/INV_2  ( .A(n124), .ZN(\SB1_0_20/i0_0 ) );
  INV_X1 \SB1_0_20/INV_1  ( .A(n125), .ZN(\SB1_0_20/i0[6] ) );
  INV_X1 \SB1_0_20/INV_0  ( .A(n126), .ZN(\SB1_0_20/i0[9] ) );
  INV_X1 \SB1_0_21/INV_3  ( .A(n129), .ZN(\SB1_0_21/i0[10] ) );
  INV_X1 \SB1_0_21/INV_2  ( .A(n130), .ZN(\SB1_0_21/i0_0 ) );
  INV_X1 \SB1_0_21/INV_1  ( .A(n131), .ZN(\SB1_0_21/i0[6] ) );
  INV_X1 \SB1_0_21/INV_0  ( .A(n132), .ZN(\SB1_0_21/i0[9] ) );
  BUF_X1 \SB1_0_21/BUF_1  ( .A(n131), .Z(\SB1_0_21/i1_7 ) );
  INV_X1 \SB1_0_22/INV_4  ( .A(n134), .ZN(\SB1_0_22/i0_4 ) );
  INV_X1 \SB1_0_22/INV_3  ( .A(n135), .ZN(\SB1_0_22/i0[10] ) );
  INV_X1 \SB1_0_22/INV_2  ( .A(n136), .ZN(\SB1_0_22/i0_0 ) );
  INV_X1 \SB1_0_22/INV_1  ( .A(n137), .ZN(\SB1_0_22/i0[6] ) );
  INV_X1 \SB1_0_22/INV_0  ( .A(n138), .ZN(\SB1_0_22/i0[9] ) );
  BUF_X1 \SB1_0_22/BUF_1  ( .A(n137), .Z(\SB1_0_22/i1_7 ) );
  INV_X1 \SB1_0_23/INV_1  ( .A(n143), .ZN(\SB1_0_23/i0[6] ) );
  INV_X1 \SB1_0_24/INV_4  ( .A(n146), .ZN(\SB1_0_24/i0_4 ) );
  INV_X1 \SB1_0_24/INV_3  ( .A(n147), .ZN(\SB1_0_24/i0[10] ) );
  INV_X1 \SB1_0_24/INV_2  ( .A(n148), .ZN(\SB1_0_24/i0_0 ) );
  INV_X1 \SB1_0_24/INV_1  ( .A(n149), .ZN(\SB1_0_24/i0[6] ) );
  INV_X1 \SB1_0_24/INV_0  ( .A(n150), .ZN(\SB1_0_24/i0[9] ) );
  INV_X1 \SB1_0_25/INV_3  ( .A(n153), .ZN(\SB1_0_25/i0[10] ) );
  INV_X1 \SB1_0_25/INV_1  ( .A(n155), .ZN(\SB1_0_25/i0[6] ) );
  INV_X1 \SB1_0_25/INV_0  ( .A(n156), .ZN(\SB1_0_25/i0[9] ) );
  BUF_X1 \SB1_0_25/BUF_5  ( .A(n151), .Z(\SB1_0_25/i1_5 ) );
  BUF_X1 \SB1_0_25/BUF_1  ( .A(n155), .Z(\SB1_0_25/i1_7 ) );
  INV_X1 \SB1_0_26/INV_3  ( .A(n159), .ZN(\SB1_0_26/i0[10] ) );
  INV_X1 \SB1_0_26/INV_2  ( .A(n160), .ZN(\SB1_0_26/i0_0 ) );
  INV_X1 \SB1_0_26/INV_1  ( .A(n161), .ZN(\SB1_0_26/i0[6] ) );
  INV_X1 \SB1_0_26/INV_0  ( .A(n162), .ZN(\SB1_0_26/i0[9] ) );
  INV_X1 \SB1_0_27/INV_4  ( .A(n164), .ZN(\SB1_0_27/i0_4 ) );
  INV_X1 \SB1_0_27/INV_3  ( .A(n165), .ZN(\SB1_0_27/i0[10] ) );
  INV_X1 \SB1_0_27/INV_2  ( .A(n166), .ZN(\SB1_0_27/i0_0 ) );
  INV_X1 \SB1_0_27/INV_1  ( .A(n167), .ZN(\SB1_0_27/i0[6] ) );
  INV_X1 \SB1_0_27/INV_0  ( .A(n168), .ZN(\SB1_0_27/i0[9] ) );
  BUF_X1 \SB1_0_27/BUF_1  ( .A(n167), .Z(\SB1_0_27/i1_7 ) );
  INV_X1 \SB1_0_28/INV_4  ( .A(n170), .ZN(\SB1_0_28/i0_4 ) );
  INV_X1 \SB1_0_28/INV_2  ( .A(n172), .ZN(\SB1_0_28/i0_0 ) );
  INV_X1 \SB1_0_28/INV_1  ( .A(n173), .ZN(\SB1_0_28/i0[6] ) );
  INV_X1 \SB1_0_28/INV_0  ( .A(n174), .ZN(\SB1_0_28/i0[9] ) );
  BUF_X1 \SB1_0_28/BUF_5  ( .A(n169), .Z(\SB1_0_28/i1_5 ) );
  INV_X1 \SB1_0_29/INV_3  ( .A(n177), .ZN(\SB1_0_29/i0[10] ) );
  INV_X1 \SB1_0_29/INV_2  ( .A(n178), .ZN(\SB1_0_29/i0_0 ) );
  INV_X1 \SB1_0_29/INV_1  ( .A(n179), .ZN(\SB1_0_29/i0[6] ) );
  INV_X1 \SB1_0_29/INV_0  ( .A(n180), .ZN(\SB1_0_29/i0[9] ) );
  BUF_X1 \SB1_0_29/BUF_1  ( .A(n179), .Z(\SB1_0_29/i1_7 ) );
  INV_X1 \SB1_0_30/INV_4  ( .A(n182), .ZN(\SB1_0_30/i0_4 ) );
  INV_X1 \SB1_0_30/INV_3  ( .A(n183), .ZN(\SB1_0_30/i0[10] ) );
  INV_X1 \SB1_0_30/INV_2  ( .A(n184), .ZN(\SB1_0_30/i0_0 ) );
  INV_X1 \SB1_0_30/INV_1  ( .A(n185), .ZN(\SB1_0_30/i0[6] ) );
  INV_X1 \SB1_0_30/INV_0  ( .A(n186), .ZN(\SB1_0_30/i0[9] ) );
  INV_X1 \SB1_0_31/INV_4  ( .A(n188), .ZN(\SB1_0_31/i0_4 ) );
  INV_X1 \SB1_0_31/INV_3  ( .A(n189), .ZN(\SB1_0_31/i0[10] ) );
  INV_X1 \SB1_0_31/INV_2  ( .A(n190), .ZN(\SB1_0_31/i0_0 ) );
  INV_X1 \SB1_0_31/INV_1  ( .A(n191), .ZN(\SB1_0_31/i0[6] ) );
  INV_X1 \SB1_0_31/INV_0  ( .A(n192), .ZN(\SB1_0_31/i0[9] ) );
  BUF_X1 \SB1_0_31/BUF_1  ( .A(n191), .Z(\SB1_0_31/i1_7 ) );
  INV_X1 \SB1_1_0/INV_4  ( .A(\RI1[1][190] ), .ZN(\SB1_1_0/i0_4 ) );
  INV_X1 \SB1_1_0/INV_3  ( .A(\RI1[1][189] ), .ZN(\SB1_1_0/i0[10] ) );
  INV_X1 \SB1_1_0/INV_2  ( .A(\RI1[1][188] ), .ZN(\SB1_1_0/i0_0 ) );
  INV_X1 \SB1_1_0/INV_1  ( .A(\RI1[1][187] ), .ZN(\SB1_1_0/i0[6] ) );
  INV_X1 \SB1_1_1/INV_4  ( .A(\RI1[1][184] ), .ZN(\SB1_1_1/i0_4 ) );
  INV_X1 \SB1_1_1/INV_3  ( .A(\RI1[1][183] ), .ZN(\SB1_1_1/i0[10] ) );
  INV_X1 \SB1_1_1/INV_2  ( .A(\RI1[1][182] ), .ZN(\SB1_1_1/i0_0 ) );
  INV_X1 \SB1_1_1/INV_1  ( .A(\RI1[1][181] ), .ZN(\SB1_1_1/i0[6] ) );
  INV_X1 \SB1_1_1/INV_0  ( .A(\RI1[1][180] ), .ZN(\SB1_1_1/i0[9] ) );
  BUF_X1 \SB1_1_1/BUF_5  ( .A(\RI1[1][185] ), .Z(\SB1_1_1/i1_5 ) );
  INV_X1 \SB1_1_2/INV_4  ( .A(\RI1[1][178] ), .ZN(\SB1_1_2/i0_4 ) );
  INV_X1 \SB1_1_2/INV_3  ( .A(\RI1[1][177] ), .ZN(\SB1_1_2/i0[10] ) );
  INV_X1 \SB1_1_2/INV_2  ( .A(\RI1[1][176] ), .ZN(\SB1_1_2/i0_0 ) );
  INV_X1 \SB1_1_2/INV_1  ( .A(\RI1[1][175] ), .ZN(\SB1_1_2/i0[6] ) );
  INV_X1 \SB1_1_2/INV_0  ( .A(\RI1[1][174] ), .ZN(\SB1_1_2/i0[9] ) );
  INV_X1 \SB1_1_3/INV_2  ( .A(\RI1[1][170] ), .ZN(\SB1_1_3/i0_0 ) );
  INV_X1 \SB1_1_3/INV_1  ( .A(\RI1[1][169] ), .ZN(\SB1_1_3/i0[6] ) );
  BUF_X1 \SB1_1_3/BUF_5  ( .A(\RI1[1][173] ), .Z(\SB1_1_3/i1_5 ) );
  INV_X1 \SB1_1_4/INV_4  ( .A(\RI1[1][166] ), .ZN(\SB1_1_4/i0_4 ) );
  INV_X1 \SB1_1_4/INV_3  ( .A(\RI1[1][165] ), .ZN(\SB1_1_4/i0[10] ) );
  INV_X1 \SB1_1_4/INV_2  ( .A(\RI1[1][164] ), .ZN(\SB1_1_4/i0_0 ) );
  BUF_X1 \SB1_1_4/BUF_5  ( .A(\RI1[1][167] ), .Z(\SB1_1_4/i1_5 ) );
  INV_X1 \SB1_1_5/INV_4  ( .A(\RI1[1][160] ), .ZN(\SB1_1_5/i0_4 ) );
  INV_X1 \SB1_1_5/INV_3  ( .A(\RI1[1][159] ), .ZN(\SB1_1_5/i0[10] ) );
  INV_X1 \SB1_1_5/INV_2  ( .A(\RI1[1][158] ), .ZN(\SB1_1_5/i0_0 ) );
  INV_X1 \SB1_1_5/INV_1  ( .A(\RI1[1][157] ), .ZN(\SB1_1_5/i0[6] ) );
  BUF_X1 \SB1_1_5/BUF_5  ( .A(\RI1[1][161] ), .Z(\SB1_1_5/i1_5 ) );
  INV_X1 \SB1_1_6/INV_3  ( .A(\RI1[1][153] ), .ZN(\SB1_1_6/i0[10] ) );
  INV_X1 \SB1_1_6/INV_2  ( .A(\RI1[1][152] ), .ZN(\SB1_1_6/i0_0 ) );
  INV_X1 \SB1_1_6/INV_1  ( .A(\RI1[1][151] ), .ZN(\SB1_1_6/i0[6] ) );
  INV_X1 \SB1_1_6/INV_0  ( .A(\RI1[1][150] ), .ZN(\SB1_1_6/i0[9] ) );
  BUF_X1 \SB1_1_6/BUF_5  ( .A(\RI1[1][155] ), .Z(\SB1_1_6/i1_5 ) );
  INV_X1 \SB1_1_7/INV_4  ( .A(\RI1[1][148] ), .ZN(\SB1_1_7/i0_4 ) );
  INV_X1 \SB1_1_7/INV_3  ( .A(\RI1[1][147] ), .ZN(\SB1_1_7/i0[10] ) );
  INV_X1 \SB1_1_7/INV_2  ( .A(\RI1[1][146] ), .ZN(\SB1_1_7/i0_0 ) );
  INV_X1 \SB1_1_7/INV_1  ( .A(\RI1[1][145] ), .ZN(\SB1_1_7/i0[6] ) );
  INV_X1 \SB1_1_7/INV_0  ( .A(\RI1[1][144] ), .ZN(\SB1_1_7/i0[9] ) );
  INV_X1 \SB1_1_8/INV_2  ( .A(\RI1[1][140] ), .ZN(\SB1_1_8/i0_0 ) );
  INV_X1 \SB1_1_8/INV_1  ( .A(\RI1[1][139] ), .ZN(\SB1_1_8/i0[6] ) );
  BUF_X1 \SB1_1_8/BUF_5  ( .A(\RI1[1][143] ), .Z(\SB1_1_8/i1_5 ) );
  INV_X1 \SB1_1_9/INV_4  ( .A(\RI1[1][136] ), .ZN(\SB1_1_9/i0_4 ) );
  INV_X1 \SB1_1_9/INV_2  ( .A(\RI1[1][134] ), .ZN(\SB1_1_9/i0_0 ) );
  INV_X1 \SB1_1_9/INV_1  ( .A(\RI1[1][133] ), .ZN(\SB1_1_9/i0[6] ) );
  INV_X1 \SB1_1_10/INV_4  ( .A(\RI1[1][130] ), .ZN(\SB1_1_10/i0_4 ) );
  INV_X1 \SB1_1_10/INV_3  ( .A(\RI1[1][129] ), .ZN(\SB1_1_10/i0[10] ) );
  INV_X1 \SB1_1_10/INV_2  ( .A(\RI1[1][128] ), .ZN(\SB1_1_10/i0_0 ) );
  INV_X1 \SB1_1_10/INV_1  ( .A(\RI1[1][127] ), .ZN(\SB1_1_10/i0[6] ) );
  INV_X1 \SB1_1_11/INV_3  ( .A(\RI1[1][123] ), .ZN(\SB1_1_11/i0[10] ) );
  INV_X1 \SB1_1_11/INV_2  ( .A(\RI1[1][122] ), .ZN(\SB1_1_11/i0_0 ) );
  INV_X1 \SB1_1_11/INV_1  ( .A(\RI1[1][121] ), .ZN(\SB1_1_11/i0[6] ) );
  BUF_X1 \SB1_1_11/BUF_5  ( .A(\RI1[1][125] ), .Z(\SB1_1_11/i1_5 ) );
  INV_X1 \SB1_1_12/INV_4  ( .A(\RI1[1][118] ), .ZN(\SB1_1_12/i0_4 ) );
  INV_X1 \SB1_1_12/INV_3  ( .A(\RI1[1][117] ), .ZN(\SB1_1_12/i0[10] ) );
  INV_X1 \SB1_1_12/INV_2  ( .A(\RI1[1][116] ), .ZN(\SB1_1_12/i0_0 ) );
  INV_X1 \SB1_1_12/INV_1  ( .A(\RI1[1][115] ), .ZN(\SB1_1_12/i0[6] ) );
  INV_X1 \SB1_1_12/INV_0  ( .A(\RI1[1][114] ), .ZN(\SB1_1_12/i0[9] ) );
  BUF_X1 \SB1_1_12/BUF_5  ( .A(\RI1[1][119] ), .Z(\SB1_1_12/i1_5 ) );
  INV_X1 \SB1_1_13/INV_4  ( .A(\RI1[1][112] ), .ZN(\SB1_1_13/i0_4 ) );
  INV_X1 \SB1_1_13/INV_3  ( .A(\RI1[1][111] ), .ZN(\SB1_1_13/i0[10] ) );
  INV_X1 \SB1_1_13/INV_2  ( .A(\RI1[1][110] ), .ZN(\SB1_1_13/i0_0 ) );
  INV_X1 \SB1_1_13/INV_1  ( .A(\RI1[1][109] ), .ZN(\SB1_1_13/i0[6] ) );
  INV_X1 \SB1_1_14/INV_4  ( .A(\RI1[1][106] ), .ZN(\SB1_1_14/i0_4 ) );
  INV_X1 \SB1_1_14/INV_3  ( .A(\RI1[1][105] ), .ZN(\SB1_1_14/i0[10] ) );
  INV_X1 \SB1_1_14/INV_1  ( .A(\RI1[1][103] ), .ZN(\SB1_1_14/i0[6] ) );
  BUF_X1 \SB1_1_14/BUF_5  ( .A(\RI1[1][107] ), .Z(\SB1_1_14/i1_5 ) );
  INV_X1 \SB1_1_15/INV_4  ( .A(\RI1[1][100] ), .ZN(\SB1_1_15/i0_4 ) );
  INV_X1 \SB1_1_15/INV_3  ( .A(\RI1[1][99] ), .ZN(\SB1_1_15/i0[10] ) );
  INV_X1 \SB1_1_15/INV_2  ( .A(\RI1[1][98] ), .ZN(\SB1_1_15/i0_0 ) );
  INV_X1 \SB1_1_15/INV_1  ( .A(\RI1[1][97] ), .ZN(\SB1_1_15/i0[6] ) );
  BUF_X1 \SB1_1_15/BUF_5  ( .A(\RI1[1][101] ), .Z(\SB1_1_15/i1_5 ) );
  BUF_X1 \SB1_1_15/BUF_1  ( .A(\RI1[1][97] ), .Z(\SB1_1_15/i1_7 ) );
  INV_X1 \SB1_1_16/INV_3  ( .A(\RI1[1][93] ), .ZN(\SB1_1_16/i0[10] ) );
  INV_X1 \SB1_1_16/INV_1  ( .A(\RI1[1][91] ), .ZN(\SB1_1_16/i0[6] ) );
  INV_X1 \SB1_1_16/INV_0  ( .A(\RI1[1][90] ), .ZN(\SB1_1_16/i0[9] ) );
  BUF_X1 \SB1_1_16/BUF_5  ( .A(\RI1[1][95] ), .Z(\SB1_1_16/i1_5 ) );
  INV_X1 \SB1_1_17/INV_4  ( .A(\RI1[1][88] ), .ZN(\SB1_1_17/i0_4 ) );
  INV_X1 \SB1_1_17/INV_3  ( .A(\RI1[1][87] ), .ZN(\SB1_1_17/i0[10] ) );
  INV_X1 \SB1_1_17/INV_2  ( .A(\RI1[1][86] ), .ZN(\SB1_1_17/i0_0 ) );
  INV_X1 \SB1_1_17/INV_1  ( .A(\RI1[1][85] ), .ZN(\SB1_1_17/i0[6] ) );
  INV_X1 \SB1_1_17/INV_0  ( .A(\RI1[1][84] ), .ZN(\SB1_1_17/i0[9] ) );
  BUF_X1 \SB1_1_17/BUF_5  ( .A(\RI1[1][89] ), .Z(\SB1_1_17/i1_5 ) );
  INV_X1 \SB1_1_18/INV_4  ( .A(\RI1[1][82] ), .ZN(\SB1_1_18/i0_4 ) );
  INV_X1 \SB1_1_18/INV_3  ( .A(\RI1[1][81] ), .ZN(\SB1_1_18/i0[10] ) );
  INV_X1 \SB1_1_18/INV_2  ( .A(\RI1[1][80] ), .ZN(\SB1_1_18/i0_0 ) );
  INV_X1 \SB1_1_18/INV_1  ( .A(\RI1[1][79] ), .ZN(\SB1_1_18/i0[6] ) );
  BUF_X1 \SB1_1_18/BUF_5  ( .A(\RI1[1][83] ), .Z(\SB1_1_18/i1_5 ) );
  INV_X1 \SB1_1_19/INV_4  ( .A(\RI1[1][76] ), .ZN(\SB1_1_19/i0_4 ) );
  INV_X1 \SB1_1_19/INV_3  ( .A(\RI1[1][75] ), .ZN(\SB1_1_19/i0[10] ) );
  INV_X1 \SB1_1_19/INV_2  ( .A(\RI1[1][74] ), .ZN(\SB1_1_19/i0_0 ) );
  INV_X1 \SB1_1_19/INV_1  ( .A(\RI1[1][73] ), .ZN(\SB1_1_19/i0[6] ) );
  BUF_X1 \SB1_1_19/BUF_5  ( .A(\RI1[1][77] ), .Z(\SB1_1_19/i1_5 ) );
  INV_X1 \SB1_1_20/INV_4  ( .A(\RI1[1][70] ), .ZN(\SB1_1_20/i0_4 ) );
  INV_X1 \SB1_1_20/INV_2  ( .A(\RI1[1][68] ), .ZN(\SB1_1_20/i0_0 ) );
  BUF_X1 \SB1_1_20/BUF_5  ( .A(\RI1[1][71] ), .Z(\SB1_1_20/i1_5 ) );
  INV_X1 \SB1_1_21/INV_3  ( .A(\RI1[1][63] ), .ZN(\SB1_1_21/i0[10] ) );
  INV_X1 \SB1_1_21/INV_2  ( .A(\RI1[1][62] ), .ZN(\SB1_1_21/i0_0 ) );
  INV_X1 \SB1_1_21/INV_1  ( .A(\RI1[1][61] ), .ZN(\SB1_1_21/i0[6] ) );
  BUF_X1 \SB1_1_21/BUF_5  ( .A(\RI1[1][65] ), .Z(\SB1_1_21/i1_5 ) );
  BUF_X1 \SB1_1_21/BUF_1  ( .A(\RI1[1][61] ), .Z(\SB1_1_21/i1_7 ) );
  INV_X1 \SB1_1_22/INV_4  ( .A(\RI1[1][58] ), .ZN(\SB1_1_22/i0_4 ) );
  INV_X1 \SB1_1_22/INV_3  ( .A(\RI1[1][57] ), .ZN(\SB1_1_22/i0[10] ) );
  INV_X1 \SB1_1_22/INV_2  ( .A(\RI1[1][56] ), .ZN(\SB1_1_22/i0_0 ) );
  INV_X1 \SB1_1_22/INV_1  ( .A(\RI1[1][55] ), .ZN(\SB1_1_22/i0[6] ) );
  INV_X1 \SB1_1_22/INV_0  ( .A(\RI1[1][54] ), .ZN(\SB1_1_22/i0[9] ) );
  BUF_X1 \SB1_1_22/BUF_5  ( .A(\RI1[1][59] ), .Z(\SB1_1_22/i1_5 ) );
  INV_X1 \SB1_1_23/INV_4  ( .A(\RI1[1][52] ), .ZN(\SB1_1_23/i0_4 ) );
  INV_X1 \SB1_1_23/INV_3  ( .A(\RI1[1][51] ), .ZN(\SB1_1_23/i0[10] ) );
  INV_X1 \SB1_1_23/INV_2  ( .A(\RI1[1][50] ), .ZN(\SB1_1_23/i0_0 ) );
  INV_X1 \SB1_1_23/INV_1  ( .A(\RI1[1][49] ), .ZN(\SB1_1_23/i0[6] ) );
  INV_X1 \SB1_1_23/INV_0  ( .A(\RI1[1][48] ), .ZN(\SB1_1_23/i0[9] ) );
  BUF_X1 \SB1_1_23/BUF_5  ( .A(\RI1[1][53] ), .Z(\SB1_1_23/i1_5 ) );
  INV_X1 \SB1_1_24/INV_4  ( .A(\RI1[1][46] ), .ZN(\SB1_1_24/i0_4 ) );
  INV_X1 \SB1_1_24/INV_3  ( .A(\RI1[1][45] ), .ZN(\SB1_1_24/i0[10] ) );
  INV_X1 \SB1_1_24/INV_2  ( .A(\RI1[1][44] ), .ZN(\SB1_1_24/i0_0 ) );
  INV_X1 \SB1_1_24/INV_1  ( .A(\RI1[1][43] ), .ZN(\SB1_1_24/i0[6] ) );
  INV_X1 \SB1_1_25/INV_4  ( .A(\RI1[1][40] ), .ZN(\SB1_1_25/i0_4 ) );
  INV_X1 \SB1_1_25/INV_3  ( .A(\RI1[1][39] ), .ZN(\SB1_1_25/i0[10] ) );
  INV_X1 \SB1_1_25/INV_2  ( .A(\RI1[1][38] ), .ZN(\SB1_1_25/i0_0 ) );
  INV_X1 \SB1_1_25/INV_1  ( .A(\RI1[1][37] ), .ZN(\SB1_1_25/i0[6] ) );
  BUF_X1 \SB1_1_25/BUF_5  ( .A(\RI1[1][41] ), .Z(\SB1_1_25/i1_5 ) );
  INV_X1 \SB1_1_26/INV_3  ( .A(\RI1[1][33] ), .ZN(\SB1_1_26/i0[10] ) );
  INV_X1 \SB1_1_26/INV_2  ( .A(\RI1[1][32] ), .ZN(\SB1_1_26/i0_0 ) );
  INV_X1 \SB1_1_26/INV_1  ( .A(\RI1[1][31] ), .ZN(\SB1_1_26/i0[6] ) );
  BUF_X1 \SB1_1_26/BUF_5  ( .A(\RI1[1][35] ), .Z(\SB1_1_26/i1_5 ) );
  INV_X1 \SB1_1_27/INV_3  ( .A(\RI1[1][27] ), .ZN(\SB1_1_27/i0[10] ) );
  INV_X1 \SB1_1_27/INV_2  ( .A(\RI1[1][26] ), .ZN(\SB1_1_27/i0_0 ) );
  INV_X1 \SB1_1_27/INV_1  ( .A(\RI1[1][25] ), .ZN(\SB1_1_27/i0[6] ) );
  BUF_X1 \SB1_1_27/BUF_1  ( .A(\RI1[1][25] ), .Z(\SB1_1_27/i1_7 ) );
  INV_X1 \SB1_1_28/INV_4  ( .A(\RI1[1][22] ), .ZN(\SB1_1_28/i0_4 ) );
  INV_X1 \SB1_1_28/INV_3  ( .A(\RI1[1][21] ), .ZN(\SB1_1_28/i0[10] ) );
  INV_X1 \SB1_1_28/INV_2  ( .A(\RI1[1][20] ), .ZN(\SB1_1_28/i0_0 ) );
  INV_X1 \SB1_1_28/INV_1  ( .A(\RI1[1][19] ), .ZN(\SB1_1_28/i0[6] ) );
  INV_X1 \SB1_1_28/INV_0  ( .A(\RI1[1][18] ), .ZN(\SB1_1_28/i0[9] ) );
  BUF_X1 \SB1_1_28/BUF_5  ( .A(\RI1[1][23] ), .Z(\SB1_1_28/i1_5 ) );
  INV_X1 \SB1_1_29/INV_4  ( .A(\RI1[1][16] ), .ZN(\SB1_1_29/i0_4 ) );
  INV_X1 \SB1_1_29/INV_3  ( .A(\RI1[1][15] ), .ZN(\SB1_1_29/i0[10] ) );
  INV_X1 \SB1_1_29/INV_2  ( .A(\RI1[1][14] ), .ZN(\SB1_1_29/i0_0 ) );
  INV_X1 \SB1_1_29/INV_1  ( .A(\RI1[1][13] ), .ZN(\SB1_1_29/i0[6] ) );
  BUF_X1 \SB1_1_29/BUF_5  ( .A(\RI1[1][17] ), .Z(\SB1_1_29/i1_5 ) );
  INV_X1 \SB1_1_30/INV_3  ( .A(\RI1[1][9] ), .ZN(\SB1_1_30/i0[10] ) );
  INV_X1 \SB1_1_30/INV_2  ( .A(\RI1[1][8] ), .ZN(\SB1_1_30/i0_0 ) );
  INV_X1 \SB1_1_30/INV_1  ( .A(\RI1[1][7] ), .ZN(\SB1_1_30/i0[6] ) );
  BUF_X1 \SB1_1_30/BUF_5  ( .A(\RI1[1][11] ), .Z(\SB1_1_30/i1_5 ) );
  INV_X1 \SB1_1_31/INV_3  ( .A(\RI1[1][3] ), .ZN(\SB1_1_31/i0[10] ) );
  INV_X1 \SB1_1_31/INV_2  ( .A(\RI1[1][2] ), .ZN(\SB1_1_31/i0_0 ) );
  INV_X1 \SB1_1_31/INV_1  ( .A(\RI1[1][1] ), .ZN(\SB1_1_31/i0[6] ) );
  BUF_X1 \SB1_1_31/BUF_5  ( .A(\RI1[1][5] ), .Z(\SB1_1_31/i1_5 ) );
  INV_X1 \SB1_2_0/INV_4  ( .A(\RI1[2][190] ), .ZN(\SB1_2_0/i0_4 ) );
  INV_X1 \SB1_2_0/INV_3  ( .A(\RI1[2][189] ), .ZN(\SB1_2_0/i0[10] ) );
  INV_X1 \SB1_2_0/INV_2  ( .A(\RI1[2][188] ), .ZN(\SB1_2_0/i0_0 ) );
  INV_X1 \SB1_2_0/INV_1  ( .A(\RI1[2][187] ), .ZN(\SB1_2_0/i0[6] ) );
  INV_X1 \SB1_2_1/INV_3  ( .A(\RI1[2][183] ), .ZN(\SB1_2_1/i0[10] ) );
  INV_X1 \SB1_2_1/INV_2  ( .A(\RI1[2][182] ), .ZN(\SB1_2_1/i0_0 ) );
  INV_X1 \SB1_2_1/INV_1  ( .A(\RI1[2][181] ), .ZN(\SB1_2_1/i0[6] ) );
  INV_X1 \SB1_2_1/INV_0  ( .A(\RI1[2][180] ), .ZN(\SB1_2_1/i0[9] ) );
  BUF_X1 \SB1_2_1/BUF_5  ( .A(\RI1[2][185] ), .Z(\SB1_2_1/i1_5 ) );
  INV_X1 \SB1_2_2/INV_3  ( .A(\RI1[2][177] ), .ZN(\SB1_2_2/i0[10] ) );
  INV_X1 \SB1_2_2/INV_2  ( .A(\RI1[2][176] ), .ZN(\SB1_2_2/i0_0 ) );
  INV_X1 \SB1_2_2/INV_1  ( .A(\RI1[2][175] ), .ZN(\SB1_2_2/i0[6] ) );
  INV_X1 \SB1_2_3/INV_3  ( .A(\RI1[2][171] ), .ZN(\SB1_2_3/i0[10] ) );
  INV_X1 \SB1_2_3/INV_2  ( .A(\RI1[2][170] ), .ZN(\SB1_2_3/i0_0 ) );
  INV_X1 \SB1_2_3/INV_1  ( .A(\RI1[2][169] ), .ZN(\SB1_2_3/i0[6] ) );
  BUF_X1 \SB1_2_3/BUF_5  ( .A(\RI1[2][173] ), .Z(\SB1_2_3/i1_5 ) );
  INV_X1 \SB1_2_4/INV_3  ( .A(\RI1[2][165] ), .ZN(\SB1_2_4/i0[10] ) );
  INV_X1 \SB1_2_4/INV_2  ( .A(\RI1[2][164] ), .ZN(\SB1_2_4/i0_0 ) );
  INV_X1 \SB1_2_4/INV_1  ( .A(\RI1[2][163] ), .ZN(\SB1_2_4/i0[6] ) );
  BUF_X1 \SB1_2_4/BUF_5  ( .A(\RI1[2][167] ), .Z(\SB1_2_4/i1_5 ) );
  INV_X1 \SB1_2_5/INV_4  ( .A(\RI1[2][160] ), .ZN(\SB1_2_5/i0_4 ) );
  INV_X1 \SB1_2_5/INV_3  ( .A(\RI1[2][159] ), .ZN(\SB1_2_5/i0[10] ) );
  INV_X1 \SB1_2_5/INV_1  ( .A(\RI1[2][157] ), .ZN(\SB1_2_5/i0[6] ) );
  BUF_X1 \SB1_2_5/BUF_5  ( .A(\RI1[2][161] ), .Z(\SB1_2_5/i1_5 ) );
  INV_X1 \SB1_2_6/INV_2  ( .A(\RI1[2][152] ), .ZN(\SB1_2_6/i0_0 ) );
  INV_X1 \SB1_2_6/INV_1  ( .A(\RI1[2][151] ), .ZN(\SB1_2_6/i0[6] ) );
  BUF_X1 \SB1_2_6/BUF_5  ( .A(\RI1[2][155] ), .Z(\SB1_2_6/i1_5 ) );
  INV_X1 \SB1_2_7/INV_3  ( .A(\RI1[2][147] ), .ZN(\SB1_2_7/i0[10] ) );
  INV_X1 \SB1_2_7/INV_2  ( .A(\RI1[2][146] ), .ZN(\SB1_2_7/i0_0 ) );
  INV_X1 \SB1_2_7/INV_1  ( .A(\RI1[2][145] ), .ZN(\SB1_2_7/i0[6] ) );
  BUF_X1 \SB1_2_7/BUF_5  ( .A(\RI1[2][149] ), .Z(\SB1_2_7/i1_5 ) );
  INV_X1 \SB1_2_8/INV_4  ( .A(\RI1[2][142] ), .ZN(\SB1_2_8/i0_4 ) );
  INV_X1 \SB1_2_8/INV_3  ( .A(\RI1[2][141] ), .ZN(\SB1_2_8/i0[10] ) );
  INV_X1 \SB1_2_8/INV_2  ( .A(\RI1[2][140] ), .ZN(\SB1_2_8/i0_0 ) );
  INV_X1 \SB1_2_8/INV_1  ( .A(\RI1[2][139] ), .ZN(\SB1_2_8/i0[6] ) );
  BUF_X1 \SB1_2_8/BUF_5  ( .A(\RI1[2][143] ), .Z(\SB1_2_8/i1_5 ) );
  INV_X1 \SB1_2_9/INV_4  ( .A(\RI1[2][136] ), .ZN(\SB1_2_9/i0_4 ) );
  INV_X1 \SB1_2_9/INV_3  ( .A(\RI1[2][135] ), .ZN(\SB1_2_9/i0[10] ) );
  INV_X1 \SB1_2_9/INV_2  ( .A(\RI1[2][134] ), .ZN(\SB1_2_9/i0_0 ) );
  INV_X1 \SB1_2_9/INV_1  ( .A(\RI1[2][133] ), .ZN(\SB1_2_9/i0[6] ) );
  INV_X1 \SB1_2_9/INV_0  ( .A(\RI1[2][132] ), .ZN(\SB1_2_9/i0[9] ) );
  BUF_X1 \SB1_2_9/BUF_5  ( .A(\RI1[2][137] ), .Z(\SB1_2_9/i1_5 ) );
  INV_X1 \SB1_2_10/INV_3  ( .A(\RI1[2][129] ), .ZN(\SB1_2_10/i0[10] ) );
  INV_X1 \SB1_2_10/INV_2  ( .A(\RI1[2][128] ), .ZN(\SB1_2_10/i0_0 ) );
  INV_X1 \SB1_2_10/INV_1  ( .A(\RI1[2][127] ), .ZN(\SB1_2_10/i0[6] ) );
  INV_X1 \SB1_2_10/INV_0  ( .A(\RI1[2][126] ), .ZN(\SB1_2_10/i0[9] ) );
  BUF_X1 \SB1_2_10/BUF_5  ( .A(\RI1[2][131] ), .Z(\SB1_2_10/i1_5 ) );
  INV_X1 \SB1_2_11/INV_4  ( .A(\RI1[2][124] ), .ZN(\SB1_2_11/i0_4 ) );
  INV_X1 \SB1_2_11/INV_3  ( .A(\RI1[2][123] ), .ZN(\SB1_2_11/i0[10] ) );
  INV_X1 \SB1_2_11/INV_2  ( .A(\RI1[2][122] ), .ZN(\SB1_2_11/i0_0 ) );
  INV_X1 \SB1_2_11/INV_1  ( .A(\RI1[2][121] ), .ZN(\SB1_2_11/i0[6] ) );
  BUF_X1 \SB1_2_11/BUF_5  ( .A(\RI1[2][125] ), .Z(\SB1_2_11/i1_5 ) );
  INV_X1 \SB1_2_12/INV_3  ( .A(\RI1[2][117] ), .ZN(\SB1_2_12/i0[10] ) );
  INV_X1 \SB1_2_12/INV_2  ( .A(\RI1[2][116] ), .ZN(\SB1_2_12/i0_0 ) );
  BUF_X1 \SB1_2_12/BUF_5  ( .A(\RI1[2][119] ), .Z(\SB1_2_12/i1_5 ) );
  INV_X1 \SB1_2_13/INV_3  ( .A(\RI1[2][111] ), .ZN(\SB1_2_13/i0[10] ) );
  INV_X1 \SB1_2_13/INV_1  ( .A(\RI1[2][109] ), .ZN(\SB1_2_13/i0[6] ) );
  BUF_X1 \SB1_2_13/BUF_5  ( .A(\RI1[2][113] ), .Z(\SB1_2_13/i1_5 ) );
  INV_X1 \SB1_2_14/INV_3  ( .A(\RI1[2][105] ), .ZN(\SB1_2_14/i0[10] ) );
  INV_X1 \SB1_2_14/INV_2  ( .A(\RI1[2][104] ), .ZN(\SB1_2_14/i0_0 ) );
  INV_X1 \SB1_2_14/INV_1  ( .A(\RI1[2][103] ), .ZN(\SB1_2_14/i0[6] ) );
  INV_X1 \SB1_2_14/INV_0  ( .A(\RI1[2][102] ), .ZN(\SB1_2_14/i0[9] ) );
  BUF_X1 \SB1_2_14/BUF_5  ( .A(\RI1[2][107] ), .Z(\SB1_2_14/i1_5 ) );
  INV_X1 \SB1_2_15/INV_3  ( .A(\RI1[2][99] ), .ZN(\SB1_2_15/i0[10] ) );
  INV_X1 \SB1_2_15/INV_2  ( .A(\RI1[2][98] ), .ZN(\SB1_2_15/i0_0 ) );
  INV_X1 \SB1_2_15/INV_1  ( .A(\RI1[2][97] ), .ZN(\SB1_2_15/i0[6] ) );
  INV_X1 \SB1_2_15/INV_0  ( .A(\RI1[2][96] ), .ZN(\SB1_2_15/i0[9] ) );
  BUF_X1 \SB1_2_15/BUF_5  ( .A(\RI1[2][101] ), .Z(\SB1_2_15/i1_5 ) );
  INV_X1 \SB1_2_16/INV_4  ( .A(\RI1[2][94] ), .ZN(\SB1_2_16/i0_4 ) );
  INV_X1 \SB1_2_16/INV_3  ( .A(\RI1[2][93] ), .ZN(\SB1_2_16/i0[10] ) );
  INV_X1 \SB1_2_16/INV_2  ( .A(\RI1[2][92] ), .ZN(\SB1_2_16/i0_0 ) );
  BUF_X1 \SB1_2_16/BUF_5  ( .A(\RI1[2][95] ), .Z(\SB1_2_16/i1_5 ) );
  INV_X1 \SB1_2_17/INV_3  ( .A(\RI1[2][87] ), .ZN(\SB1_2_17/i0[10] ) );
  INV_X1 \SB1_2_17/INV_2  ( .A(\RI1[2][86] ), .ZN(\SB1_2_17/i0_0 ) );
  INV_X1 \SB1_2_17/INV_1  ( .A(\RI1[2][85] ), .ZN(\SB1_2_17/i0[6] ) );
  BUF_X1 \SB1_2_17/BUF_5  ( .A(\RI1[2][89] ), .Z(\SB1_2_17/i1_5 ) );
  INV_X1 \SB1_2_18/INV_4  ( .A(\RI1[2][82] ), .ZN(\SB1_2_18/i0_4 ) );
  INV_X1 \SB1_2_18/INV_3  ( .A(\RI1[2][81] ), .ZN(\SB1_2_18/i0[10] ) );
  INV_X1 \SB1_2_18/INV_2  ( .A(\RI1[2][80] ), .ZN(\SB1_2_18/i0_0 ) );
  INV_X1 \SB1_2_18/INV_1  ( .A(\RI1[2][79] ), .ZN(\SB1_2_18/i0[6] ) );
  BUF_X1 \SB1_2_18/BUF_5  ( .A(\RI1[2][83] ), .Z(\SB1_2_18/i1_5 ) );
  INV_X1 \SB1_2_19/INV_4  ( .A(\RI1[2][76] ), .ZN(\SB1_2_19/i0_4 ) );
  INV_X1 \SB1_2_19/INV_3  ( .A(\RI1[2][75] ), .ZN(\SB1_2_19/i0[10] ) );
  INV_X1 \SB1_2_19/INV_2  ( .A(\RI1[2][74] ), .ZN(\SB1_2_19/i0_0 ) );
  INV_X1 \SB1_2_19/INV_1  ( .A(\RI1[2][73] ), .ZN(\SB1_2_19/i0[6] ) );
  BUF_X1 \SB1_2_19/BUF_5  ( .A(\RI1[2][77] ), .Z(\SB1_2_19/i1_5 ) );
  INV_X1 \SB1_2_20/INV_4  ( .A(\RI1[2][70] ), .ZN(\SB1_2_20/i0_4 ) );
  INV_X1 \SB1_2_20/INV_3  ( .A(\RI1[2][69] ), .ZN(\SB1_2_20/i0[10] ) );
  INV_X1 \SB1_2_20/INV_2  ( .A(\RI1[2][68] ), .ZN(\SB1_2_20/i0_0 ) );
  INV_X1 \SB1_2_20/INV_1  ( .A(\RI1[2][67] ), .ZN(\SB1_2_20/i0[6] ) );
  BUF_X1 \SB1_2_20/BUF_5  ( .A(\RI1[2][71] ), .Z(\SB1_2_20/i1_5 ) );
  INV_X1 \SB1_2_21/INV_4  ( .A(\RI1[2][64] ), .ZN(\SB1_2_21/i0_4 ) );
  INV_X1 \SB1_2_21/INV_3  ( .A(\RI1[2][63] ), .ZN(\SB1_2_21/i0[10] ) );
  INV_X1 \SB1_2_21/INV_2  ( .A(\RI1[2][62] ), .ZN(\SB1_2_21/i0_0 ) );
  INV_X1 \SB1_2_21/INV_1  ( .A(\RI1[2][61] ), .ZN(\SB1_2_21/i0[6] ) );
  INV_X1 \SB1_2_21/INV_0  ( .A(\RI1[2][60] ), .ZN(\SB1_2_21/i0[9] ) );
  BUF_X1 \SB1_2_21/BUF_5  ( .A(\RI1[2][65] ), .Z(\SB1_2_21/i1_5 ) );
  INV_X1 \SB1_2_22/INV_3  ( .A(\RI1[2][57] ), .ZN(\SB1_2_22/i0[10] ) );
  INV_X1 \SB1_2_22/INV_2  ( .A(\RI1[2][56] ), .ZN(\SB1_2_22/i0_0 ) );
  INV_X1 \SB1_2_22/INV_1  ( .A(\RI1[2][55] ), .ZN(\SB1_2_22/i0[6] ) );
  BUF_X1 \SB1_2_22/BUF_5  ( .A(\RI1[2][59] ), .Z(\SB1_2_22/i1_5 ) );
  INV_X1 \SB1_2_23/INV_4  ( .A(\RI1[2][52] ), .ZN(\SB1_2_23/i0_4 ) );
  INV_X1 \SB1_2_23/INV_3  ( .A(\RI1[2][51] ), .ZN(\SB1_2_23/i0[10] ) );
  INV_X1 \SB1_2_23/INV_2  ( .A(\RI1[2][50] ), .ZN(\SB1_2_23/i0_0 ) );
  INV_X1 \SB1_2_23/INV_1  ( .A(\RI1[2][49] ), .ZN(\SB1_2_23/i0[6] ) );
  BUF_X1 \SB1_2_23/BUF_5  ( .A(\RI1[2][53] ), .Z(\SB1_2_23/i1_5 ) );
  INV_X1 \SB1_2_24/INV_3  ( .A(\RI1[2][45] ), .ZN(\SB1_2_24/i0[10] ) );
  INV_X1 \SB1_2_24/INV_2  ( .A(\RI1[2][44] ), .ZN(\SB1_2_24/i0_0 ) );
  INV_X1 \SB1_2_24/INV_1  ( .A(\RI1[2][43] ), .ZN(\SB1_2_24/i0[6] ) );
  BUF_X1 \SB1_2_24/BUF_5  ( .A(\RI1[2][47] ), .Z(\SB1_2_24/i1_5 ) );
  INV_X1 \SB1_2_25/INV_3  ( .A(\RI1[2][39] ), .ZN(\SB1_2_25/i0[10] ) );
  INV_X1 \SB1_2_25/INV_2  ( .A(\RI1[2][38] ), .ZN(\SB1_2_25/i0_0 ) );
  INV_X1 \SB1_2_25/INV_1  ( .A(\RI1[2][37] ), .ZN(\SB1_2_25/i0[6] ) );
  INV_X1 \SB1_2_25/INV_0  ( .A(\RI1[2][36] ), .ZN(\SB1_2_25/i0[9] ) );
  BUF_X1 \SB1_2_25/BUF_5  ( .A(\RI1[2][41] ), .Z(\SB1_2_25/i1_5 ) );
  INV_X1 \SB1_2_26/INV_3  ( .A(\RI1[2][33] ), .ZN(\SB1_2_26/i0[10] ) );
  INV_X1 \SB1_2_26/INV_2  ( .A(\RI1[2][32] ), .ZN(\SB1_2_26/i0_0 ) );
  INV_X1 \SB1_2_26/INV_1  ( .A(\RI1[2][31] ), .ZN(\SB1_2_26/i0[6] ) );
  BUF_X1 \SB1_2_26/BUF_5  ( .A(\RI1[2][35] ), .Z(\SB1_2_26/i1_5 ) );
  INV_X1 \SB1_2_27/INV_4  ( .A(\RI1[2][28] ), .ZN(\SB1_2_27/i0_4 ) );
  INV_X1 \SB1_2_27/INV_3  ( .A(\RI1[2][27] ), .ZN(\SB1_2_27/i0[10] ) );
  INV_X1 \SB1_2_27/INV_2  ( .A(\RI1[2][26] ), .ZN(\SB1_2_27/i0_0 ) );
  INV_X1 \SB1_2_27/INV_1  ( .A(\RI1[2][25] ), .ZN(\SB1_2_27/i0[6] ) );
  BUF_X1 \SB1_2_27/BUF_5  ( .A(\RI1[2][29] ), .Z(\SB1_2_27/i1_5 ) );
  INV_X1 \SB1_2_28/INV_4  ( .A(\RI1[2][22] ), .ZN(\SB1_2_28/i0_4 ) );
  INV_X1 \SB1_2_28/INV_3  ( .A(\RI1[2][21] ), .ZN(\SB1_2_28/i0[10] ) );
  INV_X1 \SB1_2_28/INV_2  ( .A(\RI1[2][20] ), .ZN(\SB1_2_28/i0_0 ) );
  INV_X1 \SB1_2_28/INV_1  ( .A(\RI1[2][19] ), .ZN(\SB1_2_28/i0[6] ) );
  BUF_X1 \SB1_2_28/BUF_5  ( .A(\RI1[2][23] ), .Z(\SB1_2_28/i1_5 ) );
  INV_X1 \SB1_2_29/INV_4  ( .A(\RI1[2][16] ), .ZN(\SB1_2_29/i0_4 ) );
  INV_X1 \SB1_2_29/INV_2  ( .A(\RI1[2][14] ), .ZN(\SB1_2_29/i0_0 ) );
  INV_X1 \SB1_2_29/INV_1  ( .A(\RI1[2][13] ), .ZN(\SB1_2_29/i0[6] ) );
  INV_X1 \SB1_2_29/INV_0  ( .A(\RI1[2][12] ), .ZN(\SB1_2_29/i0[9] ) );
  INV_X1 \SB1_2_30/INV_3  ( .A(\RI1[2][9] ), .ZN(\SB1_2_30/i0[10] ) );
  INV_X1 \SB1_2_30/INV_2  ( .A(\RI1[2][8] ), .ZN(\SB1_2_30/i0_0 ) );
  INV_X1 \SB1_2_30/INV_1  ( .A(\RI1[2][7] ), .ZN(\SB1_2_30/i0[6] ) );
  BUF_X1 \SB1_2_30/BUF_5  ( .A(\RI1[2][11] ), .Z(\SB1_2_30/i1_5 ) );
  INV_X1 \SB1_2_31/INV_4  ( .A(\RI1[2][4] ), .ZN(\SB1_2_31/i0_4 ) );
  INV_X1 \SB1_2_31/INV_2  ( .A(\RI1[2][2] ), .ZN(\SB1_2_31/i0_0 ) );
  INV_X1 \SB1_2_31/INV_0  ( .A(\RI1[2][0] ), .ZN(\SB1_2_31/i0[9] ) );
  BUF_X1 \SB1_2_31/BUF_5  ( .A(\RI1[2][5] ), .Z(\SB1_2_31/i1_5 ) );
  INV_X1 \SB1_3_0/INV_3  ( .A(\RI1[3][189] ), .ZN(\SB1_3_0/i0[10] ) );
  INV_X1 \SB1_3_0/INV_2  ( .A(\RI1[3][188] ), .ZN(\SB1_3_0/i0_0 ) );
  INV_X1 \SB1_3_0/INV_1  ( .A(\RI1[3][187] ), .ZN(\SB1_3_0/i0[6] ) );
  INV_X1 \SB1_3_0/INV_0  ( .A(\RI1[3][186] ), .ZN(\SB1_3_0/i0[9] ) );
  BUF_X1 \SB1_3_0/BUF_5  ( .A(\RI1[3][191] ), .Z(\SB1_3_0/i1_5 ) );
  INV_X1 \SB1_3_1/INV_3  ( .A(\RI1[3][183] ), .ZN(\SB1_3_1/i0[10] ) );
  INV_X1 \SB1_3_1/INV_2  ( .A(\RI1[3][182] ), .ZN(\SB1_3_1/i0_0 ) );
  INV_X1 \SB1_3_1/INV_1  ( .A(\RI1[3][181] ), .ZN(\SB1_3_1/i0[6] ) );
  INV_X1 \SB1_3_2/INV_3  ( .A(\RI1[3][177] ), .ZN(\SB1_3_2/i0[10] ) );
  INV_X1 \SB1_3_2/INV_2  ( .A(\RI1[3][176] ), .ZN(\SB1_3_2/i0_0 ) );
  INV_X1 \SB1_3_2/INV_1  ( .A(\RI1[3][175] ), .ZN(\SB1_3_2/i0[6] ) );
  INV_X1 \SB1_3_2/INV_0  ( .A(\RI1[3][174] ), .ZN(\SB1_3_2/i0[9] ) );
  BUF_X1 \SB1_3_2/BUF_5  ( .A(\RI1[3][179] ), .Z(\SB1_3_2/i1_5 ) );
  INV_X1 \SB1_3_3/INV_3  ( .A(\RI1[3][171] ), .ZN(\SB1_3_3/i0[10] ) );
  INV_X1 \SB1_3_3/INV_2  ( .A(\RI1[3][170] ), .ZN(\SB1_3_3/i0_0 ) );
  INV_X1 \SB1_3_3/INV_1  ( .A(\RI1[3][169] ), .ZN(\SB1_3_3/i0[6] ) );
  INV_X1 \SB1_3_3/INV_0  ( .A(\RI1[3][168] ), .ZN(\SB1_3_3/i0[9] ) );
  BUF_X1 \SB1_3_3/BUF_5  ( .A(\RI1[3][173] ), .Z(\SB1_3_3/i1_5 ) );
  INV_X1 \SB1_3_4/INV_3  ( .A(\RI1[3][165] ), .ZN(\SB1_3_4/i0[10] ) );
  INV_X1 \SB1_3_4/INV_2  ( .A(\RI1[3][164] ), .ZN(\SB1_3_4/i0_0 ) );
  INV_X1 \SB1_3_4/INV_1  ( .A(\RI1[3][163] ), .ZN(\SB1_3_4/i0[6] ) );
  INV_X1 \SB1_3_4/INV_0  ( .A(\RI1[3][162] ), .ZN(\SB1_3_4/i0[9] ) );
  BUF_X1 \SB1_3_4/BUF_5  ( .A(\RI1[3][167] ), .Z(\SB1_3_4/i1_5 ) );
  INV_X1 \SB1_3_5/INV_4  ( .A(\RI1[3][160] ), .ZN(\SB1_3_5/i0_4 ) );
  INV_X1 \SB1_3_5/INV_3  ( .A(\RI1[3][159] ), .ZN(\SB1_3_5/i0[10] ) );
  INV_X1 \SB1_3_5/INV_2  ( .A(\RI1[3][158] ), .ZN(\SB1_3_5/i0_0 ) );
  INV_X1 \SB1_3_5/INV_1  ( .A(\RI1[3][157] ), .ZN(\SB1_3_5/i0[6] ) );
  INV_X1 \SB1_3_5/INV_0  ( .A(\RI1[3][156] ), .ZN(\SB1_3_5/i0[9] ) );
  BUF_X1 \SB1_3_5/BUF_5  ( .A(\RI1[3][161] ), .Z(\SB1_3_5/i1_5 ) );
  INV_X1 \SB1_3_6/INV_4  ( .A(\RI1[3][154] ), .ZN(\SB1_3_6/i0_4 ) );
  INV_X1 \SB1_3_6/INV_3  ( .A(\RI1[3][153] ), .ZN(\SB1_3_6/i0[10] ) );
  INV_X1 \SB1_3_6/INV_2  ( .A(\RI1[3][152] ), .ZN(\SB1_3_6/i0_0 ) );
  INV_X1 \SB1_3_6/INV_1  ( .A(\RI1[3][151] ), .ZN(\SB1_3_6/i0[6] ) );
  INV_X1 \SB1_3_6/INV_0  ( .A(\RI1[3][150] ), .ZN(\SB1_3_6/i0[9] ) );
  BUF_X1 \SB1_3_6/BUF_5  ( .A(\RI1[3][155] ), .Z(\SB1_3_6/i1_5 ) );
  INV_X1 \SB1_3_7/INV_3  ( .A(\RI1[3][147] ), .ZN(\SB1_3_7/i0[10] ) );
  INV_X1 \SB1_3_7/INV_2  ( .A(\RI1[3][146] ), .ZN(\SB1_3_7/i0_0 ) );
  INV_X1 \SB1_3_7/INV_1  ( .A(\RI1[3][145] ), .ZN(\SB1_3_7/i0[6] ) );
  INV_X1 \SB1_3_7/INV_0  ( .A(\RI1[3][144] ), .ZN(\SB1_3_7/i0[9] ) );
  BUF_X1 \SB1_3_7/BUF_5  ( .A(\RI1[3][149] ), .Z(\SB1_3_7/i1_5 ) );
  INV_X1 \SB1_3_8/INV_3  ( .A(\RI1[3][141] ), .ZN(\SB1_3_8/i0[10] ) );
  INV_X1 \SB1_3_8/INV_2  ( .A(\RI1[3][140] ), .ZN(\SB1_3_8/i0_0 ) );
  INV_X1 \SB1_3_8/INV_1  ( .A(\RI1[3][139] ), .ZN(\SB1_3_8/i0[6] ) );
  INV_X1 \SB1_3_8/INV_0  ( .A(\RI1[3][138] ), .ZN(\SB1_3_8/i0[9] ) );
  BUF_X1 \SB1_3_8/BUF_5  ( .A(\RI1[3][143] ), .Z(\SB1_3_8/i1_5 ) );
  INV_X1 \SB1_3_9/INV_4  ( .A(\RI1[3][136] ), .ZN(\SB1_3_9/i0_4 ) );
  INV_X1 \SB1_3_9/INV_3  ( .A(\RI1[3][135] ), .ZN(\SB1_3_9/i0[10] ) );
  INV_X1 \SB1_3_9/INV_2  ( .A(\RI1[3][134] ), .ZN(\SB1_3_9/i0_0 ) );
  INV_X1 \SB1_3_9/INV_1  ( .A(\RI1[3][133] ), .ZN(\SB1_3_9/i0[6] ) );
  INV_X1 \SB1_3_9/INV_0  ( .A(\RI1[3][132] ), .ZN(\SB1_3_9/i0[9] ) );
  BUF_X1 \SB1_3_9/BUF_5  ( .A(\RI1[3][137] ), .Z(\SB1_3_9/i1_5 ) );
  INV_X1 \SB1_3_10/INV_4  ( .A(\RI1[3][130] ), .ZN(\SB1_3_10/i0_4 ) );
  INV_X1 \SB1_3_10/INV_3  ( .A(\RI1[3][129] ), .ZN(\SB1_3_10/i0[10] ) );
  INV_X1 \SB1_3_10/INV_2  ( .A(\RI1[3][128] ), .ZN(\SB1_3_10/i0_0 ) );
  INV_X1 \SB1_3_10/INV_1  ( .A(\RI1[3][127] ), .ZN(\SB1_3_10/i0[6] ) );
  BUF_X1 \SB1_3_10/BUF_5  ( .A(\RI1[3][131] ), .Z(\SB1_3_10/i1_5 ) );
  INV_X1 \SB1_3_11/INV_3  ( .A(\RI1[3][123] ), .ZN(\SB1_3_11/i0[10] ) );
  INV_X1 \SB1_3_11/INV_2  ( .A(\RI1[3][122] ), .ZN(\SB1_3_11/i0_0 ) );
  INV_X1 \SB1_3_11/INV_1  ( .A(\RI1[3][121] ), .ZN(\SB1_3_11/i0[6] ) );
  BUF_X1 \SB1_3_11/BUF_5  ( .A(\RI1[3][125] ), .Z(\SB1_3_11/i1_5 ) );
  INV_X1 \SB1_3_12/INV_3  ( .A(\RI1[3][117] ), .ZN(\SB1_3_12/i0[10] ) );
  INV_X1 \SB1_3_12/INV_2  ( .A(\RI1[3][116] ), .ZN(\SB1_3_12/i0_0 ) );
  INV_X1 \SB1_3_12/INV_1  ( .A(\RI1[3][115] ), .ZN(\SB1_3_12/i0[6] ) );
  INV_X1 \SB1_3_12/INV_0  ( .A(\RI1[3][114] ), .ZN(\SB1_3_12/i0[9] ) );
  BUF_X1 \SB1_3_12/BUF_5  ( .A(\RI1[3][119] ), .Z(\SB1_3_12/i1_5 ) );
  INV_X1 \SB1_3_13/INV_4  ( .A(\RI1[3][112] ), .ZN(\SB1_3_13/i0_4 ) );
  INV_X1 \SB1_3_13/INV_3  ( .A(\RI1[3][111] ), .ZN(\SB1_3_13/i0[10] ) );
  INV_X1 \SB1_3_13/INV_2  ( .A(\RI1[3][110] ), .ZN(\SB1_3_13/i0_0 ) );
  INV_X1 \SB1_3_13/INV_1  ( .A(\RI1[3][109] ), .ZN(\SB1_3_13/i0[6] ) );
  INV_X1 \SB1_3_13/INV_0  ( .A(\RI1[3][108] ), .ZN(\SB1_3_13/i0[9] ) );
  BUF_X1 \SB1_3_13/BUF_5  ( .A(\RI1[3][113] ), .Z(\SB1_3_13/i1_5 ) );
  INV_X1 \SB1_3_14/INV_3  ( .A(\RI1[3][105] ), .ZN(\SB1_3_14/i0[10] ) );
  INV_X1 \SB1_3_14/INV_2  ( .A(\RI1[3][104] ), .ZN(\SB1_3_14/i0_0 ) );
  INV_X1 \SB1_3_14/INV_1  ( .A(\RI1[3][103] ), .ZN(\SB1_3_14/i0[6] ) );
  BUF_X1 \SB1_3_14/BUF_5  ( .A(\RI1[3][107] ), .Z(\SB1_3_14/i1_5 ) );
  INV_X1 \SB1_3_15/INV_4  ( .A(\RI1[3][100] ), .ZN(\SB1_3_15/i0_4 ) );
  INV_X1 \SB1_3_15/INV_2  ( .A(\RI1[3][98] ), .ZN(\SB1_3_15/i0_0 ) );
  INV_X1 \SB1_3_15/INV_1  ( .A(\RI1[3][97] ), .ZN(\SB1_3_15/i0[6] ) );
  BUF_X1 \SB1_3_15/BUF_5  ( .A(\RI1[3][101] ), .Z(\SB1_3_15/i1_5 ) );
  INV_X1 \SB1_3_16/INV_3  ( .A(\RI1[3][93] ), .ZN(\SB1_3_16/i0[10] ) );
  INV_X1 \SB1_3_16/INV_2  ( .A(\RI1[3][92] ), .ZN(\SB1_3_16/i0_0 ) );
  INV_X1 \SB1_3_16/INV_1  ( .A(\RI1[3][91] ), .ZN(\SB1_3_16/i0[6] ) );
  BUF_X1 \SB1_3_16/BUF_5  ( .A(\RI1[3][95] ), .Z(\SB1_3_16/i1_5 ) );
  INV_X1 \SB1_3_17/INV_3  ( .A(\RI1[3][87] ), .ZN(\SB1_3_17/i0[10] ) );
  INV_X1 \SB1_3_17/INV_2  ( .A(\RI1[3][86] ), .ZN(\SB1_3_17/i0_0 ) );
  INV_X1 \SB1_3_17/INV_1  ( .A(\RI1[3][85] ), .ZN(\SB1_3_17/i0[6] ) );
  INV_X1 \SB1_3_17/INV_0  ( .A(\RI1[3][84] ), .ZN(\SB1_3_17/i0[9] ) );
  BUF_X1 \SB1_3_17/BUF_5  ( .A(\RI1[3][89] ), .Z(\SB1_3_17/i1_5 ) );
  INV_X1 \SB1_3_18/INV_3  ( .A(\RI1[3][81] ), .ZN(\SB1_3_18/i0[10] ) );
  INV_X1 \SB1_3_18/INV_2  ( .A(\RI1[3][80] ), .ZN(\SB1_3_18/i0_0 ) );
  INV_X1 \SB1_3_18/INV_1  ( .A(\RI1[3][79] ), .ZN(\SB1_3_18/i0[6] ) );
  BUF_X1 \SB1_3_18/BUF_5  ( .A(\RI1[3][83] ), .Z(\SB1_3_18/i1_5 ) );
  INV_X1 \SB1_3_19/INV_3  ( .A(\RI1[3][75] ), .ZN(\SB1_3_19/i0[10] ) );
  INV_X1 \SB1_3_19/INV_2  ( .A(\RI1[3][74] ), .ZN(\SB1_3_19/i0_0 ) );
  INV_X1 \SB1_3_19/INV_1  ( .A(\RI1[3][73] ), .ZN(\SB1_3_19/i0[6] ) );
  INV_X1 \SB1_3_19/INV_0  ( .A(\RI1[3][72] ), .ZN(\SB1_3_19/i0[9] ) );
  BUF_X1 \SB1_3_19/BUF_5  ( .A(\RI1[3][77] ), .Z(\SB1_3_19/i1_5 ) );
  INV_X1 \SB1_3_20/INV_4  ( .A(\RI1[3][70] ), .ZN(\SB1_3_20/i0_4 ) );
  INV_X1 \SB1_3_20/INV_3  ( .A(\RI1[3][69] ), .ZN(\SB1_3_20/i0[10] ) );
  INV_X1 \SB1_3_20/INV_2  ( .A(\RI1[3][68] ), .ZN(\SB1_3_20/i0_0 ) );
  INV_X1 \SB1_3_20/INV_1  ( .A(\RI1[3][67] ), .ZN(\SB1_3_20/i0[6] ) );
  BUF_X1 \SB1_3_20/BUF_5  ( .A(\RI1[3][71] ), .Z(\SB1_3_20/i1_5 ) );
  INV_X1 \SB1_3_21/INV_4  ( .A(\RI1[3][64] ), .ZN(\SB1_3_21/i0_4 ) );
  INV_X1 \SB1_3_21/INV_3  ( .A(\RI1[3][63] ), .ZN(\SB1_3_21/i0[10] ) );
  INV_X1 \SB1_3_21/INV_1  ( .A(\RI1[3][61] ), .ZN(\SB1_3_21/i0[6] ) );
  INV_X1 \SB1_3_21/INV_0  ( .A(\RI1[3][60] ), .ZN(\SB1_3_21/i0[9] ) );
  BUF_X1 \SB1_3_21/BUF_5  ( .A(\RI1[3][65] ), .Z(\SB1_3_21/i1_5 ) );
  INV_X1 \SB1_3_22/INV_3  ( .A(\RI1[3][57] ), .ZN(\SB1_3_22/i0[10] ) );
  INV_X1 \SB1_3_22/INV_2  ( .A(\RI1[3][56] ), .ZN(\SB1_3_22/i0_0 ) );
  INV_X1 \SB1_3_22/INV_1  ( .A(\RI1[3][55] ), .ZN(\SB1_3_22/i0[6] ) );
  INV_X1 \SB1_3_22/INV_0  ( .A(\RI1[3][54] ), .ZN(\SB1_3_22/i0[9] ) );
  BUF_X1 \SB1_3_22/BUF_5  ( .A(\RI1[3][59] ), .Z(\SB1_3_22/i1_5 ) );
  INV_X1 \SB1_3_23/INV_4  ( .A(\RI1[3][52] ), .ZN(\SB1_3_23/i0_4 ) );
  INV_X1 \SB1_3_23/INV_3  ( .A(\RI1[3][51] ), .ZN(\SB1_3_23/i0[10] ) );
  INV_X1 \SB1_3_23/INV_2  ( .A(\RI1[3][50] ), .ZN(\SB1_3_23/i0_0 ) );
  INV_X1 \SB1_3_23/INV_1  ( .A(\RI1[3][49] ), .ZN(\SB1_3_23/i0[6] ) );
  INV_X1 \SB1_3_24/INV_3  ( .A(\RI1[3][45] ), .ZN(\SB1_3_24/i0[10] ) );
  INV_X1 \SB1_3_24/INV_2  ( .A(\RI1[3][44] ), .ZN(\SB1_3_24/i0_0 ) );
  INV_X1 \SB1_3_24/INV_1  ( .A(\RI1[3][43] ), .ZN(\SB1_3_24/i0[6] ) );
  INV_X1 \SB1_3_24/INV_0  ( .A(\RI1[3][42] ), .ZN(\SB1_3_24/i0[9] ) );
  BUF_X1 \SB1_3_24/BUF_5  ( .A(\RI1[3][47] ), .Z(\SB1_3_24/i1_5 ) );
  INV_X1 \SB1_3_25/INV_3  ( .A(\RI1[3][39] ), .ZN(\SB1_3_25/i0[10] ) );
  INV_X1 \SB1_3_25/INV_1  ( .A(\RI1[3][37] ), .ZN(\SB1_3_25/i0[6] ) );
  INV_X1 \SB1_3_25/INV_0  ( .A(\RI1[3][36] ), .ZN(\SB1_3_25/i0[9] ) );
  BUF_X1 \SB1_3_25/BUF_5  ( .A(\RI1[3][41] ), .Z(\SB1_3_25/i1_5 ) );
  INV_X1 \SB1_3_26/INV_3  ( .A(\RI1[3][33] ), .ZN(\SB1_3_26/i0[10] ) );
  INV_X1 \SB1_3_26/INV_2  ( .A(\RI1[3][32] ), .ZN(\SB1_3_26/i0_0 ) );
  INV_X1 \SB1_3_26/INV_1  ( .A(\RI1[3][31] ), .ZN(\SB1_3_26/i0[6] ) );
  BUF_X1 \SB1_3_26/BUF_5  ( .A(\RI1[3][35] ), .Z(\SB1_3_26/i1_5 ) );
  INV_X1 \SB1_3_27/INV_4  ( .A(\RI1[3][28] ), .ZN(\SB1_3_27/i0_4 ) );
  INV_X1 \SB1_3_27/INV_3  ( .A(\RI1[3][27] ), .ZN(\SB1_3_27/i0[10] ) );
  INV_X1 \SB1_3_27/INV_2  ( .A(\RI1[3][26] ), .ZN(\SB1_3_27/i0_0 ) );
  INV_X1 \SB1_3_27/INV_1  ( .A(\RI1[3][25] ), .ZN(\SB1_3_27/i0[6] ) );
  INV_X1 \SB1_3_27/INV_0  ( .A(\RI1[3][24] ), .ZN(\SB1_3_27/i0[9] ) );
  BUF_X1 \SB1_3_27/BUF_5  ( .A(\RI1[3][29] ), .Z(\SB1_3_27/i1_5 ) );
  INV_X1 \SB1_3_28/INV_3  ( .A(\RI1[3][21] ), .ZN(\SB1_3_28/i0[10] ) );
  INV_X1 \SB1_3_28/INV_2  ( .A(\RI1[3][20] ), .ZN(\SB1_3_28/i0_0 ) );
  INV_X1 \SB1_3_28/INV_1  ( .A(\RI1[3][19] ), .ZN(\SB1_3_28/i0[6] ) );
  INV_X1 \SB1_3_28/INV_0  ( .A(\RI1[3][18] ), .ZN(\SB1_3_28/i0[9] ) );
  BUF_X1 \SB1_3_28/BUF_5  ( .A(\RI1[3][23] ), .Z(\SB1_3_28/i1_5 ) );
  INV_X1 \SB1_3_29/INV_3  ( .A(\RI1[3][15] ), .ZN(\SB1_3_29/i0[10] ) );
  INV_X1 \SB1_3_29/INV_2  ( .A(\RI1[3][14] ), .ZN(\SB1_3_29/i0_0 ) );
  INV_X1 \SB1_3_29/INV_1  ( .A(\RI1[3][13] ), .ZN(\SB1_3_29/i0[6] ) );
  INV_X1 \SB1_3_29/INV_0  ( .A(\RI1[3][12] ), .ZN(\SB1_3_29/i0[9] ) );
  BUF_X1 \SB1_3_29/BUF_5  ( .A(\RI1[3][17] ), .Z(\SB1_3_29/i1_5 ) );
  INV_X1 \SB1_3_30/INV_3  ( .A(\RI1[3][9] ), .ZN(\SB1_3_30/i0[10] ) );
  INV_X1 \SB1_3_30/INV_2  ( .A(\RI1[3][8] ), .ZN(\SB1_3_30/i0_0 ) );
  INV_X1 \SB1_3_30/INV_1  ( .A(\RI1[3][7] ), .ZN(\SB1_3_30/i0[6] ) );
  BUF_X1 \SB1_3_30/BUF_5  ( .A(\RI1[3][11] ), .Z(\SB1_3_30/i1_5 ) );
  INV_X1 \SB1_3_31/INV_3  ( .A(\RI1[3][3] ), .ZN(\SB1_3_31/i0[10] ) );
  INV_X1 \SB1_3_31/INV_2  ( .A(\RI1[3][2] ), .ZN(\SB1_3_31/i0_0 ) );
  INV_X1 \SB1_3_31/INV_1  ( .A(\RI1[3][1] ), .ZN(\SB1_3_31/i0[6] ) );
  INV_X1 \SB1_3_31/INV_0  ( .A(\RI1[3][0] ), .ZN(\SB1_3_31/i0[9] ) );
  BUF_X1 \SB1_3_31/BUF_5  ( .A(\RI1[3][5] ), .Z(\SB1_3_31/i1_5 ) );
  INV_X1 \SB3_0/INV_3  ( .A(\RI1[4][189] ), .ZN(\SB3_0/i0[10] ) );
  INV_X1 \SB3_0/INV_2  ( .A(\RI1[4][188] ), .ZN(\SB3_0/i0_0 ) );
  INV_X1 \SB3_0/INV_1  ( .A(\RI1[4][187] ), .ZN(\SB3_0/i0[6] ) );
  INV_X1 \SB3_0/INV_0  ( .A(\RI1[4][186] ), .ZN(\SB3_0/i0[9] ) );
  BUF_X1 \SB3_0/BUF_1  ( .A(\RI1[4][187] ), .Z(\SB3_0/i1_7 ) );
  INV_X1 \SB3_1/INV_4  ( .A(\RI1[4][184] ), .ZN(\SB3_1/i0_4 ) );
  INV_X1 \SB3_1/INV_3  ( .A(\RI1[4][183] ), .ZN(\SB3_1/i0[10] ) );
  INV_X1 \SB3_1/INV_2  ( .A(\RI1[4][182] ), .ZN(\SB3_1/i0_0 ) );
  INV_X1 \SB3_1/INV_1  ( .A(\RI1[4][181] ), .ZN(\SB3_1/i0[6] ) );
  INV_X1 \SB3_1/INV_0  ( .A(\RI1[4][180] ), .ZN(\SB3_1/i0[9] ) );
  BUF_X1 \SB3_1/BUF_5  ( .A(\RI1[4][185] ), .Z(\SB3_1/i1_5 ) );
  BUF_X1 \SB3_1/BUF_2  ( .A(\RI1[4][182] ), .Z(\SB3_1/i1[9] ) );
  BUF_X1 \SB3_1/BUF_1  ( .A(\RI1[4][181] ), .Z(\SB3_1/i1_7 ) );
  INV_X1 \SB3_2/INV_3  ( .A(\RI1[4][177] ), .ZN(\SB3_2/i0[10] ) );
  INV_X1 \SB3_2/INV_2  ( .A(\RI1[4][176] ), .ZN(\SB3_2/i0_0 ) );
  INV_X1 \SB3_2/INV_1  ( .A(\RI1[4][175] ), .ZN(\SB3_2/i0[6] ) );
  INV_X1 \SB3_2/INV_0  ( .A(\RI1[4][174] ), .ZN(\SB3_2/i0[9] ) );
  BUF_X1 \SB3_2/BUF_1  ( .A(\RI1[4][175] ), .Z(\SB3_2/i1_7 ) );
  BUF_X1 \SB3_2/BUF_0  ( .A(\RI1[4][174] ), .Z(\SB3_2/i3[0] ) );
  INV_X1 \SB3_3/INV_4  ( .A(\RI1[4][172] ), .ZN(\SB3_3/i0_4 ) );
  INV_X1 \SB3_3/INV_3  ( .A(\RI1[4][171] ), .ZN(\SB3_3/i0[10] ) );
  INV_X1 \SB3_3/INV_2  ( .A(\RI1[4][170] ), .ZN(\SB3_3/i0_0 ) );
  INV_X1 \SB3_3/INV_1  ( .A(\RI1[4][169] ), .ZN(\SB3_3/i0[6] ) );
  INV_X1 \SB3_3/INV_0  ( .A(\RI1[4][168] ), .ZN(\SB3_3/i0[9] ) );
  BUF_X1 \SB3_3/BUF_1  ( .A(\RI1[4][169] ), .Z(\SB3_3/i1_7 ) );
  INV_X1 \SB3_4/INV_4  ( .A(\RI1[4][166] ), .ZN(\SB3_4/i0_4 ) );
  INV_X1 \SB3_4/INV_3  ( .A(\RI1[4][165] ), .ZN(\SB3_4/i0[10] ) );
  INV_X1 \SB3_4/INV_2  ( .A(\RI1[4][164] ), .ZN(\SB3_4/i0_0 ) );
  INV_X1 \SB3_4/INV_1  ( .A(\RI1[4][163] ), .ZN(\SB3_4/i0[6] ) );
  INV_X1 \SB3_4/INV_0  ( .A(\RI1[4][162] ), .ZN(\SB3_4/i0[9] ) );
  BUF_X1 \SB3_4/BUF_5  ( .A(\RI1[4][167] ), .Z(\SB3_4/i1_5 ) );
  BUF_X1 \SB3_4/BUF_1  ( .A(\RI1[4][163] ), .Z(\SB3_4/i1_7 ) );
  INV_X1 \SB3_5/INV_3  ( .A(\RI1[4][159] ), .ZN(\SB3_5/i0[10] ) );
  INV_X1 \SB3_5/INV_2  ( .A(\RI1[4][158] ), .ZN(\SB3_5/i0_0 ) );
  INV_X1 \SB3_5/INV_1  ( .A(\RI1[4][157] ), .ZN(\SB3_5/i0[6] ) );
  INV_X1 \SB3_5/INV_0  ( .A(\RI1[4][156] ), .ZN(\SB3_5/i0[9] ) );
  BUF_X1 \SB3_5/BUF_1  ( .A(\RI1[4][157] ), .Z(\SB3_5/i1_7 ) );
  INV_X1 \SB3_6/INV_4  ( .A(\RI1[4][154] ), .ZN(\SB3_6/i0_4 ) );
  INV_X1 \SB3_6/INV_3  ( .A(\RI1[4][153] ), .ZN(\SB3_6/i0[10] ) );
  INV_X1 \SB3_6/INV_2  ( .A(\RI1[4][152] ), .ZN(\SB3_6/i0_0 ) );
  INV_X1 \SB3_6/INV_1  ( .A(\RI1[4][151] ), .ZN(\SB3_6/i0[6] ) );
  INV_X1 \SB3_6/INV_0  ( .A(\RI1[4][150] ), .ZN(\SB3_6/i0[9] ) );
  BUF_X1 \SB3_6/BUF_1  ( .A(\RI1[4][151] ), .Z(\SB3_6/i1_7 ) );
  INV_X1 \SB3_7/INV_4  ( .A(\RI1[4][148] ), .ZN(\SB3_7/i0_4 ) );
  INV_X1 \SB3_7/INV_3  ( .A(\RI1[4][147] ), .ZN(\SB3_7/i0[10] ) );
  INV_X1 \SB3_7/INV_2  ( .A(\RI1[4][146] ), .ZN(\SB3_7/i0_0 ) );
  INV_X1 \SB3_7/INV_1  ( .A(\RI1[4][145] ), .ZN(\SB3_7/i0[6] ) );
  INV_X1 \SB3_7/INV_0  ( .A(\RI1[4][144] ), .ZN(\SB3_7/i0[9] ) );
  BUF_X1 \SB3_7/BUF_1  ( .A(\RI1[4][145] ), .Z(\SB3_7/i1_7 ) );
  INV_X1 \SB3_8/INV_4  ( .A(\RI1[4][142] ), .ZN(\SB3_8/i0_4 ) );
  INV_X1 \SB3_8/INV_3  ( .A(\RI1[4][141] ), .ZN(\SB3_8/i0[10] ) );
  INV_X1 \SB3_8/INV_2  ( .A(\RI1[4][140] ), .ZN(\SB3_8/i0_0 ) );
  INV_X1 \SB3_8/INV_1  ( .A(\RI1[4][139] ), .ZN(\SB3_8/i0[6] ) );
  INV_X1 \SB3_8/INV_0  ( .A(\RI1[4][138] ), .ZN(\SB3_8/i0[9] ) );
  BUF_X1 \SB3_8/BUF_1  ( .A(\RI1[4][139] ), .Z(\SB3_8/i1_7 ) );
  INV_X1 \SB3_9/INV_4  ( .A(\RI1[4][136] ), .ZN(\SB3_9/i0_4 ) );
  INV_X1 \SB3_9/INV_3  ( .A(\RI1[4][135] ), .ZN(\SB3_9/i0[10] ) );
  INV_X1 \SB3_9/INV_2  ( .A(\RI1[4][134] ), .ZN(\SB3_9/i0_0 ) );
  INV_X1 \SB3_9/INV_1  ( .A(\RI1[4][133] ), .ZN(\SB3_9/i0[6] ) );
  INV_X1 \SB3_9/INV_0  ( .A(\RI1[4][132] ), .ZN(\SB3_9/i0[9] ) );
  BUF_X1 \SB3_9/BUF_1  ( .A(\RI1[4][133] ), .Z(\SB3_9/i1_7 ) );
  INV_X1 \SB3_10/INV_4  ( .A(\RI1[4][130] ), .ZN(\SB3_10/i0_4 ) );
  INV_X1 \SB3_10/INV_3  ( .A(\RI1[4][129] ), .ZN(\SB3_10/i0[10] ) );
  INV_X1 \SB3_10/INV_2  ( .A(\RI1[4][128] ), .ZN(\SB3_10/i0_0 ) );
  INV_X1 \SB3_10/INV_1  ( .A(\RI1[4][127] ), .ZN(\SB3_10/i0[6] ) );
  INV_X1 \SB3_10/INV_0  ( .A(\RI1[4][126] ), .ZN(\SB3_10/i0[9] ) );
  BUF_X1 \SB3_10/BUF_5  ( .A(\RI1[4][131] ), .Z(\SB3_10/i1_5 ) );
  BUF_X1 \SB3_10/BUF_4  ( .A(\RI1[4][130] ), .Z(\SB3_10/i0[7] ) );
  BUF_X1 \SB3_10/BUF_1  ( .A(\RI1[4][127] ), .Z(\SB3_10/i1_7 ) );
  INV_X1 \SB3_11/INV_3  ( .A(\RI1[4][123] ), .ZN(\SB3_11/i0[10] ) );
  INV_X1 \SB3_11/INV_2  ( .A(\RI1[4][122] ), .ZN(\SB3_11/i0_0 ) );
  INV_X1 \SB3_11/INV_1  ( .A(\RI1[4][121] ), .ZN(\SB3_11/i0[6] ) );
  INV_X1 \SB3_11/INV_0  ( .A(\RI1[4][120] ), .ZN(\SB3_11/i0[9] ) );
  BUF_X1 \SB3_11/BUF_5  ( .A(\RI1[4][125] ), .Z(\SB3_11/i1_5 ) );
  BUF_X1 \SB3_11/BUF_1  ( .A(\RI1[4][121] ), .Z(\SB3_11/i1_7 ) );
  INV_X1 \SB3_12/INV_4  ( .A(\RI1[4][118] ), .ZN(\SB3_12/i0_4 ) );
  INV_X1 \SB3_12/INV_3  ( .A(\RI1[4][117] ), .ZN(\SB3_12/i0[10] ) );
  INV_X1 \SB3_12/INV_2  ( .A(\RI1[4][116] ), .ZN(\SB3_12/i0_0 ) );
  INV_X1 \SB3_12/INV_1  ( .A(\RI1[4][115] ), .ZN(\SB3_12/i0[6] ) );
  INV_X1 \SB3_12/INV_0  ( .A(\RI1[4][114] ), .ZN(\SB3_12/i0[9] ) );
  BUF_X1 \SB3_12/BUF_1  ( .A(\RI1[4][115] ), .Z(\SB3_12/i1_7 ) );
  INV_X1 \SB3_13/INV_4  ( .A(\RI1[4][112] ), .ZN(\SB3_13/i0_4 ) );
  INV_X1 \SB3_13/INV_3  ( .A(\RI1[4][111] ), .ZN(\SB3_13/i0[10] ) );
  INV_X1 \SB3_13/INV_2  ( .A(\RI1[4][110] ), .ZN(\SB3_13/i0_0 ) );
  INV_X1 \SB3_13/INV_1  ( .A(\RI1[4][109] ), .ZN(\SB3_13/i0[6] ) );
  INV_X1 \SB3_13/INV_0  ( .A(\RI1[4][108] ), .ZN(\SB3_13/i0[9] ) );
  BUF_X1 \SB3_13/BUF_1  ( .A(\RI1[4][109] ), .Z(\SB3_13/i1_7 ) );
  INV_X1 \SB3_14/INV_4  ( .A(\RI1[4][106] ), .ZN(\SB3_14/i0_4 ) );
  INV_X1 \SB3_14/INV_3  ( .A(\RI1[4][105] ), .ZN(\SB3_14/i0[10] ) );
  INV_X1 \SB3_14/INV_2  ( .A(\RI1[4][104] ), .ZN(\SB3_14/i0_0 ) );
  INV_X1 \SB3_14/INV_1  ( .A(\RI1[4][103] ), .ZN(\SB3_14/i0[6] ) );
  INV_X1 \SB3_14/INV_0  ( .A(\RI1[4][102] ), .ZN(\SB3_14/i0[9] ) );
  BUF_X1 \SB3_14/BUF_5  ( .A(\RI1[4][107] ), .Z(\SB3_14/i1_5 ) );
  BUF_X1 \SB3_14/BUF_1  ( .A(\RI1[4][103] ), .Z(\SB3_14/i1_7 ) );
  INV_X1 \SB3_15/INV_4  ( .A(\RI1[4][100] ), .ZN(\SB3_15/i0_4 ) );
  INV_X1 \SB3_15/INV_3  ( .A(\RI1[4][99] ), .ZN(\SB3_15/i0[10] ) );
  INV_X1 \SB3_15/INV_2  ( .A(\RI1[4][98] ), .ZN(\SB3_15/i0_0 ) );
  INV_X1 \SB3_15/INV_1  ( .A(\RI1[4][97] ), .ZN(\SB3_15/i0[6] ) );
  INV_X1 \SB3_15/INV_0  ( .A(\RI1[4][96] ), .ZN(\SB3_15/i0[9] ) );
  BUF_X1 \SB3_15/BUF_1  ( .A(\RI1[4][97] ), .Z(\SB3_15/i1_7 ) );
  INV_X1 \SB3_16/INV_4  ( .A(\RI1[4][94] ), .ZN(\SB3_16/i0_4 ) );
  INV_X1 \SB3_16/INV_3  ( .A(\RI1[4][93] ), .ZN(\SB3_16/i0[10] ) );
  INV_X1 \SB3_16/INV_2  ( .A(\RI1[4][92] ), .ZN(\SB3_16/i0_0 ) );
  INV_X1 \SB3_16/INV_1  ( .A(\RI1[4][91] ), .ZN(\SB3_16/i0[6] ) );
  INV_X1 \SB3_16/INV_0  ( .A(\RI1[4][90] ), .ZN(\SB3_16/i0[9] ) );
  BUF_X1 \SB3_16/BUF_5  ( .A(\RI1[4][95] ), .Z(\SB3_16/i1_5 ) );
  BUF_X1 \SB3_16/BUF_1  ( .A(\RI1[4][91] ), .Z(\SB3_16/i1_7 ) );
  INV_X1 \SB3_17/INV_3  ( .A(\RI1[4][87] ), .ZN(\SB3_17/i0[10] ) );
  INV_X1 \SB3_17/INV_2  ( .A(\RI1[4][86] ), .ZN(\SB3_17/i0_0 ) );
  INV_X1 \SB3_17/INV_1  ( .A(\RI1[4][85] ), .ZN(\SB3_17/i0[6] ) );
  INV_X1 \SB3_17/INV_0  ( .A(\RI1[4][84] ), .ZN(\SB3_17/i0[9] ) );
  BUF_X1 \SB3_17/BUF_5  ( .A(\RI1[4][89] ), .Z(\SB3_17/i1_5 ) );
  BUF_X1 \SB3_17/BUF_1  ( .A(\RI1[4][85] ), .Z(\SB3_17/i1_7 ) );
  INV_X1 \SB3_18/INV_4  ( .A(\RI1[4][82] ), .ZN(\SB3_18/i0_4 ) );
  INV_X1 \SB3_18/INV_3  ( .A(\RI1[4][81] ), .ZN(\SB3_18/i0[10] ) );
  INV_X1 \SB3_18/INV_2  ( .A(\RI1[4][80] ), .ZN(\SB3_18/i0_0 ) );
  INV_X1 \SB3_18/INV_1  ( .A(\RI1[4][79] ), .ZN(\SB3_18/i0[6] ) );
  INV_X1 \SB3_18/INV_0  ( .A(\RI1[4][78] ), .ZN(\SB3_18/i0[9] ) );
  BUF_X1 \SB3_18/BUF_5  ( .A(\RI1[4][83] ), .Z(\SB3_18/i1_5 ) );
  BUF_X1 \SB3_18/BUF_1  ( .A(\RI1[4][79] ), .Z(\SB3_18/i1_7 ) );
  INV_X1 \SB3_19/INV_3  ( .A(\RI1[4][75] ), .ZN(\SB3_19/i0[10] ) );
  INV_X1 \SB3_19/INV_2  ( .A(\RI1[4][74] ), .ZN(\SB3_19/i0_0 ) );
  INV_X1 \SB3_19/INV_1  ( .A(\RI1[4][73] ), .ZN(\SB3_19/i0[6] ) );
  INV_X1 \SB3_19/INV_0  ( .A(\RI1[4][72] ), .ZN(\SB3_19/i0[9] ) );
  BUF_X1 \SB3_19/BUF_1  ( .A(\RI1[4][73] ), .Z(\SB3_19/i1_7 ) );
  BUF_X1 \SB3_19/BUF_0  ( .A(\RI1[4][72] ), .Z(\SB3_19/i3[0] ) );
  INV_X1 \SB3_20/INV_3  ( .A(\RI1[4][69] ), .ZN(\SB3_20/i0[10] ) );
  INV_X1 \SB3_20/INV_2  ( .A(\RI1[4][68] ), .ZN(\SB3_20/i0_0 ) );
  INV_X1 \SB3_20/INV_1  ( .A(\RI1[4][67] ), .ZN(\SB3_20/i0[6] ) );
  INV_X1 \SB3_20/INV_0  ( .A(\RI1[4][66] ), .ZN(\SB3_20/i0[9] ) );
  BUF_X1 \SB3_20/BUF_5  ( .A(\RI1[4][71] ), .Z(\SB3_20/i1_5 ) );
  BUF_X1 \SB3_20/BUF_3  ( .A(\RI1[4][69] ), .Z(\SB3_20/i0[8] ) );
  BUF_X1 \SB3_20/BUF_1  ( .A(\RI1[4][67] ), .Z(\SB3_20/i1_7 ) );
  INV_X1 \SB3_21/INV_4  ( .A(\RI1[4][64] ), .ZN(\SB3_21/i0_4 ) );
  INV_X1 \SB3_21/INV_3  ( .A(\RI1[4][63] ), .ZN(\SB3_21/i0[10] ) );
  INV_X1 \SB3_21/INV_2  ( .A(\RI1[4][62] ), .ZN(\SB3_21/i0_0 ) );
  INV_X1 \SB3_21/INV_1  ( .A(\RI1[4][61] ), .ZN(\SB3_21/i0[6] ) );
  INV_X1 \SB3_21/INV_0  ( .A(\RI1[4][60] ), .ZN(\SB3_21/i0[9] ) );
  BUF_X1 \SB3_21/BUF_5  ( .A(\RI1[4][65] ), .Z(\SB3_21/i1_5 ) );
  BUF_X1 \SB3_21/BUF_1  ( .A(\RI1[4][61] ), .Z(\SB3_21/i1_7 ) );
  INV_X1 \SB3_22/INV_4  ( .A(\RI1[4][58] ), .ZN(\SB3_22/i0_4 ) );
  INV_X1 \SB3_22/INV_3  ( .A(\RI1[4][57] ), .ZN(\SB3_22/i0[10] ) );
  INV_X1 \SB3_22/INV_2  ( .A(\RI1[4][56] ), .ZN(\SB3_22/i0_0 ) );
  INV_X1 \SB3_22/INV_1  ( .A(\RI1[4][55] ), .ZN(\SB3_22/i0[6] ) );
  INV_X1 \SB3_22/INV_0  ( .A(\RI1[4][54] ), .ZN(\SB3_22/i0[9] ) );
  BUF_X1 \SB3_22/BUF_1  ( .A(\RI1[4][55] ), .Z(\SB3_22/i1_7 ) );
  INV_X1 \SB3_23/INV_4  ( .A(\RI1[4][52] ), .ZN(\SB3_23/i0_4 ) );
  INV_X1 \SB3_23/INV_3  ( .A(\RI1[4][51] ), .ZN(\SB3_23/i0[10] ) );
  INV_X1 \SB3_23/INV_2  ( .A(\RI1[4][50] ), .ZN(\SB3_23/i0_0 ) );
  INV_X1 \SB3_23/INV_1  ( .A(\RI1[4][49] ), .ZN(\SB3_23/i0[6] ) );
  INV_X1 \SB3_23/INV_0  ( .A(\RI1[4][48] ), .ZN(\SB3_23/i0[9] ) );
  BUF_X1 \SB3_23/BUF_5  ( .A(\RI1[4][53] ), .Z(\SB3_23/i1_5 ) );
  BUF_X1 \SB3_23/BUF_1  ( .A(\RI1[4][49] ), .Z(\SB3_23/i1_7 ) );
  INV_X1 \SB3_24/INV_4  ( .A(\RI1[4][46] ), .ZN(\SB3_24/i0_4 ) );
  INV_X1 \SB3_24/INV_3  ( .A(\RI1[4][45] ), .ZN(\SB3_24/i0[10] ) );
  INV_X1 \SB3_24/INV_2  ( .A(\RI1[4][44] ), .ZN(\SB3_24/i0_0 ) );
  INV_X1 \SB3_24/INV_1  ( .A(\RI1[4][43] ), .ZN(\SB3_24/i0[6] ) );
  INV_X1 \SB3_24/INV_0  ( .A(\RI1[4][42] ), .ZN(\SB3_24/i0[9] ) );
  BUF_X1 \SB3_24/BUF_5  ( .A(\RI1[4][47] ), .Z(\SB3_24/i1_5 ) );
  BUF_X1 \SB3_24/BUF_1  ( .A(\RI1[4][43] ), .Z(\SB3_24/i1_7 ) );
  INV_X1 \SB3_25/INV_4  ( .A(\RI1[4][40] ), .ZN(\SB3_25/i0_4 ) );
  INV_X1 \SB3_25/INV_3  ( .A(\RI1[4][39] ), .ZN(\SB3_25/i0[10] ) );
  INV_X1 \SB3_25/INV_2  ( .A(\RI1[4][38] ), .ZN(\SB3_25/i0_0 ) );
  INV_X1 \SB3_25/INV_1  ( .A(\RI1[4][37] ), .ZN(\SB3_25/i0[6] ) );
  INV_X1 \SB3_25/INV_0  ( .A(\RI1[4][36] ), .ZN(\SB3_25/i0[9] ) );
  BUF_X1 \SB3_25/BUF_5  ( .A(\RI1[4][41] ), .Z(\SB3_25/i1_5 ) );
  BUF_X1 \SB3_25/BUF_3  ( .A(\RI1[4][39] ), .Z(\SB3_25/i0[8] ) );
  BUF_X1 \SB3_25/BUF_1  ( .A(\RI1[4][37] ), .Z(\SB3_25/i1_7 ) );
  INV_X1 \SB3_26/INV_4  ( .A(\RI1[4][34] ), .ZN(\SB3_26/i0_4 ) );
  INV_X1 \SB3_26/INV_3  ( .A(\RI1[4][33] ), .ZN(\SB3_26/i0[10] ) );
  INV_X1 \SB3_26/INV_2  ( .A(\RI1[4][32] ), .ZN(\SB3_26/i0_0 ) );
  INV_X1 \SB3_26/INV_1  ( .A(\RI1[4][31] ), .ZN(\SB3_26/i0[6] ) );
  INV_X1 \SB3_26/INV_0  ( .A(\RI1[4][30] ), .ZN(\SB3_26/i0[9] ) );
  BUF_X1 \SB3_26/BUF_1  ( .A(\RI1[4][31] ), .Z(\SB3_26/i1_7 ) );
  INV_X1 \SB3_27/INV_4  ( .A(\RI1[4][28] ), .ZN(\SB3_27/i0_4 ) );
  INV_X1 \SB3_27/INV_3  ( .A(\RI1[4][27] ), .ZN(\SB3_27/i0[10] ) );
  INV_X1 \SB3_27/INV_2  ( .A(\RI1[4][26] ), .ZN(\SB3_27/i0_0 ) );
  INV_X1 \SB3_27/INV_1  ( .A(\RI1[4][25] ), .ZN(\SB3_27/i0[6] ) );
  INV_X1 \SB3_27/INV_0  ( .A(\RI1[4][24] ), .ZN(\SB3_27/i0[9] ) );
  BUF_X1 \SB3_27/BUF_5  ( .A(\RI1[4][29] ), .Z(\SB3_27/i1_5 ) );
  BUF_X1 \SB3_27/BUF_1  ( .A(\RI1[4][25] ), .Z(\SB3_27/i1_7 ) );
  INV_X1 \SB3_28/INV_4  ( .A(\RI1[4][22] ), .ZN(\SB3_28/i0_4 ) );
  INV_X1 \SB3_28/INV_3  ( .A(\RI1[4][21] ), .ZN(\SB3_28/i0[10] ) );
  INV_X1 \SB3_28/INV_2  ( .A(\RI1[4][20] ), .ZN(\SB3_28/i0_0 ) );
  INV_X1 \SB3_28/INV_1  ( .A(\RI1[4][19] ), .ZN(\SB3_28/i0[6] ) );
  INV_X1 \SB3_28/INV_0  ( .A(\RI1[4][18] ), .ZN(\SB3_28/i0[9] ) );
  BUF_X1 \SB3_28/BUF_5  ( .A(\RI1[4][23] ), .Z(\SB3_28/i1_5 ) );
  BUF_X1 \SB3_28/BUF_2  ( .A(\RI1[4][20] ), .Z(\SB3_28/i1[9] ) );
  BUF_X1 \SB3_28/BUF_1  ( .A(\RI1[4][19] ), .Z(\SB3_28/i1_7 ) );
  INV_X1 \SB3_29/INV_3  ( .A(\RI1[4][15] ), .ZN(\SB3_29/i0[10] ) );
  INV_X1 \SB3_29/INV_2  ( .A(\RI1[4][14] ), .ZN(\SB3_29/i0_0 ) );
  INV_X1 \SB3_29/INV_1  ( .A(\RI1[4][13] ), .ZN(\SB3_29/i0[6] ) );
  INV_X1 \SB3_29/INV_0  ( .A(\RI1[4][12] ), .ZN(\SB3_29/i0[9] ) );
  BUF_X1 \SB3_29/BUF_5  ( .A(\RI1[4][17] ), .Z(\SB3_29/i1_5 ) );
  BUF_X1 \SB3_29/BUF_4  ( .A(\RI1[4][16] ), .Z(\SB3_29/i0[7] ) );
  BUF_X1 \SB3_29/BUF_1  ( .A(\RI1[4][13] ), .Z(\SB3_29/i1_7 ) );
  INV_X1 \SB3_30/INV_4  ( .A(\RI1[4][10] ), .ZN(\SB3_30/i0_4 ) );
  INV_X1 \SB3_30/INV_3  ( .A(\RI1[4][9] ), .ZN(\SB3_30/i0[10] ) );
  INV_X1 \SB3_30/INV_2  ( .A(\RI1[4][8] ), .ZN(\SB3_30/i0_0 ) );
  INV_X1 \SB3_30/INV_1  ( .A(\RI1[4][7] ), .ZN(\SB3_30/i0[6] ) );
  INV_X1 \SB3_30/INV_0  ( .A(\RI1[4][6] ), .ZN(\SB3_30/i0[9] ) );
  BUF_X1 \SB3_30/BUF_1  ( .A(\RI1[4][7] ), .Z(\SB3_30/i1_7 ) );
  INV_X1 \SB3_31/INV_4  ( .A(\RI1[4][4] ), .ZN(\SB3_31/i0_4 ) );
  INV_X1 \SB3_31/INV_3  ( .A(\RI1[4][3] ), .ZN(\SB3_31/i0[10] ) );
  INV_X1 \SB3_31/INV_2  ( .A(\RI1[4][2] ), .ZN(\SB3_31/i0_0 ) );
  INV_X1 \SB3_31/INV_1  ( .A(\RI1[4][1] ), .ZN(\SB3_31/i0[6] ) );
  INV_X1 \SB3_31/INV_0  ( .A(\RI1[4][0] ), .ZN(\SB3_31/i0[9] ) );
  BUF_X1 \SB3_31/BUF_5  ( .A(\RI1[4][5] ), .Z(\SB3_31/i1_5 ) );
  BUF_X1 \SB3_31/BUF_1  ( .A(\RI1[4][1] ), .Z(\SB3_31/i1_7 ) );
  INV_X1 \SB2_0_0/INV_5  ( .A(\RI3[0][191] ), .ZN(\SB2_0_0/i1_5 ) );
  INV_X1 \SB2_0_0/INV_4  ( .A(\RI3[0][190] ), .ZN(\SB2_0_0/i0[7] ) );
  INV_X1 \SB2_0_0/INV_3  ( .A(\RI3[0][189] ), .ZN(\SB2_0_0/i0[8] ) );
  INV_X1 \SB2_0_0/INV_2  ( .A(\RI3[0][188] ), .ZN(\SB2_0_0/i1[9] ) );
  INV_X1 \SB2_0_0/INV_1  ( .A(\RI3[0][187] ), .ZN(\SB2_0_0/i1_7 ) );
  INV_X1 \SB2_0_0/INV_0  ( .A(\RI3[0][186] ), .ZN(\SB2_0_0/i3[0] ) );
  INV_X1 \SB2_0_1/INV_5  ( .A(\RI3[0][185] ), .ZN(\SB2_0_1/i1_5 ) );
  INV_X1 \SB2_0_1/INV_4  ( .A(\RI3[0][184] ), .ZN(\SB2_0_1/i0[7] ) );
  INV_X1 \SB2_0_1/INV_3  ( .A(\RI3[0][183] ), .ZN(\SB2_0_1/i0[8] ) );
  INV_X1 \SB2_0_1/INV_1  ( .A(\RI3[0][181] ), .ZN(\SB2_0_1/i1_7 ) );
  INV_X1 \SB2_0_1/INV_0  ( .A(\RI3[0][180] ), .ZN(\SB2_0_1/i3[0] ) );
  INV_X1 \SB2_0_2/INV_5  ( .A(\RI3[0][179] ), .ZN(\SB2_0_2/i1_5 ) );
  INV_X1 \SB2_0_2/INV_4  ( .A(\RI3[0][178] ), .ZN(\SB2_0_2/i0[7] ) );
  INV_X1 \SB2_0_2/INV_3  ( .A(\RI3[0][177] ), .ZN(\SB2_0_2/i0[8] ) );
  INV_X1 \SB2_0_2/INV_2  ( .A(\RI3[0][176] ), .ZN(\SB2_0_2/i1[9] ) );
  INV_X1 \SB2_0_2/INV_1  ( .A(\RI3[0][175] ), .ZN(\SB2_0_2/i1_7 ) );
  INV_X1 \SB2_0_2/INV_0  ( .A(\RI3[0][174] ), .ZN(\SB2_0_2/i3[0] ) );
  INV_X1 \SB2_0_3/INV_5  ( .A(\RI3[0][173] ), .ZN(\SB2_0_3/i1_5 ) );
  INV_X1 \SB2_0_3/INV_4  ( .A(\SB2_0_3/i0_4 ), .ZN(\SB2_0_3/i0[7] ) );
  INV_X1 \SB2_0_3/INV_3  ( .A(\RI3[0][171] ), .ZN(\SB2_0_3/i0[8] ) );
  INV_X1 \SB2_0_3/INV_2  ( .A(\RI3[0][170] ), .ZN(\SB2_0_3/i1[9] ) );
  INV_X1 \SB2_0_3/INV_1  ( .A(\RI3[0][169] ), .ZN(\SB2_0_3/i1_7 ) );
  INV_X1 \SB2_0_3/INV_0  ( .A(\RI3[0][168] ), .ZN(\SB2_0_3/i3[0] ) );
  INV_X1 \SB2_0_4/INV_5  ( .A(\RI3[0][167] ), .ZN(\SB2_0_4/i1_5 ) );
  INV_X1 \SB2_0_4/INV_4  ( .A(\RI3[0][166] ), .ZN(\SB2_0_4/i0[7] ) );
  INV_X1 \SB2_0_4/INV_3  ( .A(\RI3[0][165] ), .ZN(\SB2_0_4/i0[8] ) );
  INV_X1 \SB2_0_4/INV_2  ( .A(\RI3[0][164] ), .ZN(\SB2_0_4/i1[9] ) );
  INV_X1 \SB2_0_4/INV_1  ( .A(\RI3[0][163] ), .ZN(\SB2_0_4/i1_7 ) );
  INV_X1 \SB2_0_4/INV_0  ( .A(\RI3[0][162] ), .ZN(\SB2_0_4/i3[0] ) );
  INV_X1 \SB2_0_5/INV_5  ( .A(\RI3[0][161] ), .ZN(\SB2_0_5/i1_5 ) );
  INV_X1 \SB2_0_5/INV_4  ( .A(\RI3[0][160] ), .ZN(\SB2_0_5/i0[7] ) );
  INV_X1 \SB2_0_5/INV_3  ( .A(\RI3[0][159] ), .ZN(\SB2_0_5/i0[8] ) );
  INV_X1 \SB2_0_5/INV_2  ( .A(\RI3[0][158] ), .ZN(\SB2_0_5/i1[9] ) );
  INV_X1 \SB2_0_5/INV_1  ( .A(\RI3[0][157] ), .ZN(\SB2_0_5/i1_7 ) );
  INV_X1 \SB2_0_5/INV_0  ( .A(\RI3[0][156] ), .ZN(\SB2_0_5/i3[0] ) );
  INV_X1 \SB2_0_6/INV_5  ( .A(\RI3[0][155] ), .ZN(\SB2_0_6/i1_5 ) );
  INV_X1 \SB2_0_6/INV_4  ( .A(\RI3[0][154] ), .ZN(\SB2_0_6/i0[7] ) );
  INV_X1 \SB2_0_6/INV_3  ( .A(\RI3[0][153] ), .ZN(\SB2_0_6/i0[8] ) );
  INV_X1 \SB2_0_6/INV_2  ( .A(\RI3[0][152] ), .ZN(\SB2_0_6/i1[9] ) );
  INV_X1 \SB2_0_6/INV_1  ( .A(\RI3[0][151] ), .ZN(\SB2_0_6/i1_7 ) );
  INV_X1 \SB2_0_6/INV_0  ( .A(\RI3[0][150] ), .ZN(\SB2_0_6/i3[0] ) );
  INV_X1 \SB2_0_7/INV_5  ( .A(\RI3[0][149] ), .ZN(\SB2_0_7/i1_5 ) );
  INV_X1 \SB2_0_7/INV_4  ( .A(\RI3[0][148] ), .ZN(\SB2_0_7/i0[7] ) );
  INV_X1 \SB2_0_7/INV_3  ( .A(\RI3[0][147] ), .ZN(\SB2_0_7/i0[8] ) );
  INV_X1 \SB2_0_7/INV_2  ( .A(\RI3[0][146] ), .ZN(\SB2_0_7/i1[9] ) );
  INV_X1 \SB2_0_7/INV_1  ( .A(\RI3[0][145] ), .ZN(\SB2_0_7/i1_7 ) );
  INV_X1 \SB2_0_7/INV_0  ( .A(\RI3[0][144] ), .ZN(\SB2_0_7/i3[0] ) );
  INV_X1 \SB2_0_8/INV_5  ( .A(\RI3[0][143] ), .ZN(\SB2_0_8/i1_5 ) );
  INV_X1 \SB2_0_8/INV_4  ( .A(\RI3[0][142] ), .ZN(\SB2_0_8/i0[7] ) );
  INV_X1 \SB2_0_8/INV_3  ( .A(\RI3[0][141] ), .ZN(\SB2_0_8/i0[8] ) );
  INV_X1 \SB2_0_8/INV_1  ( .A(\RI3[0][139] ), .ZN(\SB2_0_8/i1_7 ) );
  INV_X1 \SB2_0_8/INV_0  ( .A(\RI3[0][138] ), .ZN(\SB2_0_8/i3[0] ) );
  INV_X1 \SB2_0_9/INV_5  ( .A(\RI3[0][137] ), .ZN(\SB2_0_9/i1_5 ) );
  INV_X1 \SB2_0_9/INV_4  ( .A(\RI3[0][136] ), .ZN(\SB2_0_9/i0[7] ) );
  INV_X1 \SB2_0_9/INV_3  ( .A(\RI3[0][135] ), .ZN(\SB2_0_9/i0[8] ) );
  INV_X1 \SB2_0_9/INV_2  ( .A(\RI3[0][134] ), .ZN(\SB2_0_9/i1[9] ) );
  INV_X1 \SB2_0_9/INV_1  ( .A(\RI3[0][133] ), .ZN(\SB2_0_9/i1_7 ) );
  INV_X1 \SB2_0_9/INV_0  ( .A(\RI3[0][132] ), .ZN(\SB2_0_9/i3[0] ) );
  INV_X1 \SB2_0_10/INV_5  ( .A(\RI3[0][131] ), .ZN(\SB2_0_10/i1_5 ) );
  INV_X1 \SB2_0_10/INV_4  ( .A(\RI3[0][130] ), .ZN(\SB2_0_10/i0[7] ) );
  INV_X1 \SB2_0_10/INV_3  ( .A(\RI3[0][129] ), .ZN(\SB2_0_10/i0[8] ) );
  INV_X1 \SB2_0_10/INV_1  ( .A(\RI3[0][127] ), .ZN(\SB2_0_10/i1_7 ) );
  INV_X1 \SB2_0_10/INV_0  ( .A(\RI3[0][126] ), .ZN(\SB2_0_10/i3[0] ) );
  INV_X1 \SB2_0_11/INV_5  ( .A(\RI3[0][125] ), .ZN(\SB2_0_11/i1_5 ) );
  INV_X1 \SB2_0_11/INV_4  ( .A(\RI3[0][124] ), .ZN(\SB2_0_11/i0[7] ) );
  INV_X1 \SB2_0_11/INV_3  ( .A(\RI3[0][123] ), .ZN(\SB2_0_11/i0[8] ) );
  INV_X1 \SB2_0_11/INV_2  ( .A(\RI3[0][122] ), .ZN(\SB2_0_11/i1[9] ) );
  INV_X1 \SB2_0_11/INV_1  ( .A(\RI3[0][121] ), .ZN(\SB2_0_11/i1_7 ) );
  INV_X1 \SB2_0_11/INV_0  ( .A(\RI3[0][120] ), .ZN(\SB2_0_11/i3[0] ) );
  BUF_X1 \SB2_0_11/BUF_1  ( .A(\RI3[0][121] ), .Z(\SB2_0_11/i0[6] ) );
  INV_X1 \SB2_0_12/INV_5  ( .A(\RI3[0][119] ), .ZN(\SB2_0_12/i1_5 ) );
  INV_X1 \SB2_0_12/INV_4  ( .A(\RI3[0][118] ), .ZN(\SB2_0_12/i0[7] ) );
  INV_X1 \SB2_0_12/INV_3  ( .A(\RI3[0][117] ), .ZN(\SB2_0_12/i0[8] ) );
  INV_X1 \SB2_0_12/INV_1  ( .A(\RI3[0][115] ), .ZN(\SB2_0_12/i1_7 ) );
  INV_X1 \SB2_0_12/INV_0  ( .A(\RI3[0][114] ), .ZN(\SB2_0_12/i3[0] ) );
  BUF_X1 \SB2_0_12/BUF_0  ( .A(\RI3[0][114] ), .Z(\SB2_0_12/i0[9] ) );
  INV_X1 \SB2_0_13/INV_5  ( .A(\RI3[0][113] ), .ZN(\SB2_0_13/i1_5 ) );
  INV_X1 \SB2_0_13/INV_4  ( .A(\RI3[0][112] ), .ZN(\SB2_0_13/i0[7] ) );
  INV_X1 \SB2_0_13/INV_3  ( .A(\RI3[0][111] ), .ZN(\SB2_0_13/i0[8] ) );
  INV_X1 \SB2_0_13/INV_1  ( .A(\RI3[0][109] ), .ZN(\SB2_0_13/i1_7 ) );
  INV_X1 \SB2_0_13/INV_0  ( .A(\RI3[0][108] ), .ZN(\SB2_0_13/i3[0] ) );
  INV_X1 \SB2_0_14/INV_5  ( .A(\RI3[0][107] ), .ZN(\SB2_0_14/i1_5 ) );
  INV_X1 \SB2_0_14/INV_4  ( .A(\RI3[0][106] ), .ZN(\SB2_0_14/i0[7] ) );
  INV_X1 \SB2_0_14/INV_3  ( .A(\RI3[0][105] ), .ZN(\SB2_0_14/i0[8] ) );
  INV_X1 \SB2_0_14/INV_2  ( .A(\RI3[0][104] ), .ZN(\SB2_0_14/i1[9] ) );
  INV_X1 \SB2_0_14/INV_1  ( .A(\RI3[0][103] ), .ZN(\SB2_0_14/i1_7 ) );
  INV_X1 \SB2_0_14/INV_0  ( .A(\RI3[0][102] ), .ZN(\SB2_0_14/i3[0] ) );
  INV_X1 \SB2_0_15/INV_5  ( .A(\RI3[0][101] ), .ZN(\SB2_0_15/i1_5 ) );
  INV_X1 \SB2_0_15/INV_4  ( .A(\SB2_0_15/i0_4 ), .ZN(\SB2_0_15/i0[7] ) );
  INV_X1 \SB2_0_15/INV_3  ( .A(\RI3[0][99] ), .ZN(\SB2_0_15/i0[8] ) );
  INV_X1 \SB2_0_15/INV_2  ( .A(\RI3[0][98] ), .ZN(\SB2_0_15/i1[9] ) );
  INV_X1 \SB2_0_15/INV_1  ( .A(\RI3[0][97] ), .ZN(\SB2_0_15/i1_7 ) );
  INV_X1 \SB2_0_15/INV_0  ( .A(\RI3[0][96] ), .ZN(\SB2_0_15/i3[0] ) );
  INV_X1 \SB2_0_16/INV_5  ( .A(\RI3[0][95] ), .ZN(\SB2_0_16/i1_5 ) );
  INV_X1 \SB2_0_16/INV_4  ( .A(\RI3[0][94] ), .ZN(\SB2_0_16/i0[7] ) );
  INV_X1 \SB2_0_16/INV_3  ( .A(\RI3[0][93] ), .ZN(\SB2_0_16/i0[8] ) );
  INV_X1 \SB2_0_16/INV_2  ( .A(\RI3[0][92] ), .ZN(\SB2_0_16/i1[9] ) );
  INV_X1 \SB2_0_16/INV_1  ( .A(\RI3[0][91] ), .ZN(\SB2_0_16/i1_7 ) );
  INV_X1 \SB2_0_16/INV_0  ( .A(\RI3[0][90] ), .ZN(\SB2_0_16/i3[0] ) );
  INV_X1 \SB2_0_17/INV_5  ( .A(\RI3[0][89] ), .ZN(\SB2_0_17/i1_5 ) );
  INV_X1 \SB2_0_17/INV_4  ( .A(\RI3[0][88] ), .ZN(\SB2_0_17/i0[7] ) );
  INV_X1 \SB2_0_17/INV_3  ( .A(\RI3[0][87] ), .ZN(\SB2_0_17/i0[8] ) );
  INV_X1 \SB2_0_17/INV_2  ( .A(\RI3[0][86] ), .ZN(\SB2_0_17/i1[9] ) );
  INV_X1 \SB2_0_17/INV_1  ( .A(\RI3[0][85] ), .ZN(\SB2_0_17/i1_7 ) );
  INV_X1 \SB2_0_17/INV_0  ( .A(\RI3[0][84] ), .ZN(\SB2_0_17/i3[0] ) );
  INV_X1 \SB2_0_18/INV_4  ( .A(\RI3[0][82] ), .ZN(\SB2_0_18/i0[7] ) );
  INV_X1 \SB2_0_18/INV_3  ( .A(\RI3[0][81] ), .ZN(\SB2_0_18/i0[8] ) );
  INV_X1 \SB2_0_18/INV_1  ( .A(\RI3[0][79] ), .ZN(\SB2_0_18/i1_7 ) );
  INV_X1 \SB2_0_18/INV_0  ( .A(\RI3[0][78] ), .ZN(\SB2_0_18/i3[0] ) );
  INV_X1 \SB2_0_19/INV_5  ( .A(\RI3[0][77] ), .ZN(\SB2_0_19/i1_5 ) );
  INV_X1 \SB2_0_19/INV_4  ( .A(\RI3[0][76] ), .ZN(\SB2_0_19/i0[7] ) );
  INV_X1 \SB2_0_19/INV_3  ( .A(\RI3[0][75] ), .ZN(\SB2_0_19/i0[8] ) );
  INV_X1 \SB2_0_19/INV_2  ( .A(\RI3[0][74] ), .ZN(\SB2_0_19/i1[9] ) );
  INV_X1 \SB2_0_19/INV_1  ( .A(\RI3[0][73] ), .ZN(\SB2_0_19/i1_7 ) );
  INV_X1 \SB2_0_19/INV_0  ( .A(\RI3[0][72] ), .ZN(\SB2_0_19/i3[0] ) );
  INV_X1 \SB2_0_20/INV_5  ( .A(\RI3[0][71] ), .ZN(\SB2_0_20/i1_5 ) );
  INV_X1 \SB2_0_20/INV_4  ( .A(\RI3[0][70] ), .ZN(\SB2_0_20/i0[7] ) );
  INV_X1 \SB2_0_20/INV_3  ( .A(\RI3[0][69] ), .ZN(\SB2_0_20/i0[8] ) );
  INV_X1 \SB2_0_20/INV_1  ( .A(\RI3[0][67] ), .ZN(\SB2_0_20/i1_7 ) );
  INV_X1 \SB2_0_20/INV_0  ( .A(\RI3[0][66] ), .ZN(\SB2_0_20/i3[0] ) );
  INV_X1 \SB2_0_21/INV_5  ( .A(\RI3[0][65] ), .ZN(\SB2_0_21/i1_5 ) );
  INV_X1 \SB2_0_21/INV_4  ( .A(\RI3[0][64] ), .ZN(\SB2_0_21/i0[7] ) );
  INV_X1 \SB2_0_21/INV_3  ( .A(\RI3[0][63] ), .ZN(\SB2_0_21/i0[8] ) );
  INV_X1 \SB2_0_21/INV_1  ( .A(\RI3[0][61] ), .ZN(\SB2_0_21/i1_7 ) );
  INV_X1 \SB2_0_21/INV_0  ( .A(\RI3[0][60] ), .ZN(\SB2_0_21/i3[0] ) );
  INV_X1 \SB2_0_22/INV_5  ( .A(\RI3[0][59] ), .ZN(\SB2_0_22/i1_5 ) );
  INV_X1 \SB2_0_22/INV_4  ( .A(\RI3[0][58] ), .ZN(\SB2_0_22/i0[7] ) );
  INV_X1 \SB2_0_22/INV_3  ( .A(\RI3[0][57] ), .ZN(\SB2_0_22/i0[8] ) );
  INV_X1 \SB2_0_22/INV_2  ( .A(\RI3[0][56] ), .ZN(\SB2_0_22/i1[9] ) );
  INV_X1 \SB2_0_22/INV_1  ( .A(\RI3[0][55] ), .ZN(\SB2_0_22/i1_7 ) );
  INV_X1 \SB2_0_22/INV_0  ( .A(\RI3[0][54] ), .ZN(\SB2_0_22/i3[0] ) );
  INV_X1 \SB2_0_23/INV_4  ( .A(\SB2_0_23/i0_4 ), .ZN(\SB2_0_23/i0[7] ) );
  INV_X1 \SB2_0_23/INV_3  ( .A(\RI3[0][51] ), .ZN(\SB2_0_23/i0[8] ) );
  INV_X1 \SB2_0_23/INV_1  ( .A(\RI3[0][49] ), .ZN(\SB2_0_23/i1_7 ) );
  INV_X1 \SB2_0_23/INV_0  ( .A(\RI3[0][48] ), .ZN(\SB2_0_23/i3[0] ) );
  INV_X1 \SB2_0_24/INV_5  ( .A(\RI3[0][47] ), .ZN(\SB2_0_24/i1_5 ) );
  INV_X1 \SB2_0_24/INV_4  ( .A(\RI3[0][46] ), .ZN(\SB2_0_24/i0[7] ) );
  INV_X1 \SB2_0_24/INV_3  ( .A(\RI3[0][45] ), .ZN(\SB2_0_24/i0[8] ) );
  INV_X1 \SB2_0_24/INV_2  ( .A(\RI3[0][44] ), .ZN(\SB2_0_24/i1[9] ) );
  INV_X1 \SB2_0_24/INV_1  ( .A(\RI3[0][43] ), .ZN(\SB2_0_24/i1_7 ) );
  INV_X1 \SB2_0_24/INV_0  ( .A(\RI3[0][42] ), .ZN(\SB2_0_24/i3[0] ) );
  INV_X1 \SB2_0_25/INV_5  ( .A(\RI3[0][41] ), .ZN(\SB2_0_25/i1_5 ) );
  INV_X1 \SB2_0_25/INV_4  ( .A(\RI3[0][40] ), .ZN(\SB2_0_25/i0[7] ) );
  INV_X1 \SB2_0_25/INV_3  ( .A(\RI3[0][39] ), .ZN(\SB2_0_25/i0[8] ) );
  INV_X1 \SB2_0_25/INV_2  ( .A(\RI3[0][38] ), .ZN(\SB2_0_25/i1[9] ) );
  INV_X1 \SB2_0_25/INV_1  ( .A(\RI3[0][37] ), .ZN(\SB2_0_25/i1_7 ) );
  INV_X1 \SB2_0_25/INV_0  ( .A(\RI3[0][36] ), .ZN(\SB2_0_25/i3[0] ) );
  INV_X1 \SB2_0_26/INV_5  ( .A(\RI3[0][35] ), .ZN(\SB2_0_26/i1_5 ) );
  INV_X1 \SB2_0_26/INV_4  ( .A(\RI3[0][34] ), .ZN(\SB2_0_26/i0[7] ) );
  INV_X1 \SB2_0_26/INV_3  ( .A(\RI3[0][33] ), .ZN(\SB2_0_26/i0[8] ) );
  INV_X1 \SB2_0_26/INV_2  ( .A(\RI3[0][32] ), .ZN(\SB2_0_26/i1[9] ) );
  INV_X1 \SB2_0_26/INV_1  ( .A(\RI3[0][31] ), .ZN(\SB2_0_26/i1_7 ) );
  INV_X1 \SB2_0_26/INV_0  ( .A(\RI3[0][30] ), .ZN(\SB2_0_26/i3[0] ) );
  INV_X1 \SB2_0_27/INV_5  ( .A(\RI3[0][29] ), .ZN(\SB2_0_27/i1_5 ) );
  INV_X1 \SB2_0_27/INV_4  ( .A(\RI3[0][28] ), .ZN(\SB2_0_27/i0[7] ) );
  INV_X1 \SB2_0_27/INV_3  ( .A(\RI3[0][27] ), .ZN(\SB2_0_27/i0[8] ) );
  INV_X1 \SB2_0_27/INV_2  ( .A(\RI3[0][26] ), .ZN(\SB2_0_27/i1[9] ) );
  INV_X1 \SB2_0_27/INV_1  ( .A(\RI3[0][25] ), .ZN(\SB2_0_27/i1_7 ) );
  INV_X1 \SB2_0_27/INV_0  ( .A(\RI3[0][24] ), .ZN(\SB2_0_27/i3[0] ) );
  INV_X1 \SB2_0_28/INV_5  ( .A(\RI3[0][23] ), .ZN(\SB2_0_28/i1_5 ) );
  INV_X1 \SB2_0_28/INV_4  ( .A(\RI3[0][22] ), .ZN(\SB2_0_28/i0[7] ) );
  INV_X1 \SB2_0_28/INV_3  ( .A(\RI3[0][21] ), .ZN(\SB2_0_28/i0[8] ) );
  INV_X1 \SB2_0_28/INV_2  ( .A(\RI3[0][20] ), .ZN(\SB2_0_28/i1[9] ) );
  INV_X1 \SB2_0_28/INV_1  ( .A(\RI3[0][19] ), .ZN(\SB2_0_28/i1_7 ) );
  INV_X1 \SB2_0_28/INV_0  ( .A(\RI3[0][18] ), .ZN(\SB2_0_28/i3[0] ) );
  INV_X1 \SB2_0_29/INV_5  ( .A(\RI3[0][17] ), .ZN(\SB2_0_29/i1_5 ) );
  INV_X1 \SB2_0_29/INV_4  ( .A(\RI3[0][16] ), .ZN(\SB2_0_29/i0[7] ) );
  INV_X1 \SB2_0_29/INV_3  ( .A(\RI3[0][15] ), .ZN(\SB2_0_29/i0[8] ) );
  INV_X1 \SB2_0_29/INV_2  ( .A(\RI3[0][14] ), .ZN(\SB2_0_29/i1[9] ) );
  INV_X1 \SB2_0_29/INV_1  ( .A(\RI3[0][13] ), .ZN(\SB2_0_29/i1_7 ) );
  INV_X1 \SB2_0_29/INV_0  ( .A(\RI3[0][12] ), .ZN(\SB2_0_29/i3[0] ) );
  INV_X1 \SB2_0_30/INV_5  ( .A(\RI3[0][11] ), .ZN(\SB2_0_30/i1_5 ) );
  INV_X1 \SB2_0_30/INV_4  ( .A(\RI3[0][10] ), .ZN(\SB2_0_30/i0[7] ) );
  INV_X1 \SB2_0_30/INV_3  ( .A(\RI3[0][9] ), .ZN(\SB2_0_30/i0[8] ) );
  INV_X1 \SB2_0_30/INV_2  ( .A(\RI3[0][8] ), .ZN(\SB2_0_30/i1[9] ) );
  INV_X1 \SB2_0_30/INV_1  ( .A(\RI3[0][7] ), .ZN(\SB2_0_30/i1_7 ) );
  INV_X1 \SB2_0_30/INV_0  ( .A(\RI3[0][6] ), .ZN(\SB2_0_30/i3[0] ) );
  INV_X1 \SB2_0_31/INV_5  ( .A(\RI3[0][5] ), .ZN(\SB2_0_31/i1_5 ) );
  INV_X1 \SB2_0_31/INV_4  ( .A(\RI3[0][4] ), .ZN(\SB2_0_31/i0[7] ) );
  INV_X1 \SB2_0_31/INV_3  ( .A(\RI3[0][3] ), .ZN(\SB2_0_31/i0[8] ) );
  INV_X1 \SB2_0_31/INV_2  ( .A(\RI3[0][2] ), .ZN(\SB2_0_31/i1[9] ) );
  INV_X1 \SB2_0_31/INV_1  ( .A(\RI3[0][1] ), .ZN(\SB2_0_31/i1_7 ) );
  INV_X1 \SB2_0_31/INV_0  ( .A(\RI3[0][0] ), .ZN(\SB2_0_31/i3[0] ) );
  INV_X1 \SB2_1_0/INV_5  ( .A(\RI3[1][191] ), .ZN(\SB2_1_0/i1_5 ) );
  INV_X1 \SB2_1_0/INV_4  ( .A(\RI3[1][190] ), .ZN(\SB2_1_0/i0[7] ) );
  INV_X1 \SB2_1_0/INV_3  ( .A(\RI3[1][189] ), .ZN(\SB2_1_0/i0[8] ) );
  INV_X1 \SB2_1_0/INV_2  ( .A(\RI3[1][188] ), .ZN(\SB2_1_0/i1[9] ) );
  INV_X1 \SB2_1_0/INV_1  ( .A(\RI3[1][187] ), .ZN(\SB2_1_0/i1_7 ) );
  INV_X1 \SB2_1_0/INV_0  ( .A(\RI3[1][186] ), .ZN(\SB2_1_0/i3[0] ) );
  INV_X1 \SB2_1_1/INV_5  ( .A(\RI3[1][185] ), .ZN(\SB2_1_1/i1_5 ) );
  INV_X1 \SB2_1_1/INV_4  ( .A(\RI3[1][184] ), .ZN(\SB2_1_1/i0[7] ) );
  INV_X1 \SB2_1_1/INV_3  ( .A(\RI3[1][183] ), .ZN(\SB2_1_1/i0[8] ) );
  INV_X1 \SB2_1_1/INV_2  ( .A(\RI3[1][182] ), .ZN(\SB2_1_1/i1[9] ) );
  INV_X1 \SB2_1_1/INV_1  ( .A(\RI3[1][181] ), .ZN(\SB2_1_1/i1_7 ) );
  INV_X1 \SB2_1_1/INV_0  ( .A(\RI3[1][180] ), .ZN(\SB2_1_1/i3[0] ) );
  INV_X1 \SB2_1_2/INV_4  ( .A(\RI3[1][178] ), .ZN(\SB2_1_2/i0[7] ) );
  INV_X1 \SB2_1_2/INV_3  ( .A(\RI3[1][177] ), .ZN(\SB2_1_2/i0[8] ) );
  INV_X1 \SB2_1_2/INV_2  ( .A(\RI3[1][176] ), .ZN(\SB2_1_2/i1[9] ) );
  INV_X1 \SB2_1_2/INV_1  ( .A(\RI3[1][175] ), .ZN(\SB2_1_2/i1_7 ) );
  INV_X1 \SB2_1_2/INV_0  ( .A(\RI3[1][174] ), .ZN(\SB2_1_2/i3[0] ) );
  INV_X1 \SB2_1_3/INV_5  ( .A(\RI3[1][173] ), .ZN(\SB2_1_3/i1_5 ) );
  INV_X1 \SB2_1_3/INV_4  ( .A(\RI3[1][172] ), .ZN(\SB2_1_3/i0[7] ) );
  INV_X1 \SB2_1_3/INV_3  ( .A(\RI3[1][171] ), .ZN(\SB2_1_3/i0[8] ) );
  INV_X1 \SB2_1_3/INV_2  ( .A(\RI3[1][170] ), .ZN(\SB2_1_3/i1[9] ) );
  INV_X1 \SB2_1_3/INV_1  ( .A(\RI3[1][169] ), .ZN(\SB2_1_3/i1_7 ) );
  INV_X1 \SB2_1_3/INV_0  ( .A(\RI3[1][168] ), .ZN(\SB2_1_3/i3[0] ) );
  INV_X1 \SB2_1_4/INV_5  ( .A(\RI3[1][167] ), .ZN(\SB2_1_4/i1_5 ) );
  INV_X1 \SB2_1_4/INV_4  ( .A(\RI3[1][166] ), .ZN(\SB2_1_4/i0[7] ) );
  INV_X1 \SB2_1_4/INV_3  ( .A(\RI3[1][165] ), .ZN(\SB2_1_4/i0[8] ) );
  INV_X1 \SB2_1_4/INV_2  ( .A(\RI3[1][164] ), .ZN(\SB2_1_4/i1[9] ) );
  INV_X1 \SB2_1_4/INV_1  ( .A(\RI3[1][163] ), .ZN(\SB2_1_4/i1_7 ) );
  INV_X1 \SB2_1_4/INV_0  ( .A(\RI3[1][162] ), .ZN(\SB2_1_4/i3[0] ) );
  INV_X1 \SB2_1_5/INV_5  ( .A(\RI3[1][161] ), .ZN(\SB2_1_5/i1_5 ) );
  INV_X1 \SB2_1_5/INV_4  ( .A(\RI3[1][160] ), .ZN(\SB2_1_5/i0[7] ) );
  INV_X1 \SB2_1_5/INV_3  ( .A(\RI3[1][159] ), .ZN(\SB2_1_5/i0[8] ) );
  INV_X1 \SB2_1_5/INV_2  ( .A(\RI3[1][158] ), .ZN(\SB2_1_5/i1[9] ) );
  INV_X1 \SB2_1_5/INV_1  ( .A(\RI3[1][157] ), .ZN(\SB2_1_5/i1_7 ) );
  INV_X1 \SB2_1_5/INV_0  ( .A(\RI3[1][156] ), .ZN(\SB2_1_5/i3[0] ) );
  INV_X1 \SB2_1_6/INV_5  ( .A(\RI3[1][155] ), .ZN(\SB2_1_6/i1_5 ) );
  INV_X1 \SB2_1_6/INV_4  ( .A(\RI3[1][154] ), .ZN(\SB2_1_6/i0[7] ) );
  INV_X1 \SB2_1_6/INV_3  ( .A(\RI3[1][153] ), .ZN(\SB2_1_6/i0[8] ) );
  INV_X1 \SB2_1_6/INV_1  ( .A(\RI3[1][151] ), .ZN(\SB2_1_6/i1_7 ) );
  INV_X1 \SB2_1_6/INV_0  ( .A(\RI3[1][150] ), .ZN(\SB2_1_6/i3[0] ) );
  INV_X1 \SB2_1_7/INV_5  ( .A(\RI3[1][149] ), .ZN(\SB2_1_7/i1_5 ) );
  INV_X1 \SB2_1_7/INV_4  ( .A(\SB2_1_7/i0_4 ), .ZN(\SB2_1_7/i0[7] ) );
  INV_X1 \SB2_1_7/INV_3  ( .A(\RI3[1][147] ), .ZN(\SB2_1_7/i0[8] ) );
  INV_X1 \SB2_1_7/INV_2  ( .A(\RI3[1][146] ), .ZN(\SB2_1_7/i1[9] ) );
  INV_X1 \SB2_1_7/INV_1  ( .A(\RI3[1][145] ), .ZN(\SB2_1_7/i1_7 ) );
  INV_X1 \SB2_1_7/INV_0  ( .A(\RI3[1][144] ), .ZN(\SB2_1_7/i3[0] ) );
  INV_X1 \SB2_1_8/INV_5  ( .A(\RI3[1][143] ), .ZN(\SB2_1_8/i1_5 ) );
  INV_X1 \SB2_1_8/INV_4  ( .A(\RI3[1][142] ), .ZN(\SB2_1_8/i0[7] ) );
  INV_X1 \SB2_1_8/INV_3  ( .A(\RI3[1][141] ), .ZN(\SB2_1_8/i0[8] ) );
  INV_X1 \SB2_1_8/INV_2  ( .A(\RI3[1][140] ), .ZN(\SB2_1_8/i1[9] ) );
  INV_X1 \SB2_1_8/INV_1  ( .A(\RI3[1][139] ), .ZN(\SB2_1_8/i1_7 ) );
  INV_X1 \SB2_1_8/INV_0  ( .A(\RI3[1][138] ), .ZN(\SB2_1_8/i3[0] ) );
  INV_X1 \SB2_1_9/INV_5  ( .A(\RI3[1][137] ), .ZN(\SB2_1_9/i1_5 ) );
  INV_X1 \SB2_1_9/INV_4  ( .A(\RI3[1][136] ), .ZN(\SB2_1_9/i0[7] ) );
  INV_X1 \SB2_1_9/INV_3  ( .A(\RI3[1][135] ), .ZN(\SB2_1_9/i0[8] ) );
  INV_X1 \SB2_1_9/INV_2  ( .A(\RI3[1][134] ), .ZN(\SB2_1_9/i1[9] ) );
  INV_X1 \SB2_1_9/INV_1  ( .A(\RI3[1][133] ), .ZN(\SB2_1_9/i1_7 ) );
  INV_X1 \SB2_1_9/INV_0  ( .A(\RI3[1][132] ), .ZN(\SB2_1_9/i3[0] ) );
  INV_X1 \SB2_1_10/INV_5  ( .A(\RI3[1][131] ), .ZN(\SB2_1_10/i1_5 ) );
  INV_X1 \SB2_1_10/INV_4  ( .A(\RI3[1][130] ), .ZN(\SB2_1_10/i0[7] ) );
  INV_X1 \SB2_1_10/INV_3  ( .A(\RI3[1][129] ), .ZN(\SB2_1_10/i0[8] ) );
  INV_X1 \SB2_1_10/INV_2  ( .A(\RI3[1][128] ), .ZN(\SB2_1_10/i1[9] ) );
  INV_X1 \SB2_1_10/INV_1  ( .A(\RI3[1][127] ), .ZN(\SB2_1_10/i1_7 ) );
  INV_X1 \SB2_1_10/INV_0  ( .A(\RI3[1][126] ), .ZN(\SB2_1_10/i3[0] ) );
  INV_X1 \SB2_1_11/INV_5  ( .A(\RI3[1][125] ), .ZN(\SB2_1_11/i1_5 ) );
  INV_X1 \SB2_1_11/INV_4  ( .A(\RI3[1][124] ), .ZN(\SB2_1_11/i0[7] ) );
  INV_X1 \SB2_1_11/INV_3  ( .A(\RI3[1][123] ), .ZN(\SB2_1_11/i0[8] ) );
  INV_X1 \SB2_1_11/INV_2  ( .A(\RI3[1][122] ), .ZN(\SB2_1_11/i1[9] ) );
  INV_X1 \SB2_1_11/INV_1  ( .A(\RI3[1][121] ), .ZN(\SB2_1_11/i1_7 ) );
  INV_X1 \SB2_1_11/INV_0  ( .A(\RI3[1][120] ), .ZN(\SB2_1_11/i3[0] ) );
  INV_X1 \SB2_1_12/INV_5  ( .A(\RI3[1][119] ), .ZN(\SB2_1_12/i1_5 ) );
  INV_X1 \SB2_1_12/INV_4  ( .A(\RI3[1][118] ), .ZN(\SB2_1_12/i0[7] ) );
  INV_X1 \SB2_1_12/INV_3  ( .A(\RI3[1][117] ), .ZN(\SB2_1_12/i0[8] ) );
  INV_X1 \SB2_1_12/INV_2  ( .A(\RI3[1][116] ), .ZN(\SB2_1_12/i1[9] ) );
  INV_X1 \SB2_1_12/INV_1  ( .A(\RI3[1][115] ), .ZN(\SB2_1_12/i1_7 ) );
  INV_X1 \SB2_1_12/INV_0  ( .A(\RI3[1][114] ), .ZN(\SB2_1_12/i3[0] ) );
  INV_X1 \SB2_1_13/INV_5  ( .A(\RI3[1][113] ), .ZN(\SB2_1_13/i1_5 ) );
  INV_X1 \SB2_1_13/INV_4  ( .A(\RI3[1][112] ), .ZN(\SB2_1_13/i0[7] ) );
  INV_X1 \SB2_1_13/INV_3  ( .A(\RI3[1][111] ), .ZN(\SB2_1_13/i0[8] ) );
  INV_X1 \SB2_1_13/INV_2  ( .A(\RI3[1][110] ), .ZN(\SB2_1_13/i1[9] ) );
  INV_X1 \SB2_1_13/INV_1  ( .A(\RI3[1][109] ), .ZN(\SB2_1_13/i1_7 ) );
  INV_X1 \SB2_1_13/INV_0  ( .A(\RI3[1][108] ), .ZN(\SB2_1_13/i3[0] ) );
  INV_X1 \SB2_1_14/INV_5  ( .A(\RI3[1][107] ), .ZN(\SB2_1_14/i1_5 ) );
  INV_X1 \SB2_1_14/INV_4  ( .A(\RI3[1][106] ), .ZN(\SB2_1_14/i0[7] ) );
  INV_X1 \SB2_1_14/INV_3  ( .A(\RI3[1][105] ), .ZN(\SB2_1_14/i0[8] ) );
  INV_X1 \SB2_1_14/INV_1  ( .A(\RI3[1][103] ), .ZN(\SB2_1_14/i1_7 ) );
  INV_X1 \SB2_1_14/INV_0  ( .A(\RI3[1][102] ), .ZN(\SB2_1_14/i3[0] ) );
  INV_X1 \SB2_1_15/INV_5  ( .A(\RI3[1][101] ), .ZN(\SB2_1_15/i1_5 ) );
  INV_X1 \SB2_1_15/INV_4  ( .A(\RI3[1][100] ), .ZN(\SB2_1_15/i0[7] ) );
  INV_X1 \SB2_1_15/INV_3  ( .A(\RI3[1][99] ), .ZN(\SB2_1_15/i0[8] ) );
  INV_X1 \SB2_1_15/INV_1  ( .A(\RI3[1][97] ), .ZN(\SB2_1_15/i1_7 ) );
  INV_X1 \SB2_1_15/INV_0  ( .A(\RI3[1][96] ), .ZN(\SB2_1_15/i3[0] ) );
  INV_X1 \SB2_1_16/INV_5  ( .A(\RI3[1][95] ), .ZN(\SB2_1_16/i1_5 ) );
  INV_X1 \SB2_1_16/INV_4  ( .A(\RI3[1][94] ), .ZN(\SB2_1_16/i0[7] ) );
  INV_X1 \SB2_1_16/INV_3  ( .A(\RI3[1][93] ), .ZN(\SB2_1_16/i0[8] ) );
  INV_X1 \SB2_1_16/INV_2  ( .A(\RI3[1][92] ), .ZN(\SB2_1_16/i1[9] ) );
  INV_X1 \SB2_1_16/INV_1  ( .A(\RI3[1][91] ), .ZN(\SB2_1_16/i1_7 ) );
  INV_X1 \SB2_1_16/INV_0  ( .A(\RI3[1][90] ), .ZN(\SB2_1_16/i3[0] ) );
  INV_X1 \SB2_1_17/INV_5  ( .A(\RI3[1][89] ), .ZN(\SB2_1_17/i1_5 ) );
  INV_X1 \SB2_1_17/INV_4  ( .A(\RI3[1][88] ), .ZN(\SB2_1_17/i0[7] ) );
  INV_X1 \SB2_1_17/INV_3  ( .A(\RI3[1][87] ), .ZN(\SB2_1_17/i0[8] ) );
  INV_X1 \SB2_1_17/INV_1  ( .A(\RI3[1][85] ), .ZN(\SB2_1_17/i1_7 ) );
  INV_X1 \SB2_1_17/INV_0  ( .A(\RI3[1][84] ), .ZN(\SB2_1_17/i3[0] ) );
  INV_X1 \SB2_1_18/INV_5  ( .A(\RI3[1][83] ), .ZN(\SB2_1_18/i1_5 ) );
  INV_X1 \SB2_1_18/INV_4  ( .A(\RI3[1][82] ), .ZN(\SB2_1_18/i0[7] ) );
  INV_X1 \SB2_1_18/INV_3  ( .A(\RI3[1][81] ), .ZN(\SB2_1_18/i0[8] ) );
  INV_X1 \SB2_1_18/INV_2  ( .A(\RI3[1][80] ), .ZN(\SB2_1_18/i1[9] ) );
  INV_X1 \SB2_1_18/INV_1  ( .A(\RI3[1][79] ), .ZN(\SB2_1_18/i1_7 ) );
  INV_X1 \SB2_1_18/INV_0  ( .A(\RI3[1][78] ), .ZN(\SB2_1_18/i3[0] ) );
  INV_X1 \SB2_1_19/INV_5  ( .A(\RI3[1][77] ), .ZN(\SB2_1_19/i1_5 ) );
  INV_X1 \SB2_1_19/INV_4  ( .A(\RI3[1][76] ), .ZN(\SB2_1_19/i0[7] ) );
  INV_X1 \SB2_1_19/INV_3  ( .A(\RI3[1][75] ), .ZN(\SB2_1_19/i0[8] ) );
  INV_X1 \SB2_1_19/INV_2  ( .A(\RI3[1][74] ), .ZN(\SB2_1_19/i1[9] ) );
  INV_X1 \SB2_1_19/INV_1  ( .A(\RI3[1][73] ), .ZN(\SB2_1_19/i1_7 ) );
  INV_X1 \SB2_1_19/INV_0  ( .A(\RI3[1][72] ), .ZN(\SB2_1_19/i3[0] ) );
  INV_X1 \SB2_1_20/INV_5  ( .A(\RI3[1][71] ), .ZN(\SB2_1_20/i1_5 ) );
  INV_X1 \SB2_1_20/INV_4  ( .A(\RI3[1][70] ), .ZN(\SB2_1_20/i0[7] ) );
  INV_X1 \SB2_1_20/INV_3  ( .A(\RI3[1][69] ), .ZN(\SB2_1_20/i0[8] ) );
  INV_X1 \SB2_1_20/INV_2  ( .A(\RI3[1][68] ), .ZN(\SB2_1_20/i1[9] ) );
  INV_X1 \SB2_1_20/INV_1  ( .A(\RI3[1][67] ), .ZN(\SB2_1_20/i1_7 ) );
  INV_X1 \SB2_1_20/INV_0  ( .A(\RI3[1][66] ), .ZN(\SB2_1_20/i3[0] ) );
  INV_X1 \SB2_1_21/INV_5  ( .A(\RI3[1][65] ), .ZN(\SB2_1_21/i1_5 ) );
  INV_X1 \SB2_1_21/INV_4  ( .A(\RI3[1][64] ), .ZN(\SB2_1_21/i0[7] ) );
  INV_X1 \SB2_1_21/INV_3  ( .A(\RI3[1][63] ), .ZN(\SB2_1_21/i0[8] ) );
  INV_X1 \SB2_1_21/INV_2  ( .A(\RI3[1][62] ), .ZN(\SB2_1_21/i1[9] ) );
  INV_X1 \SB2_1_21/INV_1  ( .A(\RI3[1][61] ), .ZN(\SB2_1_21/i1_7 ) );
  INV_X1 \SB2_1_21/INV_0  ( .A(\RI3[1][60] ), .ZN(\SB2_1_21/i3[0] ) );
  INV_X1 \SB2_1_22/INV_5  ( .A(\RI3[1][59] ), .ZN(\SB2_1_22/i1_5 ) );
  INV_X1 \SB2_1_22/INV_4  ( .A(\RI3[1][58] ), .ZN(\SB2_1_22/i0[7] ) );
  INV_X1 \SB2_1_22/INV_3  ( .A(\RI3[1][57] ), .ZN(\SB2_1_22/i0[8] ) );
  INV_X1 \SB2_1_22/INV_2  ( .A(\RI3[1][56] ), .ZN(\SB2_1_22/i1[9] ) );
  INV_X1 \SB2_1_22/INV_1  ( .A(\RI3[1][55] ), .ZN(\SB2_1_22/i1_7 ) );
  INV_X1 \SB2_1_22/INV_0  ( .A(\RI3[1][54] ), .ZN(\SB2_1_22/i3[0] ) );
  INV_X1 \SB2_1_23/INV_5  ( .A(\RI3[1][53] ), .ZN(\SB2_1_23/i1_5 ) );
  INV_X1 \SB2_1_23/INV_4  ( .A(\RI3[1][52] ), .ZN(\SB2_1_23/i0[7] ) );
  INV_X1 \SB2_1_23/INV_3  ( .A(\RI3[1][51] ), .ZN(\SB2_1_23/i0[8] ) );
  INV_X1 \SB2_1_23/INV_2  ( .A(\RI3[1][50] ), .ZN(\SB2_1_23/i1[9] ) );
  INV_X1 \SB2_1_23/INV_1  ( .A(\RI3[1][49] ), .ZN(\SB2_1_23/i1_7 ) );
  INV_X1 \SB2_1_23/INV_0  ( .A(\RI3[1][48] ), .ZN(\SB2_1_23/i3[0] ) );
  BUF_X1 \SB2_1_23/BUF_0  ( .A(\RI3[1][48] ), .Z(\SB2_1_23/i0[9] ) );
  INV_X1 \SB2_1_24/INV_5  ( .A(\RI3[1][47] ), .ZN(\SB2_1_24/i1_5 ) );
  INV_X1 \SB2_1_24/INV_4  ( .A(\RI3[1][46] ), .ZN(\SB2_1_24/i0[7] ) );
  INV_X1 \SB2_1_24/INV_3  ( .A(\RI3[1][45] ), .ZN(\SB2_1_24/i0[8] ) );
  INV_X1 \SB2_1_24/INV_2  ( .A(\RI3[1][44] ), .ZN(\SB2_1_24/i1[9] ) );
  INV_X1 \SB2_1_24/INV_1  ( .A(\RI3[1][43] ), .ZN(\SB2_1_24/i1_7 ) );
  INV_X1 \SB2_1_24/INV_0  ( .A(\RI3[1][42] ), .ZN(\SB2_1_24/i3[0] ) );
  INV_X1 \SB2_1_25/INV_5  ( .A(\RI3[1][41] ), .ZN(\SB2_1_25/i1_5 ) );
  INV_X1 \SB2_1_25/INV_4  ( .A(\RI3[1][40] ), .ZN(\SB2_1_25/i0[7] ) );
  INV_X1 \SB2_1_25/INV_3  ( .A(\RI3[1][39] ), .ZN(\SB2_1_25/i0[8] ) );
  INV_X1 \SB2_1_25/INV_2  ( .A(\RI3[1][38] ), .ZN(\SB2_1_25/i1[9] ) );
  INV_X1 \SB2_1_25/INV_1  ( .A(\RI3[1][37] ), .ZN(\SB2_1_25/i1_7 ) );
  INV_X1 \SB2_1_25/INV_0  ( .A(\RI3[1][36] ), .ZN(\SB2_1_25/i3[0] ) );
  INV_X1 \SB2_1_26/INV_5  ( .A(\RI3[1][35] ), .ZN(\SB2_1_26/i1_5 ) );
  INV_X1 \SB2_1_26/INV_4  ( .A(\RI3[1][34] ), .ZN(\SB2_1_26/i0[7] ) );
  INV_X1 \SB2_1_26/INV_3  ( .A(\RI3[1][33] ), .ZN(\SB2_1_26/i0[8] ) );
  INV_X1 \SB2_1_26/INV_2  ( .A(\RI3[1][32] ), .ZN(\SB2_1_26/i1[9] ) );
  INV_X1 \SB2_1_26/INV_1  ( .A(\RI3[1][31] ), .ZN(\SB2_1_26/i1_7 ) );
  INV_X1 \SB2_1_26/INV_0  ( .A(\RI3[1][30] ), .ZN(\SB2_1_26/i3[0] ) );
  INV_X1 \SB2_1_27/INV_5  ( .A(\RI3[1][29] ), .ZN(\SB2_1_27/i1_5 ) );
  INV_X1 \SB2_1_27/INV_4  ( .A(\RI3[1][28] ), .ZN(\SB2_1_27/i0[7] ) );
  INV_X1 \SB2_1_27/INV_3  ( .A(\RI3[1][27] ), .ZN(\SB2_1_27/i0[8] ) );
  INV_X1 \SB2_1_27/INV_2  ( .A(\RI3[1][26] ), .ZN(\SB2_1_27/i1[9] ) );
  INV_X1 \SB2_1_27/INV_1  ( .A(\RI3[1][25] ), .ZN(\SB2_1_27/i1_7 ) );
  INV_X1 \SB2_1_27/INV_0  ( .A(\RI3[1][24] ), .ZN(\SB2_1_27/i3[0] ) );
  INV_X1 \SB2_1_28/INV_5  ( .A(\RI3[1][23] ), .ZN(\SB2_1_28/i1_5 ) );
  INV_X1 \SB2_1_28/INV_4  ( .A(\RI3[1][22] ), .ZN(\SB2_1_28/i0[7] ) );
  INV_X1 \SB2_1_28/INV_3  ( .A(\RI3[1][21] ), .ZN(\SB2_1_28/i0[8] ) );
  INV_X1 \SB2_1_28/INV_2  ( .A(\RI3[1][20] ), .ZN(\SB2_1_28/i1[9] ) );
  INV_X1 \SB2_1_28/INV_1  ( .A(\RI3[1][19] ), .ZN(\SB2_1_28/i1_7 ) );
  INV_X1 \SB2_1_28/INV_0  ( .A(\RI3[1][18] ), .ZN(\SB2_1_28/i3[0] ) );
  INV_X1 \SB2_1_29/INV_5  ( .A(\RI3[1][17] ), .ZN(\SB2_1_29/i1_5 ) );
  INV_X1 \SB2_1_29/INV_4  ( .A(\RI3[1][16] ), .ZN(\SB2_1_29/i0[7] ) );
  INV_X1 \SB2_1_29/INV_3  ( .A(\RI3[1][15] ), .ZN(\SB2_1_29/i0[8] ) );
  INV_X1 \SB2_1_29/INV_2  ( .A(\RI3[1][14] ), .ZN(\SB2_1_29/i1[9] ) );
  INV_X1 \SB2_1_29/INV_1  ( .A(\RI3[1][13] ), .ZN(\SB2_1_29/i1_7 ) );
  INV_X1 \SB2_1_29/INV_0  ( .A(\RI3[1][12] ), .ZN(\SB2_1_29/i3[0] ) );
  INV_X1 \SB2_1_30/INV_5  ( .A(\RI3[1][11] ), .ZN(\SB2_1_30/i1_5 ) );
  INV_X1 \SB2_1_30/INV_4  ( .A(\RI3[1][10] ), .ZN(\SB2_1_30/i0[7] ) );
  INV_X1 \SB2_1_30/INV_3  ( .A(\RI3[1][9] ), .ZN(\SB2_1_30/i0[8] ) );
  INV_X1 \SB2_1_30/INV_2  ( .A(\RI3[1][8] ), .ZN(\SB2_1_30/i1[9] ) );
  INV_X1 \SB2_1_30/INV_1  ( .A(\RI3[1][7] ), .ZN(\SB2_1_30/i1_7 ) );
  INV_X1 \SB2_1_30/INV_0  ( .A(\RI3[1][6] ), .ZN(\SB2_1_30/i3[0] ) );
  INV_X1 \SB2_1_31/INV_5  ( .A(\RI3[1][5] ), .ZN(\SB2_1_31/i1_5 ) );
  INV_X1 \SB2_1_31/INV_4  ( .A(\RI3[1][4] ), .ZN(\SB2_1_31/i0[7] ) );
  INV_X1 \SB2_1_31/INV_3  ( .A(\RI3[1][3] ), .ZN(\SB2_1_31/i0[8] ) );
  INV_X1 \SB2_1_31/INV_1  ( .A(\RI3[1][1] ), .ZN(\SB2_1_31/i1_7 ) );
  INV_X1 \SB2_1_31/INV_0  ( .A(\RI3[1][0] ), .ZN(\SB2_1_31/i3[0] ) );
  INV_X1 \SB2_2_0/INV_5  ( .A(\RI3[2][191] ), .ZN(\SB2_2_0/i1_5 ) );
  INV_X1 \SB2_2_0/INV_4  ( .A(\RI3[2][190] ), .ZN(\SB2_2_0/i0[7] ) );
  INV_X1 \SB2_2_0/INV_3  ( .A(\RI3[2][189] ), .ZN(\SB2_2_0/i0[8] ) );
  INV_X1 \SB2_2_0/INV_2  ( .A(\RI3[2][188] ), .ZN(\SB2_2_0/i1[9] ) );
  INV_X1 \SB2_2_0/INV_1  ( .A(\RI3[2][187] ), .ZN(\SB2_2_0/i1_7 ) );
  INV_X1 \SB2_2_0/INV_0  ( .A(\RI3[2][186] ), .ZN(\SB2_2_0/i3[0] ) );
  INV_X1 \SB2_2_1/INV_5  ( .A(\RI3[2][185] ), .ZN(\SB2_2_1/i1_5 ) );
  INV_X1 \SB2_2_1/INV_4  ( .A(\RI3[2][184] ), .ZN(\SB2_2_1/i0[7] ) );
  INV_X1 \SB2_2_1/INV_3  ( .A(\RI3[2][183] ), .ZN(\SB2_2_1/i0[8] ) );
  INV_X1 \SB2_2_1/INV_1  ( .A(\RI3[2][181] ), .ZN(\SB2_2_1/i1_7 ) );
  INV_X1 \SB2_2_1/INV_0  ( .A(\RI3[2][180] ), .ZN(\SB2_2_1/i3[0] ) );
  BUF_X1 \SB2_2_1/BUF_0  ( .A(\RI3[2][180] ), .Z(\SB2_2_1/i0[9] ) );
  INV_X1 \SB2_2_2/INV_5  ( .A(\RI3[2][179] ), .ZN(\SB2_2_2/i1_5 ) );
  INV_X1 \SB2_2_2/INV_4  ( .A(\RI3[2][178] ), .ZN(\SB2_2_2/i0[7] ) );
  INV_X1 \SB2_2_2/INV_3  ( .A(\RI3[2][177] ), .ZN(\SB2_2_2/i0[8] ) );
  INV_X1 \SB2_2_2/INV_1  ( .A(\RI3[2][175] ), .ZN(\SB2_2_2/i1_7 ) );
  INV_X1 \SB2_2_2/INV_0  ( .A(\RI3[2][174] ), .ZN(\SB2_2_2/i3[0] ) );
  INV_X1 \SB2_2_3/INV_5  ( .A(\RI3[2][173] ), .ZN(\SB2_2_3/i1_5 ) );
  INV_X1 \SB2_2_3/INV_4  ( .A(\RI3[2][172] ), .ZN(\SB2_2_3/i0[7] ) );
  INV_X1 \SB2_2_3/INV_3  ( .A(\RI3[2][171] ), .ZN(\SB2_2_3/i0[8] ) );
  INV_X1 \SB2_2_3/INV_2  ( .A(\RI3[2][170] ), .ZN(\SB2_2_3/i1[9] ) );
  INV_X1 \SB2_2_3/INV_1  ( .A(\RI3[2][169] ), .ZN(\SB2_2_3/i1_7 ) );
  INV_X1 \SB2_2_3/INV_0  ( .A(\RI3[2][168] ), .ZN(\SB2_2_3/i3[0] ) );
  BUF_X1 \SB2_2_3/BUF_1  ( .A(\RI3[2][169] ), .Z(\SB2_2_3/i0[6] ) );
  INV_X1 \SB2_2_4/INV_5  ( .A(\RI3[2][167] ), .ZN(\SB2_2_4/i1_5 ) );
  INV_X1 \SB2_2_4/INV_4  ( .A(\RI3[2][166] ), .ZN(\SB2_2_4/i0[7] ) );
  INV_X1 \SB2_2_4/INV_3  ( .A(\RI3[2][165] ), .ZN(\SB2_2_4/i0[8] ) );
  INV_X1 \SB2_2_4/INV_2  ( .A(\RI3[2][164] ), .ZN(\SB2_2_4/i1[9] ) );
  INV_X1 \SB2_2_4/INV_1  ( .A(\RI3[2][163] ), .ZN(\SB2_2_4/i1_7 ) );
  INV_X1 \SB2_2_4/INV_0  ( .A(\RI3[2][162] ), .ZN(\SB2_2_4/i3[0] ) );
  INV_X1 \SB2_2_5/INV_5  ( .A(\RI3[2][161] ), .ZN(\SB2_2_5/i1_5 ) );
  INV_X1 \SB2_2_5/INV_4  ( .A(\RI3[2][160] ), .ZN(\SB2_2_5/i0[7] ) );
  INV_X1 \SB2_2_5/INV_3  ( .A(\RI3[2][159] ), .ZN(\SB2_2_5/i0[8] ) );
  INV_X1 \SB2_2_5/INV_1  ( .A(\RI3[2][157] ), .ZN(\SB2_2_5/i1_7 ) );
  INV_X1 \SB2_2_5/INV_0  ( .A(\RI3[2][156] ), .ZN(\SB2_2_5/i3[0] ) );
  INV_X1 \SB2_2_6/INV_5  ( .A(\RI3[2][155] ), .ZN(\SB2_2_6/i1_5 ) );
  INV_X1 \SB2_2_6/INV_4  ( .A(\RI3[2][154] ), .ZN(\SB2_2_6/i0[7] ) );
  INV_X1 \SB2_2_6/INV_3  ( .A(\RI3[2][153] ), .ZN(\SB2_2_6/i0[8] ) );
  INV_X1 \SB2_2_6/INV_1  ( .A(\RI3[2][151] ), .ZN(\SB2_2_6/i1_7 ) );
  INV_X1 \SB2_2_6/INV_0  ( .A(\RI3[2][150] ), .ZN(\SB2_2_6/i3[0] ) );
  INV_X1 \SB2_2_7/INV_5  ( .A(\RI3[2][149] ), .ZN(\SB2_2_7/i1_5 ) );
  INV_X1 \SB2_2_7/INV_4  ( .A(\RI3[2][148] ), .ZN(\SB2_2_7/i0[7] ) );
  INV_X1 \SB2_2_7/INV_3  ( .A(\RI3[2][147] ), .ZN(\SB2_2_7/i0[8] ) );
  INV_X1 \SB2_2_7/INV_1  ( .A(\RI3[2][145] ), .ZN(\SB2_2_7/i1_7 ) );
  INV_X1 \SB2_2_7/INV_0  ( .A(\RI3[2][144] ), .ZN(\SB2_2_7/i3[0] ) );
  INV_X1 \SB2_2_8/INV_5  ( .A(\RI3[2][143] ), .ZN(\SB2_2_8/i1_5 ) );
  INV_X1 \SB2_2_8/INV_4  ( .A(\RI3[2][142] ), .ZN(\SB2_2_8/i0[7] ) );
  INV_X1 \SB2_2_8/INV_3  ( .A(\RI3[2][141] ), .ZN(\SB2_2_8/i0[8] ) );
  INV_X1 \SB2_2_8/INV_2  ( .A(\RI3[2][140] ), .ZN(\SB2_2_8/i1[9] ) );
  INV_X1 \SB2_2_8/INV_1  ( .A(\RI3[2][139] ), .ZN(\SB2_2_8/i1_7 ) );
  INV_X1 \SB2_2_8/INV_0  ( .A(\RI3[2][138] ), .ZN(\SB2_2_8/i3[0] ) );
  INV_X1 \SB2_2_9/INV_5  ( .A(\RI3[2][137] ), .ZN(\SB2_2_9/i1_5 ) );
  INV_X1 \SB2_2_9/INV_4  ( .A(\RI3[2][136] ), .ZN(\SB2_2_9/i0[7] ) );
  INV_X1 \SB2_2_9/INV_3  ( .A(\RI3[2][135] ), .ZN(\SB2_2_9/i0[8] ) );
  INV_X1 \SB2_2_9/INV_2  ( .A(\RI3[2][134] ), .ZN(\SB2_2_9/i1[9] ) );
  INV_X1 \SB2_2_9/INV_1  ( .A(\RI3[2][133] ), .ZN(\SB2_2_9/i1_7 ) );
  INV_X1 \SB2_2_9/INV_0  ( .A(\RI3[2][132] ), .ZN(\SB2_2_9/i3[0] ) );
  INV_X1 \SB2_2_10/INV_5  ( .A(\RI3[2][131] ), .ZN(\SB2_2_10/i1_5 ) );
  INV_X1 \SB2_2_10/INV_4  ( .A(\RI3[2][130] ), .ZN(\SB2_2_10/i0[7] ) );
  INV_X1 \SB2_2_10/INV_3  ( .A(\RI3[2][129] ), .ZN(\SB2_2_10/i0[8] ) );
  INV_X1 \SB2_2_10/INV_2  ( .A(\RI3[2][128] ), .ZN(\SB2_2_10/i1[9] ) );
  INV_X1 \SB2_2_10/INV_1  ( .A(\RI3[2][127] ), .ZN(\SB2_2_10/i1_7 ) );
  INV_X1 \SB2_2_10/INV_0  ( .A(\RI3[2][126] ), .ZN(\SB2_2_10/i3[0] ) );
  INV_X1 \SB2_2_11/INV_5  ( .A(\RI3[2][125] ), .ZN(\SB2_2_11/i1_5 ) );
  INV_X1 \SB2_2_11/INV_4  ( .A(\RI3[2][124] ), .ZN(\SB2_2_11/i0[7] ) );
  INV_X1 \SB2_2_11/INV_3  ( .A(\RI3[2][123] ), .ZN(\SB2_2_11/i0[8] ) );
  INV_X1 \SB2_2_11/INV_2  ( .A(\RI3[2][122] ), .ZN(\SB2_2_11/i1[9] ) );
  INV_X1 \SB2_2_11/INV_1  ( .A(\RI3[2][121] ), .ZN(\SB2_2_11/i1_7 ) );
  INV_X1 \SB2_2_11/INV_0  ( .A(\RI3[2][120] ), .ZN(\SB2_2_11/i3[0] ) );
  INV_X1 \SB2_2_12/INV_5  ( .A(\RI3[2][119] ), .ZN(\SB2_2_12/i1_5 ) );
  INV_X1 \SB2_2_12/INV_4  ( .A(\RI3[2][118] ), .ZN(\SB2_2_12/i0[7] ) );
  INV_X1 \SB2_2_12/INV_3  ( .A(\RI3[2][117] ), .ZN(\SB2_2_12/i0[8] ) );
  INV_X1 \SB2_2_12/INV_2  ( .A(\RI3[2][116] ), .ZN(\SB2_2_12/i1[9] ) );
  INV_X1 \SB2_2_12/INV_1  ( .A(\RI3[2][115] ), .ZN(\SB2_2_12/i1_7 ) );
  INV_X1 \SB2_2_12/INV_0  ( .A(\RI3[2][114] ), .ZN(\SB2_2_12/i3[0] ) );
  INV_X1 \SB2_2_13/INV_5  ( .A(\RI3[2][113] ), .ZN(\SB2_2_13/i1_5 ) );
  INV_X1 \SB2_2_13/INV_4  ( .A(\RI3[2][112] ), .ZN(\SB2_2_13/i0[7] ) );
  INV_X1 \SB2_2_13/INV_3  ( .A(\RI3[2][111] ), .ZN(\SB2_2_13/i0[8] ) );
  INV_X1 \SB2_2_13/INV_2  ( .A(\RI3[2][110] ), .ZN(\SB2_2_13/i1[9] ) );
  INV_X1 \SB2_2_13/INV_1  ( .A(\RI3[2][109] ), .ZN(\SB2_2_13/i1_7 ) );
  INV_X1 \SB2_2_13/INV_0  ( .A(\RI3[2][108] ), .ZN(\SB2_2_13/i3[0] ) );
  INV_X1 \SB2_2_14/INV_5  ( .A(\RI3[2][107] ), .ZN(\SB2_2_14/i1_5 ) );
  INV_X1 \SB2_2_14/INV_4  ( .A(\RI3[2][106] ), .ZN(\SB2_2_14/i0[7] ) );
  INV_X1 \SB2_2_14/INV_3  ( .A(\RI3[2][105] ), .ZN(\SB2_2_14/i0[8] ) );
  INV_X1 \SB2_2_14/INV_2  ( .A(\RI3[2][104] ), .ZN(\SB2_2_14/i1[9] ) );
  INV_X1 \SB2_2_14/INV_1  ( .A(\RI3[2][103] ), .ZN(\SB2_2_14/i1_7 ) );
  INV_X1 \SB2_2_14/INV_0  ( .A(\RI3[2][102] ), .ZN(\SB2_2_14/i3[0] ) );
  INV_X1 \SB2_2_15/INV_5  ( .A(\RI3[2][101] ), .ZN(\SB2_2_15/i1_5 ) );
  INV_X1 \SB2_2_15/INV_4  ( .A(\RI3[2][100] ), .ZN(\SB2_2_15/i0[7] ) );
  INV_X1 \SB2_2_15/INV_3  ( .A(\RI3[2][99] ), .ZN(\SB2_2_15/i0[8] ) );
  INV_X1 \SB2_2_15/INV_2  ( .A(\RI3[2][98] ), .ZN(\SB2_2_15/i1[9] ) );
  INV_X1 \SB2_2_15/INV_1  ( .A(\RI3[2][97] ), .ZN(\SB2_2_15/i1_7 ) );
  INV_X1 \SB2_2_15/INV_0  ( .A(\RI3[2][96] ), .ZN(\SB2_2_15/i3[0] ) );
  INV_X1 \SB2_2_16/INV_5  ( .A(\RI3[2][95] ), .ZN(\SB2_2_16/i1_5 ) );
  INV_X1 \SB2_2_16/INV_4  ( .A(\RI3[2][94] ), .ZN(\SB2_2_16/i0[7] ) );
  INV_X1 \SB2_2_16/INV_3  ( .A(\RI3[2][93] ), .ZN(\SB2_2_16/i0[8] ) );
  INV_X1 \SB2_2_16/INV_2  ( .A(\RI3[2][92] ), .ZN(\SB2_2_16/i1[9] ) );
  INV_X1 \SB2_2_16/INV_1  ( .A(\RI3[2][91] ), .ZN(\SB2_2_16/i1_7 ) );
  INV_X1 \SB2_2_16/INV_0  ( .A(\RI3[2][90] ), .ZN(\SB2_2_16/i3[0] ) );
  INV_X1 \SB2_2_17/INV_5  ( .A(\RI3[2][89] ), .ZN(\SB2_2_17/i1_5 ) );
  INV_X1 \SB2_2_17/INV_4  ( .A(\RI3[2][88] ), .ZN(\SB2_2_17/i0[7] ) );
  INV_X1 \SB2_2_17/INV_3  ( .A(\RI3[2][87] ), .ZN(\SB2_2_17/i0[8] ) );
  INV_X1 \SB2_2_17/INV_2  ( .A(\RI3[2][86] ), .ZN(\SB2_2_17/i1[9] ) );
  INV_X1 \SB2_2_17/INV_1  ( .A(\RI3[2][85] ), .ZN(\SB2_2_17/i1_7 ) );
  INV_X1 \SB2_2_17/INV_0  ( .A(\RI3[2][84] ), .ZN(\SB2_2_17/i3[0] ) );
  INV_X1 \SB2_2_18/INV_5  ( .A(\RI3[2][83] ), .ZN(\SB2_2_18/i1_5 ) );
  INV_X1 \SB2_2_18/INV_4  ( .A(\RI3[2][82] ), .ZN(\SB2_2_18/i0[7] ) );
  INV_X1 \SB2_2_18/INV_3  ( .A(\RI3[2][81] ), .ZN(\SB2_2_18/i0[8] ) );
  INV_X1 \SB2_2_18/INV_2  ( .A(\RI3[2][80] ), .ZN(\SB2_2_18/i1[9] ) );
  INV_X1 \SB2_2_18/INV_1  ( .A(\RI3[2][79] ), .ZN(\SB2_2_18/i1_7 ) );
  INV_X1 \SB2_2_18/INV_0  ( .A(\RI3[2][78] ), .ZN(\SB2_2_18/i3[0] ) );
  INV_X1 \SB2_2_19/INV_5  ( .A(\RI3[2][77] ), .ZN(\SB2_2_19/i1_5 ) );
  INV_X1 \SB2_2_19/INV_4  ( .A(\RI3[2][76] ), .ZN(\SB2_2_19/i0[7] ) );
  INV_X1 \SB2_2_19/INV_3  ( .A(\RI3[2][75] ), .ZN(\SB2_2_19/i0[8] ) );
  INV_X1 \SB2_2_19/INV_2  ( .A(\RI3[2][74] ), .ZN(\SB2_2_19/i1[9] ) );
  INV_X1 \SB2_2_19/INV_1  ( .A(\RI3[2][73] ), .ZN(\SB2_2_19/i1_7 ) );
  INV_X1 \SB2_2_19/INV_0  ( .A(\RI3[2][72] ), .ZN(\SB2_2_19/i3[0] ) );
  INV_X1 \SB2_2_20/INV_5  ( .A(\RI3[2][71] ), .ZN(\SB2_2_20/i1_5 ) );
  INV_X1 \SB2_2_20/INV_4  ( .A(\RI3[2][70] ), .ZN(\SB2_2_20/i0[7] ) );
  INV_X1 \SB2_2_20/INV_3  ( .A(\RI3[2][69] ), .ZN(\SB2_2_20/i0[8] ) );
  INV_X1 \SB2_2_20/INV_2  ( .A(\RI3[2][68] ), .ZN(\SB2_2_20/i1[9] ) );
  INV_X1 \SB2_2_20/INV_1  ( .A(\RI3[2][67] ), .ZN(\SB2_2_20/i1_7 ) );
  INV_X1 \SB2_2_20/INV_0  ( .A(\RI3[2][66] ), .ZN(\SB2_2_20/i3[0] ) );
  INV_X1 \SB2_2_21/INV_5  ( .A(\RI3[2][65] ), .ZN(\SB2_2_21/i1_5 ) );
  INV_X1 \SB2_2_21/INV_4  ( .A(\RI3[2][64] ), .ZN(\SB2_2_21/i0[7] ) );
  INV_X1 \SB2_2_21/INV_3  ( .A(\RI3[2][63] ), .ZN(\SB2_2_21/i0[8] ) );
  INV_X1 \SB2_2_21/INV_2  ( .A(\RI3[2][62] ), .ZN(\SB2_2_21/i1[9] ) );
  INV_X1 \SB2_2_21/INV_1  ( .A(\RI3[2][61] ), .ZN(\SB2_2_21/i1_7 ) );
  INV_X1 \SB2_2_21/INV_0  ( .A(\RI3[2][60] ), .ZN(\SB2_2_21/i3[0] ) );
  INV_X1 \SB2_2_22/INV_5  ( .A(\RI3[2][59] ), .ZN(\SB2_2_22/i1_5 ) );
  INV_X1 \SB2_2_22/INV_4  ( .A(\RI3[2][58] ), .ZN(\SB2_2_22/i0[7] ) );
  INV_X1 \SB2_2_22/INV_3  ( .A(\RI3[2][57] ), .ZN(\SB2_2_22/i0[8] ) );
  INV_X1 \SB2_2_22/INV_1  ( .A(\RI3[2][55] ), .ZN(\SB2_2_22/i1_7 ) );
  INV_X1 \SB2_2_22/INV_0  ( .A(\RI3[2][54] ), .ZN(\SB2_2_22/i3[0] ) );
  INV_X1 \SB2_2_23/INV_5  ( .A(\RI3[2][53] ), .ZN(\SB2_2_23/i1_5 ) );
  INV_X1 \SB2_2_23/INV_4  ( .A(\RI3[2][52] ), .ZN(\SB2_2_23/i0[7] ) );
  INV_X1 \SB2_2_23/INV_3  ( .A(\RI3[2][51] ), .ZN(\SB2_2_23/i0[8] ) );
  INV_X1 \SB2_2_23/INV_2  ( .A(\RI3[2][50] ), .ZN(\SB2_2_23/i1[9] ) );
  INV_X1 \SB2_2_23/INV_1  ( .A(\RI3[2][49] ), .ZN(\SB2_2_23/i1_7 ) );
  INV_X1 \SB2_2_23/INV_0  ( .A(\RI3[2][48] ), .ZN(\SB2_2_23/i3[0] ) );
  INV_X1 \SB2_2_24/INV_5  ( .A(\RI3[2][47] ), .ZN(\SB2_2_24/i1_5 ) );
  INV_X1 \SB2_2_24/INV_4  ( .A(\RI3[2][46] ), .ZN(\SB2_2_24/i0[7] ) );
  INV_X1 \SB2_2_24/INV_3  ( .A(\RI3[2][45] ), .ZN(\SB2_2_24/i0[8] ) );
  INV_X1 \SB2_2_24/INV_2  ( .A(\RI3[2][44] ), .ZN(\SB2_2_24/i1[9] ) );
  INV_X1 \SB2_2_24/INV_1  ( .A(\RI3[2][43] ), .ZN(\SB2_2_24/i1_7 ) );
  INV_X1 \SB2_2_24/INV_0  ( .A(\RI3[2][42] ), .ZN(\SB2_2_24/i3[0] ) );
  INV_X1 \SB2_2_25/INV_5  ( .A(\RI3[2][41] ), .ZN(\SB2_2_25/i1_5 ) );
  INV_X1 \SB2_2_25/INV_4  ( .A(\RI3[2][40] ), .ZN(\SB2_2_25/i0[7] ) );
  INV_X1 \SB2_2_25/INV_3  ( .A(\RI3[2][39] ), .ZN(\SB2_2_25/i0[8] ) );
  INV_X1 \SB2_2_25/INV_2  ( .A(\RI3[2][38] ), .ZN(\SB2_2_25/i1[9] ) );
  INV_X1 \SB2_2_25/INV_1  ( .A(\RI3[2][37] ), .ZN(\SB2_2_25/i1_7 ) );
  INV_X1 \SB2_2_25/INV_0  ( .A(\RI3[2][36] ), .ZN(\SB2_2_25/i3[0] ) );
  INV_X1 \SB2_2_26/INV_5  ( .A(\RI3[2][35] ), .ZN(\SB2_2_26/i1_5 ) );
  INV_X1 \SB2_2_26/INV_4  ( .A(\RI3[2][34] ), .ZN(\SB2_2_26/i0[7] ) );
  INV_X1 \SB2_2_26/INV_3  ( .A(\RI3[2][33] ), .ZN(\SB2_2_26/i0[8] ) );
  INV_X1 \SB2_2_26/INV_2  ( .A(\RI3[2][32] ), .ZN(\SB2_2_26/i1[9] ) );
  INV_X1 \SB2_2_26/INV_1  ( .A(\RI3[2][31] ), .ZN(\SB2_2_26/i1_7 ) );
  INV_X1 \SB2_2_26/INV_0  ( .A(\RI3[2][30] ), .ZN(\SB2_2_26/i3[0] ) );
  INV_X1 \SB2_2_27/INV_5  ( .A(\RI3[2][29] ), .ZN(\SB2_2_27/i1_5 ) );
  INV_X1 \SB2_2_27/INV_4  ( .A(\RI3[2][28] ), .ZN(\SB2_2_27/i0[7] ) );
  INV_X1 \SB2_2_27/INV_2  ( .A(\RI3[2][26] ), .ZN(\SB2_2_27/i1[9] ) );
  INV_X1 \SB2_2_27/INV_1  ( .A(\RI3[2][25] ), .ZN(\SB2_2_27/i1_7 ) );
  INV_X1 \SB2_2_27/INV_0  ( .A(\RI3[2][24] ), .ZN(\SB2_2_27/i3[0] ) );
  INV_X1 \SB2_2_28/INV_5  ( .A(\RI3[2][23] ), .ZN(\SB2_2_28/i1_5 ) );
  INV_X1 \SB2_2_28/INV_4  ( .A(\RI3[2][22] ), .ZN(\SB2_2_28/i0[7] ) );
  INV_X1 \SB2_2_28/INV_3  ( .A(\RI3[2][21] ), .ZN(\SB2_2_28/i0[8] ) );
  INV_X1 \SB2_2_28/INV_1  ( .A(\RI3[2][19] ), .ZN(\SB2_2_28/i1_7 ) );
  INV_X1 \SB2_2_28/INV_0  ( .A(\RI3[2][18] ), .ZN(\SB2_2_28/i3[0] ) );
  INV_X1 \SB2_2_29/INV_5  ( .A(\RI3[2][17] ), .ZN(\SB2_2_29/i1_5 ) );
  INV_X1 \SB2_2_29/INV_4  ( .A(\RI3[2][16] ), .ZN(\SB2_2_29/i0[7] ) );
  INV_X1 \SB2_2_29/INV_3  ( .A(\RI3[2][15] ), .ZN(\SB2_2_29/i0[8] ) );
  INV_X1 \SB2_2_29/INV_2  ( .A(\RI3[2][14] ), .ZN(\SB2_2_29/i1[9] ) );
  INV_X1 \SB2_2_29/INV_1  ( .A(\RI3[2][13] ), .ZN(\SB2_2_29/i1_7 ) );
  INV_X1 \SB2_2_29/INV_0  ( .A(\RI3[2][12] ), .ZN(\SB2_2_29/i3[0] ) );
  INV_X1 \SB2_2_30/INV_5  ( .A(\RI3[2][11] ), .ZN(\SB2_2_30/i1_5 ) );
  INV_X1 \SB2_2_30/INV_4  ( .A(\RI3[2][10] ), .ZN(\SB2_2_30/i0[7] ) );
  INV_X1 \SB2_2_30/INV_3  ( .A(\RI3[2][9] ), .ZN(\SB2_2_30/i0[8] ) );
  INV_X1 \SB2_2_30/INV_1  ( .A(\RI3[2][7] ), .ZN(\SB2_2_30/i1_7 ) );
  INV_X1 \SB2_2_30/INV_0  ( .A(\RI3[2][6] ), .ZN(\SB2_2_30/i3[0] ) );
  INV_X1 \SB2_2_31/INV_5  ( .A(\RI3[2][5] ), .ZN(\SB2_2_31/i1_5 ) );
  INV_X1 \SB2_2_31/INV_4  ( .A(\RI3[2][4] ), .ZN(\SB2_2_31/i0[7] ) );
  INV_X1 \SB2_2_31/INV_3  ( .A(\RI3[2][3] ), .ZN(\SB2_2_31/i0[8] ) );
  INV_X1 \SB2_2_31/INV_2  ( .A(\RI3[2][2] ), .ZN(\SB2_2_31/i1[9] ) );
  INV_X1 \SB2_2_31/INV_1  ( .A(\RI3[2][1] ), .ZN(\SB2_2_31/i1_7 ) );
  INV_X1 \SB2_2_31/INV_0  ( .A(\RI3[2][0] ), .ZN(\SB2_2_31/i3[0] ) );
  INV_X1 \SB2_3_0/INV_5  ( .A(\RI3[3][191] ), .ZN(\SB2_3_0/i1_5 ) );
  INV_X1 \SB2_3_0/INV_4  ( .A(\RI3[3][190] ), .ZN(\SB2_3_0/i0[7] ) );
  INV_X1 \SB2_3_0/INV_3  ( .A(\RI3[3][189] ), .ZN(\SB2_3_0/i0[8] ) );
  INV_X1 \SB2_3_0/INV_2  ( .A(\RI3[3][188] ), .ZN(\SB2_3_0/i1[9] ) );
  INV_X1 \SB2_3_0/INV_1  ( .A(\RI3[3][187] ), .ZN(\SB2_3_0/i1_7 ) );
  INV_X1 \SB2_3_0/INV_0  ( .A(\RI3[3][186] ), .ZN(\SB2_3_0/i3[0] ) );
  BUF_X1 \SB2_3_0/BUF_0  ( .A(\RI3[3][186] ), .Z(\SB2_3_0/i0[9] ) );
  INV_X1 \SB2_3_1/INV_5  ( .A(\RI3[3][185] ), .ZN(\SB2_3_1/i1_5 ) );
  INV_X1 \SB2_3_1/INV_4  ( .A(\RI3[3][184] ), .ZN(\SB2_3_1/i0[7] ) );
  INV_X1 \SB2_3_1/INV_3  ( .A(\RI3[3][183] ), .ZN(\SB2_3_1/i0[8] ) );
  INV_X1 \SB2_3_1/INV_2  ( .A(\RI3[3][182] ), .ZN(\SB2_3_1/i1[9] ) );
  INV_X1 \SB2_3_1/INV_1  ( .A(\RI3[3][181] ), .ZN(\SB2_3_1/i1_7 ) );
  INV_X1 \SB2_3_1/INV_0  ( .A(\RI3[3][180] ), .ZN(\SB2_3_1/i3[0] ) );
  INV_X1 \SB2_3_2/INV_5  ( .A(\RI3[3][179] ), .ZN(\SB2_3_2/i1_5 ) );
  INV_X1 \SB2_3_2/INV_4  ( .A(\RI3[3][178] ), .ZN(\SB2_3_2/i0[7] ) );
  INV_X1 \SB2_3_2/INV_3  ( .A(\RI3[3][177] ), .ZN(\SB2_3_2/i0[8] ) );
  INV_X1 \SB2_3_2/INV_2  ( .A(\RI3[3][176] ), .ZN(\SB2_3_2/i1[9] ) );
  INV_X1 \SB2_3_2/INV_1  ( .A(\RI3[3][175] ), .ZN(\SB2_3_2/i1_7 ) );
  INV_X1 \SB2_3_2/INV_0  ( .A(\RI3[3][174] ), .ZN(\SB2_3_2/i3[0] ) );
  INV_X1 \SB2_3_3/INV_5  ( .A(\RI3[3][173] ), .ZN(\SB2_3_3/i1_5 ) );
  INV_X1 \SB2_3_3/INV_4  ( .A(\RI3[3][172] ), .ZN(\SB2_3_3/i0[7] ) );
  INV_X1 \SB2_3_3/INV_3  ( .A(\RI3[3][171] ), .ZN(\SB2_3_3/i0[8] ) );
  INV_X1 \SB2_3_3/INV_2  ( .A(\RI3[3][170] ), .ZN(\SB2_3_3/i1[9] ) );
  INV_X1 \SB2_3_3/INV_1  ( .A(\RI3[3][169] ), .ZN(\SB2_3_3/i1_7 ) );
  INV_X1 \SB2_3_3/INV_0  ( .A(\RI3[3][168] ), .ZN(\SB2_3_3/i3[0] ) );
  INV_X1 \SB2_3_4/INV_5  ( .A(\RI3[3][167] ), .ZN(\SB2_3_4/i1_5 ) );
  INV_X1 \SB2_3_4/INV_4  ( .A(\SB2_3_4/i0_4 ), .ZN(\SB2_3_4/i0[7] ) );
  INV_X1 \SB2_3_4/INV_3  ( .A(\RI3[3][165] ), .ZN(\SB2_3_4/i0[8] ) );
  INV_X1 \SB2_3_4/INV_1  ( .A(\RI3[3][163] ), .ZN(\SB2_3_4/i1_7 ) );
  INV_X1 \SB2_3_4/INV_0  ( .A(\RI3[3][162] ), .ZN(\SB2_3_4/i3[0] ) );
  INV_X1 \SB2_3_5/INV_5  ( .A(\RI3[3][161] ), .ZN(\SB2_3_5/i1_5 ) );
  INV_X1 \SB2_3_5/INV_4  ( .A(\SB2_3_5/i0_4 ), .ZN(\SB2_3_5/i0[7] ) );
  INV_X1 \SB2_3_5/INV_3  ( .A(\RI3[3][159] ), .ZN(\SB2_3_5/i0[8] ) );
  INV_X1 \SB2_3_5/INV_2  ( .A(\RI3[3][158] ), .ZN(\SB2_3_5/i1[9] ) );
  INV_X1 \SB2_3_5/INV_1  ( .A(\RI3[3][157] ), .ZN(\SB2_3_5/i1_7 ) );
  INV_X1 \SB2_3_5/INV_0  ( .A(\RI3[3][156] ), .ZN(\SB2_3_5/i3[0] ) );
  INV_X1 \SB2_3_6/INV_5  ( .A(\RI3[3][155] ), .ZN(\SB2_3_6/i1_5 ) );
  INV_X1 \SB2_3_6/INV_4  ( .A(\RI3[3][154] ), .ZN(\SB2_3_6/i0[7] ) );
  INV_X1 \SB2_3_6/INV_3  ( .A(\RI3[3][153] ), .ZN(\SB2_3_6/i0[8] ) );
  INV_X1 \SB2_3_6/INV_1  ( .A(\RI3[3][151] ), .ZN(\SB2_3_6/i1_7 ) );
  INV_X1 \SB2_3_6/INV_0  ( .A(\RI3[3][150] ), .ZN(\SB2_3_6/i3[0] ) );
  BUF_X1 \SB2_3_6/BUF_0  ( .A(\RI3[3][150] ), .Z(\SB2_3_6/i0[9] ) );
  INV_X1 \SB2_3_7/INV_5  ( .A(\RI3[3][149] ), .ZN(\SB2_3_7/i1_5 ) );
  INV_X1 \SB2_3_7/INV_4  ( .A(\RI3[3][148] ), .ZN(\SB2_3_7/i0[7] ) );
  INV_X1 \SB2_3_7/INV_3  ( .A(\RI3[3][147] ), .ZN(\SB2_3_7/i0[8] ) );
  INV_X1 \SB2_3_7/INV_1  ( .A(\RI3[3][145] ), .ZN(\SB2_3_7/i1_7 ) );
  INV_X1 \SB2_3_7/INV_0  ( .A(\RI3[3][144] ), .ZN(\SB2_3_7/i3[0] ) );
  INV_X1 \SB2_3_8/INV_5  ( .A(\RI3[3][143] ), .ZN(\SB2_3_8/i1_5 ) );
  INV_X1 \SB2_3_8/INV_4  ( .A(\SB2_3_8/i0_4 ), .ZN(\SB2_3_8/i0[7] ) );
  INV_X1 \SB2_3_8/INV_3  ( .A(\RI3[3][141] ), .ZN(\SB2_3_8/i0[8] ) );
  INV_X1 \SB2_3_8/INV_2  ( .A(\RI3[3][140] ), .ZN(\SB2_3_8/i1[9] ) );
  INV_X1 \SB2_3_8/INV_1  ( .A(\RI3[3][139] ), .ZN(\SB2_3_8/i1_7 ) );
  INV_X1 \SB2_3_8/INV_0  ( .A(\RI3[3][138] ), .ZN(\SB2_3_8/i3[0] ) );
  INV_X1 \SB2_3_9/INV_5  ( .A(\RI3[3][137] ), .ZN(\SB2_3_9/i1_5 ) );
  INV_X1 \SB2_3_9/INV_4  ( .A(\RI3[3][136] ), .ZN(\SB2_3_9/i0[7] ) );
  INV_X1 \SB2_3_9/INV_3  ( .A(\RI3[3][135] ), .ZN(\SB2_3_9/i0[8] ) );
  INV_X1 \SB2_3_9/INV_1  ( .A(\RI3[3][133] ), .ZN(\SB2_3_9/i1_7 ) );
  INV_X1 \SB2_3_9/INV_0  ( .A(\RI3[3][132] ), .ZN(\SB2_3_9/i3[0] ) );
  INV_X1 \SB2_3_10/INV_5  ( .A(\RI3[3][131] ), .ZN(\SB2_3_10/i1_5 ) );
  INV_X1 \SB2_3_10/INV_4  ( .A(\RI3[3][130] ), .ZN(\SB2_3_10/i0[7] ) );
  INV_X1 \SB2_3_10/INV_3  ( .A(\RI3[3][129] ), .ZN(\SB2_3_10/i0[8] ) );
  INV_X1 \SB2_3_10/INV_2  ( .A(\RI3[3][128] ), .ZN(\SB2_3_10/i1[9] ) );
  INV_X1 \SB2_3_10/INV_1  ( .A(\RI3[3][127] ), .ZN(\SB2_3_10/i1_7 ) );
  INV_X1 \SB2_3_10/INV_0  ( .A(\RI3[3][126] ), .ZN(\SB2_3_10/i3[0] ) );
  BUF_X1 \SB2_3_10/BUF_1  ( .A(\RI3[3][127] ), .Z(\SB2_3_10/i0[6] ) );
  INV_X1 \SB2_3_11/INV_5  ( .A(\RI3[3][125] ), .ZN(\SB2_3_11/i1_5 ) );
  INV_X1 \SB2_3_11/INV_4  ( .A(\RI3[3][124] ), .ZN(\SB2_3_11/i0[7] ) );
  INV_X1 \SB2_3_11/INV_3  ( .A(\RI3[3][123] ), .ZN(\SB2_3_11/i0[8] ) );
  INV_X1 \SB2_3_11/INV_2  ( .A(\RI3[3][122] ), .ZN(\SB2_3_11/i1[9] ) );
  INV_X1 \SB2_3_11/INV_1  ( .A(\RI3[3][121] ), .ZN(\SB2_3_11/i1_7 ) );
  INV_X1 \SB2_3_11/INV_0  ( .A(\RI3[3][120] ), .ZN(\SB2_3_11/i3[0] ) );
  INV_X1 \SB2_3_12/INV_5  ( .A(\RI3[3][119] ), .ZN(\SB2_3_12/i1_5 ) );
  INV_X1 \SB2_3_12/INV_4  ( .A(\RI3[3][118] ), .ZN(\SB2_3_12/i0[7] ) );
  INV_X1 \SB2_3_12/INV_3  ( .A(\RI3[3][117] ), .ZN(\SB2_3_12/i0[8] ) );
  INV_X1 \SB2_3_12/INV_2  ( .A(\RI3[3][116] ), .ZN(\SB2_3_12/i1[9] ) );
  INV_X1 \SB2_3_12/INV_1  ( .A(\RI3[3][115] ), .ZN(\SB2_3_12/i1_7 ) );
  INV_X1 \SB2_3_12/INV_0  ( .A(\RI3[3][114] ), .ZN(\SB2_3_12/i3[0] ) );
  BUF_X1 \SB2_3_12/BUF_0  ( .A(\RI3[3][114] ), .Z(\SB2_3_12/i0[9] ) );
  INV_X1 \SB2_3_13/INV_5  ( .A(\RI3[3][113] ), .ZN(\SB2_3_13/i1_5 ) );
  INV_X1 \SB2_3_13/INV_4  ( .A(\SB2_3_13/i0_4 ), .ZN(\SB2_3_13/i0[7] ) );
  INV_X1 \SB2_3_13/INV_3  ( .A(\RI3[3][111] ), .ZN(\SB2_3_13/i0[8] ) );
  INV_X1 \SB2_3_13/INV_1  ( .A(\RI3[3][109] ), .ZN(\SB2_3_13/i1_7 ) );
  INV_X1 \SB2_3_13/INV_0  ( .A(\RI3[3][108] ), .ZN(\SB2_3_13/i3[0] ) );
  INV_X1 \SB2_3_14/INV_5  ( .A(\RI3[3][107] ), .ZN(\SB2_3_14/i1_5 ) );
  INV_X1 \SB2_3_14/INV_4  ( .A(\RI3[3][106] ), .ZN(\SB2_3_14/i0[7] ) );
  INV_X1 \SB2_3_14/INV_3  ( .A(\RI3[3][105] ), .ZN(\SB2_3_14/i0[8] ) );
  INV_X1 \SB2_3_14/INV_2  ( .A(\RI3[3][104] ), .ZN(\SB2_3_14/i1[9] ) );
  INV_X1 \SB2_3_14/INV_1  ( .A(\RI3[3][103] ), .ZN(\SB2_3_14/i1_7 ) );
  INV_X1 \SB2_3_14/INV_0  ( .A(\RI3[3][102] ), .ZN(\SB2_3_14/i3[0] ) );
  BUF_X1 \SB2_3_14/BUF_1  ( .A(\RI3[3][103] ), .Z(\SB2_3_14/i0[6] ) );
  INV_X1 \SB2_3_15/INV_5  ( .A(\RI3[3][101] ), .ZN(\SB2_3_15/i1_5 ) );
  INV_X1 \SB2_3_15/INV_4  ( .A(\SB2_3_15/i0_4 ), .ZN(\SB2_3_15/i0[7] ) );
  INV_X1 \SB2_3_15/INV_3  ( .A(\RI3[3][99] ), .ZN(\SB2_3_15/i0[8] ) );
  INV_X1 \SB2_3_15/INV_2  ( .A(\RI3[3][98] ), .ZN(\SB2_3_15/i1[9] ) );
  INV_X1 \SB2_3_15/INV_0  ( .A(\RI3[3][96] ), .ZN(\SB2_3_15/i3[0] ) );
  INV_X1 \SB2_3_16/INV_5  ( .A(\RI3[3][95] ), .ZN(\SB2_3_16/i1_5 ) );
  INV_X1 \SB2_3_16/INV_3  ( .A(\RI3[3][93] ), .ZN(\SB2_3_16/i0[8] ) );
  INV_X1 \SB2_3_16/INV_2  ( .A(\RI3[3][92] ), .ZN(\SB2_3_16/i1[9] ) );
  INV_X1 \SB2_3_16/INV_1  ( .A(\RI3[3][91] ), .ZN(\SB2_3_16/i1_7 ) );
  INV_X1 \SB2_3_16/INV_0  ( .A(\RI3[3][90] ), .ZN(\SB2_3_16/i3[0] ) );
  INV_X1 \SB2_3_17/INV_5  ( .A(\RI3[3][89] ), .ZN(\SB2_3_17/i1_5 ) );
  INV_X1 \SB2_3_17/INV_4  ( .A(\RI3[3][88] ), .ZN(\SB2_3_17/i0[7] ) );
  INV_X1 \SB2_3_17/INV_3  ( .A(\RI3[3][87] ), .ZN(\SB2_3_17/i0[8] ) );
  INV_X1 \SB2_3_17/INV_1  ( .A(\RI3[3][85] ), .ZN(\SB2_3_17/i1_7 ) );
  INV_X1 \SB2_3_17/INV_0  ( .A(\RI3[3][84] ), .ZN(\SB2_3_17/i3[0] ) );
  BUF_X1 \SB2_3_17/BUF_0  ( .A(\RI3[3][84] ), .Z(\SB2_3_17/i0[9] ) );
  INV_X1 \SB2_3_18/INV_5  ( .A(\RI3[3][83] ), .ZN(\SB2_3_18/i1_5 ) );
  INV_X1 \SB2_3_18/INV_4  ( .A(\SB2_3_18/i0_4 ), .ZN(\SB2_3_18/i0[7] ) );
  INV_X1 \SB2_3_18/INV_3  ( .A(\RI3[3][81] ), .ZN(\SB2_3_18/i0[8] ) );
  INV_X1 \SB2_3_18/INV_2  ( .A(\RI3[3][80] ), .ZN(\SB2_3_18/i1[9] ) );
  INV_X1 \SB2_3_18/INV_1  ( .A(\RI3[3][79] ), .ZN(\SB2_3_18/i1_7 ) );
  INV_X1 \SB2_3_18/INV_0  ( .A(\RI3[3][78] ), .ZN(\SB2_3_18/i3[0] ) );
  BUF_X1 \SB2_3_18/BUF_0  ( .A(\RI3[3][78] ), .Z(\SB2_3_18/i0[9] ) );
  INV_X1 \SB2_3_19/INV_5  ( .A(\RI3[3][77] ), .ZN(\SB2_3_19/i1_5 ) );
  INV_X1 \SB2_3_19/INV_4  ( .A(\RI3[3][76] ), .ZN(\SB2_3_19/i0[7] ) );
  INV_X1 \SB2_3_19/INV_3  ( .A(\RI3[3][75] ), .ZN(\SB2_3_19/i0[8] ) );
  INV_X1 \SB2_3_19/INV_2  ( .A(\RI3[3][74] ), .ZN(\SB2_3_19/i1[9] ) );
  INV_X1 \SB2_3_19/INV_1  ( .A(\RI3[3][73] ), .ZN(\SB2_3_19/i1_7 ) );
  INV_X1 \SB2_3_19/INV_0  ( .A(\RI3[3][72] ), .ZN(\SB2_3_19/i3[0] ) );
  INV_X1 \SB2_3_20/INV_5  ( .A(\RI3[3][71] ), .ZN(\SB2_3_20/i1_5 ) );
  INV_X1 \SB2_3_20/INV_4  ( .A(\SB2_3_20/i0_4 ), .ZN(\SB2_3_20/i0[7] ) );
  INV_X1 \SB2_3_20/INV_3  ( .A(\RI3[3][69] ), .ZN(\SB2_3_20/i0[8] ) );
  INV_X1 \SB2_3_20/INV_2  ( .A(\RI3[3][68] ), .ZN(\SB2_3_20/i1[9] ) );
  INV_X1 \SB2_3_20/INV_1  ( .A(\RI3[3][67] ), .ZN(\SB2_3_20/i1_7 ) );
  INV_X1 \SB2_3_20/INV_0  ( .A(\RI3[3][66] ), .ZN(\SB2_3_20/i3[0] ) );
  INV_X1 \SB2_3_21/INV_5  ( .A(\RI3[3][65] ), .ZN(\SB2_3_21/i1_5 ) );
  INV_X1 \SB2_3_21/INV_4  ( .A(\RI3[3][64] ), .ZN(\SB2_3_21/i0[7] ) );
  INV_X1 \SB2_3_21/INV_3  ( .A(\RI3[3][63] ), .ZN(\SB2_3_21/i0[8] ) );
  INV_X1 \SB2_3_21/INV_1  ( .A(\RI3[3][61] ), .ZN(\SB2_3_21/i1_7 ) );
  INV_X1 \SB2_3_21/INV_0  ( .A(\RI3[3][60] ), .ZN(\SB2_3_21/i3[0] ) );
  INV_X1 \SB2_3_22/INV_5  ( .A(\RI3[3][59] ), .ZN(\SB2_3_22/i1_5 ) );
  INV_X1 \SB2_3_22/INV_4  ( .A(\SB2_3_22/i0_4 ), .ZN(\SB2_3_22/i0[7] ) );
  INV_X1 \SB2_3_22/INV_3  ( .A(\RI3[3][57] ), .ZN(\SB2_3_22/i0[8] ) );
  INV_X1 \SB2_3_22/INV_2  ( .A(\RI3[3][56] ), .ZN(\SB2_3_22/i1[9] ) );
  INV_X1 \SB2_3_22/INV_1  ( .A(\RI3[3][55] ), .ZN(\SB2_3_22/i1_7 ) );
  INV_X1 \SB2_3_22/INV_0  ( .A(\RI3[3][54] ), .ZN(\SB2_3_22/i3[0] ) );
  INV_X1 \SB2_3_23/INV_5  ( .A(\RI3[3][53] ), .ZN(\SB2_3_23/i1_5 ) );
  INV_X1 \SB2_3_23/INV_4  ( .A(\SB2_3_23/i0_4 ), .ZN(\SB2_3_23/i0[7] ) );
  INV_X1 \SB2_3_23/INV_3  ( .A(\RI3[3][51] ), .ZN(\SB2_3_23/i0[8] ) );
  INV_X1 \SB2_3_23/INV_2  ( .A(\RI3[3][50] ), .ZN(\SB2_3_23/i1[9] ) );
  INV_X1 \SB2_3_23/INV_1  ( .A(\RI3[3][49] ), .ZN(\SB2_3_23/i1_7 ) );
  INV_X1 \SB2_3_23/INV_0  ( .A(\RI3[3][48] ), .ZN(\SB2_3_23/i3[0] ) );
  INV_X1 \SB2_3_24/INV_5  ( .A(\RI3[3][47] ), .ZN(\SB2_3_24/i1_5 ) );
  INV_X1 \SB2_3_24/INV_4  ( .A(\RI3[3][46] ), .ZN(\SB2_3_24/i0[7] ) );
  INV_X1 \SB2_3_24/INV_3  ( .A(\RI3[3][45] ), .ZN(\SB2_3_24/i0[8] ) );
  INV_X1 \SB2_3_24/INV_2  ( .A(\RI3[3][44] ), .ZN(\SB2_3_24/i1[9] ) );
  INV_X1 \SB2_3_24/INV_1  ( .A(\RI3[3][43] ), .ZN(\SB2_3_24/i1_7 ) );
  INV_X1 \SB2_3_24/INV_0  ( .A(\RI3[3][42] ), .ZN(\SB2_3_24/i3[0] ) );
  INV_X1 \SB2_3_25/INV_5  ( .A(\RI3[3][41] ), .ZN(\SB2_3_25/i1_5 ) );
  INV_X1 \SB2_3_25/INV_4  ( .A(\SB2_3_25/i0_4 ), .ZN(\SB2_3_25/i0[7] ) );
  INV_X1 \SB2_3_25/INV_3  ( .A(\RI3[3][39] ), .ZN(\SB2_3_25/i0[8] ) );
  INV_X1 \SB2_3_25/INV_1  ( .A(\RI3[3][37] ), .ZN(\SB2_3_25/i1_7 ) );
  INV_X1 \SB2_3_25/INV_0  ( .A(\RI3[3][36] ), .ZN(\SB2_3_25/i3[0] ) );
  INV_X1 \SB2_3_26/INV_5  ( .A(\RI3[3][35] ), .ZN(\SB2_3_26/i1_5 ) );
  INV_X1 \SB2_3_26/INV_4  ( .A(\SB2_3_26/i0_4 ), .ZN(\SB2_3_26/i0[7] ) );
  INV_X1 \SB2_3_26/INV_3  ( .A(\RI3[3][33] ), .ZN(\SB2_3_26/i0[8] ) );
  INV_X1 \SB2_3_26/INV_2  ( .A(\RI3[3][32] ), .ZN(\SB2_3_26/i1[9] ) );
  INV_X1 \SB2_3_26/INV_1  ( .A(\RI3[3][31] ), .ZN(\SB2_3_26/i1_7 ) );
  INV_X1 \SB2_3_26/INV_0  ( .A(\RI3[3][30] ), .ZN(\SB2_3_26/i3[0] ) );
  INV_X1 \SB2_3_27/INV_4  ( .A(\RI3[3][28] ), .ZN(\SB2_3_27/i0[7] ) );
  INV_X1 \SB2_3_27/INV_3  ( .A(\RI3[3][27] ), .ZN(\SB2_3_27/i0[8] ) );
  INV_X1 \SB2_3_27/INV_2  ( .A(\RI3[3][26] ), .ZN(\SB2_3_27/i1[9] ) );
  INV_X1 \SB2_3_27/INV_1  ( .A(\RI3[3][25] ), .ZN(\SB2_3_27/i1_7 ) );
  INV_X1 \SB2_3_27/INV_0  ( .A(\RI3[3][24] ), .ZN(\SB2_3_27/i3[0] ) );
  INV_X1 \SB2_3_28/INV_5  ( .A(\RI3[3][23] ), .ZN(\SB2_3_28/i1_5 ) );
  INV_X1 \SB2_3_28/INV_4  ( .A(\SB2_3_28/i0_4 ), .ZN(\SB2_3_28/i0[7] ) );
  INV_X1 \SB2_3_28/INV_3  ( .A(\RI3[3][21] ), .ZN(\SB2_3_28/i0[8] ) );
  INV_X1 \SB2_3_28/INV_2  ( .A(\RI3[3][20] ), .ZN(\SB2_3_28/i1[9] ) );
  INV_X1 \SB2_3_28/INV_1  ( .A(\RI3[3][19] ), .ZN(\SB2_3_28/i1_7 ) );
  INV_X1 \SB2_3_28/INV_0  ( .A(\RI3[3][18] ), .ZN(\SB2_3_28/i3[0] ) );
  INV_X1 \SB2_3_29/INV_5  ( .A(\RI3[3][17] ), .ZN(\SB2_3_29/i1_5 ) );
  INV_X1 \SB2_3_29/INV_4  ( .A(\RI3[3][16] ), .ZN(\SB2_3_29/i0[7] ) );
  INV_X1 \SB2_3_29/INV_3  ( .A(\RI3[3][15] ), .ZN(\SB2_3_29/i0[8] ) );
  INV_X1 \SB2_3_29/INV_2  ( .A(\RI3[3][14] ), .ZN(\SB2_3_29/i1[9] ) );
  INV_X1 \SB2_3_29/INV_1  ( .A(\RI3[3][13] ), .ZN(\SB2_3_29/i1_7 ) );
  INV_X1 \SB2_3_29/INV_0  ( .A(\RI3[3][12] ), .ZN(\SB2_3_29/i3[0] ) );
  INV_X1 \SB2_3_30/INV_5  ( .A(\RI3[3][11] ), .ZN(\SB2_3_30/i1_5 ) );
  INV_X1 \SB2_3_30/INV_4  ( .A(\RI3[3][10] ), .ZN(\SB2_3_30/i0[7] ) );
  INV_X1 \SB2_3_30/INV_3  ( .A(\RI3[3][9] ), .ZN(\SB2_3_30/i0[8] ) );
  INV_X1 \SB2_3_30/INV_2  ( .A(\RI3[3][8] ), .ZN(\SB2_3_30/i1[9] ) );
  INV_X1 \SB2_3_30/INV_1  ( .A(\RI3[3][7] ), .ZN(\SB2_3_30/i1_7 ) );
  INV_X1 \SB2_3_30/INV_0  ( .A(\RI3[3][6] ), .ZN(\SB2_3_30/i3[0] ) );
  INV_X1 \SB2_3_31/INV_5  ( .A(\RI3[3][5] ), .ZN(\SB2_3_31/i1_5 ) );
  INV_X1 \SB2_3_31/INV_3  ( .A(\RI3[3][3] ), .ZN(\SB2_3_31/i0[8] ) );
  INV_X1 \SB2_3_31/INV_1  ( .A(\RI3[3][1] ), .ZN(\SB2_3_31/i1_7 ) );
  INV_X1 \SB2_3_31/INV_0  ( .A(\RI3[3][0] ), .ZN(\SB2_3_31/i3[0] ) );
  INV_X1 \SB4_0/INV_5  ( .A(\RI3[4][191] ), .ZN(\SB4_0/i1_5 ) );
  INV_X1 \SB4_0/INV_4  ( .A(\RI3[4][190] ), .ZN(\SB4_0/i0[7] ) );
  INV_X1 \SB4_0/INV_3  ( .A(\RI3[4][189] ), .ZN(\SB4_0/i0[8] ) );
  INV_X1 \SB4_0/INV_2  ( .A(\RI3[4][188] ), .ZN(\SB4_0/i1[9] ) );
  INV_X1 \SB4_0/INV_1  ( .A(\RI3[4][187] ), .ZN(\SB4_0/i1_7 ) );
  INV_X1 \SB4_0/INV_0  ( .A(\RI3[4][186] ), .ZN(\SB4_0/i3[0] ) );
  INV_X1 \SB4_1/INV_5  ( .A(\RI3[4][185] ), .ZN(\SB4_1/i1_5 ) );
  INV_X1 \SB4_1/INV_4  ( .A(\RI3[4][184] ), .ZN(\SB4_1/i0[7] ) );
  INV_X1 \SB4_1/INV_3  ( .A(\RI3[4][183] ), .ZN(\SB4_1/i0[8] ) );
  INV_X1 \SB4_1/INV_2  ( .A(\RI3[4][182] ), .ZN(\SB4_1/i1[9] ) );
  INV_X1 \SB4_1/INV_1  ( .A(\RI3[4][181] ), .ZN(\SB4_1/i1_7 ) );
  INV_X1 \SB4_1/INV_0  ( .A(\RI3[4][180] ), .ZN(\SB4_1/i3[0] ) );
  INV_X1 \SB4_2/INV_5  ( .A(\RI3[4][179] ), .ZN(\SB4_2/i1_5 ) );
  INV_X1 \SB4_2/INV_4  ( .A(\RI3[4][178] ), .ZN(\SB4_2/i0[7] ) );
  INV_X1 \SB4_2/INV_3  ( .A(\RI3[4][177] ), .ZN(\SB4_2/i0[8] ) );
  INV_X1 \SB4_2/INV_2  ( .A(\RI3[4][176] ), .ZN(\SB4_2/i1[9] ) );
  INV_X1 \SB4_2/INV_1  ( .A(\RI3[4][175] ), .ZN(\SB4_2/i1_7 ) );
  INV_X1 \SB4_3/INV_5  ( .A(\RI3[4][173] ), .ZN(\SB4_3/i1_5 ) );
  INV_X1 \SB4_3/INV_4  ( .A(\RI3[4][172] ), .ZN(\SB4_3/i0[7] ) );
  INV_X1 \SB4_3/INV_3  ( .A(\RI3[4][171] ), .ZN(\SB4_3/i0[8] ) );
  INV_X1 \SB4_3/INV_2  ( .A(\RI3[4][170] ), .ZN(\SB4_3/i1[9] ) );
  INV_X1 \SB4_3/INV_1  ( .A(\RI3[4][169] ), .ZN(\SB4_3/i1_7 ) );
  INV_X1 \SB4_3/INV_0  ( .A(\RI3[4][168] ), .ZN(\SB4_3/i3[0] ) );
  INV_X1 \SB4_4/INV_5  ( .A(\RI3[4][167] ), .ZN(\SB4_4/i1_5 ) );
  INV_X1 \SB4_4/INV_4  ( .A(\RI3[4][166] ), .ZN(\SB4_4/i0[7] ) );
  INV_X1 \SB4_4/INV_3  ( .A(\RI3[4][165] ), .ZN(\SB4_4/i0[8] ) );
  INV_X1 \SB4_4/INV_2  ( .A(\RI3[4][164] ), .ZN(\SB4_4/i1[9] ) );
  INV_X1 \SB4_4/INV_1  ( .A(\RI3[4][163] ), .ZN(\SB4_4/i1_7 ) );
  INV_X1 \SB4_4/INV_0  ( .A(\RI3[4][162] ), .ZN(\SB4_4/i3[0] ) );
  INV_X1 \SB4_5/INV_5  ( .A(\RI3[4][161] ), .ZN(\SB4_5/i1_5 ) );
  INV_X1 \SB4_5/INV_3  ( .A(\RI3[4][159] ), .ZN(\SB4_5/i0[8] ) );
  INV_X1 \SB4_5/INV_2  ( .A(\RI3[4][158] ), .ZN(\SB4_5/i1[9] ) );
  INV_X1 \SB4_5/INV_1  ( .A(\RI3[4][157] ), .ZN(\SB4_5/i1_7 ) );
  INV_X1 \SB4_5/INV_0  ( .A(\RI3[4][156] ), .ZN(\SB4_5/i3[0] ) );
  INV_X1 \SB4_6/INV_5  ( .A(\RI3[4][155] ), .ZN(\SB4_6/i1_5 ) );
  INV_X1 \SB4_6/INV_4  ( .A(\RI3[4][154] ), .ZN(\SB4_6/i0[7] ) );
  INV_X1 \SB4_6/INV_3  ( .A(\RI3[4][153] ), .ZN(\SB4_6/i0[8] ) );
  INV_X1 \SB4_6/INV_2  ( .A(\RI3[4][152] ), .ZN(\SB4_6/i1[9] ) );
  INV_X1 \SB4_6/INV_1  ( .A(\RI3[4][151] ), .ZN(\SB4_6/i1_7 ) );
  INV_X1 \SB4_6/INV_0  ( .A(\RI3[4][150] ), .ZN(\SB4_6/i3[0] ) );
  INV_X1 \SB4_7/INV_5  ( .A(\RI3[4][149] ), .ZN(\SB4_7/i1_5 ) );
  INV_X1 \SB4_7/INV_4  ( .A(\RI3[4][148] ), .ZN(\SB4_7/i0[7] ) );
  INV_X1 \SB4_7/INV_3  ( .A(\RI3[4][147] ), .ZN(\SB4_7/i0[8] ) );
  INV_X1 \SB4_7/INV_2  ( .A(\RI3[4][146] ), .ZN(\SB4_7/i1[9] ) );
  INV_X1 \SB4_7/INV_1  ( .A(\RI3[4][145] ), .ZN(\SB4_7/i1_7 ) );
  INV_X1 \SB4_7/INV_0  ( .A(\RI3[4][144] ), .ZN(\SB4_7/i3[0] ) );
  INV_X1 \SB4_8/INV_5  ( .A(\RI3[4][143] ), .ZN(\SB4_8/i1_5 ) );
  INV_X1 \SB4_8/INV_3  ( .A(\RI3[4][141] ), .ZN(\SB4_8/i0[8] ) );
  INV_X1 \SB4_8/INV_2  ( .A(\RI3[4][140] ), .ZN(\SB4_8/i1[9] ) );
  INV_X1 \SB4_8/INV_1  ( .A(\RI3[4][139] ), .ZN(\SB4_8/i1_7 ) );
  INV_X1 \SB4_8/INV_0  ( .A(\RI3[4][138] ), .ZN(\SB4_8/i3[0] ) );
  INV_X1 \SB4_9/INV_5  ( .A(\RI3[4][137] ), .ZN(\SB4_9/i1_5 ) );
  INV_X1 \SB4_9/INV_3  ( .A(\RI3[4][135] ), .ZN(\SB4_9/i0[8] ) );
  INV_X1 \SB4_9/INV_2  ( .A(\RI3[4][134] ), .ZN(\SB4_9/i1[9] ) );
  INV_X1 \SB4_9/INV_1  ( .A(\RI3[4][133] ), .ZN(\SB4_9/i1_7 ) );
  INV_X1 \SB4_9/INV_0  ( .A(\RI3[4][132] ), .ZN(\SB4_9/i3[0] ) );
  INV_X1 \SB4_10/INV_5  ( .A(\RI3[4][131] ), .ZN(\SB4_10/i1_5 ) );
  INV_X1 \SB4_10/INV_4  ( .A(\RI3[4][130] ), .ZN(\SB4_10/i0[7] ) );
  INV_X1 \SB4_10/INV_3  ( .A(\RI3[4][129] ), .ZN(\SB4_10/i0[8] ) );
  INV_X1 \SB4_10/INV_2  ( .A(\RI3[4][128] ), .ZN(\SB4_10/i1[9] ) );
  INV_X1 \SB4_10/INV_1  ( .A(\RI3[4][127] ), .ZN(\SB4_10/i1_7 ) );
  INV_X1 \SB4_10/INV_0  ( .A(\RI3[4][126] ), .ZN(\SB4_10/i3[0] ) );
  BUF_X1 \SB4_10/BUF_1  ( .A(\RI3[4][127] ), .Z(\SB4_10/i0[6] ) );
  INV_X1 \SB4_11/INV_5  ( .A(\RI3[4][125] ), .ZN(\SB4_11/i1_5 ) );
  INV_X1 \SB4_11/INV_3  ( .A(\RI3[4][123] ), .ZN(\SB4_11/i0[8] ) );
  INV_X1 \SB4_11/INV_2  ( .A(\RI3[4][122] ), .ZN(\SB4_11/i1[9] ) );
  INV_X1 \SB4_11/INV_1  ( .A(\RI3[4][121] ), .ZN(\SB4_11/i1_7 ) );
  INV_X1 \SB4_11/INV_0  ( .A(\RI3[4][120] ), .ZN(\SB4_11/i3[0] ) );
  INV_X1 \SB4_12/INV_5  ( .A(\RI3[4][119] ), .ZN(\SB4_12/i1_5 ) );
  INV_X1 \SB4_12/INV_4  ( .A(\RI3[4][118] ), .ZN(\SB4_12/i0[7] ) );
  INV_X1 \SB4_12/INV_3  ( .A(\RI3[4][117] ), .ZN(\SB4_12/i0[8] ) );
  INV_X1 \SB4_12/INV_2  ( .A(\RI3[4][116] ), .ZN(\SB4_12/i1[9] ) );
  INV_X1 \SB4_12/INV_1  ( .A(\RI3[4][115] ), .ZN(\SB4_12/i1_7 ) );
  INV_X1 \SB4_12/INV_0  ( .A(\RI3[4][114] ), .ZN(\SB4_12/i3[0] ) );
  INV_X1 \SB4_13/INV_5  ( .A(\RI3[4][113] ), .ZN(\SB4_13/i1_5 ) );
  INV_X1 \SB4_13/INV_4  ( .A(\RI3[4][112] ), .ZN(\SB4_13/i0[7] ) );
  INV_X1 \SB4_13/INV_3  ( .A(\RI3[4][111] ), .ZN(\SB4_13/i0[8] ) );
  INV_X1 \SB4_13/INV_2  ( .A(\RI3[4][110] ), .ZN(\SB4_13/i1[9] ) );
  INV_X1 \SB4_13/INV_1  ( .A(\RI3[4][109] ), .ZN(\SB4_13/i1_7 ) );
  INV_X1 \SB4_13/INV_0  ( .A(\RI3[4][108] ), .ZN(\SB4_13/i3[0] ) );
  INV_X1 \SB4_14/INV_5  ( .A(\RI3[4][107] ), .ZN(\SB4_14/i1_5 ) );
  INV_X1 \SB4_14/INV_3  ( .A(\RI3[4][105] ), .ZN(\SB4_14/i0[8] ) );
  INV_X1 \SB4_14/INV_2  ( .A(\RI3[4][104] ), .ZN(\SB4_14/i1[9] ) );
  INV_X1 \SB4_14/INV_1  ( .A(\RI3[4][103] ), .ZN(\SB4_14/i1_7 ) );
  INV_X1 \SB4_14/INV_0  ( .A(\RI3[4][102] ), .ZN(\SB4_14/i3[0] ) );
  INV_X1 \SB4_15/INV_5  ( .A(\RI3[4][101] ), .ZN(\SB4_15/i1_5 ) );
  INV_X1 \SB4_15/INV_4  ( .A(\RI3[4][100] ), .ZN(\SB4_15/i0[7] ) );
  INV_X1 \SB4_15/INV_3  ( .A(\RI3[4][99] ), .ZN(\SB4_15/i0[8] ) );
  INV_X1 \SB4_15/INV_2  ( .A(\RI3[4][98] ), .ZN(\SB4_15/i1[9] ) );
  INV_X1 \SB4_15/INV_1  ( .A(\RI3[4][97] ), .ZN(\SB4_15/i1_7 ) );
  INV_X1 \SB4_15/INV_0  ( .A(\RI3[4][96] ), .ZN(\SB4_15/i3[0] ) );
  INV_X1 \SB4_16/INV_5  ( .A(\RI3[4][95] ), .ZN(\SB4_16/i1_5 ) );
  INV_X1 \SB4_16/INV_4  ( .A(\RI3[4][94] ), .ZN(\SB4_16/i0[7] ) );
  INV_X1 \SB4_16/INV_3  ( .A(\RI3[4][93] ), .ZN(\SB4_16/i0[8] ) );
  INV_X1 \SB4_16/INV_2  ( .A(\RI3[4][92] ), .ZN(\SB4_16/i1[9] ) );
  INV_X1 \SB4_16/INV_1  ( .A(\RI3[4][91] ), .ZN(\SB4_16/i1_7 ) );
  INV_X1 \SB4_16/INV_0  ( .A(\RI3[4][90] ), .ZN(\SB4_16/i3[0] ) );
  INV_X1 \SB4_17/INV_5  ( .A(\RI3[4][89] ), .ZN(\SB4_17/i1_5 ) );
  INV_X1 \SB4_17/INV_4  ( .A(\RI3[4][88] ), .ZN(\SB4_17/i0[7] ) );
  INV_X1 \SB4_17/INV_3  ( .A(\RI3[4][87] ), .ZN(\SB4_17/i0[8] ) );
  INV_X1 \SB4_17/INV_1  ( .A(\RI3[4][85] ), .ZN(\SB4_17/i1_7 ) );
  INV_X1 \SB4_17/INV_0  ( .A(\RI3[4][84] ), .ZN(\SB4_17/i3[0] ) );
  INV_X1 \SB4_18/INV_5  ( .A(\RI3[4][83] ), .ZN(\SB4_18/i1_5 ) );
  INV_X1 \SB4_18/INV_4  ( .A(\RI3[4][82] ), .ZN(\SB4_18/i0[7] ) );
  INV_X1 \SB4_18/INV_3  ( .A(\RI3[4][81] ), .ZN(\SB4_18/i0[8] ) );
  INV_X1 \SB4_18/INV_1  ( .A(\RI3[4][79] ), .ZN(\SB4_18/i1_7 ) );
  INV_X1 \SB4_18/INV_0  ( .A(\RI3[4][78] ), .ZN(\SB4_18/i3[0] ) );
  INV_X1 \SB4_19/INV_5  ( .A(\RI3[4][77] ), .ZN(\SB4_19/i1_5 ) );
  INV_X1 \SB4_19/INV_4  ( .A(\RI3[4][76] ), .ZN(\SB4_19/i0[7] ) );
  INV_X1 \SB4_19/INV_3  ( .A(\RI3[4][75] ), .ZN(\SB4_19/i0[8] ) );
  INV_X1 \SB4_19/INV_2  ( .A(\RI3[4][74] ), .ZN(\SB4_19/i1[9] ) );
  INV_X1 \SB4_19/INV_1  ( .A(\RI3[4][73] ), .ZN(\SB4_19/i1_7 ) );
  INV_X1 \SB4_19/INV_0  ( .A(\RI3[4][72] ), .ZN(\SB4_19/i3[0] ) );
  INV_X1 \SB4_20/INV_5  ( .A(\RI3[4][71] ), .ZN(\SB4_20/i1_5 ) );
  INV_X1 \SB4_20/INV_3  ( .A(\RI3[4][69] ), .ZN(\SB4_20/i0[8] ) );
  INV_X1 \SB4_20/INV_2  ( .A(\RI3[4][68] ), .ZN(\SB4_20/i1[9] ) );
  INV_X1 \SB4_20/INV_1  ( .A(\RI3[4][67] ), .ZN(\SB4_20/i1_7 ) );
  INV_X1 \SB4_20/INV_0  ( .A(\RI3[4][66] ), .ZN(\SB4_20/i3[0] ) );
  INV_X1 \SB4_21/INV_5  ( .A(\RI3[4][65] ), .ZN(\SB4_21/i1_5 ) );
  INV_X1 \SB4_21/INV_4  ( .A(\RI3[4][64] ), .ZN(\SB4_21/i0[7] ) );
  INV_X1 \SB4_21/INV_3  ( .A(\RI3[4][63] ), .ZN(\SB4_21/i0[8] ) );
  INV_X1 \SB4_21/INV_1  ( .A(\RI3[4][61] ), .ZN(\SB4_21/i1_7 ) );
  INV_X1 \SB4_21/INV_0  ( .A(\RI3[4][60] ), .ZN(\SB4_21/i3[0] ) );
  INV_X1 \SB4_22/INV_5  ( .A(\RI3[4][59] ), .ZN(\SB4_22/i1_5 ) );
  INV_X1 \SB4_22/INV_4  ( .A(\RI3[4][58] ), .ZN(\SB4_22/i0[7] ) );
  INV_X1 \SB4_22/INV_3  ( .A(\RI3[4][57] ), .ZN(\SB4_22/i0[8] ) );
  INV_X1 \SB4_22/INV_1  ( .A(\RI3[4][55] ), .ZN(\SB4_22/i1_7 ) );
  INV_X1 \SB4_23/INV_5  ( .A(\RI3[4][53] ), .ZN(\SB4_23/i1_5 ) );
  INV_X1 \SB4_23/INV_4  ( .A(\RI3[4][52] ), .ZN(\SB4_23/i0[7] ) );
  INV_X1 \SB4_23/INV_3  ( .A(\RI3[4][51] ), .ZN(\SB4_23/i0[8] ) );
  INV_X1 \SB4_23/INV_2  ( .A(\RI3[4][50] ), .ZN(\SB4_23/i1[9] ) );
  INV_X1 \SB4_23/INV_1  ( .A(\RI3[4][49] ), .ZN(\SB4_23/i1_7 ) );
  INV_X1 \SB4_23/INV_0  ( .A(\RI3[4][48] ), .ZN(\SB4_23/i3[0] ) );
  INV_X1 \SB4_24/INV_5  ( .A(\RI3[4][47] ), .ZN(\SB4_24/i1_5 ) );
  INV_X1 \SB4_24/INV_4  ( .A(\RI3[4][46] ), .ZN(\SB4_24/i0[7] ) );
  INV_X1 \SB4_24/INV_3  ( .A(\RI3[4][45] ), .ZN(\SB4_24/i0[8] ) );
  INV_X1 \SB4_24/INV_2  ( .A(\RI3[4][44] ), .ZN(\SB4_24/i1[9] ) );
  INV_X1 \SB4_24/INV_1  ( .A(\RI3[4][43] ), .ZN(\SB4_24/i1_7 ) );
  INV_X1 \SB4_24/INV_0  ( .A(\RI3[4][42] ), .ZN(\SB4_24/i3[0] ) );
  BUF_X1 \SB4_24/BUF_1  ( .A(\RI3[4][43] ), .Z(\SB4_24/i0[6] ) );
  INV_X1 \SB4_25/INV_5  ( .A(\RI3[4][41] ), .ZN(\SB4_25/i1_5 ) );
  INV_X1 \SB4_25/INV_3  ( .A(\RI3[4][39] ), .ZN(\SB4_25/i0[8] ) );
  INV_X1 \SB4_25/INV_2  ( .A(\RI3[4][38] ), .ZN(\SB4_25/i1[9] ) );
  INV_X1 \SB4_25/INV_1  ( .A(\RI3[4][37] ), .ZN(\SB4_25/i1_7 ) );
  INV_X1 \SB4_25/INV_0  ( .A(\RI3[4][36] ), .ZN(\SB4_25/i3[0] ) );
  INV_X1 \SB4_26/INV_5  ( .A(\RI3[4][35] ), .ZN(\SB4_26/i1_5 ) );
  INV_X1 \SB4_26/INV_4  ( .A(\RI3[4][34] ), .ZN(\SB4_26/i0[7] ) );
  INV_X1 \SB4_26/INV_3  ( .A(\RI3[4][33] ), .ZN(\SB4_26/i0[8] ) );
  INV_X1 \SB4_26/INV_2  ( .A(\RI3[4][32] ), .ZN(\SB4_26/i1[9] ) );
  INV_X1 \SB4_26/INV_1  ( .A(\RI3[4][31] ), .ZN(\SB4_26/i1_7 ) );
  INV_X1 \SB4_26/INV_0  ( .A(\RI3[4][30] ), .ZN(\SB4_26/i3[0] ) );
  INV_X1 \SB4_27/INV_5  ( .A(\RI3[4][29] ), .ZN(\SB4_27/i1_5 ) );
  INV_X1 \SB4_27/INV_3  ( .A(\RI3[4][27] ), .ZN(\SB4_27/i0[8] ) );
  INV_X1 \SB4_27/INV_2  ( .A(\RI3[4][26] ), .ZN(\SB4_27/i1[9] ) );
  INV_X1 \SB4_27/INV_1  ( .A(\RI3[4][25] ), .ZN(\SB4_27/i1_7 ) );
  INV_X1 \SB4_27/INV_0  ( .A(\RI3[4][24] ), .ZN(\SB4_27/i3[0] ) );
  INV_X1 \SB4_28/INV_5  ( .A(\RI3[4][23] ), .ZN(\SB4_28/i1_5 ) );
  INV_X1 \SB4_28/INV_4  ( .A(\RI3[4][22] ), .ZN(\SB4_28/i0[7] ) );
  INV_X1 \SB4_28/INV_3  ( .A(\RI3[4][21] ), .ZN(\SB4_28/i0[8] ) );
  INV_X1 \SB4_28/INV_2  ( .A(\RI3[4][20] ), .ZN(\SB4_28/i1[9] ) );
  INV_X1 \SB4_28/INV_1  ( .A(\RI3[4][19] ), .ZN(\SB4_28/i1_7 ) );
  INV_X1 \SB4_28/INV_0  ( .A(\RI3[4][18] ), .ZN(\SB4_28/i3[0] ) );
  INV_X1 \SB4_29/INV_5  ( .A(\RI3[4][17] ), .ZN(\SB4_29/i1_5 ) );
  INV_X1 \SB4_29/INV_3  ( .A(\RI3[4][15] ), .ZN(\SB4_29/i0[8] ) );
  INV_X1 \SB4_29/INV_2  ( .A(\RI3[4][14] ), .ZN(\SB4_29/i1[9] ) );
  INV_X1 \SB4_30/INV_5  ( .A(\RI3[4][11] ), .ZN(\SB4_30/i1_5 ) );
  INV_X1 \SB4_30/INV_4  ( .A(\RI3[4][10] ), .ZN(\SB4_30/i0[7] ) );
  INV_X1 \SB4_30/INV_3  ( .A(\RI3[4][9] ), .ZN(\SB4_30/i0[8] ) );
  INV_X1 \SB4_30/INV_2  ( .A(\RI3[4][8] ), .ZN(\SB4_30/i1[9] ) );
  INV_X1 \SB4_30/INV_1  ( .A(\RI3[4][7] ), .ZN(\SB4_30/i1_7 ) );
  INV_X1 \SB4_30/INV_0  ( .A(\RI3[4][6] ), .ZN(\SB4_30/i3[0] ) );
  INV_X1 \SB4_31/INV_4  ( .A(\RI3[4][4] ), .ZN(\SB4_31/i0[7] ) );
  INV_X1 \SB4_31/INV_3  ( .A(\RI3[4][3] ), .ZN(\SB4_31/i0[8] ) );
  INV_X1 \SB4_31/INV_2  ( .A(\RI3[4][2] ), .ZN(\SB4_31/i1[9] ) );
  INV_X1 \SB4_31/INV_1  ( .A(\RI3[4][1] ), .ZN(\SB4_31/i1_7 ) );
  INV_X1 \SB4_31/INV_0  ( .A(\RI3[4][0] ), .ZN(\SB4_31/i3[0] ) );
  NAND4_X1 \SB1_0_0/Component_Function_2/N5  ( .A1(
        \SB1_0_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_0/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][14] ) );
  NAND4_X1 \SB1_0_0/Component_Function_3/N5  ( .A1(
        \SB1_0_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_0/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][9] ) );
  NAND4_X1 \SB1_0_0/Component_Function_4/N5  ( .A1(
        \SB1_0_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_0/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][4] ) );
  NAND4_X1 \SB1_0_1/Component_Function_3/N5  ( .A1(
        \SB1_0_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][3] ) );
  NAND4_X1 \SB1_0_1/Component_Function_4/N5  ( .A1(
        \SB1_0_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][190] ) );
  NAND4_X1 \SB1_0_2/Component_Function_2/N5  ( .A1(
        \SB1_0_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_2/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][2] ) );
  NAND4_X1 \SB1_0_2/Component_Function_3/N5  ( .A1(
        \SB1_0_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_2/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][189] ) );
  NAND4_X1 \SB1_0_2/Component_Function_4/N5  ( .A1(
        \SB1_0_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_2/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][184] ) );
  NAND4_X1 \SB1_0_3/Component_Function_2/N5  ( .A1(
        \SB1_0_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_3/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][188] ) );
  NAND4_X1 \SB1_0_3/Component_Function_3/N5  ( .A1(
        \SB1_0_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][183] ) );
  NAND4_X1 \SB1_0_3/Component_Function_4/N5  ( .A1(
        \SB1_0_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][178] ) );
  NAND4_X1 \SB1_0_4/Component_Function_3/N5  ( .A1(
        \SB1_0_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][177] ) );
  NAND4_X1 \SB1_0_5/Component_Function_2/N5  ( .A1(
        \SB1_0_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_5/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_5/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_5/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][176] ) );
  NAND4_X1 \SB1_0_5/Component_Function_3/N5  ( .A1(
        \SB1_0_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][171] ) );
  NAND4_X1 \SB1_0_5/Component_Function_4/N5  ( .A1(
        \SB1_0_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_5/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][166] ) );
  NAND4_X1 \SB1_0_6/Component_Function_2/N5  ( .A1(
        \SB1_0_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_6/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_6/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][170] ) );
  NAND4_X1 \SB1_0_6/Component_Function_3/N5  ( .A1(
        \SB1_0_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][165] ) );
  NAND4_X1 \SB1_0_6/Component_Function_4/N5  ( .A1(
        \SB1_0_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_6/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][160] ) );
  NAND4_X1 \SB1_0_7/Component_Function_2/N5  ( .A1(
        \SB1_0_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_7/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][164] ) );
  NAND4_X1 \SB1_0_7/Component_Function_3/N5  ( .A1(
        \SB1_0_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][159] ) );
  NAND4_X1 \SB1_0_7/Component_Function_4/N5  ( .A1(
        \SB1_0_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_7/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][154] ) );
  NAND4_X1 \SB1_0_9/Component_Function_2/N5  ( .A1(
        \SB1_0_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][152] ) );
  NAND4_X1 \SB1_0_9/Component_Function_3/N5  ( .A1(
        \SB1_0_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][147] ) );
  NAND4_X1 \SB1_0_9/Component_Function_4/N5  ( .A1(
        \SB1_0_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][142] ) );
  NAND4_X1 \SB1_0_10/Component_Function_2/N5  ( .A1(
        \SB1_0_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][146] ) );
  NAND4_X1 \SB1_0_10/Component_Function_3/N5  ( .A1(
        \SB1_0_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][141] ) );
  NAND4_X1 \SB1_0_10/Component_Function_4/N5  ( .A1(
        \SB1_0_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][136] ) );
  NAND4_X1 \SB1_0_11/Component_Function_2/N5  ( .A1(
        \SB1_0_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_11/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][140] ) );
  NAND4_X1 \SB1_0_11/Component_Function_3/N5  ( .A1(
        \SB1_0_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][135] ) );
  NAND4_X1 \SB1_0_11/Component_Function_4/N5  ( .A1(
        \SB1_0_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][130] ) );
  NAND4_X1 \SB1_0_12/Component_Function_2/N5  ( .A1(
        \SB1_0_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_12/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][134] ) );
  NAND4_X1 \SB1_0_12/Component_Function_3/N5  ( .A1(
        \SB1_0_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_12/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][129] ) );
  NAND4_X1 \SB1_0_12/Component_Function_4/N5  ( .A1(
        \SB1_0_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_12/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][124] ) );
  NAND4_X1 \SB1_0_13/Component_Function_3/N5  ( .A1(
        \SB1_0_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][123] ) );
  NAND4_X1 \SB1_0_13/Component_Function_4/N5  ( .A1(
        \SB1_0_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][118] ) );
  NAND4_X1 \SB1_0_14/Component_Function_2/N5  ( .A1(
        \SB1_0_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][122] ) );
  NAND4_X1 \SB1_0_14/Component_Function_3/N5  ( .A1(
        \SB1_0_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][117] ) );
  NAND4_X1 \SB1_0_14/Component_Function_4/N5  ( .A1(
        \SB1_0_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][112] ) );
  NAND4_X1 \SB1_0_15/Component_Function_3/N5  ( .A1(
        \SB1_0_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][111] ) );
  NAND4_X1 \SB1_0_15/Component_Function_4/N5  ( .A1(
        \SB1_0_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_15/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][106] ) );
  NAND4_X1 \SB1_0_16/Component_Function_3/N5  ( .A1(
        \SB1_0_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_16/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][105] ) );
  NAND4_X1 \SB1_0_17/Component_Function_2/N5  ( .A1(
        \SB1_0_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_17/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][104] ) );
  NAND4_X1 \SB1_0_17/Component_Function_3/N5  ( .A1(
        \SB1_0_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_17/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][99] ) );
  NAND4_X1 \SB1_0_17/Component_Function_4/N5  ( .A1(
        \SB1_0_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][94] ) );
  NAND4_X1 \SB1_0_18/Component_Function_2/N5  ( .A1(
        \SB1_0_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_18/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_18/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_18/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][98] ) );
  NAND4_X1 \SB1_0_18/Component_Function_3/N5  ( .A1(
        \SB1_0_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][93] ) );
  NAND4_X1 \SB1_0_19/Component_Function_2/N5  ( .A1(
        \SB1_0_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_19/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_19/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][92] ) );
  NAND4_X1 \SB1_0_19/Component_Function_4/N5  ( .A1(
        \SB1_0_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_19/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][82] ) );
  NAND4_X1 \SB1_0_20/Component_Function_2/N5  ( .A1(
        \SB1_0_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_20/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_20/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][86] ) );
  NAND4_X1 \SB1_0_20/Component_Function_3/N5  ( .A1(
        \SB1_0_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_20/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][81] ) );
  NAND4_X1 \SB1_0_20/Component_Function_4/N5  ( .A1(
        \SB1_0_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_20/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][76] ) );
  NAND4_X1 \SB1_0_21/Component_Function_3/N5  ( .A1(
        \SB1_0_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_21/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][75] ) );
  NAND4_X1 \SB1_0_21/Component_Function_4/N5  ( .A1(
        \SB1_0_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_21/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][70] ) );
  NAND4_X1 \SB1_0_22/Component_Function_2/N5  ( .A1(
        \SB1_0_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_22/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][74] ) );
  NAND4_X1 \SB1_0_22/Component_Function_3/N5  ( .A1(
        \SB1_0_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_22/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][69] ) );
  NAND4_X1 \SB1_0_22/Component_Function_4/N5  ( .A1(
        \SB1_0_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_22/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][64] ) );
  NAND4_X1 \SB1_0_23/Component_Function_2/N5  ( .A1(
        \SB1_0_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][68] ) );
  NAND4_X1 \SB1_0_23/Component_Function_3/N5  ( .A1(
        \SB1_0_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][63] ) );
  NAND4_X1 \SB1_0_24/Component_Function_2/N5  ( .A1(
        \SB1_0_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_24/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][62] ) );
  NAND4_X1 \SB1_0_24/Component_Function_3/N5  ( .A1(
        \SB1_0_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_24/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][57] ) );
  NAND4_X1 \SB1_0_25/Component_Function_2/N5  ( .A1(
        \SB1_0_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_25/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_25/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][56] ) );
  NAND4_X1 \SB1_0_25/Component_Function_3/N5  ( .A1(
        \SB1_0_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_25/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][51] ) );
  NAND4_X1 \SB1_0_25/Component_Function_4/N5  ( .A1(
        \SB1_0_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_25/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_25/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][46] ) );
  NAND4_X1 \SB1_0_26/Component_Function_3/N5  ( .A1(
        \SB1_0_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_26/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][45] ) );
  NAND4_X1 \SB1_0_26/Component_Function_4/N5  ( .A1(
        \SB1_0_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_26/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][40] ) );
  NAND4_X1 \SB1_0_27/Component_Function_2/N5  ( .A1(
        \SB1_0_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][44] ) );
  NAND4_X1 \SB1_0_27/Component_Function_3/N5  ( .A1(
        \SB1_0_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][39] ) );
  NAND4_X1 \SB1_0_28/Component_Function_2/N5  ( .A1(
        \SB1_0_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_28/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][38] ) );
  NAND4_X1 \SB1_0_28/Component_Function_3/N5  ( .A1(
        \SB1_0_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_28/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][33] ) );
  NAND4_X1 \SB1_0_28/Component_Function_4/N5  ( .A1(
        \SB1_0_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_28/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][28] ) );
  NAND4_X1 \SB1_0_29/Component_Function_2/N5  ( .A1(
        \SB1_0_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_29/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][32] ) );
  NAND4_X1 \SB1_0_29/Component_Function_3/N5  ( .A1(
        \SB1_0_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_29/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][27] ) );
  NAND4_X1 \SB1_0_29/Component_Function_4/N5  ( .A1(
        \SB1_0_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_29/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][22] ) );
  NAND4_X1 \SB1_0_30/Component_Function_2/N5  ( .A1(
        \SB1_0_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][26] ) );
  NAND4_X1 \SB1_0_30/Component_Function_4/N5  ( .A1(
        \SB1_0_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][16] ) );
  NAND4_X1 \SB1_0_31/Component_Function_3/N5  ( .A1(
        \SB1_0_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][15] ) );
  NAND4_X1 \SB1_0_31/Component_Function_4/N5  ( .A1(
        \SB1_0_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][10] ) );
  NAND4_X1 \SB2_0_5/Component_Function_2/N5  ( .A1(
        \SB2_0_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_5/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_5/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[0][176] ) );
  NAND4_X1 \SB2_0_5/Component_Function_4/N5  ( .A1(
        \SB2_0_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_5/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][166] ) );
  NAND4_X1 \SB2_0_10/Component_Function_4/N5  ( .A1(
        \SB2_0_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_10/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][136] ) );
  NAND4_X1 \SB2_0_12/Component_Function_2/N5  ( .A1(
        \SB2_0_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[0][134] ) );
  NAND4_X1 \SB2_0_12/Component_Function_4/N5  ( .A1(
        \SB2_0_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][124] ) );
  NAND4_X1 \SB2_0_13/Component_Function_4/N5  ( .A1(
        \SB2_0_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_13/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][118] ) );
  NAND4_X1 \SB2_0_15/Component_Function_4/N5  ( .A1(
        \SB2_0_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_15/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][106] ) );
  NAND4_X1 \SB2_0_17/Component_Function_3/N5  ( .A1(
        \SB2_0_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_17/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[0][99] ) );
  NAND4_X1 \SB2_0_17/Component_Function_4/N5  ( .A1(
        \SB2_0_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][94] ) );
  NAND4_X1 \SB2_0_18/Component_Function_4/N5  ( .A1(
        \SB2_0_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_18/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][88] ) );
  NAND4_X1 \SB2_0_19/Component_Function_3/N5  ( .A1(
        \SB2_0_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_19/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[0][87] ) );
  NAND4_X1 \SB2_0_19/Component_Function_4/N5  ( .A1(
        \SB2_0_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_19/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][82] ) );
  NAND4_X1 \SB2_0_28/Component_Function_4/N5  ( .A1(
        \SB2_0_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_28/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][28] ) );
  NAND4_X1 \SB2_0_29/Component_Function_3/N5  ( .A1(
        \SB2_0_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[0][27] ) );
  NAND4_X1 \SB2_0_29/Component_Function_4/N5  ( .A1(
        \SB2_0_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][22] ) );
  NAND4_X1 \SB1_1_0/Component_Function_2/N5  ( .A1(
        \SB1_1_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_0/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_0/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_0/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][14] ) );
  NAND4_X1 \SB1_1_0/Component_Function_3/N5  ( .A1(
        \SB1_1_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_0/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][9] ) );
  NAND4_X1 \SB1_1_0/Component_Function_4/N5  ( .A1(
        \SB1_1_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_0/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][4] ) );
  NAND4_X1 \SB1_1_1/Component_Function_3/N5  ( .A1(
        \SB1_1_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_1/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_1/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][3] ) );
  NAND4_X1 \SB1_1_1/Component_Function_4/N5  ( .A1(
        \SB1_1_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_1/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][190] ) );
  NAND4_X1 \SB1_1_2/Component_Function_2/N5  ( .A1(
        \SB1_1_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_2/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_2/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][2] ) );
  NAND4_X1 \SB1_1_2/Component_Function_3/N5  ( .A1(
        \SB1_1_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_2/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][189] ) );
  NAND4_X1 \SB1_1_3/Component_Function_3/N5  ( .A1(
        \SB1_1_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][183] ) );
  NAND4_X1 \SB1_1_3/Component_Function_4/N5  ( .A1(
        \SB1_1_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][178] ) );
  NAND4_X1 \SB1_1_4/Component_Function_3/N5  ( .A1(
        \SB1_1_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][177] ) );
  NAND4_X1 \SB1_1_5/Component_Function_2/N5  ( .A1(
        \SB1_1_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][176] ) );
  NAND4_X1 \SB1_1_5/Component_Function_3/N5  ( .A1(
        \SB1_1_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][171] ) );
  NAND4_X1 \SB1_1_5/Component_Function_4/N5  ( .A1(
        \SB1_1_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][166] ) );
  NAND4_X1 \SB1_1_6/Component_Function_3/N5  ( .A1(
        \SB1_1_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][165] ) );
  NAND4_X1 \SB1_1_6/Component_Function_4/N5  ( .A1(
        \SB1_1_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_6/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][160] ) );
  NAND4_X1 \SB1_1_8/Component_Function_2/N5  ( .A1(
        \SB1_1_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_8/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_8/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][158] ) );
  NAND4_X1 \SB1_1_9/Component_Function_2/N5  ( .A1(
        \SB1_1_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][152] ) );
  NAND4_X1 \SB1_1_9/Component_Function_3/N5  ( .A1(
        \SB1_1_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][147] ) );
  NAND4_X1 \SB1_1_9/Component_Function_4/N5  ( .A1(
        \SB1_1_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][142] ) );
  NAND4_X1 \SB1_1_10/Component_Function_3/N5  ( .A1(
        \SB1_1_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_10/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][141] ) );
  NAND4_X1 \SB1_1_10/Component_Function_4/N5  ( .A1(
        \SB1_1_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_10/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][136] ) );
  NAND4_X1 \SB1_1_11/Component_Function_3/N5  ( .A1(
        \SB1_1_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_11/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][135] ) );
  NAND4_X1 \SB1_1_11/Component_Function_4/N5  ( .A1(
        \SB1_1_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_11/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][130] ) );
  NAND4_X1 \SB1_1_12/Component_Function_3/N5  ( .A1(
        \SB1_1_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_12/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][129] ) );
  NAND4_X1 \SB1_1_13/Component_Function_3/N5  ( .A1(
        \SB1_1_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][123] ) );
  NAND4_X1 \SB1_1_13/Component_Function_4/N5  ( .A1(
        \SB1_1_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_13/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][118] ) );
  NAND4_X1 \SB1_1_14/Component_Function_2/N5  ( .A1(
        \SB1_1_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][122] ) );
  NAND4_X1 \SB1_1_14/Component_Function_3/N5  ( .A1(
        \SB1_1_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][117] ) );
  NAND4_X1 \SB1_1_14/Component_Function_4/N5  ( .A1(
        \SB1_1_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][112] ) );
  NAND4_X1 \SB1_1_15/Component_Function_2/N5  ( .A1(
        \SB1_1_15/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_15/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_15/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][116] ) );
  NAND4_X1 \SB1_1_15/Component_Function_3/N5  ( .A1(
        \SB1_1_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][111] ) );
  NAND4_X1 \SB1_1_15/Component_Function_4/N5  ( .A1(
        \SB1_1_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_15/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][106] ) );
  NAND4_X1 \SB1_1_16/Component_Function_2/N5  ( .A1(
        \SB1_1_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_16/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_16/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][110] ) );
  NAND4_X1 \SB1_1_16/Component_Function_3/N5  ( .A1(
        \SB1_1_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_16/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][105] ) );
  NAND4_X1 \SB1_1_17/Component_Function_3/N5  ( .A1(
        \SB1_1_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_17/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_17/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][99] ) );
  NAND4_X1 \SB1_1_17/Component_Function_4/N5  ( .A1(
        \SB1_1_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][94] ) );
  NAND4_X1 \SB1_1_18/Component_Function_2/N5  ( .A1(
        \SB1_1_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_18/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][98] ) );
  NAND4_X1 \SB1_1_18/Component_Function_3/N5  ( .A1(
        \SB1_1_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][93] ) );
  NAND4_X1 \SB1_1_18/Component_Function_4/N5  ( .A1(
        \SB1_1_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_18/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][88] ) );
  NAND4_X1 \SB1_1_19/Component_Function_2/N5  ( .A1(
        \SB1_1_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][92] ) );
  NAND4_X1 \SB1_1_19/Component_Function_3/N5  ( .A1(
        \SB1_1_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][87] ) );
  NAND4_X1 \SB1_1_19/Component_Function_4/N5  ( .A1(
        \SB1_1_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][82] ) );
  NAND4_X1 \SB1_1_20/Component_Function_4/N5  ( .A1(
        \SB1_1_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_20/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][76] ) );
  NAND4_X1 \SB1_1_21/Component_Function_2/N5  ( .A1(
        \SB1_1_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_21/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][80] ) );
  NAND4_X1 \SB1_1_21/Component_Function_3/N5  ( .A1(
        \SB1_1_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_21/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][75] ) );
  NAND4_X1 \SB1_1_21/Component_Function_4/N5  ( .A1(
        \SB1_1_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_21/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][70] ) );
  NAND4_X1 \SB1_1_22/Component_Function_3/N5  ( .A1(
        \SB1_1_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_22/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][69] ) );
  NAND4_X1 \SB1_1_22/Component_Function_4/N5  ( .A1(
        \SB1_1_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_22/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][64] ) );
  NAND4_X1 \SB1_1_23/Component_Function_2/N5  ( .A1(
        \SB1_1_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_23/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_23/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][68] ) );
  NAND4_X1 \SB1_1_23/Component_Function_3/N5  ( .A1(
        \SB1_1_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][63] ) );
  NAND4_X1 \SB1_1_23/Component_Function_4/N5  ( .A1(
        \SB1_1_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_23/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][58] ) );
  NAND4_X1 \SB1_1_24/Component_Function_3/N5  ( .A1(
        \SB1_1_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_24/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][57] ) );
  NAND4_X1 \SB1_1_24/Component_Function_4/N5  ( .A1(
        \SB1_1_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_24/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][52] ) );
  NAND4_X1 \SB1_1_25/Component_Function_3/N5  ( .A1(
        \SB1_1_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_25/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][51] ) );
  NAND4_X1 \SB1_1_25/Component_Function_4/N5  ( .A1(
        \SB1_1_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_25/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][46] ) );
  NAND4_X1 \SB1_1_26/Component_Function_2/N5  ( .A1(
        \SB1_1_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_26/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_26/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][50] ) );
  NAND4_X1 \SB1_1_26/Component_Function_3/N5  ( .A1(
        \SB1_1_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_26/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][45] ) );
  NAND4_X1 \SB1_1_26/Component_Function_4/N5  ( .A1(
        \SB1_1_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_26/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][40] ) );
  NAND4_X1 \SB1_1_27/Component_Function_3/N5  ( .A1(
        \SB1_1_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][39] ) );
  NAND4_X1 \SB1_1_27/Component_Function_4/N5  ( .A1(
        \SB1_1_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_27/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][34] ) );
  NAND4_X1 \SB1_1_28/Component_Function_3/N5  ( .A1(
        \SB1_1_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_28/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][33] ) );
  NAND4_X1 \SB1_1_29/Component_Function_2/N5  ( .A1(
        \SB1_1_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][32] ) );
  NAND4_X1 \SB1_1_29/Component_Function_3/N5  ( .A1(
        \SB1_1_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][27] ) );
  NAND4_X1 \SB1_1_29/Component_Function_4/N5  ( .A1(
        \SB1_1_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][22] ) );
  NAND4_X1 \SB1_1_30/Component_Function_3/N5  ( .A1(
        \SB1_1_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_30/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][21] ) );
  NAND4_X1 \SB1_1_30/Component_Function_4/N5  ( .A1(
        \SB1_1_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_30/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[1][16] ) );
  NAND4_X1 \SB1_1_31/Component_Function_2/N5  ( .A1(
        \SB1_1_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_31/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][20] ) );
  NAND4_X1 \SB1_1_31/Component_Function_3/N5  ( .A1(
        \SB1_1_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_31/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[1][15] ) );
  NAND4_X1 \SB2_1_0/Component_Function_4/N5  ( .A1(
        \SB2_1_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_0/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][4] ) );
  NAND4_X1 \SB2_1_1/Component_Function_3/N5  ( .A1(
        \SB2_1_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_1/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_1/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][3] ) );
  NAND4_X1 \SB2_1_1/Component_Function_4/N5  ( .A1(
        \SB2_1_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_1/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][190] ) );
  NAND4_X1 \SB2_1_2/Component_Function_4/N5  ( .A1(
        \SB2_1_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_2/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][184] ) );
  NAND4_X1 \SB2_1_4/Component_Function_2/N5  ( .A1(
        \SB2_1_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_1_4/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[1][182] ) );
  NAND4_X1 \SB2_1_4/Component_Function_4/N5  ( .A1(
        \SB2_1_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_4/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][172] ) );
  NAND4_X1 \SB2_1_9/Component_Function_4/N5  ( .A1(
        \SB2_1_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_9/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][142] ) );
  NAND4_X1 \SB2_1_10/Component_Function_4/N5  ( .A1(
        \SB2_1_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_10/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][136] ) );
  NAND4_X1 \SB2_1_12/Component_Function_4/N5  ( .A1(
        \SB2_1_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_12/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][124] ) );
  NAND4_X1 \SB2_1_13/Component_Function_2/N5  ( .A1(
        \SB2_1_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_1_13/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[1][128] ) );
  NAND4_X1 \SB2_1_13/Component_Function_4/N5  ( .A1(
        \SB2_1_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_13/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][118] ) );
  NAND4_X1 \SB2_1_15/Component_Function_3/N5  ( .A1(
        \SB2_1_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][111] ) );
  NAND4_X1 \SB2_1_16/Component_Function_4/N5  ( .A1(
        \SB2_1_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_16/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_16/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][100] ) );
  NAND4_X1 \SB2_1_17/Component_Function_4/N5  ( .A1(
        \SB2_1_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][94] ) );
  NAND4_X1 \SB2_1_18/Component_Function_4/N5  ( .A1(
        \SB2_1_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][88] ) );
  NAND4_X1 \SB2_1_21/Component_Function_4/N5  ( .A1(
        \SB2_1_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_21/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][70] ) );
  NAND4_X1 \SB2_1_23/Component_Function_3/N5  ( .A1(
        \SB2_1_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][63] ) );
  NAND4_X1 \SB2_1_23/Component_Function_4/N5  ( .A1(
        \SB2_1_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_23/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][58] ) );
  NAND4_X1 \SB2_1_24/Component_Function_4/N5  ( .A1(
        \SB2_1_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_24/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][52] ) );
  NAND4_X1 \SB2_1_25/Component_Function_4/N5  ( .A1(
        \SB2_1_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_25/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][46] ) );
  NAND4_X1 \SB2_1_26/Component_Function_4/N5  ( .A1(
        \SB2_1_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_26/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[1][40] ) );
  NAND4_X1 \SB2_1_27/Component_Function_2/N5  ( .A1(
        \SB2_1_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_27/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_1_27/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[1][44] ) );
  NAND4_X1 \SB2_1_27/Component_Function_3/N5  ( .A1(
        \SB2_1_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][39] ) );
  NAND4_X1 \SB2_1_28/Component_Function_3/N5  ( .A1(
        \SB2_1_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_28/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][33] ) );
  NAND4_X1 \SB2_1_30/Component_Function_3/N5  ( .A1(
        \SB2_1_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_30/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][21] ) );
  NAND4_X1 \SB1_2_0/Component_Function_3/N5  ( .A1(
        \SB1_2_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_0/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][9] ) );
  NAND4_X1 \SB1_2_0/Component_Function_4/N5  ( .A1(
        \SB1_2_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_0/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][4] ) );
  NAND4_X1 \SB1_2_1/Component_Function_4/N5  ( .A1(
        \SB1_2_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_1/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][190] ) );
  NAND4_X1 \SB1_2_2/Component_Function_2/N5  ( .A1(
        \SB1_2_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_2/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_2/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[2][2] ) );
  NAND4_X1 \SB1_2_2/Component_Function_3/N5  ( .A1(
        \SB1_2_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_2/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][189] ) );
  NAND4_X1 \SB1_2_2/Component_Function_4/N5  ( .A1(
        \SB1_2_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_2/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][184] ) );
  NAND4_X1 \SB1_2_3/Component_Function_3/N5  ( .A1(
        \SB1_2_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_3/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][183] ) );
  NAND4_X1 \SB1_2_3/Component_Function_4/N5  ( .A1(
        \SB1_2_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_3/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][178] ) );
  NAND4_X1 \SB1_2_4/Component_Function_3/N5  ( .A1(
        \SB1_2_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][177] ) );
  NAND4_X1 \SB1_2_4/Component_Function_4/N5  ( .A1(
        \SB1_2_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_4/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][172] ) );
  NAND4_X1 \SB1_2_5/Component_Function_3/N5  ( .A1(
        \SB1_2_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][171] ) );
  NAND4_X1 \SB1_2_5/Component_Function_4/N5  ( .A1(
        \SB1_2_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_5/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][166] ) );
  NAND4_X1 \SB1_2_6/Component_Function_3/N5  ( .A1(
        \SB1_2_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][165] ) );
  NAND4_X1 \SB1_2_6/Component_Function_4/N5  ( .A1(
        \SB1_2_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_6/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][160] ) );
  NAND4_X1 \SB1_2_7/Component_Function_3/N5  ( .A1(
        \SB1_2_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_7/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][159] ) );
  NAND4_X1 \SB1_2_7/Component_Function_4/N5  ( .A1(
        \SB1_2_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_7/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_7/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][154] ) );
  NAND4_X1 \SB1_2_8/Component_Function_3/N5  ( .A1(
        \SB1_2_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_8/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_8/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][153] ) );
  NAND4_X1 \SB1_2_8/Component_Function_4/N5  ( .A1(
        \SB1_2_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_8/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_8/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][148] ) );
  NAND4_X1 \SB1_2_9/Component_Function_3/N5  ( .A1(
        \SB1_2_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_9/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][147] ) );
  NAND4_X1 \SB1_2_9/Component_Function_4/N5  ( .A1(
        \SB1_2_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_9/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][142] ) );
  NAND4_X1 \SB1_2_10/Component_Function_3/N5  ( .A1(
        \SB1_2_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_10/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_10/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][141] ) );
  NAND4_X1 \SB1_2_10/Component_Function_4/N5  ( .A1(
        \SB1_2_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_10/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][136] ) );
  NAND4_X1 \SB1_2_11/Component_Function_3/N5  ( .A1(
        \SB1_2_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_11/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][135] ) );
  NAND4_X1 \SB1_2_11/Component_Function_4/N5  ( .A1(
        \SB1_2_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_11/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][130] ) );
  NAND4_X1 \SB1_2_12/Component_Function_2/N5  ( .A1(
        \SB1_2_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_12/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[2][134] ) );
  NAND4_X1 \SB1_2_12/Component_Function_3/N5  ( .A1(
        \SB1_2_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_12/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][129] ) );
  NAND4_X1 \SB1_2_12/Component_Function_4/N5  ( .A1(
        \SB1_2_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_12/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][124] ) );
  NAND4_X1 \SB1_2_13/Component_Function_3/N5  ( .A1(
        \SB1_2_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][123] ) );
  NAND4_X1 \SB1_2_13/Component_Function_4/N5  ( .A1(
        \SB1_2_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_13/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][118] ) );
  NAND4_X1 \SB1_2_14/Component_Function_3/N5  ( .A1(
        \SB1_2_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][117] ) );
  NAND4_X1 \SB1_2_15/Component_Function_3/N5  ( .A1(
        \SB1_2_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][111] ) );
  NAND4_X1 \SB1_2_15/Component_Function_4/N5  ( .A1(
        \SB1_2_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_15/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][106] ) );
  NAND4_X1 \SB1_2_16/Component_Function_3/N5  ( .A1(
        \SB1_2_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_16/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][105] ) );
  NAND4_X1 \SB1_2_16/Component_Function_4/N5  ( .A1(
        \SB1_2_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_16/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][100] ) );
  NAND4_X1 \SB1_2_17/Component_Function_2/N5  ( .A1(
        \SB1_2_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_17/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[2][104] ) );
  NAND4_X1 \SB1_2_17/Component_Function_3/N5  ( .A1(
        \SB1_2_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_17/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][99] ) );
  NAND4_X1 \SB1_2_17/Component_Function_4/N5  ( .A1(
        \SB1_2_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][94] ) );
  NAND4_X1 \SB1_2_18/Component_Function_3/N5  ( .A1(
        \SB1_2_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][93] ) );
  NAND4_X1 \SB1_2_18/Component_Function_4/N5  ( .A1(
        \SB1_2_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_18/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][88] ) );
  NAND4_X1 \SB1_2_19/Component_Function_3/N5  ( .A1(
        \SB1_2_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_19/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][87] ) );
  NAND4_X1 \SB1_2_20/Component_Function_2/N5  ( .A1(
        \SB1_2_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_2_20/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[2][86] ) );
  NAND4_X1 \SB1_2_20/Component_Function_3/N5  ( .A1(
        \SB1_2_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][81] ) );
  NAND4_X1 \SB1_2_20/Component_Function_4/N5  ( .A1(
        \SB1_2_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][76] ) );
  NAND4_X1 \SB1_2_21/Component_Function_3/N5  ( .A1(
        \SB1_2_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_21/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][75] ) );
  NAND4_X1 \SB1_2_21/Component_Function_4/N5  ( .A1(
        \SB1_2_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_21/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][70] ) );
  NAND4_X1 \SB1_2_22/Component_Function_2/N5  ( .A1(
        \SB1_2_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_22/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_22/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[2][74] ) );
  NAND4_X1 \SB1_2_22/Component_Function_3/N5  ( .A1(
        \SB1_2_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_22/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][69] ) );
  NAND4_X1 \SB1_2_23/Component_Function_3/N5  ( .A1(
        \SB1_2_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][63] ) );
  NAND4_X1 \SB1_2_23/Component_Function_4/N5  ( .A1(
        \SB1_2_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_23/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][58] ) );
  NAND4_X1 \SB1_2_24/Component_Function_3/N5  ( .A1(
        \SB1_2_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_24/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][57] ) );
  NAND4_X1 \SB1_2_25/Component_Function_3/N5  ( .A1(
        \SB1_2_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_25/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][51] ) );
  NAND4_X1 \SB1_2_26/Component_Function_3/N5  ( .A1(
        \SB1_2_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_26/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][45] ) );
  NAND4_X1 \SB1_2_26/Component_Function_4/N5  ( .A1(
        \SB1_2_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_26/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][40] ) );
  NAND4_X1 \SB1_2_27/Component_Function_3/N5  ( .A1(
        \SB1_2_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][39] ) );
  NAND4_X1 \SB1_2_27/Component_Function_4/N5  ( .A1(
        \SB1_2_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_27/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_27/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][34] ) );
  NAND4_X1 \SB1_2_28/Component_Function_3/N5  ( .A1(
        \SB1_2_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_28/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][33] ) );
  NAND4_X1 \SB1_2_28/Component_Function_4/N5  ( .A1(
        \SB1_2_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_28/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][28] ) );
  NAND4_X1 \SB1_2_29/Component_Function_2/N5  ( .A1(
        \SB1_2_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_29/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[2][32] ) );
  NAND4_X1 \SB1_2_29/Component_Function_3/N5  ( .A1(
        \SB1_2_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_29/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][27] ) );
  NAND4_X1 \SB1_2_29/Component_Function_4/N5  ( .A1(
        \SB1_2_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_29/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][22] ) );
  NAND4_X1 \SB1_2_30/Component_Function_3/N5  ( .A1(
        \SB1_2_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_30/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[2][21] ) );
  NAND4_X1 \SB1_2_30/Component_Function_4/N5  ( .A1(
        \SB1_2_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_30/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][16] ) );
  NAND4_X1 \SB1_2_31/Component_Function_4/N5  ( .A1(
        \SB1_2_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_31/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_31/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[2][10] ) );
  NAND4_X1 \SB2_2_0/Component_Function_3/N5  ( .A1(
        \SB2_2_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_0/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][9] ) );
  NAND4_X1 \SB2_2_3/Component_Function_3/N5  ( .A1(
        \SB2_2_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_3/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][183] ) );
  NAND4_X1 \SB2_2_4/Component_Function_2/N5  ( .A1(
        \SB2_2_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][182] ) );
  NAND4_X1 \SB2_2_6/Component_Function_3/N5  ( .A1(
        \SB2_2_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][165] ) );
  NAND4_X1 \SB2_2_7/Component_Function_2/N5  ( .A1(
        \SB2_2_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_7/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_7/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][164] ) );
  NAND4_X1 \SB2_2_7/Component_Function_4/N5  ( .A1(
        \SB2_2_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_7/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_7/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[2][154] ) );
  NAND4_X1 \SB2_2_12/Component_Function_2/N5  ( .A1(
        \SB2_2_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_12/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][134] ) );
  NAND4_X1 \SB2_2_12/Component_Function_3/N5  ( .A1(
        \SB2_2_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_12/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][129] ) );
  NAND4_X1 \SB2_2_13/Component_Function_2/N5  ( .A1(
        \SB2_2_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][128] ) );
  NAND4_X1 \SB2_2_14/Component_Function_2/N5  ( .A1(
        \SB2_2_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_14/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][122] ) );
  NAND4_X1 \SB2_2_15/Component_Function_3/N5  ( .A1(
        \SB2_2_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][111] ) );
  NAND4_X1 \SB2_2_16/Component_Function_2/N5  ( .A1(
        \SB2_2_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_16/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_16/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][110] ) );
  NAND4_X1 \SB2_2_16/Component_Function_4/N5  ( .A1(
        \SB2_2_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_16/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_16/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[2][100] ) );
  NAND4_X1 \SB2_2_19/Component_Function_2/N5  ( .A1(
        \SB2_2_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_19/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][92] ) );
  NAND4_X1 \SB2_2_21/Component_Function_3/N5  ( .A1(
        \SB2_2_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_21/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][75] ) );
  NAND4_X1 \SB2_2_22/Component_Function_2/N5  ( .A1(
        \SB2_2_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_22/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_22/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][74] ) );
  NAND4_X1 \SB2_2_24/Component_Function_4/N5  ( .A1(
        \SB2_2_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_24/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[2][52] ) );
  NAND4_X1 \SB2_2_28/Component_Function_3/N5  ( .A1(
        \SB2_2_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_28/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][33] ) );
  NAND4_X1 \SB2_2_30/Component_Function_2/N5  ( .A1(
        \SB2_2_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_30/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_30/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[2][26] ) );
  NAND4_X1 \SB2_2_30/Component_Function_4/N5  ( .A1(
        \SB2_2_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_30/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[2][16] ) );
  NAND4_X1 \SB2_2_31/Component_Function_4/N5  ( .A1(
        \SB2_2_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_31/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_31/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[2][10] ) );
  NAND4_X1 \SB1_3_0/Component_Function_2/N5  ( .A1(
        \SB1_3_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][14] ) );
  NAND4_X1 \SB1_3_0/Component_Function_3/N5  ( .A1(
        \SB1_3_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][9] ) );
  NAND4_X1 \SB1_3_1/Component_Function_2/N5  ( .A1(
        \SB1_3_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_1/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_1/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][8] ) );
  NAND4_X1 \SB1_3_1/Component_Function_4/N5  ( .A1(
        \SB1_3_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_1/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][190] ) );
  NAND4_X1 \SB1_3_2/Component_Function_3/N5  ( .A1(
        \SB1_3_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_2/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][189] ) );
  NAND4_X1 \SB1_3_3/Component_Function_3/N5  ( .A1(
        \SB1_3_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_3/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][183] ) );
  NAND4_X1 \SB1_3_3/Component_Function_4/N5  ( .A1(
        \SB1_3_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_3/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][178] ) );
  NAND4_X1 \SB1_3_4/Component_Function_2/N5  ( .A1(
        \SB1_3_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_4/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_4/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][182] ) );
  NAND4_X1 \SB1_3_4/Component_Function_3/N5  ( .A1(
        \SB1_3_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][177] ) );
  NAND4_X1 \SB1_3_4/Component_Function_4/N5  ( .A1(
        \SB1_3_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_4/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][172] ) );
  NAND4_X1 \SB1_3_5/Component_Function_3/N5  ( .A1(
        \SB1_3_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][171] ) );
  NAND4_X1 \SB1_3_6/Component_Function_2/N5  ( .A1(
        \SB1_3_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_6/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][170] ) );
  NAND4_X1 \SB1_3_6/Component_Function_3/N5  ( .A1(
        \SB1_3_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][165] ) );
  NAND4_X1 \SB1_3_7/Component_Function_3/N5  ( .A1(
        \SB1_3_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_7/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][159] ) );
  NAND4_X1 \SB1_3_8/Component_Function_3/N5  ( .A1(
        \SB1_3_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_8/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_8/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][153] ) );
  NAND4_X1 \SB1_3_8/Component_Function_4/N5  ( .A1(
        \SB1_3_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_8/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_8/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][148] ) );
  NAND4_X1 \SB1_3_10/Component_Function_2/N5  ( .A1(
        \SB1_3_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][146] ) );
  NAND4_X1 \SB1_3_10/Component_Function_3/N5  ( .A1(
        \SB1_3_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][141] ) );
  NAND4_X1 \SB1_3_10/Component_Function_4/N5  ( .A1(
        \SB1_3_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][136] ) );
  NAND4_X1 \SB1_3_11/Component_Function_2/N5  ( .A1(
        \SB1_3_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_11/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_11/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][140] ) );
  NAND4_X1 \SB1_3_11/Component_Function_4/N5  ( .A1(
        \SB1_3_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_11/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][130] ) );
  NAND4_X1 \SB1_3_12/Component_Function_2/N5  ( .A1(
        \SB1_3_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_12/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][134] ) );
  NAND4_X1 \SB1_3_13/Component_Function_2/N5  ( .A1(
        \SB1_3_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][128] ) );
  NAND4_X1 \SB1_3_13/Component_Function_3/N5  ( .A1(
        \SB1_3_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][123] ) );
  NAND4_X1 \SB1_3_14/Component_Function_2/N5  ( .A1(
        \SB1_3_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_14/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_14/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][122] ) );
  NAND4_X1 \SB1_3_14/Component_Function_3/N5  ( .A1(
        \SB1_3_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][117] ) );
  NAND4_X1 \SB1_3_15/Component_Function_3/N5  ( .A1(
        \SB1_3_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][111] ) );
  NAND4_X1 \SB1_3_15/Component_Function_4/N5  ( .A1(
        \SB1_3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][106] ) );
  NAND4_X1 \SB1_3_16/Component_Function_2/N5  ( .A1(
        \SB1_3_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_16/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][110] ) );
  NAND4_X1 \SB1_3_16/Component_Function_3/N5  ( .A1(
        \SB1_3_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_16/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][105] ) );
  NAND4_X1 \SB1_3_17/Component_Function_2/N5  ( .A1(
        \SB1_3_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_17/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_17/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][104] ) );
  NAND4_X1 \SB1_3_17/Component_Function_3/N5  ( .A1(
        \SB1_3_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_17/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_17/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][99] ) );
  NAND4_X1 \SB1_3_18/Component_Function_3/N5  ( .A1(
        \SB1_3_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][93] ) );
  NAND4_X1 \SB1_3_18/Component_Function_4/N5  ( .A1(
        \SB1_3_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][88] ) );
  NAND4_X1 \SB1_3_19/Component_Function_2/N5  ( .A1(
        \SB1_3_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_19/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][92] ) );
  NAND4_X1 \SB1_3_20/Component_Function_3/N5  ( .A1(
        \SB1_3_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_20/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][81] ) );
  NAND4_X1 \SB1_3_20/Component_Function_4/N5  ( .A1(
        \SB1_3_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_20/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][76] ) );
  NAND4_X1 \SB1_3_21/Component_Function_2/N5  ( .A1(
        \SB1_3_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_21/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][80] ) );
  NAND4_X1 \SB1_3_21/Component_Function_3/N5  ( .A1(
        \SB1_3_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_21/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][75] ) );
  NAND4_X1 \SB1_3_22/Component_Function_2/N5  ( .A1(
        \SB1_3_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_22/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][74] ) );
  NAND4_X1 \SB1_3_22/Component_Function_3/N5  ( .A1(
        \SB1_3_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_22/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][69] ) );
  NAND4_X1 \SB1_3_23/Component_Function_2/N5  ( .A1(
        \SB1_3_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_23/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_23/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][68] ) );
  NAND4_X1 \SB1_3_23/Component_Function_3/N5  ( .A1(
        \SB1_3_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][63] ) );
  NAND4_X1 \SB1_3_24/Component_Function_3/N5  ( .A1(
        \SB1_3_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][57] ) );
  NAND4_X1 \SB1_3_25/Component_Function_3/N5  ( .A1(
        \SB1_3_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_25/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][51] ) );
  NAND4_X1 \SB1_3_26/Component_Function_3/N5  ( .A1(
        \SB1_3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_26/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][45] ) );
  NAND4_X1 \SB1_3_27/Component_Function_3/N5  ( .A1(
        \SB1_3_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][39] ) );
  NAND4_X1 \SB1_3_28/Component_Function_3/N5  ( .A1(
        \SB1_3_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_28/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][33] ) );
  NAND4_X1 \SB1_3_28/Component_Function_4/N5  ( .A1(
        \SB1_3_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_28/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][28] ) );
  NAND4_X1 \SB1_3_29/Component_Function_2/N5  ( .A1(
        \SB1_3_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_29/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_29/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[3][32] ) );
  NAND4_X1 \SB1_3_29/Component_Function_3/N5  ( .A1(
        \SB1_3_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_29/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_29/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][27] ) );
  NAND4_X1 \SB1_3_30/Component_Function_4/N5  ( .A1(
        \SB1_3_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_30/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][16] ) );
  NAND4_X1 \SB1_3_31/Component_Function_3/N5  ( .A1(
        \SB1_3_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_31/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[3][15] ) );
  NAND4_X1 \SB2_3_4/Component_Function_4/N5  ( .A1(
        \SB2_3_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_4/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][172] ) );
  NAND4_X1 \SB2_3_7/Component_Function_4/N5  ( .A1(
        \SB2_3_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_7/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][154] ) );
  NAND4_X1 \SB2_3_8/Component_Function_2/N5  ( .A1(
        \SB2_3_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_8/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_8/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[3][158] ) );
  NAND4_X1 \SB2_3_8/Component_Function_4/N5  ( .A1(
        \SB2_3_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_8/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_8/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][148] ) );
  NAND4_X1 \SB2_3_10/Component_Function_3/N5  ( .A1(
        \SB2_3_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_10/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_10/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][141] ) );
  NAND4_X1 \SB2_3_14/Component_Function_3/N5  ( .A1(
        \SB2_3_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][117] ) );
  NAND4_X1 \SB2_3_15/Component_Function_3/N5  ( .A1(
        \SB2_3_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][111] ) );
  NAND4_X1 \SB2_3_18/Component_Function_4/N5  ( .A1(
        \SB2_3_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_18/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][88] ) );
  NAND4_X1 \SB2_3_20/Component_Function_4/N5  ( .A1(
        \SB2_3_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_20/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][76] ) );
  NAND4_X1 \SB2_3_22/Component_Function_4/N5  ( .A1(
        \SB2_3_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][64] ) );
  NAND4_X1 \SB2_3_23/Component_Function_2/N5  ( .A1(
        \SB2_3_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_23/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[3][68] ) );
  NAND4_X1 \SB2_3_26/Component_Function_4/N5  ( .A1(
        \SB2_3_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_26/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][40] ) );
  NAND4_X1 \SB2_3_30/Component_Function_3/N5  ( .A1(
        \SB2_3_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_30/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_30/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][21] ) );
  NAND4_X1 \SB2_3_30/Component_Function_4/N5  ( .A1(
        \SB2_3_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_30/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][16] ) );
  NAND4_X1 \SB3_1/Component_Function_2/N5  ( .A1(
        \SB3_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_1/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][8] ) );
  NAND4_X1 \SB3_1/Component_Function_3/N5  ( .A1(
        \SB3_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_1/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][3] ) );
  NAND4_X1 \SB3_1/Component_Function_4/N5  ( .A1(
        \SB3_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_1/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][190] ) );
  NAND4_X1 \SB3_2/Component_Function_3/N5  ( .A1(
        \SB3_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_2/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][189] ) );
  NAND4_X1 \SB3_3/Component_Function_3/N5  ( .A1(
        \SB3_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_3/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][183] ) );
  NAND4_X1 \SB3_3/Component_Function_4/N5  ( .A1(
        \SB3_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_3/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][178] ) );
  NAND4_X1 \SB3_4/Component_Function_3/N5  ( .A1(
        \SB3_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][177] ) );
  NAND4_X1 \SB3_4/Component_Function_4/N5  ( .A1(
        \SB3_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_4/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][172] ) );
  NAND4_X1 \SB3_5/Component_Function_2/N5  ( .A1(
        \SB3_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_5/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][176] ) );
  NAND4_X1 \SB3_5/Component_Function_4/N5  ( .A1(
        \SB3_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_5/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][166] ) );
  NAND4_X1 \SB3_6/Component_Function_2/N5  ( .A1(
        \SB3_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][170] ) );
  NAND4_X1 \SB3_6/Component_Function_3/N5  ( .A1(
        \SB3_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][165] ) );
  NAND4_X1 \SB3_7/Component_Function_2/N5  ( .A1(
        \SB3_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_7/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_7/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][164] ) );
  NAND4_X1 \SB3_7/Component_Function_4/N5  ( .A1(
        \SB3_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_7/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_7/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][154] ) );
  NAND4_X1 \SB3_8/Component_Function_2/N5  ( .A1(
        \SB3_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][158] ) );
  NAND4_X1 \SB3_8/Component_Function_3/N5  ( .A1(
        \SB3_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][153] ) );
  NAND4_X1 \SB3_9/Component_Function_2/N5  ( .A1(
        \SB3_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][152] ) );
  NAND4_X1 \SB3_9/Component_Function_3/N5  ( .A1(
        \SB3_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][147] ) );
  NAND4_X1 \SB3_10/Component_Function_2/N5  ( .A1(
        \SB3_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_10/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][146] ) );
  NAND4_X1 \SB3_10/Component_Function_3/N5  ( .A1(
        \SB3_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_10/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][141] ) );
  NAND4_X1 \SB3_11/Component_Function_2/N5  ( .A1(
        \SB3_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_11/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][140] ) );
  NAND4_X1 \SB3_11/Component_Function_4/N5  ( .A1(
        \SB3_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_11/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][130] ) );
  NAND4_X1 \SB3_12/Component_Function_3/N5  ( .A1(
        \SB3_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_12/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][129] ) );
  NAND4_X1 \SB3_13/Component_Function_2/N5  ( .A1(
        \SB3_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_13/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][128] ) );
  NAND4_X1 \SB3_13/Component_Function_3/N5  ( .A1(
        \SB3_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][123] ) );
  NAND4_X1 \SB3_13/Component_Function_4/N5  ( .A1(
        \SB3_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_13/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][118] ) );
  NAND4_X1 \SB3_14/Component_Function_2/N5  ( .A1(
        \SB3_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_14/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][122] ) );
  NAND4_X1 \SB3_14/Component_Function_4/N5  ( .A1(
        \SB3_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_14/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][112] ) );
  NAND4_X1 \SB3_15/Component_Function_3/N5  ( .A1(
        \SB3_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_15/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][111] ) );
  NAND4_X1 \SB3_16/Component_Function_2/N5  ( .A1(
        \SB3_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_16/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][110] ) );
  NAND4_X1 \SB3_16/Component_Function_3/N5  ( .A1(
        \SB3_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_16/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][105] ) );
  NAND4_X1 \SB3_17/Component_Function_2/N5  ( .A1(
        \SB3_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_17/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][104] ) );
  NAND4_X1 \SB3_17/Component_Function_3/N5  ( .A1(
        \SB3_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_17/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][99] ) );
  NAND4_X1 \SB3_17/Component_Function_4/N5  ( .A1(
        \SB3_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][94] ) );
  NAND4_X1 \SB3_18/Component_Function_2/N5  ( .A1(
        \SB3_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][98] ) );
  NAND4_X1 \SB3_18/Component_Function_3/N5  ( .A1(
        \SB3_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][93] ) );
  NAND4_X1 \SB3_18/Component_Function_4/N5  ( .A1(
        \SB3_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][88] ) );
  NAND4_X1 \SB3_19/Component_Function_2/N5  ( .A1(
        \SB3_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][92] ) );
  NAND4_X1 \SB3_19/Component_Function_3/N5  ( .A1(
        \SB3_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][87] ) );
  NAND4_X1 \SB3_19/Component_Function_4/N5  ( .A1(
        \SB3_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][82] ) );
  NAND4_X1 \SB3_20/Component_Function_4/N5  ( .A1(
        \SB3_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_20/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][76] ) );
  NAND4_X1 \SB3_21/Component_Function_2/N5  ( .A1(
        \SB3_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][80] ) );
  NAND4_X1 \SB3_21/Component_Function_3/N5  ( .A1(
        \SB3_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][75] ) );
  NAND4_X1 \SB3_22/Component_Function_3/N5  ( .A1(
        \SB3_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][69] ) );
  NAND4_X1 \SB3_22/Component_Function_4/N5  ( .A1(
        \SB3_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][64] ) );
  NAND4_X1 \SB3_23/Component_Function_2/N5  ( .A1(
        \SB3_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_23/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_23/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][68] ) );
  NAND4_X1 \SB3_24/Component_Function_2/N5  ( .A1(
        \SB3_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_24/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][62] ) );
  NAND4_X1 \SB3_24/Component_Function_4/N5  ( .A1(
        \SB3_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_24/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][52] ) );
  NAND4_X1 \SB3_25/Component_Function_2/N5  ( .A1(
        \SB3_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_25/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][56] ) );
  NAND4_X1 \SB3_25/Component_Function_3/N5  ( .A1(
        \SB3_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_25/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][51] ) );
  NAND4_X1 \SB3_25/Component_Function_4/N5  ( .A1(
        \SB3_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_25/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][46] ) );
  NAND4_X1 \SB3_26/Component_Function_3/N5  ( .A1(
        \SB3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][45] ) );
  NAND4_X1 \SB3_26/Component_Function_4/N5  ( .A1(
        \SB3_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][40] ) );
  NAND4_X1 \SB3_27/Component_Function_2/N5  ( .A1(
        \SB3_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_27/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_27/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][44] ) );
  NAND4_X1 \SB3_27/Component_Function_3/N5  ( .A1(
        \SB3_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][39] ) );
  NAND4_X1 \SB3_27/Component_Function_4/N5  ( .A1(
        \SB3_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_27/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][34] ) );
  NAND4_X1 \SB3_28/Component_Function_2/N5  ( .A1(
        \SB3_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_28/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[4][38] ) );
  NAND4_X1 \SB3_29/Component_Function_4/N5  ( .A1(
        \SB3_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_29/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][22] ) );
  NAND4_X1 \SB3_30/Component_Function_3/N5  ( .A1(
        \SB3_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_30/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_30/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][21] ) );
  NAND4_X1 \SB3_31/Component_Function_3/N5  ( .A1(
        \SB3_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[4][15] ) );
  NAND4_X1 \SB3_31/Component_Function_4/N5  ( .A1(
        \SB3_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[4][10] ) );
  NAND4_X1 \SB4_5/Component_Function_3/N5  ( .A1(
        \SB4_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI4[4][159] ) );
  NAND4_X1 \SB4_14/Component_Function_3/N5  ( .A1(
        \SB4_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI4[4][105] ) );
  NAND4_X1 \SB4_18/Component_Function_3/N5  ( .A1(
        \SB4_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI4[4][81] ) );
  NAND4_X1 \SB4_19/Component_Function_3/N5  ( .A1(
        \SB4_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_19/Component_Function_3/NAND4_in[3] ), .ZN(\RI4[4][75] ) );
  NAND4_X1 \SB4_23/Component_Function_3/N5  ( .A1(
        \SB4_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI4[4][51] ) );
  NAND4_X1 \SB4_31/Component_Function_3/N5  ( .A1(
        \SB4_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_31/Component_Function_3/NAND4_in[3] ), .ZN(\RI4[4][3] ) );
  NAND4_X1 \SB1_0_0/Component_Function_0/N5  ( .A1(
        \SB1_0_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][24] ) );
  NAND4_X1 \SB1_0_0/Component_Function_1/N5  ( .A1(
        \SB1_0_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][19] ) );
  NAND4_X1 \SB1_0_0/Component_Function_5/N5  ( .A1(
        \SB1_0_0/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_0/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][191] ) );
  NAND4_X1 \SB1_0_1/Component_Function_0/N5  ( .A1(
        \SB1_0_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][18] ) );
  NAND4_X1 \SB1_0_1/Component_Function_5/N5  ( .A1(
        \SB1_0_1/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][185] ) );
  NAND4_X1 \SB1_0_2/Component_Function_0/N5  ( .A1(
        \SB1_0_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_2/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][12] ) );
  NAND4_X1 \SB1_0_2/Component_Function_1/N5  ( .A1(
        \SB1_0_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_2/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][7] ) );
  NAND4_X1 \SB1_0_3/Component_Function_1/N5  ( .A1(
        \SB1_0_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][1] ) );
  NAND4_X1 \SB1_0_3/Component_Function_5/N5  ( .A1(
        \SB1_0_3/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_3/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][173] ) );
  NAND4_X1 \SB1_0_4/Component_Function_0/N5  ( .A1(
        \SB1_0_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][0] ) );
  NAND4_X1 \SB1_0_4/Component_Function_1/N5  ( .A1(
        \SB1_0_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][187] ) );
  NAND4_X1 \SB1_0_4/Component_Function_5/N5  ( .A1(
        \SB1_0_4/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][167] ) );
  NAND4_X1 \SB1_0_5/Component_Function_0/N5  ( .A1(
        \SB1_0_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_5/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][186] ) );
  NAND4_X1 \SB1_0_5/Component_Function_1/N5  ( .A1(
        \SB1_0_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][181] ) );
  NAND4_X1 \SB1_0_6/Component_Function_0/N5  ( .A1(
        \SB1_0_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_6/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][180] ) );
  NAND4_X1 \SB1_0_6/Component_Function_1/N5  ( .A1(
        \SB1_0_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][175] ) );
  NAND4_X1 \SB1_0_7/Component_Function_0/N5  ( .A1(
        \SB1_0_7/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][174] ) );
  NAND4_X1 \SB1_0_7/Component_Function_1/N5  ( .A1(
        \SB1_0_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][169] ) );
  NAND4_X1 \SB1_0_7/Component_Function_5/N5  ( .A1(
        \SB1_0_7/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_7/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][149] ) );
  NAND4_X1 \SB1_0_8/Component_Function_0/N5  ( .A1(
        \SB1_0_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_8/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][168] ) );
  NAND4_X1 \SB1_0_8/Component_Function_1/N5  ( .A1(
        \SB1_0_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][163] ) );
  NAND4_X1 \SB1_0_9/Component_Function_0/N5  ( .A1(
        \SB1_0_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][162] ) );
  NAND4_X1 \SB1_0_9/Component_Function_1/N5  ( .A1(
        \SB1_0_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][157] ) );
  NAND4_X1 \SB1_0_9/Component_Function_5/N5  ( .A1(
        \SB1_0_9/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][137] ) );
  NAND4_X1 \SB1_0_10/Component_Function_0/N5  ( .A1(
        \SB1_0_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][156] ) );
  NAND4_X1 \SB1_0_10/Component_Function_1/N5  ( .A1(
        \SB1_0_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][151] ) );
  NAND4_X1 \SB1_0_10/Component_Function_5/N5  ( .A1(
        \SB1_0_10/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][131] ) );
  NAND4_X1 \SB1_0_11/Component_Function_0/N5  ( .A1(
        \SB1_0_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][150] ) );
  NAND4_X1 \SB1_0_11/Component_Function_1/N5  ( .A1(
        \SB1_0_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][145] ) );
  NAND4_X1 \SB1_0_12/Component_Function_0/N5  ( .A1(
        \SB1_0_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_12/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][144] ) );
  NAND4_X1 \SB1_0_12/Component_Function_1/N5  ( .A1(
        \SB1_0_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_12/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][139] ) );
  NAND4_X1 \SB1_0_12/Component_Function_5/N5  ( .A1(
        \SB1_0_12/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_12/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_12/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][119] ) );
  NAND4_X1 \SB1_0_13/Component_Function_0/N5  ( .A1(
        \SB1_0_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][138] ) );
  NAND4_X1 \SB1_0_13/Component_Function_1/N5  ( .A1(
        \SB1_0_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][133] ) );
  NAND4_X1 \SB1_0_13/Component_Function_5/N5  ( .A1(
        \SB1_0_13/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][113] ) );
  NAND4_X1 \SB1_0_14/Component_Function_0/N5  ( .A1(
        \SB1_0_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][132] ) );
  NAND4_X1 \SB1_0_14/Component_Function_1/N5  ( .A1(
        \SB1_0_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][127] ) );
  NAND4_X1 \SB1_0_14/Component_Function_5/N5  ( .A1(
        \SB1_0_14/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][107] ) );
  NAND4_X1 \SB1_0_15/Component_Function_0/N5  ( .A1(
        \SB1_0_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_15/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][126] ) );
  NAND4_X1 \SB1_0_15/Component_Function_1/N5  ( .A1(
        \SB1_0_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][121] ) );
  NAND4_X1 \SB1_0_16/Component_Function_1/N5  ( .A1(
        \SB1_0_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_16/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][115] ) );
  NAND4_X1 \SB1_0_17/Component_Function_0/N5  ( .A1(
        \SB1_0_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][114] ) );
  NAND4_X1 \SB1_0_17/Component_Function_1/N5  ( .A1(
        \SB1_0_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][109] ) );
  NAND4_X1 \SB1_0_17/Component_Function_5/N5  ( .A1(
        \SB1_0_17/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_17/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][89] ) );
  NAND4_X1 \SB1_0_18/Component_Function_1/N5  ( .A1(
        \SB1_0_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_18/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][103] ) );
  NAND4_X1 \SB1_0_19/Component_Function_0/N5  ( .A1(
        \SB1_0_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][102] ) );
  NAND4_X1 \SB1_0_19/Component_Function_5/N5  ( .A1(
        \SB1_0_19/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_19/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_19/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][77] ) );
  NAND4_X1 \SB1_0_20/Component_Function_0/N5  ( .A1(
        \SB1_0_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_20/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][96] ) );
  NAND4_X1 \SB1_0_20/Component_Function_1/N5  ( .A1(
        \SB1_0_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_20/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][91] ) );
  NAND4_X1 \SB1_0_21/Component_Function_0/N5  ( .A1(
        \SB1_0_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_21/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][90] ) );
  NAND4_X1 \SB1_0_21/Component_Function_1/N5  ( .A1(
        \SB1_0_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_21/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][85] ) );
  NAND4_X1 \SB1_0_22/Component_Function_0/N5  ( .A1(
        \SB1_0_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][84] ) );
  NAND4_X1 \SB1_0_22/Component_Function_5/N5  ( .A1(
        \SB1_0_22/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_22/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_22/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][59] ) );
  NAND4_X1 \SB1_0_23/Component_Function_0/N5  ( .A1(
        \SB1_0_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][78] ) );
  NAND4_X1 \SB1_0_23/Component_Function_1/N5  ( .A1(
        \SB1_0_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][73] ) );
  NAND4_X1 \SB1_0_24/Component_Function_0/N5  ( .A1(
        \SB1_0_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_24/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][72] ) );
  NAND4_X1 \SB1_0_24/Component_Function_1/N5  ( .A1(
        \SB1_0_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][67] ) );
  NAND4_X1 \SB1_0_25/Component_Function_1/N5  ( .A1(
        \SB1_0_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][61] ) );
  NAND4_X1 \SB1_0_26/Component_Function_0/N5  ( .A1(
        \SB1_0_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_26/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][60] ) );
  NAND4_X1 \SB1_0_26/Component_Function_1/N5  ( .A1(
        \SB1_0_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][55] ) );
  NAND4_X1 \SB1_0_27/Component_Function_0/N5  ( .A1(
        \SB1_0_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][54] ) );
  NAND4_X1 \SB1_0_27/Component_Function_1/N5  ( .A1(
        \SB1_0_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][49] ) );
  NAND4_X1 \SB1_0_27/Component_Function_5/N5  ( .A1(
        \SB1_0_27/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][29] ) );
  NAND4_X1 \SB1_0_28/Component_Function_0/N5  ( .A1(
        \SB1_0_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][48] ) );
  NAND4_X1 \SB1_0_28/Component_Function_1/N5  ( .A1(
        \SB1_0_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][43] ) );
  NAND4_X1 \SB1_0_28/Component_Function_5/N5  ( .A1(
        \SB1_0_28/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_28/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][23] ) );
  NAND4_X1 \SB1_0_29/Component_Function_0/N5  ( .A1(
        \SB1_0_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][42] ) );
  NAND4_X1 \SB1_0_29/Component_Function_1/N5  ( .A1(
        \SB1_0_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][37] ) );
  NAND4_X1 \SB1_0_30/Component_Function_0/N5  ( .A1(
        \SB1_0_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][36] ) );
  NAND4_X1 \SB1_0_30/Component_Function_1/N5  ( .A1(
        \SB1_0_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][31] ) );
  NAND4_X1 \SB1_0_30/Component_Function_5/N5  ( .A1(
        \SB1_0_30/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][11] ) );
  NAND4_X1 \SB1_0_31/Component_Function_0/N5  ( .A1(
        \SB1_0_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[0][30] ) );
  NAND4_X1 \SB1_0_31/Component_Function_1/N5  ( .A1(
        \SB1_0_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][25] ) );
  NAND4_X1 \SB1_0_31/Component_Function_5/N5  ( .A1(
        \SB1_0_31/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][5] ) );
  NAND4_X1 \SB2_0_0/Component_Function_0/N5  ( .A1(
        \SB2_0_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][24] ) );
  NAND4_X1 \SB2_0_0/Component_Function_1/N5  ( .A1(
        \SB2_0_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][19] ) );
  NAND4_X1 \SB2_0_1/Component_Function_0/N5  ( .A1(
        \SB2_0_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_1/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][18] ) );
  NAND4_X1 \SB2_0_1/Component_Function_1/N5  ( .A1(
        \SB2_0_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_1/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][13] ) );
  NAND4_X1 \SB2_0_2/Component_Function_0/N5  ( .A1(
        \SB2_0_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_2/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][12] ) );
  NAND4_X1 \SB2_0_2/Component_Function_1/N5  ( .A1(
        \SB2_0_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_2/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][7] ) );
  NAND4_X1 \SB2_0_4/Component_Function_0/N5  ( .A1(
        \SB2_0_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_4/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][0] ) );
  NAND4_X1 \SB2_0_4/Component_Function_1/N5  ( .A1(
        \SB2_0_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][187] ) );
  NAND4_X1 \SB2_0_5/Component_Function_0/N5  ( .A1(
        \SB2_0_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_5/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][186] ) );
  NAND4_X1 \SB2_0_5/Component_Function_1/N5  ( .A1(
        \SB2_0_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][181] ) );
  NAND4_X1 \SB2_0_6/Component_Function_0/N5  ( .A1(
        \SB2_0_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][180] ) );
  NAND4_X1 \SB2_0_6/Component_Function_1/N5  ( .A1(
        \SB2_0_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][175] ) );
  NAND4_X1 \SB2_0_8/Component_Function_0/N5  ( .A1(
        \SB2_0_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_8/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][168] ) );
  NAND4_X1 \SB2_0_9/Component_Function_0/N5  ( .A1(
        \SB2_0_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][162] ) );
  NAND4_X1 \SB2_0_10/Component_Function_1/N5  ( .A1(
        \SB2_0_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][151] ) );
  NAND4_X1 \SB2_0_12/Component_Function_0/N5  ( .A1(
        \SB2_0_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][144] ) );
  NAND4_X1 \SB2_0_12/Component_Function_1/N5  ( .A1(
        \SB2_0_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][139] ) );
  NAND4_X1 \SB2_0_13/Component_Function_0/N5  ( .A1(
        \SB2_0_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][138] ) );
  NAND4_X1 \SB2_0_13/Component_Function_1/N5  ( .A1(
        \SB2_0_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][133] ) );
  NAND4_X1 \SB2_0_14/Component_Function_0/N5  ( .A1(
        \SB2_0_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_14/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][132] ) );
  NAND4_X1 \SB2_0_14/Component_Function_1/N5  ( .A1(
        \SB2_0_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_14/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][127] ) );
  NAND4_X1 \SB2_0_15/Component_Function_1/N5  ( .A1(
        \SB2_0_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][121] ) );
  NAND4_X1 \SB2_0_16/Component_Function_0/N5  ( .A1(
        \SB2_0_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_16/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][120] ) );
  NAND4_X1 \SB2_0_16/Component_Function_1/N5  ( .A1(
        \SB2_0_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_16/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][115] ) );
  NAND4_X1 \SB2_0_17/Component_Function_0/N5  ( .A1(
        \SB2_0_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][114] ) );
  NAND4_X1 \SB2_0_17/Component_Function_1/N5  ( .A1(
        \SB2_0_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][109] ) );
  NAND4_X1 \SB2_0_18/Component_Function_0/N5  ( .A1(
        \SB2_0_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_18/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][108] ) );
  NAND4_X1 \SB2_0_18/Component_Function_1/N5  ( .A1(
        \SB2_0_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_18/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][103] ) );
  NAND4_X1 \SB2_0_19/Component_Function_0/N5  ( .A1(
        \SB2_0_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][102] ) );
  NAND4_X1 \SB2_0_19/Component_Function_1/N5  ( .A1(
        \SB2_0_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_19/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][97] ) );
  NAND4_X1 \SB2_0_20/Component_Function_0/N5  ( .A1(
        \SB2_0_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][96] ) );
  NAND4_X1 \SB2_0_20/Component_Function_1/N5  ( .A1(
        \SB2_0_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][91] ) );
  NAND4_X1 \SB2_0_21/Component_Function_0/N5  ( .A1(
        \SB2_0_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_21/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][90] ) );
  NAND4_X1 \SB2_0_22/Component_Function_0/N5  ( .A1(
        \SB2_0_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][84] ) );
  NAND4_X1 \SB2_0_22/Component_Function_1/N5  ( .A1(
        \SB2_0_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][79] ) );
  NAND4_X1 \SB2_0_23/Component_Function_1/N5  ( .A1(
        \SB2_0_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][73] ) );
  NAND4_X1 \SB2_0_24/Component_Function_0/N5  ( .A1(
        \SB2_0_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_24/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][72] ) );
  NAND4_X1 \SB2_0_24/Component_Function_1/N5  ( .A1(
        \SB2_0_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][67] ) );
  NAND4_X1 \SB2_0_25/Component_Function_1/N5  ( .A1(
        \SB2_0_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][61] ) );
  NAND4_X1 \SB2_0_26/Component_Function_1/N5  ( .A1(
        \SB2_0_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][55] ) );
  NAND4_X1 \SB2_0_27/Component_Function_0/N5  ( .A1(
        \SB2_0_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_27/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][54] ) );
  NAND4_X1 \SB2_0_27/Component_Function_1/N5  ( .A1(
        \SB2_0_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][49] ) );
  NAND4_X1 \SB2_0_28/Component_Function_0/N5  ( .A1(
        \SB2_0_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][48] ) );
  NAND4_X1 \SB2_0_28/Component_Function_1/N5  ( .A1(
        \SB2_0_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][43] ) );
  NAND4_X1 \SB2_0_29/Component_Function_0/N5  ( .A1(
        \SB2_0_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][42] ) );
  NAND4_X1 \SB2_0_29/Component_Function_1/N5  ( .A1(
        \SB2_0_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][37] ) );
  NAND4_X1 \SB2_0_30/Component_Function_0/N5  ( .A1(
        \SB2_0_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][36] ) );
  NAND4_X1 \SB2_0_30/Component_Function_1/N5  ( .A1(
        \SB2_0_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_30/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][31] ) );
  NAND4_X1 \SB2_0_31/Component_Function_0/N5  ( .A1(
        \SB2_0_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][30] ) );
  NAND4_X1 \SB2_0_31/Component_Function_1/N5  ( .A1(
        \SB2_0_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_31/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][25] ) );
  NAND4_X1 \SB1_1_0/Component_Function_0/N5  ( .A1(
        \SB1_1_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][24] ) );
  NAND4_X1 \SB1_1_0/Component_Function_1/N5  ( .A1(
        \SB1_1_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][19] ) );
  NAND4_X1 \SB1_1_1/Component_Function_1/N5  ( .A1(
        \SB1_1_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_1/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][13] ) );
  NAND4_X1 \SB1_1_2/Component_Function_0/N5  ( .A1(
        \SB1_1_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_2/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][12] ) );
  NAND4_X1 \SB1_1_3/Component_Function_0/N5  ( .A1(
        \SB1_1_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][6] ) );
  NAND4_X1 \SB1_1_3/Component_Function_1/N5  ( .A1(
        \SB1_1_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][1] ) );
  NAND4_X1 \SB1_1_4/Component_Function_0/N5  ( .A1(
        \SB1_1_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_4/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][0] ) );
  NAND4_X1 \SB1_1_4/Component_Function_1/N5  ( .A1(
        \SB1_1_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][187] ) );
  NAND4_X1 \SB1_1_5/Component_Function_0/N5  ( .A1(
        \SB1_1_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][186] ) );
  NAND4_X1 \SB1_1_5/Component_Function_1/N5  ( .A1(
        \SB1_1_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][181] ) );
  NAND4_X1 \SB1_1_6/Component_Function_0/N5  ( .A1(
        \SB1_1_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_6/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][180] ) );
  NAND4_X1 \SB1_1_6/Component_Function_1/N5  ( .A1(
        \SB1_1_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][175] ) );
  NAND4_X1 \SB1_1_7/Component_Function_0/N5  ( .A1(
        \SB1_1_7/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_7/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][174] ) );
  NAND4_X1 \SB1_1_7/Component_Function_1/N5  ( .A1(
        \SB1_1_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][169] ) );
  NAND4_X1 \SB1_1_8/Component_Function_0/N5  ( .A1(
        \SB1_1_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_8/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][168] ) );
  NAND4_X1 \SB1_1_8/Component_Function_1/N5  ( .A1(
        \SB1_1_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][163] ) );
  NAND4_X1 \SB1_1_9/Component_Function_0/N5  ( .A1(
        \SB1_1_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][162] ) );
  NAND4_X1 \SB1_1_9/Component_Function_1/N5  ( .A1(
        \SB1_1_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][157] ) );
  NAND4_X1 \SB1_1_10/Component_Function_0/N5  ( .A1(
        \SB1_1_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_10/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][156] ) );
  NAND4_X1 \SB1_1_10/Component_Function_1/N5  ( .A1(
        \SB1_1_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][151] ) );
  NAND4_X1 \SB1_1_11/Component_Function_0/N5  ( .A1(
        \SB1_1_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][150] ) );
  NAND4_X1 \SB1_1_11/Component_Function_1/N5  ( .A1(
        \SB1_1_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][145] ) );
  NAND4_X1 \SB1_1_13/Component_Function_0/N5  ( .A1(
        \SB1_1_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][138] ) );
  NAND4_X1 \SB1_1_13/Component_Function_1/N5  ( .A1(
        \SB1_1_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][133] ) );
  NAND4_X1 \SB1_1_14/Component_Function_0/N5  ( .A1(
        \SB1_1_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][132] ) );
  NAND4_X1 \SB1_1_14/Component_Function_1/N5  ( .A1(
        \SB1_1_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][127] ) );
  NAND4_X1 \SB1_1_15/Component_Function_1/N5  ( .A1(
        \SB1_1_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][121] ) );
  NAND4_X1 \SB1_1_16/Component_Function_0/N5  ( .A1(
        \SB1_1_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_16/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][120] ) );
  NAND4_X1 \SB1_1_16/Component_Function_1/N5  ( .A1(
        \SB1_1_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_16/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][115] ) );
  NAND4_X1 \SB1_1_17/Component_Function_0/N5  ( .A1(
        \SB1_1_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][114] ) );
  NAND4_X1 \SB1_1_17/Component_Function_1/N5  ( .A1(
        \SB1_1_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][109] ) );
  NAND4_X1 \SB1_1_18/Component_Function_0/N5  ( .A1(
        \SB1_1_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_18/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][108] ) );
  NAND4_X1 \SB1_1_19/Component_Function_0/N5  ( .A1(
        \SB1_1_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][102] ) );
  NAND4_X1 \SB1_1_19/Component_Function_1/N5  ( .A1(
        \SB1_1_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][97] ) );
  NAND4_X1 \SB1_1_20/Component_Function_0/N5  ( .A1(
        \SB1_1_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_20/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][96] ) );
  NAND4_X1 \SB1_1_20/Component_Function_1/N5  ( .A1(
        \SB1_1_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_20/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][91] ) );
  NAND4_X1 \SB1_1_21/Component_Function_0/N5  ( .A1(
        \SB1_1_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_21/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][90] ) );
  NAND4_X1 \SB1_1_22/Component_Function_0/N5  ( .A1(
        \SB1_1_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][84] ) );
  NAND4_X1 \SB1_1_22/Component_Function_1/N5  ( .A1(
        \SB1_1_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][79] ) );
  NAND4_X1 \SB1_1_23/Component_Function_0/N5  ( .A1(
        \SB1_1_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_23/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][78] ) );
  NAND4_X1 \SB1_1_23/Component_Function_1/N5  ( .A1(
        \SB1_1_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][73] ) );
  NAND4_X1 \SB1_1_24/Component_Function_0/N5  ( .A1(
        \SB1_1_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_24/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][72] ) );
  NAND4_X1 \SB1_1_25/Component_Function_0/N5  ( .A1(
        \SB1_1_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_25/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][66] ) );
  NAND4_X1 \SB1_1_25/Component_Function_1/N5  ( .A1(
        \SB1_1_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][61] ) );
  NAND4_X1 \SB1_1_26/Component_Function_0/N5  ( .A1(
        \SB1_1_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_26/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][60] ) );
  NAND4_X1 \SB1_1_26/Component_Function_1/N5  ( .A1(
        \SB1_1_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][55] ) );
  NAND4_X1 \SB1_1_27/Component_Function_0/N5  ( .A1(
        \SB1_1_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_27/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][54] ) );
  NAND4_X1 \SB1_1_27/Component_Function_1/N5  ( .A1(
        \SB1_1_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][49] ) );
  NAND4_X1 \SB1_1_28/Component_Function_0/N5  ( .A1(
        \SB1_1_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][48] ) );
  NAND4_X1 \SB1_1_28/Component_Function_1/N5  ( .A1(
        \SB1_1_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][43] ) );
  NAND4_X1 \SB1_1_29/Component_Function_0/N5  ( .A1(
        \SB1_1_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][42] ) );
  NAND4_X1 \SB1_1_29/Component_Function_1/N5  ( .A1(
        \SB1_1_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][37] ) );
  NAND4_X1 \SB1_1_30/Component_Function_0/N5  ( .A1(
        \SB1_1_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][36] ) );
  NAND4_X1 \SB1_1_31/Component_Function_0/N5  ( .A1(
        \SB1_1_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[1][30] ) );
  NAND4_X1 \SB1_1_31/Component_Function_1/N5  ( .A1(
        \SB1_1_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_31/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[1][25] ) );
  NAND4_X1 \SB2_1_0/Component_Function_0/N5  ( .A1(
        \SB2_1_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][24] ) );
  NAND4_X1 \SB2_1_0/Component_Function_1/N5  ( .A1(
        \SB2_1_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][19] ) );
  NAND4_X1 \SB2_1_1/Component_Function_0/N5  ( .A1(
        \SB2_1_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_1/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][18] ) );
  NAND4_X1 \SB2_1_1/Component_Function_1/N5  ( .A1(
        \SB2_1_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_1/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][13] ) );
  NAND4_X1 \SB2_1_2/Component_Function_0/N5  ( .A1(
        \SB2_1_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_2/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][12] ) );
  NAND4_X1 \SB2_1_2/Component_Function_1/N5  ( .A1(
        \SB2_1_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_2/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][7] ) );
  NAND4_X1 \SB2_1_3/Component_Function_0/N5  ( .A1(
        \SB2_1_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_3/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][6] ) );
  NAND4_X1 \SB2_1_4/Component_Function_0/N5  ( .A1(
        \SB2_1_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_4/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][0] ) );
  NAND4_X1 \SB2_1_4/Component_Function_1/N5  ( .A1(
        \SB2_1_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][187] ) );
  NAND4_X1 \SB2_1_5/Component_Function_0/N5  ( .A1(
        \SB2_1_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_5/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][186] ) );
  NAND4_X1 \SB2_1_5/Component_Function_1/N5  ( .A1(
        \SB2_1_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][181] ) );
  NAND4_X1 \SB2_1_6/Component_Function_0/N5  ( .A1(
        \SB2_1_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_6/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][180] ) );
  NAND4_X1 \SB2_1_6/Component_Function_1/N5  ( .A1(
        \SB2_1_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][175] ) );
  NAND4_X1 \SB2_1_7/Component_Function_1/N5  ( .A1(
        \SB2_1_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][169] ) );
  NAND4_X1 \SB2_1_8/Component_Function_0/N5  ( .A1(
        \SB2_1_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_8/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][168] ) );
  NAND4_X1 \SB2_1_8/Component_Function_1/N5  ( .A1(
        \SB2_1_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][163] ) );
  NAND4_X1 \SB2_1_9/Component_Function_0/N5  ( .A1(
        \SB2_1_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][162] ) );
  NAND4_X1 \SB2_1_9/Component_Function_1/N5  ( .A1(
        \SB2_1_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][157] ) );
  NAND4_X1 \SB2_1_10/Component_Function_0/N5  ( .A1(
        \SB2_1_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_10/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][156] ) );
  NAND4_X1 \SB2_1_10/Component_Function_1/N5  ( .A1(
        \SB2_1_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][151] ) );
  NAND4_X1 \SB2_1_11/Component_Function_0/N5  ( .A1(
        \SB2_1_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][150] ) );
  NAND4_X1 \SB2_1_11/Component_Function_1/N5  ( .A1(
        \SB2_1_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][145] ) );
  NAND4_X1 \SB2_1_12/Component_Function_0/N5  ( .A1(
        \SB2_1_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_12/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][144] ) );
  NAND4_X1 \SB2_1_12/Component_Function_1/N5  ( .A1(
        \SB2_1_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_12/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][139] ) );
  NAND4_X1 \SB2_1_13/Component_Function_1/N5  ( .A1(
        \SB2_1_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][133] ) );
  NAND4_X1 \SB2_1_15/Component_Function_0/N5  ( .A1(
        \SB2_1_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_15/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][126] ) );
  NAND4_X1 \SB2_1_16/Component_Function_0/N5  ( .A1(
        \SB2_1_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_16/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][120] ) );
  NAND4_X1 \SB2_1_17/Component_Function_0/N5  ( .A1(
        \SB2_1_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][114] ) );
  NAND4_X1 \SB2_1_17/Component_Function_1/N5  ( .A1(
        \SB2_1_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][109] ) );
  NAND4_X1 \SB2_1_18/Component_Function_0/N5  ( .A1(
        \SB2_1_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][108] ) );
  NAND4_X1 \SB2_1_18/Component_Function_1/N5  ( .A1(
        \SB2_1_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][103] ) );
  NAND4_X1 \SB2_1_19/Component_Function_0/N5  ( .A1(
        \SB2_1_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][102] ) );
  NAND4_X1 \SB2_1_20/Component_Function_1/N5  ( .A1(
        \SB2_1_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_20/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][91] ) );
  NAND4_X1 \SB2_1_21/Component_Function_0/N5  ( .A1(
        \SB2_1_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_21/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][90] ) );
  NAND4_X1 \SB2_1_21/Component_Function_1/N5  ( .A1(
        \SB2_1_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_21/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][85] ) );
  NAND4_X1 \SB2_1_22/Component_Function_0/N5  ( .A1(
        \SB2_1_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][84] ) );
  NAND4_X1 \SB2_1_22/Component_Function_1/N5  ( .A1(
        \SB2_1_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][79] ) );
  NAND4_X1 \SB2_1_23/Component_Function_0/N5  ( .A1(
        \SB2_1_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_23/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][78] ) );
  NAND4_X1 \SB2_1_23/Component_Function_1/N5  ( .A1(
        \SB2_1_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][73] ) );
  NAND4_X1 \SB2_1_24/Component_Function_0/N5  ( .A1(
        \SB2_1_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_24/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][72] ) );
  NAND4_X1 \SB2_1_24/Component_Function_1/N5  ( .A1(
        \SB2_1_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][67] ) );
  NAND4_X1 \SB2_1_25/Component_Function_1/N5  ( .A1(
        \SB2_1_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][61] ) );
  NAND4_X1 \SB2_1_26/Component_Function_0/N5  ( .A1(
        \SB2_1_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_26/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][60] ) );
  NAND4_X1 \SB2_1_27/Component_Function_0/N5  ( .A1(
        \SB2_1_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_27/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][54] ) );
  NAND4_X1 \SB2_1_27/Component_Function_1/N5  ( .A1(
        \SB2_1_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][49] ) );
  NAND4_X1 \SB2_1_28/Component_Function_0/N5  ( .A1(
        \SB2_1_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][48] ) );
  NAND4_X1 \SB2_1_28/Component_Function_1/N5  ( .A1(
        \SB2_1_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][43] ) );
  NAND4_X1 \SB2_1_29/Component_Function_0/N5  ( .A1(
        \SB2_1_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][42] ) );
  NAND4_X1 \SB2_1_30/Component_Function_0/N5  ( .A1(
        \SB2_1_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][36] ) );
  NAND4_X1 \SB2_1_30/Component_Function_1/N5  ( .A1(
        \SB2_1_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_30/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[1][31] ) );
  NAND4_X1 \SB2_1_31/Component_Function_0/N5  ( .A1(
        \SB2_1_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][30] ) );
  NAND4_X1 \SB1_2_0/Component_Function_0/N5  ( .A1(
        \SB1_2_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][24] ) );
  NAND4_X1 \SB1_2_0/Component_Function_1/N5  ( .A1(
        \SB1_2_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][19] ) );
  NAND4_X1 \SB1_2_1/Component_Function_0/N5  ( .A1(
        \SB1_2_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_1/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][18] ) );
  NAND4_X1 \SB1_2_1/Component_Function_1/N5  ( .A1(
        \SB1_2_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_1/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][13] ) );
  NAND4_X1 \SB1_2_3/Component_Function_0/N5  ( .A1(
        \SB1_2_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_3/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][6] ) );
  NAND4_X1 \SB1_2_3/Component_Function_1/N5  ( .A1(
        \SB1_2_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][1] ) );
  NAND4_X1 \SB1_2_4/Component_Function_1/N5  ( .A1(
        \SB1_2_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][187] ) );
  NAND4_X1 \SB1_2_5/Component_Function_0/N5  ( .A1(
        \SB1_2_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_5/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][186] ) );
  NAND4_X1 \SB1_2_5/Component_Function_1/N5  ( .A1(
        \SB1_2_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][181] ) );
  NAND4_X1 \SB1_2_6/Component_Function_0/N5  ( .A1(
        \SB1_2_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_6/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][180] ) );
  NAND4_X1 \SB1_2_6/Component_Function_1/N5  ( .A1(
        \SB1_2_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][175] ) );
  NAND4_X1 \SB1_2_7/Component_Function_1/N5  ( .A1(
        \SB1_2_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][169] ) );
  NAND4_X1 \SB1_2_8/Component_Function_1/N5  ( .A1(
        \SB1_2_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][163] ) );
  NAND4_X1 \SB1_2_9/Component_Function_0/N5  ( .A1(
        \SB1_2_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][162] ) );
  NAND4_X1 \SB1_2_9/Component_Function_1/N5  ( .A1(
        \SB1_2_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][157] ) );
  NAND4_X1 \SB1_2_10/Component_Function_1/N5  ( .A1(
        \SB1_2_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][151] ) );
  NAND4_X1 \SB1_2_11/Component_Function_0/N5  ( .A1(
        \SB1_2_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][150] ) );
  NAND4_X1 \SB1_2_11/Component_Function_1/N5  ( .A1(
        \SB1_2_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][145] ) );
  NAND4_X1 \SB1_2_12/Component_Function_1/N5  ( .A1(
        \SB1_2_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_12/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][139] ) );
  NAND4_X1 \SB1_2_13/Component_Function_0/N5  ( .A1(
        \SB1_2_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][138] ) );
  NAND4_X1 \SB1_2_13/Component_Function_1/N5  ( .A1(
        \SB1_2_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][133] ) );
  NAND4_X1 \SB1_2_14/Component_Function_0/N5  ( .A1(
        \SB1_2_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_14/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][132] ) );
  NAND4_X1 \SB1_2_14/Component_Function_1/N5  ( .A1(
        \SB1_2_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_14/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][127] ) );
  NAND4_X1 \SB1_2_15/Component_Function_0/N5  ( .A1(
        \SB1_2_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_15/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][126] ) );
  NAND4_X1 \SB1_2_15/Component_Function_1/N5  ( .A1(
        \SB1_2_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][121] ) );
  NAND4_X1 \SB1_2_16/Component_Function_0/N5  ( .A1(
        \SB1_2_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_16/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][120] ) );
  NAND4_X1 \SB1_2_16/Component_Function_1/N5  ( .A1(
        \SB1_2_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_16/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][115] ) );
  NAND4_X1 \SB1_2_17/Component_Function_0/N5  ( .A1(
        \SB1_2_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][114] ) );
  NAND4_X1 \SB1_2_17/Component_Function_1/N5  ( .A1(
        \SB1_2_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][109] ) );
  NAND4_X1 \SB1_2_18/Component_Function_0/N5  ( .A1(
        \SB1_2_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_18/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][108] ) );
  NAND4_X1 \SB1_2_18/Component_Function_1/N5  ( .A1(
        \SB1_2_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_18/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][103] ) );
  NAND4_X1 \SB1_2_19/Component_Function_0/N5  ( .A1(
        \SB1_2_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][102] ) );
  NAND4_X1 \SB1_2_19/Component_Function_1/N5  ( .A1(
        \SB1_2_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_19/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][97] ) );
  NAND4_X1 \SB1_2_20/Component_Function_0/N5  ( .A1(
        \SB1_2_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][96] ) );
  NAND4_X1 \SB1_2_20/Component_Function_1/N5  ( .A1(
        \SB1_2_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][91] ) );
  NAND4_X1 \SB1_2_21/Component_Function_0/N5  ( .A1(
        \SB1_2_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_21/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][90] ) );
  NAND4_X1 \SB1_2_21/Component_Function_1/N5  ( .A1(
        \SB1_2_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_21/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][85] ) );
  NAND4_X1 \SB1_2_22/Component_Function_0/N5  ( .A1(
        \SB1_2_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][84] ) );
  NAND4_X1 \SB1_2_22/Component_Function_1/N5  ( .A1(
        \SB1_2_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][79] ) );
  NAND4_X1 \SB1_2_23/Component_Function_0/N5  ( .A1(
        \SB1_2_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_23/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][78] ) );
  NAND4_X1 \SB1_2_23/Component_Function_1/N5  ( .A1(
        \SB1_2_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][73] ) );
  NAND4_X1 \SB1_2_24/Component_Function_0/N5  ( .A1(
        \SB1_2_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_24/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][72] ) );
  NAND4_X1 \SB1_2_24/Component_Function_1/N5  ( .A1(
        \SB1_2_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][67] ) );
  NAND4_X1 \SB1_2_25/Component_Function_0/N5  ( .A1(
        \SB1_2_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_25/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][66] ) );
  NAND4_X1 \SB1_2_25/Component_Function_1/N5  ( .A1(
        \SB1_2_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][61] ) );
  NAND4_X1 \SB1_2_26/Component_Function_1/N5  ( .A1(
        \SB1_2_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][55] ) );
  NAND4_X1 \SB1_2_27/Component_Function_0/N5  ( .A1(
        \SB1_2_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_27/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][54] ) );
  NAND4_X1 \SB1_2_27/Component_Function_1/N5  ( .A1(
        \SB1_2_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][49] ) );
  NAND4_X1 \SB1_2_28/Component_Function_0/N5  ( .A1(
        \SB1_2_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][48] ) );
  NAND4_X1 \SB1_2_28/Component_Function_1/N5  ( .A1(
        \SB1_2_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][43] ) );
  NAND4_X1 \SB1_2_29/Component_Function_0/N5  ( .A1(
        \SB1_2_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][42] ) );
  NAND4_X1 \SB1_2_29/Component_Function_1/N5  ( .A1(
        \SB1_2_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][37] ) );
  NAND4_X1 \SB1_2_30/Component_Function_0/N5  ( .A1(
        \SB1_2_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][36] ) );
  NAND4_X1 \SB1_2_30/Component_Function_1/N5  ( .A1(
        \SB1_2_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_30/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[2][31] ) );
  NAND4_X1 \SB1_2_31/Component_Function_0/N5  ( .A1(
        \SB1_2_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[2][30] ) );
  NAND4_X1 \SB2_2_0/Component_Function_0/N5  ( .A1(
        \SB2_2_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][24] ) );
  NAND4_X1 \SB2_2_0/Component_Function_1/N5  ( .A1(
        \SB2_2_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][19] ) );
  NAND4_X1 \SB2_2_1/Component_Function_0/N5  ( .A1(
        \SB2_2_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_1/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][18] ) );
  NAND4_X1 \SB2_2_2/Component_Function_0/N5  ( .A1(
        \SB2_2_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_2/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][12] ) );
  NAND4_X1 \SB2_2_2/Component_Function_1/N5  ( .A1(
        \SB2_2_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_2/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][7] ) );
  NAND4_X1 \SB2_2_3/Component_Function_0/N5  ( .A1(
        \SB2_2_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_3/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][6] ) );
  NAND4_X1 \SB2_2_3/Component_Function_1/N5  ( .A1(
        \SB2_2_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][1] ) );
  NAND4_X1 \SB2_2_4/Component_Function_0/N5  ( .A1(
        \SB2_2_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][0] ) );
  NAND4_X1 \SB2_2_5/Component_Function_0/N5  ( .A1(
        \SB2_2_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_5/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][186] ) );
  NAND4_X1 \SB2_2_5/Component_Function_1/N5  ( .A1(
        \SB2_2_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][181] ) );
  NAND4_X1 \SB2_2_6/Component_Function_0/N5  ( .A1(
        \SB2_2_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_6/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][180] ) );
  NAND4_X1 \SB2_2_6/Component_Function_1/N5  ( .A1(
        \SB2_2_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][175] ) );
  NAND4_X1 \SB2_2_7/Component_Function_0/N5  ( .A1(
        \SB2_2_7/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_7/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][174] ) );
  NAND4_X1 \SB2_2_7/Component_Function_1/N5  ( .A1(
        \SB2_2_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][169] ) );
  NAND4_X1 \SB2_2_8/Component_Function_0/N5  ( .A1(
        \SB2_2_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_8/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][168] ) );
  NAND4_X1 \SB2_2_8/Component_Function_1/N5  ( .A1(
        \SB2_2_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][163] ) );
  NAND4_X1 \SB2_2_9/Component_Function_0/N5  ( .A1(
        \SB2_2_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][162] ) );
  NAND4_X1 \SB2_2_9/Component_Function_1/N5  ( .A1(
        \SB2_2_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][157] ) );
  NAND4_X1 \SB2_2_10/Component_Function_0/N5  ( .A1(
        \SB2_2_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_10/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][156] ) );
  NAND4_X1 \SB2_2_11/Component_Function_0/N5  ( .A1(
        \SB2_2_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][150] ) );
  NAND4_X1 \SB2_2_11/Component_Function_1/N5  ( .A1(
        \SB2_2_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][145] ) );
  NAND4_X1 \SB2_2_12/Component_Function_1/N5  ( .A1(
        \SB2_2_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_12/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][139] ) );
  NAND4_X1 \SB2_2_13/Component_Function_0/N5  ( .A1(
        \SB2_2_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][138] ) );
  NAND4_X1 \SB2_2_14/Component_Function_0/N5  ( .A1(
        \SB2_2_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_14/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][132] ) );
  NAND4_X1 \SB2_2_15/Component_Function_0/N5  ( .A1(
        \SB2_2_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_15/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][126] ) );
  NAND4_X1 \SB2_2_15/Component_Function_1/N5  ( .A1(
        \SB2_2_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][121] ) );
  NAND4_X1 \SB2_2_16/Component_Function_0/N5  ( .A1(
        \SB2_2_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_16/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][120] ) );
  NAND4_X1 \SB2_2_16/Component_Function_1/N5  ( .A1(
        \SB2_2_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_16/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][115] ) );
  NAND4_X1 \SB2_2_17/Component_Function_0/N5  ( .A1(
        \SB2_2_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][114] ) );
  NAND4_X1 \SB2_2_17/Component_Function_1/N5  ( .A1(
        \SB2_2_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][109] ) );
  NAND4_X1 \SB2_2_19/Component_Function_0/N5  ( .A1(
        \SB2_2_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][102] ) );
  NAND4_X1 \SB2_2_19/Component_Function_1/N5  ( .A1(
        \SB2_2_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_19/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][97] ) );
  NAND4_X1 \SB2_2_20/Component_Function_0/N5  ( .A1(
        \SB2_2_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_20/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][96] ) );
  NAND4_X1 \SB2_2_20/Component_Function_1/N5  ( .A1(
        \SB2_2_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_20/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][91] ) );
  NAND4_X1 \SB2_2_21/Component_Function_0/N5  ( .A1(
        \SB2_2_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_21/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][90] ) );
  NAND4_X1 \SB2_2_21/Component_Function_1/N5  ( .A1(
        \SB2_2_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_21/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][85] ) );
  NAND4_X1 \SB2_2_22/Component_Function_0/N5  ( .A1(
        \SB2_2_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][84] ) );
  NAND4_X1 \SB2_2_22/Component_Function_1/N5  ( .A1(
        \SB2_2_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][79] ) );
  NAND4_X1 \SB2_2_23/Component_Function_0/N5  ( .A1(
        \SB2_2_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_23/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][78] ) );
  NAND4_X1 \SB2_2_23/Component_Function_1/N5  ( .A1(
        \SB2_2_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][73] ) );
  NAND4_X1 \SB2_2_24/Component_Function_1/N5  ( .A1(
        \SB2_2_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][67] ) );
  NAND4_X1 \SB2_2_25/Component_Function_0/N5  ( .A1(
        \SB2_2_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_25/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][66] ) );
  NAND4_X1 \SB2_2_25/Component_Function_1/N5  ( .A1(
        \SB2_2_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][61] ) );
  NAND4_X1 \SB2_2_26/Component_Function_0/N5  ( .A1(
        \SB2_2_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_26/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][60] ) );
  NAND4_X1 \SB2_2_26/Component_Function_1/N5  ( .A1(
        \SB2_2_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][55] ) );
  NAND4_X1 \SB2_2_27/Component_Function_0/N5  ( .A1(
        \SB2_2_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_27/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][54] ) );
  NAND4_X1 \SB2_2_27/Component_Function_1/N5  ( .A1(
        \SB2_2_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][49] ) );
  NAND4_X1 \SB2_2_28/Component_Function_0/N5  ( .A1(
        \SB2_2_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][48] ) );
  NAND4_X1 \SB2_2_28/Component_Function_1/N5  ( .A1(
        \SB2_2_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][43] ) );
  NAND4_X1 \SB2_2_29/Component_Function_0/N5  ( .A1(
        \SB2_2_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][42] ) );
  NAND4_X1 \SB2_2_29/Component_Function_1/N5  ( .A1(
        \SB2_2_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][37] ) );
  NAND4_X1 \SB2_2_30/Component_Function_0/N5  ( .A1(
        \SB2_2_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][36] ) );
  NAND4_X1 \SB2_2_31/Component_Function_0/N5  ( .A1(
        \SB2_2_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][30] ) );
  NAND4_X1 \SB2_2_31/Component_Function_1/N5  ( .A1(
        \SB2_2_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_31/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][25] ) );
  NAND4_X1 \SB1_3_0/Component_Function_0/N5  ( .A1(
        \SB1_3_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][24] ) );
  NAND4_X1 \SB1_3_0/Component_Function_1/N5  ( .A1(
        \SB1_3_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][19] ) );
  NAND4_X1 \SB1_3_1/Component_Function_0/N5  ( .A1(
        \SB1_3_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_1/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][18] ) );
  NAND4_X1 \SB1_3_1/Component_Function_1/N5  ( .A1(
        \SB1_3_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_1/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][13] ) );
  NAND4_X1 \SB1_3_2/Component_Function_0/N5  ( .A1(
        \SB1_3_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_2/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][12] ) );
  NAND4_X1 \SB1_3_2/Component_Function_1/N5  ( .A1(
        \SB1_3_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_2/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][7] ) );
  NAND4_X1 \SB1_3_3/Component_Function_0/N5  ( .A1(
        \SB1_3_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_3/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][6] ) );
  NAND4_X1 \SB1_3_3/Component_Function_1/N5  ( .A1(
        \SB1_3_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][1] ) );
  NAND4_X1 \SB1_3_4/Component_Function_0/N5  ( .A1(
        \SB1_3_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_4/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][0] ) );
  NAND4_X1 \SB1_3_4/Component_Function_1/N5  ( .A1(
        \SB1_3_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][187] ) );
  NAND4_X1 \SB1_3_5/Component_Function_0/N5  ( .A1(
        \SB1_3_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][186] ) );
  NAND4_X1 \SB1_3_5/Component_Function_1/N5  ( .A1(
        \SB1_3_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][181] ) );
  NAND4_X1 \SB1_3_5/Component_Function_5/N5  ( .A1(
        \SB1_3_5/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[3][161] ) );
  NAND4_X1 \SB1_3_6/Component_Function_0/N5  ( .A1(
        \SB1_3_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_6/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][180] ) );
  NAND4_X1 \SB1_3_6/Component_Function_1/N5  ( .A1(
        \SB1_3_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][175] ) );
  NAND4_X1 \SB1_3_7/Component_Function_0/N5  ( .A1(
        \SB1_3_7/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_7/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][174] ) );
  NAND4_X1 \SB1_3_7/Component_Function_1/N5  ( .A1(
        \SB1_3_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][169] ) );
  NAND4_X1 \SB1_3_8/Component_Function_0/N5  ( .A1(
        \SB1_3_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_8/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][168] ) );
  NAND4_X1 \SB1_3_9/Component_Function_0/N5  ( .A1(
        \SB1_3_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][162] ) );
  NAND4_X1 \SB1_3_9/Component_Function_1/N5  ( .A1(
        \SB1_3_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][157] ) );
  NAND4_X1 \SB1_3_10/Component_Function_0/N5  ( .A1(
        \SB1_3_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][156] ) );
  NAND4_X1 \SB1_3_10/Component_Function_1/N5  ( .A1(
        \SB1_3_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][151] ) );
  NAND4_X1 \SB1_3_10/Component_Function_5/N5  ( .A1(
        \SB1_3_10/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[3][131] ) );
  NAND4_X1 \SB1_3_11/Component_Function_0/N5  ( .A1(
        \SB1_3_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][150] ) );
  NAND4_X1 \SB1_3_11/Component_Function_1/N5  ( .A1(
        \SB1_3_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][145] ) );
  NAND4_X1 \SB1_3_11/Component_Function_5/N5  ( .A1(
        \SB1_3_11/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_3_11/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_11/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[3][125] ) );
  NAND4_X1 \SB1_3_12/Component_Function_0/N5  ( .A1(
        \SB1_3_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_12/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][144] ) );
  NAND4_X1 \SB1_3_13/Component_Function_0/N5  ( .A1(
        \SB1_3_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][138] ) );
  NAND4_X1 \SB1_3_13/Component_Function_1/N5  ( .A1(
        \SB1_3_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][133] ) );
  NAND4_X1 \SB1_3_14/Component_Function_0/N5  ( .A1(
        \SB1_3_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_14/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][132] ) );
  NAND4_X1 \SB1_3_14/Component_Function_1/N5  ( .A1(
        \SB1_3_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_14/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][127] ) );
  NAND4_X1 \SB1_3_15/Component_Function_0/N5  ( .A1(
        \SB1_3_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][126] ) );
  NAND4_X1 \SB1_3_15/Component_Function_1/N5  ( .A1(
        \SB1_3_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][121] ) );
  NAND4_X1 \SB1_3_16/Component_Function_0/N5  ( .A1(
        \SB1_3_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_16/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][120] ) );
  NAND4_X1 \SB1_3_16/Component_Function_1/N5  ( .A1(
        \SB1_3_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_16/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][115] ) );
  NAND4_X1 \SB1_3_16/Component_Function_5/N5  ( .A1(
        \SB1_3_16/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_3_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_16/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[3][95] ) );
  NAND4_X1 \SB1_3_17/Component_Function_0/N5  ( .A1(
        \SB1_3_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][114] ) );
  NAND4_X1 \SB1_3_17/Component_Function_1/N5  ( .A1(
        \SB1_3_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][109] ) );
  NAND4_X1 \SB1_3_18/Component_Function_0/N5  ( .A1(
        \SB1_3_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][108] ) );
  NAND4_X1 \SB1_3_18/Component_Function_1/N5  ( .A1(
        \SB1_3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][103] ) );
  NAND4_X1 \SB1_3_18/Component_Function_5/N5  ( .A1(
        \SB1_3_18/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[3][83] ) );
  NAND4_X1 \SB1_3_19/Component_Function_0/N5  ( .A1(
        \SB1_3_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][102] ) );
  NAND4_X1 \SB1_3_20/Component_Function_0/N5  ( .A1(
        \SB1_3_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_20/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][96] ) );
  NAND4_X1 \SB1_3_21/Component_Function_1/N5  ( .A1(
        \SB1_3_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_21/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][85] ) );
  NAND4_X1 \SB1_3_21/Component_Function_5/N5  ( .A1(
        \SB1_3_21/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_3_21/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_21/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_21/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[3][65] ) );
  NAND4_X1 \SB1_3_22/Component_Function_0/N5  ( .A1(
        \SB1_3_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][84] ) );
  NAND4_X1 \SB1_3_22/Component_Function_1/N5  ( .A1(
        \SB1_3_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][79] ) );
  NAND4_X1 \SB1_3_23/Component_Function_0/N5  ( .A1(
        \SB1_3_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_23/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][78] ) );
  NAND4_X1 \SB1_3_24/Component_Function_0/N5  ( .A1(
        \SB1_3_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][72] ) );
  NAND4_X1 \SB1_3_24/Component_Function_1/N5  ( .A1(
        \SB1_3_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][67] ) );
  NAND4_X1 \SB1_3_25/Component_Function_0/N5  ( .A1(
        \SB1_3_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_25/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][66] ) );
  NAND4_X1 \SB1_3_26/Component_Function_0/N5  ( .A1(
        \SB1_3_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_26/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][60] ) );
  NAND4_X1 \SB1_3_26/Component_Function_1/N5  ( .A1(
        \SB1_3_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][55] ) );
  NAND4_X1 \SB1_3_27/Component_Function_1/N5  ( .A1(
        \SB1_3_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][49] ) );
  NAND4_X1 \SB1_3_28/Component_Function_0/N5  ( .A1(
        \SB1_3_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][48] ) );
  NAND4_X1 \SB1_3_28/Component_Function_1/N5  ( .A1(
        \SB1_3_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][43] ) );
  NAND4_X1 \SB1_3_29/Component_Function_0/N5  ( .A1(
        \SB1_3_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][42] ) );
  NAND4_X1 \SB1_3_29/Component_Function_1/N5  ( .A1(
        \SB1_3_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][37] ) );
  NAND4_X1 \SB1_3_30/Component_Function_0/N5  ( .A1(
        \SB1_3_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][36] ) );
  NAND4_X1 \SB1_3_30/Component_Function_1/N5  ( .A1(
        \SB1_3_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_30/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][31] ) );
  NAND4_X1 \SB1_3_31/Component_Function_0/N5  ( .A1(
        \SB1_3_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[3][30] ) );
  NAND4_X1 \SB1_3_31/Component_Function_1/N5  ( .A1(
        \SB1_3_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_31/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[3][25] ) );
  NAND4_X1 \SB2_3_2/Component_Function_0/N5  ( .A1(
        \SB2_3_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_2/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][12] ) );
  NAND4_X1 \SB2_3_7/Component_Function_0/N5  ( .A1(
        \SB2_3_7/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_7/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][174] ) );
  NAND4_X1 \SB2_3_12/Component_Function_0/N5  ( .A1(
        \SB2_3_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_12/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][144] ) );
  NAND4_X1 \SB2_3_14/Component_Function_0/N5  ( .A1(
        \SB2_3_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_14/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][132] ) );
  NAND4_X1 \SB2_3_17/Component_Function_0/N5  ( .A1(
        \SB2_3_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_17/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][114] ) );
  NAND4_X1 \SB2_3_19/Component_Function_0/N5  ( .A1(
        \SB2_3_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][102] ) );
  NAND4_X1 \SB2_3_25/Component_Function_5/N5  ( .A1(
        \SB2_3_25/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_3_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_25/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_3_25/Component_Function_5/NAND4_in[3] ), .ZN(\RI5[3][41] ) );
  NAND4_X1 \SB2_3_29/Component_Function_0/N5  ( .A1(
        \SB2_3_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_29/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][42] ) );
  NAND4_X1 \SB3_0/Component_Function_0/N5  ( .A1(
        \SB3_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][24] ) );
  NAND4_X1 \SB3_0/Component_Function_1/N5  ( .A1(
        \SB3_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_0/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][19] ) );
  NAND4_X1 \SB3_0/Component_Function_5/N5  ( .A1(
        \SB3_0/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_0/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_0/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_0/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[4][191] ) );
  NAND4_X1 \SB3_2/Component_Function_1/N5  ( .A1(
        \SB3_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_2/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][7] ) );
  NAND4_X1 \SB3_3/Component_Function_1/N5  ( .A1(
        \SB3_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][1] ) );
  NAND4_X1 \SB3_4/Component_Function_0/N5  ( .A1(
        \SB3_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_4/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][0] ) );
  NAND4_X1 \SB3_4/Component_Function_1/N5  ( .A1(
        \SB3_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][187] ) );
  NAND4_X1 \SB3_4/Component_Function_5/N5  ( .A1(
        \SB3_4/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_4/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[4][167] ) );
  NAND4_X1 \SB3_5/Component_Function_1/N5  ( .A1(
        \SB3_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][181] ) );
  NAND4_X1 \SB3_5/Component_Function_5/N5  ( .A1(
        \SB3_5/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_5/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[4][161] ) );
  NAND4_X1 \SB3_6/Component_Function_1/N5  ( .A1(
        \SB3_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][175] ) );
  NAND4_X1 \SB3_6/Component_Function_5/N5  ( .A1(
        \SB3_6/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[4][155] ) );
  NAND4_X1 \SB3_7/Component_Function_1/N5  ( .A1(
        \SB3_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][169] ) );
  NAND4_X1 \SB3_8/Component_Function_0/N5  ( .A1(
        \SB3_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][168] ) );
  NAND4_X1 \SB3_8/Component_Function_1/N5  ( .A1(
        \SB3_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][163] ) );
  NAND4_X1 \SB3_9/Component_Function_0/N5  ( .A1(
        \SB3_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][162] ) );
  NAND4_X1 \SB3_9/Component_Function_1/N5  ( .A1(
        \SB3_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][157] ) );
  NAND4_X1 \SB3_10/Component_Function_1/N5  ( .A1(
        \SB3_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][151] ) );
  NAND4_X1 \SB3_11/Component_Function_0/N5  ( .A1(
        \SB3_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][150] ) );
  NAND4_X1 \SB3_11/Component_Function_1/N5  ( .A1(
        \SB3_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][145] ) );
  NAND4_X1 \SB3_12/Component_Function_0/N5  ( .A1(
        \SB3_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_12/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][144] ) );
  NAND4_X1 \SB3_12/Component_Function_1/N5  ( .A1(
        \SB3_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_12/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][139] ) );
  NAND4_X1 \SB3_13/Component_Function_0/N5  ( .A1(
        \SB3_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][138] ) );
  NAND4_X1 \SB3_13/Component_Function_1/N5  ( .A1(
        \SB3_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][133] ) );
  NAND4_X1 \SB3_13/Component_Function_5/N5  ( .A1(
        \SB3_13/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_13/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[4][113] ) );
  NAND4_X1 \SB3_14/Component_Function_1/N5  ( .A1(
        \SB3_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_14/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][127] ) );
  NAND4_X1 \SB3_15/Component_Function_1/N5  ( .A1(
        \SB3_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][121] ) );
  NAND4_X1 \SB3_16/Component_Function_0/N5  ( .A1(
        \SB3_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_16/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][120] ) );
  NAND4_X1 \SB3_16/Component_Function_1/N5  ( .A1(
        \SB3_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_16/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][115] ) );
  NAND4_X1 \SB3_17/Component_Function_1/N5  ( .A1(
        \SB3_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][109] ) );
  NAND4_X1 \SB3_18/Component_Function_1/N5  ( .A1(
        \SB3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][103] ) );
  NAND4_X1 \SB3_19/Component_Function_0/N5  ( .A1(
        \SB3_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][102] ) );
  NAND4_X1 \SB3_19/Component_Function_1/N5  ( .A1(
        \SB3_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][97] ) );
  NAND4_X1 \SB3_20/Component_Function_0/N5  ( .A1(
        \SB3_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_20/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][96] ) );
  NAND4_X1 \SB3_20/Component_Function_1/N5  ( .A1(
        \SB3_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_20/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][91] ) );
  NAND4_X1 \SB3_21/Component_Function_0/N5  ( .A1(
        \SB3_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][90] ) );
  NAND4_X1 \SB3_22/Component_Function_1/N5  ( .A1(
        \SB3_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][79] ) );
  NAND4_X1 \SB3_22/Component_Function_5/N5  ( .A1(
        \SB3_22/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[4][59] ) );
  NAND4_X1 \SB3_23/Component_Function_0/N5  ( .A1(
        \SB3_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_23/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][78] ) );
  NAND4_X1 \SB3_23/Component_Function_1/N5  ( .A1(
        \SB3_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][73] ) );
  NAND4_X1 \SB3_24/Component_Function_1/N5  ( .A1(
        \SB3_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][67] ) );
  NAND4_X1 \SB3_25/Component_Function_0/N5  ( .A1(
        \SB3_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_25/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][66] ) );
  NAND4_X1 \SB3_25/Component_Function_1/N5  ( .A1(
        \SB3_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][61] ) );
  NAND4_X1 \SB3_26/Component_Function_1/N5  ( .A1(
        \SB3_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][55] ) );
  NAND4_X1 \SB3_27/Component_Function_1/N5  ( .A1(
        \SB3_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][49] ) );
  NAND4_X1 \SB3_28/Component_Function_0/N5  ( .A1(
        \SB3_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_28/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][48] ) );
  NAND4_X1 \SB3_28/Component_Function_1/N5  ( .A1(
        \SB3_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][43] ) );
  NAND4_X1 \SB3_29/Component_Function_1/N5  ( .A1(
        \SB3_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][37] ) );
  NAND4_X1 \SB3_30/Component_Function_0/N5  ( .A1(
        \SB3_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_30/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][36] ) );
  NAND4_X1 \SB3_30/Component_Function_1/N5  ( .A1(
        \SB3_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_30/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][31] ) );
  NAND4_X1 \SB3_31/Component_Function_0/N5  ( .A1(
        \SB3_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_0/NAND4_in[3] ), .ZN(\RI3[4][30] ) );
  NAND4_X1 \SB3_31/Component_Function_1/N5  ( .A1(
        \SB3_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[4][25] ) );
  INV_X1 \SB3_1/INV_5  ( .A(\RI1[4][185] ), .ZN(\SB3_1/i0_3 ) );
  INV_X1 \SB3_11/INV_5  ( .A(\RI1[4][125] ), .ZN(\SB3_11/i0_3 ) );
  INV_X1 \SB3_14/INV_5  ( .A(\RI1[4][107] ), .ZN(\SB3_14/i0_3 ) );
  INV_X1 \SB3_18/INV_5  ( .A(\RI1[4][83] ), .ZN(\SB3_18/i0_3 ) );
  INV_X1 \SB3_23/INV_5  ( .A(\RI1[4][53] ), .ZN(\SB3_23/i0_3 ) );
  INV_X1 \SB3_28/INV_5  ( .A(\RI1[4][23] ), .ZN(\SB3_28/i0_3 ) );
  INV_X1 \SB3_29/INV_5  ( .A(\RI1[4][17] ), .ZN(\SB3_29/i0_3 ) );
  INV_X1 \SB3_30/INV_5  ( .A(\RI1[4][11] ), .ZN(\SB3_30/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_71  ( .A(\RI5[3][71] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[71] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_5  ( .A(\RI5[3][5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[5] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_11  ( .A(\RI5[3][11] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[11] ) );
  BUF_X1 \SB3_5/BUF_3  ( .A(\RI1[4][159] ), .Z(\SB3_5/i0[8] ) );
  BUF_X1 \SB3_29/BUF_3  ( .A(\RI1[4][15] ), .Z(\SB3_29/i0[8] ) );
  BUF_X1 \SB3_8/BUF_2  ( .A(\RI1[4][140] ), .Z(\SB3_8/i1[9] ) );
  BUF_X1 \SB1_1_2/BUF_5  ( .A(\RI1[1][179] ), .Z(\SB1_1_2/i1_5 ) );
  BUF_X1 \SB3_6/BUF_2  ( .A(\RI1[4][152] ), .Z(\SB3_6/i1[9] ) );
  BUF_X1 \SB1_1_13/BUF_5  ( .A(\RI1[1][113] ), .Z(\SB1_1_13/i1_5 ) );
  BUF_X1 \SB3_21/BUF_2  ( .A(\RI1[4][62] ), .Z(\SB3_21/i1[9] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_76  ( .A(\RI5[1][76] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[76] ) );
  INV_X1 \SB3_21/INV_5  ( .A(\RI1[4][65] ), .ZN(\SB3_21/i0_3 ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X4_21_1  ( .A(\MC_ARK_ARC_1_3/buf_datainput[100] ), 
        .B(n239), .ZN(\MC_ARK_ARC_1_3/temp4[64] ) );
  INV_X1 \SB3_20/INV_4  ( .A(\RI1[4][70] ), .ZN(\SB3_20/i0_4 ) );
  XNOR2_X1 \MC_ARK_ARC_1_3/X7_20_1  ( .A(\MC_ARK_ARC_1_3/temp6[70] ), .B(
        \MC_ARK_ARC_1_3/temp5[70] ), .ZN(\RI1[4][70] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_4  ( .A(\RI5[1][4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[4] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_106  ( .A(\RI5[1][106] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[106] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_10  ( .A(\RI5[2][10] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_130  ( .A(\RI5[2][130] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[130] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_40  ( .A(\RI5[2][40] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[40] ) );
  BUF_X2 \SB2_2_9/BUF_3  ( .A(\RI3[2][135] ), .Z(\SB2_2_9/i0[10] ) );
  BUF_X2 \SB4_25/BUF_5  ( .A(\RI3[4][41] ), .Z(\SB4_25/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_116  ( .A(\RI5[3][116] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[116] ) );
  BUF_X2 \SB2_0_11/BUF_5  ( .A(\RI3[0][125] ), .Z(\SB2_0_11/i0_3 ) );
  BUF_X2 \SB2_1_12/BUF_2  ( .A(\RI3[1][116] ), .Z(\SB2_1_12/i0_0 ) );
  BUF_X2 \SB2_2_19/BUF_3  ( .A(\RI3[2][75] ), .Z(\SB2_2_19/i0[10] ) );
  BUF_X2 \SB2_1_30/BUF_3  ( .A(\RI3[1][9] ), .Z(\SB2_1_30/i0[10] ) );
  BUF_X2 \SB2_0_17/BUF_4  ( .A(\RI3[0][88] ), .Z(\SB2_0_17/i0_4 ) );
  BUF_X2 \SB4_5/BUF_5  ( .A(\RI3[4][161] ), .Z(\SB4_5/i0_3 ) );
  BUF_X2 \SB2_1_3/BUF_3  ( .A(\RI3[1][171] ), .Z(\SB2_1_3/i0[10] ) );
  BUF_X2 \SB2_1_23/BUF_3  ( .A(\RI3[1][51] ), .Z(\SB2_1_23/i0[10] ) );
  BUF_X2 \SB4_10/BUF_5  ( .A(\RI3[4][131] ), .Z(\SB4_10/i0_3 ) );
  BUF_X2 \SB2_2_9/BUF_2  ( .A(\RI3[2][134] ), .Z(\SB2_2_9/i0_0 ) );
  BUF_X2 \SB2_1_1/BUF_3  ( .A(\RI3[1][183] ), .Z(\SB2_1_1/i0[10] ) );
  BUF_X2 \SB2_2_7/BUF_3  ( .A(\RI3[2][147] ), .Z(\SB2_2_7/i0[10] ) );
  BUF_X2 \SB2_2_29/BUF_3  ( .A(\RI3[2][15] ), .Z(\SB2_2_29/i0[10] ) );
  BUF_X2 \SB2_1_9/BUF_3  ( .A(\RI3[1][135] ), .Z(\SB2_1_9/i0[10] ) );
  BUF_X2 \SB2_1_26/BUF_3  ( .A(\RI3[1][33] ), .Z(\SB2_1_26/i0[10] ) );
  BUF_X2 \SB1_1_30/BUF_3  ( .A(\RI1[1][9] ), .Z(\SB1_1_30/i0[8] ) );
  BUF_X2 \SB2_1_8/BUF_2  ( .A(\RI3[1][140] ), .Z(\SB2_1_8/i0_0 ) );
  BUF_X2 \SB2_1_13/BUF_3  ( .A(\RI3[1][111] ), .Z(\SB2_1_13/i0[10] ) );
  BUF_X2 \SB2_1_24/BUF_3  ( .A(\RI3[1][45] ), .Z(\SB2_1_24/i0[10] ) );
  BUF_X2 \SB2_1_28/BUF_3  ( .A(\RI3[1][21] ), .Z(\SB2_1_28/i0[10] ) );
  BUF_X2 \SB2_1_31/BUF_3  ( .A(\RI3[1][3] ), .Z(\SB2_1_31/i0[10] ) );
  BUF_X2 \SB2_0_19/BUF_3  ( .A(\RI3[0][75] ), .Z(\SB2_0_19/i0[10] ) );
  BUF_X2 \SB2_2_30/BUF_2  ( .A(\RI3[2][8] ), .Z(\SB2_2_30/i0_0 ) );
  BUF_X2 \SB4_20/BUF_5  ( .A(\RI3[4][71] ), .Z(\SB4_20/i0_3 ) );
  BUF_X2 \SB2_1_21/BUF_3  ( .A(\RI3[1][63] ), .Z(\SB2_1_21/i0[10] ) );
  BUF_X2 \SB2_2_1/BUF_3  ( .A(\RI3[2][183] ), .Z(\SB2_2_1/i0[10] ) );
  BUF_X2 \SB2_1_25/BUF_4  ( .A(\RI3[1][40] ), .Z(\SB2_1_25/i0_4 ) );
  BUF_X2 \SB2_2_14/BUF_2  ( .A(\RI3[2][104] ), .Z(\SB2_2_14/i0_0 ) );
  BUF_X2 \SB2_1_29/BUF_4  ( .A(\RI3[1][16] ), .Z(\SB2_1_29/i0_4 ) );
  BUF_X2 \SB4_16/BUF_5  ( .A(\RI3[4][95] ), .Z(\SB4_16/i0_3 ) );
  BUF_X2 \SB2_2_24/BUF_3  ( .A(\RI3[2][45] ), .Z(\SB2_2_24/i0[10] ) );
  BUF_X2 \SB2_2_24/BUF_4  ( .A(\RI3[2][46] ), .Z(\SB2_2_24/i0_4 ) );
  BUF_X2 \SB2_0_25/BUF_4  ( .A(\RI3[0][40] ), .Z(\SB2_0_25/i0_4 ) );
  BUF_X2 \SB2_2_2/BUF_4  ( .A(\RI3[2][178] ), .Z(\SB2_2_2/i0_4 ) );
  BUF_X2 \SB2_1_26/BUF_2  ( .A(\RI3[1][32] ), .Z(\SB2_1_26/i0_0 ) );
  BUF_X2 \SB4_29/BUF_5  ( .A(\RI3[4][17] ), .Z(\SB4_29/i0_3 ) );
  BUF_X2 \SB2_2_15/BUF_4  ( .A(\RI3[2][100] ), .Z(\SB2_2_15/i0_4 ) );
  BUF_X2 \SB4_19/BUF_5  ( .A(\RI3[4][77] ), .Z(\SB4_19/i0_3 ) );
  BUF_X2 \SB2_1_13/BUF_2  ( .A(\RI3[1][110] ), .Z(\SB2_1_13/i0_0 ) );
  BUF_X2 \SB2_3_4/BUF_2  ( .A(\RI3[3][164] ), .Z(\SB2_3_4/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_9  ( .A(\RI5[0][9] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[9] ) );
  BUF_X2 \SB4_2/BUF_5  ( .A(\RI3[4][179] ), .Z(\SB4_2/i0_3 ) );
  BUF_X2 \SB2_1_16/BUF_3  ( .A(\RI3[1][93] ), .Z(\SB2_1_16/i0[10] ) );
  BUF_X2 \SB2_3_24/BUF_4  ( .A(\RI3[3][46] ), .Z(\SB2_3_24/i0_4 ) );
  BUF_X2 \SB2_2_3/BUF_4  ( .A(\RI3[2][172] ), .Z(\SB2_2_3/i0_4 ) );
  BUF_X2 \SB2_2_13/BUF_2  ( .A(\RI3[2][110] ), .Z(\SB2_2_13/i0_0 ) );
  BUF_X2 \SB2_2_11/BUF_4  ( .A(\RI3[2][124] ), .Z(\SB2_2_11/i0_4 ) );
  BUF_X2 \SB4_19/BUF_2  ( .A(\RI3[4][74] ), .Z(\SB4_19/i0_0 ) );
  BUF_X2 \SB2_2_26/BUF_4  ( .A(\RI3[2][34] ), .Z(\SB2_2_26/i0_4 ) );
  BUF_X2 \SB4_14/BUF_5  ( .A(\RI3[4][107] ), .Z(\SB4_14/i0_3 ) );
  BUF_X2 \SB2_3_18/BUF_2  ( .A(\RI3[3][80] ), .Z(\SB2_3_18/i0_0 ) );
  BUF_X2 \SB2_0_18/BUF_4  ( .A(\RI3[0][82] ), .Z(\SB2_0_18/i0_4 ) );
  BUF_X2 \SB2_1_4/BUF_2  ( .A(\RI3[1][164] ), .Z(\SB2_1_4/i0_0 ) );
  BUF_X2 \SB2_1_1/BUF_4  ( .A(\RI3[1][184] ), .Z(\SB2_1_1/i0_4 ) );
  BUF_X2 \SB2_2_0/BUF_4  ( .A(\RI3[2][190] ), .Z(\SB2_2_0/i0_4 ) );
  BUF_X2 \SB2_0_20/BUF_2  ( .A(\RI3[0][68] ), .Z(\SB2_0_20/i0_0 ) );
  BUF_X2 \SB2_1_11/BUF_4  ( .A(\RI3[1][124] ), .Z(\SB2_1_11/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_132  ( .A(\RI5[3][132] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[132] ) );
  BUF_X2 \SB2_3_24/BUF_3  ( .A(\RI3[3][45] ), .Z(\SB2_3_24/i0[10] ) );
  BUF_X2 \SB3_28/BUF_3  ( .A(\RI1[4][21] ), .Z(\SB3_28/i0[8] ) );
  BUF_X2 \SB4_25/BUF_2  ( .A(\RI3[4][38] ), .Z(\SB4_25/i0_0 ) );
  BUF_X2 \SB2_3_17/BUF_3  ( .A(\RI3[3][87] ), .Z(\SB2_3_17/i0[10] ) );
  BUF_X2 \SB2_2_15/BUF_3  ( .A(\RI3[2][99] ), .Z(\SB2_2_15/i0[10] ) );
  BUF_X2 \SB2_1_26/BUF_4  ( .A(\RI3[1][34] ), .Z(\SB2_1_26/i0_4 ) );
  BUF_X2 \SB2_3_18/BUF_3  ( .A(\RI3[3][81] ), .Z(\SB2_3_18/i0[10] ) );
  BUF_X2 \SB2_3_12/BUF_4  ( .A(\RI3[3][118] ), .Z(\SB2_3_12/i0_4 ) );
  BUF_X2 \SB2_2_31/BUF_4  ( .A(\RI3[2][4] ), .Z(\SB2_2_31/i0_4 ) );
  BUF_X2 \SB4_8/BUF_2  ( .A(\RI3[4][140] ), .Z(\SB4_8/i0_0 ) );
  BUF_X2 \SB4_4/BUF_2  ( .A(\RI3[4][164] ), .Z(\SB4_4/i0_0 ) );
  BUF_X2 \SB2_1_3/BUF_4  ( .A(\RI3[1][172] ), .Z(\SB2_1_3/i0_4 ) );
  BUF_X2 \SB2_2_17/BUF_4  ( .A(\RI3[2][88] ), .Z(\SB2_2_17/i0_4 ) );
  BUF_X2 \SB2_1_30/BUF_4  ( .A(\RI3[1][10] ), .Z(\SB2_1_30/i0_4 ) );
  BUF_X2 \SB4_30/BUF_2  ( .A(\RI3[4][8] ), .Z(\SB4_30/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_144  ( .A(\RI5[3][144] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[144] ) );
  BUF_X2 \SB4_25/BUF_4  ( .A(\RI3[4][40] ), .Z(\SB4_25/i0_4 ) );
  BUF_X2 \SB2_3_23/BUF_2  ( .A(\RI3[3][50] ), .Z(\SB2_3_23/i0_0 ) );
  BUF_X2 \SB2_2_29/BUF_5  ( .A(\RI3[2][17] ), .Z(\SB2_2_29/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_26  ( .A(\RI5[3][26] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[26] ) );
  BUF_X2 \SB2_2_7/BUF_4  ( .A(\RI3[2][148] ), .Z(\SB2_2_7/i0_4 ) );
  BUF_X2 \SB2_3_30/BUF_4  ( .A(\RI3[3][10] ), .Z(\SB2_3_30/i0_4 ) );
  BUF_X2 \SB2_0_7/BUF_5  ( .A(\RI3[0][149] ), .Z(\SB2_0_7/i0_3 ) );
  BUF_X2 \SB2_3_20/BUF_3  ( .A(\RI3[3][69] ), .Z(\SB2_3_20/i0[10] ) );
  BUF_X2 \SB2_2_18/BUF_4  ( .A(\RI3[2][82] ), .Z(\SB2_2_18/i0_4 ) );
  BUF_X2 \SB4_1/BUF_4  ( .A(\RI3[4][184] ), .Z(\SB4_1/i0_4 ) );
  BUF_X2 \SB2_0_17/BUF_5  ( .A(\RI3[0][89] ), .Z(\SB2_0_17/i0_3 ) );
  BUF_X2 \SB2_3_22/BUF_3  ( .A(\RI3[3][57] ), .Z(\SB2_3_22/i0[10] ) );
  BUF_X2 \SB2_2_20/BUF_3  ( .A(\RI3[2][69] ), .Z(\SB2_2_20/i0[10] ) );
  BUF_X2 \SB2_2_3/BUF_2  ( .A(\RI3[2][170] ), .Z(\SB2_2_3/i0_0 ) );
  BUF_X2 \SB2_1_18/BUF_3  ( .A(\RI3[1][81] ), .Z(\SB2_1_18/i0[10] ) );
  BUF_X2 \SB2_1_28/BUF_4  ( .A(\RI3[1][22] ), .Z(\SB2_1_28/i0_4 ) );
  BUF_X2 \SB1_2_20/BUF_2  ( .A(\RI1[2][68] ), .Z(\SB1_2_20/i1[9] ) );
  BUF_X2 \SB2_2_19/BUF_4  ( .A(\RI3[2][76] ), .Z(\SB2_2_19/i0_4 ) );
  BUF_X2 \SB4_6/BUF_4  ( .A(\RI3[4][154] ), .Z(\SB4_6/i0_4 ) );
  BUF_X2 \SB4_16/BUF_4  ( .A(\RI3[4][94] ), .Z(\SB4_16/i0_4 ) );
  BUF_X2 \SB2_0_15/BUF_2  ( .A(\RI3[0][98] ), .Z(\SB2_0_15/i0_0 ) );
  BUF_X2 \SB2_1_21/BUF_4  ( .A(\RI3[1][64] ), .Z(\SB2_1_21/i0_4 ) );
  BUF_X2 \SB2_2_27/BUF_2  ( .A(\RI3[2][26] ), .Z(\SB2_2_27/i0_0 ) );
  BUF_X2 \SB4_9/BUF_3  ( .A(\RI3[4][135] ), .Z(\SB4_9/i0[10] ) );
  BUF_X2 \SB2_0_14/BUF_5  ( .A(\RI3[0][107] ), .Z(\SB2_0_14/i0_3 ) );
  BUF_X2 \SB2_1_4/BUF_4  ( .A(\RI3[1][166] ), .Z(\SB2_1_4/i0_4 ) );
  BUF_X2 \SB2_3_3/BUF_4  ( .A(\RI3[3][172] ), .Z(\SB2_3_3/i0_4 ) );
  INV_X2 \SB1_1_5/INV_5  ( .A(\RI1[1][161] ), .ZN(\SB1_1_5/i0_3 ) );
  BUF_X2 \SB4_9/BUF_2  ( .A(\RI3[4][134] ), .Z(\SB4_9/i0_0 ) );
  BUF_X2 \SB4_15/BUF_2  ( .A(\RI3[4][98] ), .Z(\SB4_15/i0_0 ) );
  BUF_X2 \SB2_2_7/BUF_5  ( .A(\RI3[2][149] ), .Z(\SB2_2_7/i0_3 ) );
  BUF_X2 \SB2_2_2/BUF_5  ( .A(\RI3[2][179] ), .Z(\SB2_2_2/i0_3 ) );
  BUF_X2 \SB2_1_19/BUF_4  ( .A(\RI3[1][76] ), .Z(\SB2_1_19/i0_4 ) );
  BUF_X2 \SB4_3/BUF_2  ( .A(\RI3[4][170] ), .Z(\SB4_3/i0_0 ) );
  BUF_X2 \SB4_13/BUF_2  ( .A(\RI3[4][110] ), .Z(\SB4_13/i0_0 ) );
  BUF_X2 \SB2_3_23/BUF_3  ( .A(\RI3[3][51] ), .Z(\SB2_3_23/i0[10] ) );
  BUF_X2 \SB2_0_6/BUF_5  ( .A(\RI3[0][155] ), .Z(\SB2_0_6/i0_3 ) );
  BUF_X2 \SB2_2_16/BUF_5  ( .A(\RI3[2][95] ), .Z(\SB2_2_16/i0_3 ) );
  BUF_X2 \SB2_1_27/BUF_3  ( .A(\RI3[1][27] ), .Z(\SB2_1_27/i0[10] ) );
  INV_X2 \SB1_1_29/INV_5  ( .A(\RI1[1][17] ), .ZN(\SB1_1_29/i0_3 ) );
  BUF_X2 \SB4_0/BUF_4  ( .A(\RI3[4][190] ), .Z(\SB4_0/i0_4 ) );
  BUF_X2 \SB2_2_4/BUF_5  ( .A(\RI3[2][167] ), .Z(\SB2_2_4/i0_3 ) );
  BUF_X2 \SB2_0_18/BUF_5  ( .A(\RI3[0][83] ), .Z(\SB2_0_18/i0_3 ) );
  INV_X2 \SB1_1_27/INV_5  ( .A(\RI1[1][29] ), .ZN(\SB1_1_27/i0_3 ) );
  BUF_X2 \SB2_2_26/BUF_2  ( .A(\RI3[2][32] ), .Z(\SB2_2_26/i0_0 ) );
  BUF_X2 \SB2_1_25/BUF_3  ( .A(\RI3[1][39] ), .Z(\SB2_1_25/i0[10] ) );
  BUF_X2 \SB4_7/BUF_4  ( .A(\RI3[4][148] ), .Z(\SB4_7/i0_4 ) );
  BUF_X2 \SB2_3_7/BUF_4  ( .A(\RI3[3][148] ), .Z(\SB2_3_7/i0_4 ) );
  BUF_X2 \SB4_24/BUF_4  ( .A(\RI3[4][46] ), .Z(\SB4_24/i0_4 ) );
  BUF_X2 \SB2_0_18/BUF_2  ( .A(\RI3[0][80] ), .Z(\SB2_0_18/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_42  ( .A(\RI5[3][42] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[42] ) );
  BUF_X2 \SB2_2_10/BUF_2  ( .A(\RI3[2][128] ), .Z(\SB2_2_10/i0_0 ) );
  BUF_X2 \SB2_3_29/BUF_4  ( .A(\RI3[3][16] ), .Z(\SB2_3_29/i0_4 ) );
  BUF_X2 \SB2_1_9/BUF_2  ( .A(\RI3[1][134] ), .Z(\SB2_1_9/i0_0 ) );
  BUF_X2 \SB2_1_9/BUF_4  ( .A(\RI3[1][136] ), .Z(\SB2_1_9/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_98  ( .A(\RI5[0][98] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[98] ) );
  BUF_X2 \SB4_15/BUF_4  ( .A(\RI3[4][100] ), .Z(\SB4_15/i0_4 ) );
  BUF_X2 \SB1_2_24/BUF_2  ( .A(\RI1[2][44] ), .Z(\SB1_2_24/i1[9] ) );
  BUF_X2 \SB2_3_15/BUF_3  ( .A(\RI3[3][99] ), .Z(\SB2_3_15/i0[10] ) );
  BUF_X2 \SB2_1_14/BUF_3  ( .A(\RI3[1][105] ), .Z(\SB2_1_14/i0[10] ) );
  BUF_X2 \SB4_31/BUF_4  ( .A(\RI3[4][4] ), .Z(\SB4_31/i0_4 ) );
  BUF_X2 \SB2_2_8/BUF_2  ( .A(\RI3[2][140] ), .Z(\SB2_2_8/i0_0 ) );
  BUF_X2 \SB2_1_10/BUF_4  ( .A(\RI3[1][130] ), .Z(\SB2_1_10/i0_4 ) );
  BUF_X2 \SB2_0_5/BUF_5  ( .A(\RI3[0][161] ), .Z(\SB2_0_5/i0_3 ) );
  BUF_X2 \SB2_2_24/BUF_5  ( .A(\RI3[2][47] ), .Z(\SB2_2_24/i0_3 ) );
  BUF_X2 \SB2_1_31/BUF_2  ( .A(\RI3[1][2] ), .Z(\SB2_1_31/i0_0 ) );
  BUF_X2 \SB4_25/BUF_3  ( .A(\RI3[4][39] ), .Z(\SB4_25/i0[10] ) );
  BUF_X2 \SB4_30/BUF_4  ( .A(\RI3[4][10] ), .Z(\SB4_30/i0_4 ) );
  BUF_X2 \SB2_2_22/BUF_4  ( .A(\RI3[2][58] ), .Z(\SB2_2_22/i0_4 ) );
  BUF_X2 \SB2_1_3/BUF_2  ( .A(\RI3[1][170] ), .Z(\SB2_1_3/i0_0 ) );
  BUF_X2 \SB2_0_2/BUF_5  ( .A(\RI3[0][179] ), .Z(\SB2_0_2/i0_3 ) );
  BUF_X2 \SB2_2_24/BUF_2  ( .A(\RI3[2][44] ), .Z(\SB2_2_24/i0_0 ) );
  BUF_X2 \SB2_1_6/BUF_4  ( .A(\RI3[1][154] ), .Z(\SB2_1_6/i0_4 ) );
  BUF_X2 \SB2_1_23/BUF_4  ( .A(\RI3[1][52] ), .Z(\SB2_1_23/i0_4 ) );
  BUF_X2 \SB2_1_30/BUF_2  ( .A(\RI3[1][8] ), .Z(\SB2_1_30/i0_0 ) );
  BUF_X2 \SB4_10/BUF_4  ( .A(\RI3[4][130] ), .Z(\SB4_10/i0_4 ) );
  BUF_X2 \SB2_1_4/BUF_5  ( .A(\RI3[1][167] ), .Z(\SB2_1_4/i0_3 ) );
  BUF_X2 \SB2_3_26/BUF_2  ( .A(\RI3[3][32] ), .Z(\SB2_3_26/i0_0 ) );
  BUF_X2 \SB2_1_16/BUF_5  ( .A(\RI3[1][95] ), .Z(\SB2_1_16/i0_3 ) );
  BUF_X2 \SB4_26/BUF_4  ( .A(\RI3[4][34] ), .Z(\SB4_26/i0_4 ) );
  BUF_X2 \SB2_1_29/BUF_3  ( .A(\RI3[1][15] ), .Z(\SB2_1_29/i0[10] ) );
  BUF_X2 \SB2_2_10/BUF_3  ( .A(\RI3[2][129] ), .Z(\SB2_2_10/i0[10] ) );
  BUF_X2 \SB4_22/BUF_4  ( .A(\RI3[4][58] ), .Z(\SB4_22/i0_4 ) );
  INV_X2 \SB1_1_31/INV_5  ( .A(\RI1[1][5] ), .ZN(\SB1_1_31/i0_3 ) );
  BUF_X2 \SB2_0_22/BUF_5  ( .A(\RI3[0][59] ), .Z(\SB2_0_22/i0_3 ) );
  BUF_X2 \SB4_19/BUF_4  ( .A(\RI3[4][76] ), .Z(\SB4_19/i0_4 ) );
  BUF_X2 \SB2_1_10/BUF_3  ( .A(\RI3[1][129] ), .Z(\SB2_1_10/i0[10] ) );
  BUF_X2 \SB2_3_8/BUF_3  ( .A(\RI3[3][141] ), .Z(\SB2_3_8/i0[10] ) );
  BUF_X2 \SB4_2/BUF_4  ( .A(\RI3[4][178] ), .Z(\SB4_2/i0_4 ) );
  BUF_X2 \SB2_3_30/BUF_3  ( .A(\RI3[3][9] ), .Z(\SB2_3_30/i0[10] ) );
  BUF_X2 \SB2_1_13/BUF_4  ( .A(\RI3[1][112] ), .Z(\SB2_1_13/i0_4 ) );
  BUF_X2 \SB2_0_23/BUF_5  ( .A(\RI3[0][53] ), .Z(\SB2_0_23/i0_3 ) );
  BUF_X2 \SB2_2_3/BUF_3  ( .A(\RI3[2][171] ), .Z(\SB2_2_3/i0[10] ) );
  BUF_X2 \SB2_3_12/BUF_5  ( .A(\RI3[3][119] ), .Z(\SB2_3_12/i0_3 ) );
  BUF_X2 \SB2_0_2/BUF_4  ( .A(\RI3[0][178] ), .Z(\SB2_0_2/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_121  ( .A(\RI5[1][121] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[121] ) );
  BUF_X2 \SB2_1_15/BUF_4  ( .A(\RI3[1][100] ), .Z(\SB2_1_15/i0_4 ) );
  BUF_X2 \SB4_18/BUF_2  ( .A(\RI3[4][80] ), .Z(\SB4_18/i0_0 ) );
  BUF_X2 \SB2_0_24/BUF_4  ( .A(\RI3[0][46] ), .Z(\SB2_0_24/i0_4 ) );
  BUF_X2 \SB2_3_7/BUF_5  ( .A(\RI3[3][149] ), .Z(\SB2_3_7/i0_3 ) );
  BUF_X2 \SB2_0_16/BUF_5  ( .A(\RI3[0][95] ), .Z(\SB2_0_16/i0_3 ) );
  BUF_X2 \SB2_2_5/BUF_2  ( .A(\RI3[2][158] ), .Z(\SB2_2_5/i0_0 ) );
  BUF_X2 \SB2_3_17/BUF_5  ( .A(\RI3[3][89] ), .Z(\SB2_3_17/i0_3 ) );
  BUF_X2 \SB2_3_6/BUF_5  ( .A(\RI3[3][155] ), .Z(\SB2_3_6/i0_3 ) );
  BUF_X2 \SB2_3_27/BUF_5  ( .A(\RI3[3][29] ), .Z(\SB2_3_27/i0_3 ) );
  BUF_X2 \SB2_1_4/BUF_3  ( .A(\RI3[1][165] ), .Z(\SB2_1_4/i0[10] ) );
  BUF_X2 \SB4_1/BUF_2  ( .A(\RI3[4][182] ), .Z(\SB4_1/i0_0 ) );
  BUF_X2 \SB2_2_6/BUF_3  ( .A(\RI3[2][153] ), .Z(\SB2_2_6/i0[10] ) );
  BUF_X2 \SB4_26/BUF_2  ( .A(\RI3[4][32] ), .Z(\SB4_26/i0_0 ) );
  BUF_X2 \SB2_3_28/BUF_5  ( .A(\RI3[3][23] ), .Z(\SB2_3_28/i0_3 ) );
  BUF_X2 \SB4_2/BUF_2  ( .A(\RI3[4][176] ), .Z(\SB4_2/i0_0 ) );
  BUF_X2 \SB2_2_25/BUF_2  ( .A(\RI3[2][38] ), .Z(\SB2_2_25/i0_0 ) );
  BUF_X2 \SB4_20/BUF_2  ( .A(\RI3[4][68] ), .Z(\SB4_20/i0_0 ) );
  BUF_X2 \SB4_23/BUF_4  ( .A(\RI3[4][52] ), .Z(\SB4_23/i0_4 ) );
  BUF_X2 \SB2_1_23/BUF_5  ( .A(\RI3[1][53] ), .Z(\SB2_1_23/i0_3 ) );
  BUF_X2 \SB2_3_22/BUF_5  ( .A(\RI3[3][59] ), .Z(\SB2_3_22/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_88  ( .A(\RI5[0][88] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[88] ) );
  BUF_X2 \SB2_2_11/BUF_2  ( .A(\RI3[2][122] ), .Z(\SB2_2_11/i0_0 ) );
  BUF_X2 \SB4_0/BUF_2  ( .A(\RI3[4][188] ), .Z(\SB4_0/i0_0 ) );
  BUF_X2 \SB4_28/BUF_2  ( .A(\RI3[4][20] ), .Z(\SB4_28/i0_0 ) );
  INV_X2 \SB1_2_14/INV_5  ( .A(\RI1[2][107] ), .ZN(\SB1_2_14/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_90  ( .A(\RI5[2][90] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[90] ) );
  BUF_X2 \SB2_0_20/BUF_5  ( .A(\RI3[0][71] ), .Z(\SB2_0_20/i0_3 ) );
  BUF_X2 \SB2_3_23/BUF_5  ( .A(\RI3[3][53] ), .Z(\SB2_3_23/i0_3 ) );
  BUF_X2 \SB2_2_2/BUF_2  ( .A(\RI3[2][176] ), .Z(\SB2_2_2/i0_0 ) );
  BUF_X2 \SB2_3_5/BUF_5  ( .A(\RI3[3][161] ), .Z(\SB2_3_5/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_84  ( .A(\RI5[2][84] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[84] ) );
  BUF_X2 \SB2_3_18/BUF_5  ( .A(\RI3[3][83] ), .Z(\SB2_3_18/i0_3 ) );
  BUF_X2 \SB2_2_22/BUF_2  ( .A(\RI3[2][56] ), .Z(\SB2_2_22/i0_0 ) );
  BUF_X2 \SB2_0_27/BUF_4  ( .A(\RI3[0][28] ), .Z(\SB2_0_27/i0_4 ) );
  BUF_X2 \SB4_11/BUF_2  ( .A(\RI3[4][122] ), .Z(\SB4_11/i0_0 ) );
  BUF_X2 \SB4_31/BUF_2  ( .A(\RI3[4][2] ), .Z(\SB4_31/i0_0 ) );
  BUF_X2 \SB4_6/BUF_2  ( .A(\RI3[4][152] ), .Z(\SB4_6/i0_0 ) );
  BUF_X2 \SB2_1_8/BUF_3  ( .A(\RI3[1][141] ), .Z(\SB2_1_8/i0[10] ) );
  BUF_X2 \SB2_2_14/BUF_3  ( .A(\RI3[2][105] ), .Z(\SB2_2_14/i0[10] ) );
  BUF_X2 \SB4_13/BUF_4  ( .A(\RI3[4][112] ), .Z(\SB4_13/i0_4 ) );
  BUF_X2 \SB2_2_15/BUF_5  ( .A(\RI3[2][101] ), .Z(\SB2_2_15/i0_3 ) );
  BUF_X2 \SB4_4/BUF_4  ( .A(\RI3[4][166] ), .Z(\SB4_4/i0_4 ) );
  BUF_X2 \SB2_0_13/BUF_5  ( .A(\RI3[0][113] ), .Z(\SB2_0_13/i0_3 ) );
  BUF_X2 \SB2_1_11/BUF_5  ( .A(\RI3[1][125] ), .Z(\SB2_1_11/i0_3 ) );
  BUF_X2 \SB2_0_6/BUF_4  ( .A(\RI3[0][154] ), .Z(\SB2_0_6/i0_4 ) );
  BUF_X2 \SB2_2_19/BUF_2  ( .A(\RI3[2][74] ), .Z(\SB2_2_19/i0_0 ) );
  INV_X2 \SB1_3_17/INV_5  ( .A(\RI1[3][89] ), .ZN(\SB1_3_17/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_160  ( .A(\RI5[0][160] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[160] ) );
  BUF_X2 \SB2_1_2/BUF_3  ( .A(\RI3[1][177] ), .Z(\SB2_1_2/i0[10] ) );
  BUF_X2 \SB2_3_1/BUF_5  ( .A(\RI3[3][185] ), .Z(\SB2_3_1/i0_3 ) );
  BUF_X2 \SB2_3_0/BUF_5  ( .A(\RI3[3][191] ), .Z(\SB2_3_0/i0_3 ) );
  BUF_X2 \SB2_2_0/BUF_2  ( .A(\RI3[2][188] ), .Z(\SB2_2_0/i0_0 ) );
  BUF_X2 \SB2_1_12/BUF_5  ( .A(\RI3[1][119] ), .Z(\SB2_1_12/i0_3 ) );
  BUF_X2 \SB4_23/BUF_2  ( .A(\RI3[4][50] ), .Z(\SB4_23/i0_0 ) );
  BUF_X2 \SB2_3_29/BUF_5  ( .A(\RI3[3][17] ), .Z(\SB2_3_29/i0_3 ) );
  BUF_X2 \SB2_1_7/BUF_5  ( .A(\RI3[1][149] ), .Z(\SB2_1_7/i0_3 ) );
  BUF_X2 \SB2_2_15/BUF_2  ( .A(\RI3[2][98] ), .Z(\SB2_2_15/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_58  ( .A(\RI5[0][58] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[58] ) );
  BUF_X2 \SB4_5/BUF_2  ( .A(\RI3[4][158] ), .Z(\SB4_5/i0_0 ) );
  BUF_X2 \SB2_0_1/BUF_5  ( .A(\RI3[0][185] ), .Z(\SB2_0_1/i0_3 ) );
  BUF_X2 \SB2_2_0/BUF_5  ( .A(\RI3[2][191] ), .Z(\SB2_2_0/i0_3 ) );
  BUF_X2 \SB2_2_31/BUF_5  ( .A(\RI3[2][5] ), .Z(\SB2_2_31/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_4  ( .A(\RI5[2][4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[4] ) );
  BUF_X2 \SB2_0_21/BUF_4  ( .A(\RI3[0][64] ), .Z(\SB2_0_21/i0_4 ) );
  BUF_X2 \SB4_21/BUF_4  ( .A(\RI3[4][64] ), .Z(\SB4_21/i0_4 ) );
  BUF_X2 \SB2_2_18/BUF_5  ( .A(\RI3[2][83] ), .Z(\SB2_2_18/i0_3 ) );
  BUF_X2 \SB2_0_29/BUF_5  ( .A(\RI3[0][17] ), .Z(\SB2_0_29/i0_3 ) );
  BUF_X2 \SB2_2_23/BUF_5  ( .A(\RI3[2][53] ), .Z(\SB2_2_23/i0_3 ) );
  BUF_X2 \SB2_1_17/BUF_4  ( .A(\RI3[1][88] ), .Z(\SB2_1_17/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_114  ( .A(\RI5[1][114] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[114] ) );
  BUF_X2 \SB2_1_19/BUF_5  ( .A(\RI3[1][77] ), .Z(\SB2_1_19/i0_3 ) );
  BUF_X2 \SB2_3_1/BUF_4  ( .A(\RI3[3][184] ), .Z(\SB2_3_1/i0_4 ) );
  INV_X2 \SB1_0_5/INV_5  ( .A(n31), .ZN(\SB1_0_5/i0_3 ) );
  BUF_X2 \SB2_3_24/BUF_5  ( .A(\RI3[3][47] ), .Z(\SB2_3_24/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_180  ( .A(\RI5[2][180] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[180] ) );
  BUF_X2 \SB4_28/BUF_4  ( .A(\RI3[4][22] ), .Z(\SB4_28/i0_4 ) );
  BUF_X2 \SB2_0_3/BUF_3  ( .A(\RI3[0][171] ), .Z(\SB2_0_3/i0[10] ) );
  BUF_X2 \SB4_12/BUF_2  ( .A(\RI3[4][116] ), .Z(\SB4_12/i0_0 ) );
  BUF_X2 \SB2_1_2/BUF_5  ( .A(\RI3[1][179] ), .Z(\SB2_1_2/i0_3 ) );
  BUF_X2 \SB4_4/BUF_3  ( .A(\RI3[4][165] ), .Z(\SB4_4/i0[10] ) );
  INV_X2 \SB1_2_13/INV_5  ( .A(\RI1[2][113] ), .ZN(\SB1_2_13/i0_3 ) );
  BUF_X2 \SB4_24/BUF_2  ( .A(\RI3[4][44] ), .Z(\SB4_24/i0_0 ) );
  BUF_X2 \SB4_2/BUF_3  ( .A(\RI3[4][177] ), .Z(\SB4_2/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_172  ( .A(\RI5[3][172] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[172] ) );
  BUF_X2 \SB2_3_15/BUF_5  ( .A(\RI3[3][101] ), .Z(\SB2_3_15/i0_3 ) );
  BUF_X2 \SB2_2_12/BUF_4  ( .A(\RI3[2][118] ), .Z(\SB2_2_12/i0_4 ) );
  BUF_X2 \SB2_3_4/BUF_5  ( .A(\RI3[3][167] ), .Z(\SB2_3_4/i0_3 ) );
  BUF_X2 \SB2_3_17/BUF_4  ( .A(\RI3[3][88] ), .Z(\SB2_3_17/i0_4 ) );
  BUF_X2 \SB2_2_19/BUF_5  ( .A(\RI3[2][77] ), .Z(\SB2_2_19/i0_3 ) );
  BUF_X2 \SB4_17/BUF_4  ( .A(\RI3[4][88] ), .Z(\SB4_17/i0_4 ) );
  BUF_X2 \SB2_2_8/BUF_5  ( .A(\RI3[2][143] ), .Z(\SB2_2_8/i0_3 ) );
  BUF_X2 \SB2_3_9/BUF_4  ( .A(\RI3[3][136] ), .Z(\SB2_3_9/i0_4 ) );
  INV_X2 \SB1_3_10/INV_5  ( .A(\RI1[3][131] ), .ZN(\SB1_3_10/i0_3 ) );
  BUF_X2 \SB2_1_12/BUF_4  ( .A(\RI3[1][118] ), .Z(\SB2_1_12/i0_4 ) );
  BUF_X2 \SB2_0_16/BUF_4  ( .A(\RI3[0][94] ), .Z(\SB2_0_16/i0_4 ) );
  INV_X2 \SB1_0_17/INV_5  ( .A(n103), .ZN(\SB1_0_17/i0_3 ) );
  BUF_X2 \SB2_2_13/BUF_4  ( .A(\RI3[2][112] ), .Z(\SB2_2_13/i0_4 ) );
  BUF_X2 \SB2_3_16/BUF_5  ( .A(\RI3[3][95] ), .Z(\SB2_3_16/i0_3 ) );
  BUF_X2 \SB2_2_27/BUF_5  ( .A(\RI3[2][29] ), .Z(\SB2_2_27/i0_3 ) );
  BUF_X2 \SB2_2_9/BUF_5  ( .A(\RI3[2][137] ), .Z(\SB2_2_9/i0_3 ) );
  BUF_X2 \SB2_0_10/BUF_5  ( .A(\RI3[0][131] ), .Z(\SB2_0_10/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_190  ( .A(\RI5[1][190] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[190] ) );
  BUF_X2 \SB4_12/BUF_4  ( .A(\RI3[4][118] ), .Z(\SB4_12/i0_4 ) );
  INV_X2 \SB1_1_9/INV_5  ( .A(\RI1[1][137] ), .ZN(\SB1_1_9/i0_3 ) );
  BUF_X2 \SB4_14/BUF_2  ( .A(\RI3[4][104] ), .Z(\SB4_14/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_34  ( .A(\RI5[2][34] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[34] ) );
  BUF_X2 \SB2_0_3/BUF_5  ( .A(\RI3[0][173] ), .Z(\SB2_0_3/i0_3 ) );
  BUF_X2 \SB2_2_25/BUF_5  ( .A(\RI3[2][41] ), .Z(\SB2_2_25/i0_3 ) );
  BUF_X2 \SB2_2_30/BUF_5  ( .A(\RI3[2][11] ), .Z(\SB2_2_30/i0_3 ) );
  BUF_X2 \SB2_1_31/BUF_5  ( .A(\RI3[1][5] ), .Z(\SB2_1_31/i0_3 ) );
  BUF_X2 \SB2_2_17/BUF_5  ( .A(\RI3[2][89] ), .Z(\SB2_2_17/i0_3 ) );
  BUF_X2 \SB2_3_11/BUF_5  ( .A(\RI3[3][125] ), .Z(\SB2_3_11/i0_3 ) );
  BUF_X2 \SB2_0_29/BUF_4  ( .A(\RI3[0][16] ), .Z(\SB2_0_29/i0_4 ) );
  BUF_X2 \SB2_1_16/BUF_4  ( .A(\RI3[1][94] ), .Z(\SB2_1_16/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_120  ( .A(\RI5[1][120] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[120] ) );
  BUF_X2 \SB2_2_8/BUF_3  ( .A(\RI3[2][141] ), .Z(\SB2_2_8/i0[10] ) );
  INV_X2 \SB1_2_10/INV_5  ( .A(\RI1[2][131] ), .ZN(\SB1_2_10/i0_3 ) );
  BUF_X2 \SB4_21/BUF_2  ( .A(\RI3[4][62] ), .Z(\SB4_21/i0_0 ) );
  BUF_X2 \SB2_1_17/BUF_5  ( .A(\RI3[1][89] ), .Z(\SB2_1_17/i0_3 ) );
  BUF_X2 \SB2_2_21/BUF_5  ( .A(\RI3[2][65] ), .Z(\SB2_2_21/i0_3 ) );
  BUF_X2 \SB2_1_21/BUF_5  ( .A(\RI3[1][65] ), .Z(\SB2_1_21/i0_3 ) );
  BUF_X2 \SB2_0_28/BUF_5  ( .A(\RI3[0][23] ), .Z(\SB2_0_28/i0_3 ) );
  BUF_X2 \SB2_3_26/BUF_5  ( .A(\RI3[3][35] ), .Z(\SB2_3_26/i0_3 ) );
  BUF_X2 \SB2_2_1/BUF_5  ( .A(\RI3[2][185] ), .Z(\SB2_2_1/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_70  ( .A(\RI5[2][70] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[70] ) );
  BUF_X2 \SB2_3_8/BUF_5  ( .A(\RI3[3][143] ), .Z(\SB2_3_8/i0_3 ) );
  BUF_X2 \SB2_2_26/BUF_3  ( .A(\RI3[2][33] ), .Z(\SB2_2_26/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_28  ( .A(\RI5[0][28] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[28] ) );
  BUF_X2 \SB2_2_30/BUF_4  ( .A(\RI3[2][10] ), .Z(\SB2_2_30/i0_4 ) );
  BUF_X2 \SB2_0_12/BUF_5  ( .A(\RI3[0][119] ), .Z(\SB2_0_12/i0_3 ) );
  BUF_X2 \SB2_0_27/BUF_5  ( .A(\RI3[0][29] ), .Z(\SB2_0_27/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_70  ( .A(\RI5[1][70] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[70] ) );
  BUF_X2 \SB2_1_9/BUF_5  ( .A(\RI3[1][137] ), .Z(\SB2_1_9/i0_3 ) );
  BUF_X2 \SB2_3_10/BUF_5  ( .A(\RI3[3][131] ), .Z(\SB2_3_10/i0_3 ) );
  BUF_X2 \SB2_0_4/BUF_4  ( .A(\RI3[0][166] ), .Z(\SB2_0_4/i0_4 ) );
  BUF_X2 \SB2_2_14/BUF_4  ( .A(\RI3[2][106] ), .Z(\SB2_2_14/i0_4 ) );
  BUF_X2 \SB4_16/BUF_2  ( .A(\RI3[4][92] ), .Z(\SB4_16/i0_0 ) );
  INV_X2 \SB1_2_15/INV_5  ( .A(\RI1[2][101] ), .ZN(\SB1_2_15/i0_3 ) );
  BUF_X2 \SB2_2_11/BUF_5  ( .A(\RI3[2][125] ), .Z(\SB2_2_11/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_32  ( .A(\RI5[1][32] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[32] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_102  ( .A(\RI5[3][102] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[102] ) );
  BUF_X2 \SB2_0_30/BUF_3  ( .A(\RI3[0][9] ), .Z(\SB2_0_30/i0[10] ) );
  BUF_X2 \SB4_29/BUF_2  ( .A(\RI3[4][14] ), .Z(\SB4_29/i0_0 ) );
  BUF_X2 \SB2_2_13/BUF_3  ( .A(\RI3[2][111] ), .Z(\SB2_2_13/i0[10] ) );
  BUF_X2 \SB2_3_21/BUF_5  ( .A(\RI3[3][65] ), .Z(\SB2_3_21/i0_3 ) );
  BUF_X2 \SB2_0_15/BUF_5  ( .A(\RI3[0][101] ), .Z(\SB2_0_15/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_52  ( .A(\RI5[0][52] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[52] ) );
  BUF_X2 \SB2_3_2/BUF_4  ( .A(\RI3[3][178] ), .Z(\SB2_3_2/i0_4 ) );
  BUF_X2 \SB2_1_24/BUF_4  ( .A(\RI3[1][46] ), .Z(\SB2_1_24/i0_4 ) );
  BUF_X2 \SB2_1_29/BUF_5  ( .A(\RI3[1][17] ), .Z(\SB2_1_29/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_88  ( .A(\RI5[1][88] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[88] ) );
  BUF_X2 \SB2_1_18/BUF_5  ( .A(\RI3[1][83] ), .Z(\SB2_1_18/i0_3 ) );
  BUF_X2 \SB2_3_13/BUF_5  ( .A(\RI3[3][113] ), .Z(\SB2_3_13/i0_3 ) );
  BUF_X2 \SB4_3/BUF_4  ( .A(\RI3[4][172] ), .Z(\SB4_3/i0_4 ) );
  BUF_X2 \SB2_2_27/BUF_4  ( .A(\RI3[2][28] ), .Z(\SB2_2_27/i0_4 ) );
  BUF_X2 \SB4_7/BUF_2  ( .A(\RI3[4][146] ), .Z(\SB4_7/i0_0 ) );
  BUF_X2 \SB2_1_7/BUF_2  ( .A(\RI3[1][146] ), .Z(\SB2_1_7/i0_0 ) );
  BUF_X2 \SB2_0_31/BUF_5  ( .A(\RI3[0][5] ), .Z(\SB2_0_31/i0_3 ) );
  BUF_X2 \SB2_1_26/BUF_5  ( .A(\RI3[1][35] ), .Z(\SB2_1_26/i0_3 ) );
  INV_X2 \SB1_2_6/INV_5  ( .A(\RI1[2][155] ), .ZN(\SB1_2_6/i0_3 ) );
  BUF_X2 \SB2_2_4/BUF_4  ( .A(\RI3[2][166] ), .Z(\SB2_2_4/i0_4 ) );
  BUF_X2 \SB2_2_14/BUF_5  ( .A(\RI3[2][107] ), .Z(\SB2_2_14/i0_3 ) );
  BUF_X2 \SB2_1_18/BUF_4  ( .A(\RI3[1][82] ), .Z(\SB2_1_18/i0_4 ) );
  BUF_X2 \SB2_2_22/BUF_5  ( .A(\RI3[2][59] ), .Z(\SB2_2_22/i0_3 ) );
  BUF_X2 \SB2_2_26/BUF_5  ( .A(\RI3[2][35] ), .Z(\SB2_2_26/i0_3 ) );
  INV_X2 \SB1_0_18/INV_5  ( .A(n109), .ZN(\SB1_0_18/i0_3 ) );
  BUF_X2 \SB2_3_9/BUF_5  ( .A(\RI3[3][137] ), .Z(\SB2_3_9/i0_3 ) );
  BUF_X2 \SB2_1_14/BUF_5  ( .A(\RI3[1][107] ), .Z(\SB2_1_14/i0_3 ) );
  BUF_X2 \SB2_3_3/BUF_3  ( .A(\RI3[3][171] ), .Z(\SB2_3_3/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_78  ( .A(\RI5[2][78] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[78] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_64  ( .A(\RI5[2][64] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[64] ) );
  INV_X2 \SB1_3_5/INV_5  ( .A(\RI1[3][161] ), .ZN(\SB1_3_5/i0_3 ) );
  BUF_X2 \SB4_11/BUF_3  ( .A(\RI3[4][123] ), .Z(\SB4_11/i0[10] ) );
  BUF_X2 \SB2_1_28/BUF_5  ( .A(\RI3[1][23] ), .Z(\SB2_1_28/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_158  ( .A(\RI5[1][158] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[158] ) );
  BUF_X2 \SB2_3_19/BUF_5  ( .A(\RI3[3][77] ), .Z(\SB2_3_19/i0_3 ) );
  INV_X2 \SB1_2_7/INV_5  ( .A(\RI1[2][149] ), .ZN(\SB1_2_7/i0_3 ) );
  BUF_X2 \SB2_2_28/BUF_5  ( .A(\RI3[2][23] ), .Z(\SB2_2_28/i0_3 ) );
  BUF_X2 \SB2_2_6/BUF_4  ( .A(\RI3[2][154] ), .Z(\SB2_2_6/i0_4 ) );
  BUF_X2 \SB2_1_8/BUF_4  ( .A(\RI3[1][142] ), .Z(\SB2_1_8/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_46  ( .A(\RI5[1][46] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[46] ) );
  BUF_X2 \SB2_3_30/BUF_5  ( .A(\RI3[3][11] ), .Z(\SB2_3_30/i0_3 ) );
  BUF_X2 \SB2_1_25/BUF_5  ( .A(\RI3[1][41] ), .Z(\SB2_1_25/i0_3 ) );
  BUF_X2 \SB2_3_31/BUF_5  ( .A(\RI3[3][5] ), .Z(\SB2_3_31/i0_3 ) );
  BUF_X2 \SB4_19/BUF_3  ( .A(\RI3[4][75] ), .Z(\SB4_19/i0[10] ) );
  BUF_X2 \SB4_8/BUF_3  ( .A(\RI3[4][141] ), .Z(\SB4_8/i0[10] ) );
  BUF_X2 \SB2_2_29/BUF_4  ( .A(\RI3[2][16] ), .Z(\SB2_2_29/i0_4 ) );
  BUF_X2 \SB4_18/BUF_3  ( .A(\RI3[4][81] ), .Z(\SB4_18/i0[10] ) );
  BUF_X2 \SB2_0_1/BUF_4  ( .A(\RI3[0][184] ), .Z(\SB2_0_1/i0_4 ) );
  BUF_X2 \SB2_1_13/BUF_5  ( .A(\RI3[1][113] ), .Z(\SB2_1_13/i0_3 ) );
  BUF_X2 \SB2_2_23/BUF_4  ( .A(\RI3[2][52] ), .Z(\SB2_2_23/i0_4 ) );
  BUF_X2 \SB2_3_20/BUF_5  ( .A(\RI3[3][71] ), .Z(\SB2_3_20/i0_3 ) );
  BUF_X2 \SB2_1_24/BUF_5  ( .A(\RI3[1][47] ), .Z(\SB2_1_24/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_73  ( .A(\RI5[2][73] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[73] ) );
  BUF_X2 \SB2_3_25/BUF_5  ( .A(\RI3[3][41] ), .Z(\SB2_3_25/i0_3 ) );
  BUF_X2 \SB2_2_1/BUF_4  ( .A(\RI3[2][184] ), .Z(\SB2_2_1/i0_4 ) );
  BUF_X2 \SB4_29/BUF_3  ( .A(\RI3[4][15] ), .Z(\SB4_29/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_166  ( .A(\RI5[0][166] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[166] ) );
  BUF_X2 \SB2_2_13/BUF_5  ( .A(\RI3[2][113] ), .Z(\SB2_2_13/i0_3 ) );
  INV_X2 \SB1_1_23/INV_5  ( .A(\RI1[1][53] ), .ZN(\SB1_1_23/i0_3 ) );
  BUF_X2 \SB2_3_2/BUF_3  ( .A(\RI3[3][177] ), .Z(\SB2_3_2/i0[10] ) );
  INV_X2 \SB1_3_4/INV_5  ( .A(\RI1[3][167] ), .ZN(\SB1_3_4/i0_3 ) );
  BUF_X2 \SB2_0_0/BUF_5  ( .A(\RI3[0][191] ), .Z(\SB2_0_0/i0_3 ) );
  BUF_X2 \SB2_1_10/BUF_5  ( .A(\RI3[1][131] ), .Z(\SB2_1_10/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_79  ( .A(\RI5[1][79] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[79] ) );
  BUF_X2 \SB2_1_22/BUF_4  ( .A(\RI3[1][58] ), .Z(\SB2_1_22/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_91  ( .A(\RI5[2][91] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[91] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_12  ( .A(\RI5[3][12] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[12] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_166  ( .A(\RI5[2][166] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[166] ) );
  BUF_X2 \SB2_2_5/BUF_5  ( .A(\RI3[2][161] ), .Z(\SB2_2_5/i0_3 ) );
  BUF_X2 \SB2_3_27/BUF_4  ( .A(\RI3[3][28] ), .Z(\SB2_3_27/i0_4 ) );
  BUF_X2 \SB2_1_15/BUF_3  ( .A(\RI3[1][99] ), .Z(\SB2_1_15/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_126  ( .A(\RI5[1][126] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[126] ) );
  BUF_X2 \SB1_1_17/BUF_2  ( .A(\RI1[1][86] ), .Z(\SB1_1_17/i1[9] ) );
  BUF_X2 \SB4_26/BUF_3  ( .A(\RI3[4][33] ), .Z(\SB4_26/i0[10] ) );
  BUF_X2 \SB4_27/BUF_3  ( .A(\RI3[4][27] ), .Z(\SB4_27/i0[10] ) );
  BUF_X2 \SB2_1_0/BUF_5  ( .A(\RI3[1][191] ), .Z(\SB2_1_0/i0_3 ) );
  BUF_X2 \SB2_3_0/BUF_4  ( .A(\RI3[3][190] ), .Z(\SB2_3_0/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_151  ( .A(\RI5[2][151] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[151] ) );
  BUF_X2 \SB4_16/BUF_3  ( .A(\RI3[4][93] ), .Z(\SB4_16/i0[10] ) );
  BUF_X2 \SB2_2_10/BUF_4  ( .A(\RI3[2][130] ), .Z(\SB2_2_10/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_16  ( .A(\RI5[1][16] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[16] ) );
  BUF_X2 \SB2_1_30/BUF_5  ( .A(\RI3[1][11] ), .Z(\SB2_1_30/i0_3 ) );
  BUF_X2 \SB2_2_20/BUF_5  ( .A(\RI3[2][71] ), .Z(\SB2_2_20/i0_3 ) );
  BUF_X2 \SB4_27/BUF_2  ( .A(\RI3[4][26] ), .Z(\SB4_27/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_34  ( .A(\RI5[1][34] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[34] ) );
  BUF_X2 \SB2_3_25/BUF_3  ( .A(\RI3[3][39] ), .Z(\SB2_3_25/i0[10] ) );
  BUF_X2 \SB2_3_1/BUF_3  ( .A(\RI3[3][183] ), .Z(\SB2_3_1/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_127  ( .A(\RI5[0][127] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[127] ) );
  BUF_X2 \SB2_2_16/BUF_4  ( .A(\RI3[2][94] ), .Z(\SB2_2_16/i0_4 ) );
  BUF_X2 \SB2_0_24/BUF_2  ( .A(\RI3[0][44] ), .Z(\SB2_0_24/i0_0 ) );
  BUF_X2 \SB2_1_8/BUF_5  ( .A(\RI3[1][143] ), .Z(\SB2_1_8/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_55  ( .A(\RI5[2][55] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[55] ) );
  BUF_X2 \SB2_3_5/BUF_3  ( .A(\RI3[3][159] ), .Z(\SB2_3_5/i0[10] ) );
  BUF_X2 \SB2_2_5/BUF_4  ( .A(\RI3[2][160] ), .Z(\SB2_2_5/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_25  ( .A(\RI5[1][25] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[25] ) );
  BUF_X2 \SB2_0_30/BUF_4  ( .A(\RI3[0][10] ), .Z(\SB2_0_30/i0_4 ) );
  BUF_X2 \SB2_0_13/BUF_4  ( .A(\RI3[0][112] ), .Z(\SB2_0_13/i0_4 ) );
  BUF_X2 \SB2_2_28/BUF_4  ( .A(\RI3[2][22] ), .Z(\SB2_2_28/i0_4 ) );
  BUF_X2 \SB2_3_28/BUF_3  ( .A(\RI3[3][21] ), .Z(\SB2_3_28/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_133  ( .A(\RI5[0][133] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[133] ) );
  BUF_X2 \SB2_1_20/BUF_5  ( .A(\RI3[1][71] ), .Z(\SB2_1_20/i0_3 ) );
  BUF_X2 \SB2_1_14/BUF_4  ( .A(\RI3[1][106] ), .Z(\SB2_1_14/i0_4 ) );
  BUF_X2 \SB2_3_31/BUF_3  ( .A(\RI3[3][3] ), .Z(\SB2_3_31/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_64  ( .A(\RI5[1][64] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[64] ) );
  BUF_X2 \SB2_2_21/BUF_4  ( .A(\RI3[2][64] ), .Z(\SB2_2_21/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_91  ( .A(\RI5[1][91] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[91] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_169  ( .A(\RI5[2][169] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[169] ) );
  BUF_X2 \SB2_1_20/BUF_4  ( .A(\RI3[1][70] ), .Z(\SB2_1_20/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_85  ( .A(\RI5[2][85] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[85] ) );
  BUF_X2 \SB2_3_19/BUF_4  ( .A(\RI3[3][76] ), .Z(\SB2_3_19/i0_4 ) );
  BUF_X2 \SB2_3_10/BUF_4  ( .A(\RI3[3][130] ), .Z(\SB2_3_10/i0_4 ) );
  BUF_X2 \SB4_31/BUF_3  ( .A(\RI3[4][3] ), .Z(\SB4_31/i0[10] ) );
  BUF_X2 \SB4_21/BUF_3  ( .A(\RI3[4][63] ), .Z(\SB4_21/i0[10] ) );
  BUF_X2 \SB2_0_9/BUF_4  ( .A(\RI3[0][136] ), .Z(\SB2_0_9/i0_4 ) );
  BUF_X2 \SB2_3_4/BUF_3  ( .A(\RI3[3][165] ), .Z(\SB2_3_4/i0[10] ) );
  BUF_X2 \SB2_1_27/BUF_4  ( .A(\RI3[1][28] ), .Z(\SB2_1_27/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_49  ( .A(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[49] ) );
  BUF_X2 \SB2_0_21/BUF_5  ( .A(\RI3[0][65] ), .Z(\SB2_0_21/i0_3 ) );
  BUF_X2 \SB2_0_0/BUF_4  ( .A(\RI3[0][190] ), .Z(\SB2_0_0/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_24  ( .A(\RI5[1][24] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[24] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_19  ( .A(\RI5[0][19] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[19] ) );
  BUF_X2 \SB2_1_0/BUF_3  ( .A(\RI3[1][189] ), .Z(\SB2_1_0/i0[10] ) );
  BUF_X2 \SB4_30/BUF_3  ( .A(\RI3[4][9] ), .Z(\SB4_30/i0[10] ) );
  BUF_X2 \SB2_3_6/BUF_3  ( .A(\RI3[3][153] ), .Z(\SB2_3_6/i0[10] ) );
  BUF_X2 \SB4_14/BUF_3  ( .A(\RI3[4][105] ), .Z(\SB4_14/i0[10] ) );
  BUF_X2 \SB2_0_28/BUF_4  ( .A(\RI3[0][22] ), .Z(\SB2_0_28/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_7  ( .A(\RI5[1][7] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[7] ) );
  BUF_X2 \SB2_3_0/BUF_3  ( .A(\RI3[3][189] ), .Z(\SB2_3_0/i0[10] ) );
  BUF_X2 \SB2_1_2/BUF_4  ( .A(\RI3[1][178] ), .Z(\SB2_1_2/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_43  ( .A(\RI5[0][43] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[43] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_73  ( .A(\RI5[1][73] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[73] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_163  ( .A(\RI5[1][163] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[163] ) );
  BUF_X2 \SB2_2_20/BUF_4  ( .A(\RI3[2][70] ), .Z(\SB2_2_20/i0_4 ) );
  BUF_X2 \SB2_2_22/BUF_3  ( .A(\RI3[2][57] ), .Z(\SB2_2_22/i0[10] ) );
  BUF_X2 \SB2_3_19/BUF_3  ( .A(\RI3[3][75] ), .Z(\SB2_3_19/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_96  ( .A(\RI5[2][96] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[96] ) );
  BUF_X2 \SB4_28/BUF_3  ( .A(\RI3[4][21] ), .Z(\SB4_28/i0[10] ) );
  BUF_X2 \SB2_1_0/BUF_4  ( .A(\RI3[1][190] ), .Z(\SB2_1_0/i0_4 ) );
  BUF_X2 \SB2_3_6/BUF_2  ( .A(\RI3[3][152] ), .Z(\SB2_3_6/i0_0 ) );
  BUF_X2 \SB2_1_5/BUF_4  ( .A(\RI3[1][160] ), .Z(\SB2_1_5/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_97  ( .A(\RI5[1][97] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[97] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_133  ( .A(\RI5[1][133] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[133] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_36  ( .A(\RI5[2][36] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[36] ) );
  BUF_X2 \SB2_2_30/BUF_3  ( .A(\RI3[2][9] ), .Z(\SB2_2_30/i0[10] ) );
  BUF_X2 \SB2_3_29/BUF_3  ( .A(\RI3[3][15] ), .Z(\SB2_3_29/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_115  ( .A(\RI5[1][115] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[115] ) );
  INV_X2 \SB1_3_18/INV_5  ( .A(\RI1[3][83] ), .ZN(\SB1_3_18/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_103  ( .A(\RI5[0][103] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[103] ) );
  BUF_X2 \SB2_2_17/BUF_3  ( .A(\RI3[2][87] ), .Z(\SB2_2_17/i0[10] ) );
  INV_X2 \SB1_0_12/INV_5  ( .A(n73), .ZN(\SB1_0_12/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_67  ( .A(\RI5[2][67] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[67] ) );
  BUF_X2 \SB2_0_11/BUF_4  ( .A(\RI3[0][124] ), .Z(\SB2_0_11/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_68  ( .A(\RI5[0][68] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[68] ) );
  INV_X2 \SB1_0_13/INV_5  ( .A(n79), .ZN(\SB1_0_13/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_139  ( .A(\RI5[0][139] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[139] ) );
  BUF_X2 \SB2_0_12/BUF_4  ( .A(\RI3[0][118] ), .Z(\SB2_0_12/i0_4 ) );
  BUF_X2 \SB2_2_18/BUF_3  ( .A(\RI3[2][81] ), .Z(\SB2_2_18/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_97  ( .A(\RI5[2][97] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[97] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_49  ( .A(\RI5[2][49] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[49] ) );
  BUF_X2 \SB2_3_16/BUF_3  ( .A(\RI3[3][93] ), .Z(\SB2_3_16/i0[10] ) );
  BUF_X2 \SB2_2_31/BUF_3  ( .A(\RI3[2][3] ), .Z(\SB2_2_31/i0[10] ) );
  BUF_X2 \SB2_2_16/BUF_3  ( .A(\RI3[2][93] ), .Z(\SB2_2_16/i0[10] ) );
  BUF_X2 \SB2_3_29/BUF_2  ( .A(\RI3[3][14] ), .Z(\SB2_3_29/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_120  ( .A(\RI5[2][120] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[120] ) );
  BUF_X2 \SB4_3/BUF_3  ( .A(\RI3[4][171] ), .Z(\SB4_3/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_94  ( .A(\RI5[0][94] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[94] ) );
  BUF_X2 \SB2_0_22/BUF_4  ( .A(\RI3[0][58] ), .Z(\SB2_0_22/i0_4 ) );
  INV_X2 \SB1_0_23/INV_5  ( .A(n139), .ZN(\SB1_0_23/i0_3 ) );
  BUF_X2 \SB2_2_2/BUF_3  ( .A(\RI3[2][177] ), .Z(\SB2_2_2/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_12  ( .A(\RI5[2][12] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[12] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_145  ( .A(\RI5[1][145] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[145] ) );
  BUF_X2 \SB2_2_11/BUF_3  ( .A(\RI3[2][123] ), .Z(\SB2_2_11/i0[10] ) );
  BUF_X2 \SB2_3_13/BUF_3  ( .A(\RI3[3][111] ), .Z(\SB2_3_13/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_150  ( .A(\RI5[2][150] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[150] ) );
  BUF_X2 \SB2_2_27/BUF_3  ( .A(\RI3[2][27] ), .Z(\SB2_2_27/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_37  ( .A(\RI5[0][37] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[37] ) );
  BUF_X2 \SB2_2_28/BUF_2  ( .A(\RI3[2][20] ), .Z(\SB2_2_28/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_54  ( .A(\RI5[2][54] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[54] ) );
  BUF_X2 \SB2_1_20/BUF_3  ( .A(\RI3[1][69] ), .Z(\SB2_1_20/i0[10] ) );
  BUF_X2 \SB2_1_5/BUF_3  ( .A(\RI3[1][159] ), .Z(\SB2_1_5/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_145  ( .A(\RI5[2][145] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[145] ) );
  BUF_X2 \SB2_3_14/BUF_3  ( .A(\RI3[3][105] ), .Z(\SB2_3_14/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_96  ( .A(\RI5[1][96] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[96] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_19  ( .A(\RI5[1][19] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[19] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_157  ( .A(\RI5[2][157] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[157] ) );
  BUF_X2 \SB2_2_4/BUF_3  ( .A(\RI3[2][165] ), .Z(\SB2_2_4/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_114  ( .A(\RI5[2][114] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[114] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_162  ( .A(\RI5[0][162] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[162] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_37  ( .A(\RI5[1][37] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[37] ) );
  INV_X2 \SB1_1_25/INV_5  ( .A(\RI1[1][41] ), .ZN(\SB1_1_25/i0_3 ) );
  BUF_X2 \SB2_2_0/BUF_3  ( .A(\RI3[2][189] ), .Z(\SB2_2_0/i0[10] ) );
  BUF_X2 \SB2_1_22/BUF_2  ( .A(\RI3[1][56] ), .Z(\SB2_1_22/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_24  ( .A(\RI5[2][24] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[24] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_84  ( .A(\RI5[1][84] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[84] ) );
  BUF_X2 \SB2_3_10/BUF_3  ( .A(\RI3[3][129] ), .Z(\SB2_3_10/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_109  ( .A(\RI5[0][109] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[109] ) );
  INV_X2 \SB1_3_29/INV_5  ( .A(\RI1[3][17] ), .ZN(\SB1_3_29/i0_3 ) );
  BUF_X2 \SB2_1_19/BUF_2  ( .A(\RI3[1][74] ), .Z(\SB2_1_19/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_102  ( .A(\RI5[1][102] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[102] ) );
  INV_X2 \SB1_1_22/INV_5  ( .A(\RI1[1][59] ), .ZN(\SB1_1_22/i0_3 ) );
  INV_X2 \SB1_3_31/INV_5  ( .A(\RI1[3][5] ), .ZN(\SB1_3_31/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_139  ( .A(\RI5[2][139] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[139] ) );
  BUF_X2 \SB4_22/BUF_2  ( .A(\RI3[4][56] ), .Z(\SB4_22/i0_0 ) );
  BUF_X2 \SB2_3_7/BUF_3  ( .A(\RI3[3][147] ), .Z(\SB2_3_7/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_103  ( .A(\RI5[2][103] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[103] ) );
  BUF_X2 \SB2_1_31/BUF_4  ( .A(\RI3[1][4] ), .Z(\SB2_1_31/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_97  ( .A(\RI5[0][97] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[97] ) );
  BUF_X2 \SB2_2_20/BUF_2  ( .A(\RI3[2][68] ), .Z(\SB2_2_20/i0_0 ) );
  BUF_X2 \SB2_0_12/BUF_3  ( .A(\RI3[0][117] ), .Z(\SB2_0_12/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_144  ( .A(\RI5[0][144] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[144] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_138  ( .A(\RI5[0][138] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[138] ) );
  BUF_X2 \SB2_2_23/BUF_3  ( .A(\RI3[2][51] ), .Z(\SB2_2_23/i0[10] ) );
  INV_X2 \SB1_2_25/INV_5  ( .A(\RI1[2][41] ), .ZN(\SB1_2_25/i0_3 ) );
  BUF_X2 \SB2_2_29/BUF_2  ( .A(\RI3[2][14] ), .Z(\SB2_2_29/i0_0 ) );
  INV_X2 \SB1_2_0/INV_5  ( .A(\RI1[2][191] ), .ZN(\SB1_2_0/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_13  ( .A(\RI5[1][13] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[13] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_121  ( .A(\RI5[2][121] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[121] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_181  ( .A(\RI5[0][181] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[181] ) );
  BUF_X2 \SB2_3_16/BUF_2  ( .A(\RI3[3][92] ), .Z(\SB2_3_16/i0_0 ) );
  BUF_X2 \SB2_3_26/BUF_3  ( .A(\RI3[3][33] ), .Z(\SB2_3_26/i0[10] ) );
  BUF_X2 \SB2_0_5/BUF_4  ( .A(\RI3[0][160] ), .Z(\SB2_0_5/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_178  ( .A(\RI5[2][178] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[178] ) );
  BUF_X2 \SB2_0_20/BUF_4  ( .A(\RI3[0][70] ), .Z(\SB2_0_20/i0_4 ) );
  INV_X2 \SB1_1_26/INV_5  ( .A(\RI1[1][35] ), .ZN(\SB1_1_26/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_4  ( .A(\RI5[0][4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[4] ) );
  BUF_X2 \SB2_0_8/BUF_4  ( .A(\RI3[0][142] ), .Z(\SB2_0_8/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_18  ( .A(\RI5[0][18] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[18] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_54  ( .A(\RI5[1][54] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[54] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_151  ( .A(\RI5[1][151] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[151] ) );
  BUF_X2 \SB4_23/BUF_3  ( .A(\RI3[4][51] ), .Z(\SB4_23/i0[10] ) );
  INV_X2 \SB1_3_7/INV_5  ( .A(\RI1[3][149] ), .ZN(\SB1_3_7/i0_3 ) );
  BUF_X2 \SB4_7/BUF_3  ( .A(\RI3[4][147] ), .Z(\SB4_7/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_115  ( .A(\RI5[0][115] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[115] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_66  ( .A(\RI5[2][66] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[66] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_1  ( .A(\RI5[1][1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[1] ) );
  BUF_X2 \SB2_3_17/BUF_2  ( .A(\RI3[3][86] ), .Z(\SB2_3_17/i0_0 ) );
  INV_X2 \SB1_3_8/INV_5  ( .A(\RI1[3][143] ), .ZN(\SB1_3_8/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_37  ( .A(\RI5[2][37] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[37] ) );
  BUF_X2 \SB2_3_21/BUF_2  ( .A(\RI3[3][62] ), .Z(\SB2_3_21/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_109  ( .A(\RI5[2][109] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[109] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_55  ( .A(\RI5[1][55] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[55] ) );
  BUF_X2 \SB4_6/BUF_3  ( .A(\RI3[4][153] ), .Z(\SB4_6/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_82  ( .A(\RI5[2][82] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[82] ) );
  BUF_X2 \SB4_12/BUF_3  ( .A(\RI3[4][117] ), .Z(\SB4_12/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_13  ( .A(\RI5[2][13] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[13] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_61  ( .A(\RI5[0][61] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[61] ) );
  BUF_X2 \SB4_20/BUF_3  ( .A(\RI3[4][69] ), .Z(\SB4_20/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_60  ( .A(\RI5[2][60] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[60] ) );
  BUF_X2 \SB2_3_13/BUF_2  ( .A(\RI3[3][110] ), .Z(\SB2_3_13/i0_0 ) );
  BUF_X2 \SB2_3_19/BUF_2  ( .A(\RI3[3][74] ), .Z(\SB2_3_19/i0_0 ) );
  BUF_X2 \SB2_2_18/BUF_2  ( .A(\RI3[2][80] ), .Z(\SB2_2_18/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_151  ( .A(\RI5[0][151] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[151] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_49  ( .A(\RI5[0][49] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[49] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_73  ( .A(\RI5[0][73] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[73] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_18  ( .A(\RI5[1][18] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[18] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_172  ( .A(\RI5[1][172] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[172] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_127  ( .A(\RI5[2][127] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[127] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_48  ( .A(\RI5[1][48] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[48] ) );
  BUF_X2 \SB2_0_26/BUF_4  ( .A(\RI3[0][34] ), .Z(\SB2_0_26/i0_4 ) );
  INV_X2 \SB1_1_28/INV_5  ( .A(\RI1[1][23] ), .ZN(\SB1_1_28/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_79  ( .A(\RI5[0][79] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[79] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_22  ( .A(\RI5[1][22] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[22] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_102  ( .A(\RI5[2][102] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[102] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_67  ( .A(\RI5[0][67] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[67] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_166  ( .A(\RI5[1][166] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[166] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_175  ( .A(\RI5[0][175] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[175] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_30  ( .A(\RI5[2][30] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[30] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_175  ( .A(\RI5[2][175] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[175] ) );
  INV_X2 \SB1_2_31/INV_5  ( .A(\RI1[2][5] ), .ZN(\SB1_2_31/i0_3 ) );
  BUF_X2 \SB2_2_7/BUF_2  ( .A(\RI3[2][146] ), .Z(\SB2_2_7/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_109  ( .A(\RI5[1][109] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[109] ) );
  BUF_X2 \SB2_1_5/BUF_2  ( .A(\RI3[1][158] ), .Z(\SB2_1_5/i0_0 ) );
  BUF_X2 \SB2_1_17/BUF_2  ( .A(\RI3[1][86] ), .Z(\SB2_1_17/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_78  ( .A(\RI5[1][78] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[78] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_7  ( .A(\RI5[2][7] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[7] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_186  ( .A(\RI5[2][186] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[186] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_174  ( .A(\RI5[2][174] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[174] ) );
  BUF_X2 \SB4_10/BUF_3  ( .A(\RI3[4][129] ), .Z(\SB4_10/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_94  ( .A(\RI5[1][94] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[94] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_18  ( .A(\RI5[2][18] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[18] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_13  ( .A(\RI5[0][13] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[13] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_85  ( .A(\RI5[1][85] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[85] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_126  ( .A(\RI5[2][126] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[126] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_124  ( .A(\RI5[0][124] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[124] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_136  ( .A(\RI5[1][136] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[136] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_72  ( .A(\RI5[0][72] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[72] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_46  ( .A(\RI5[2][46] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[46] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_6  ( .A(\RI5[2][6] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[6] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_16  ( .A(\RI5[2][16] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[16] ) );
  INV_X2 \SB1_2_3/INV_5  ( .A(\RI1[2][173] ), .ZN(\SB1_2_3/i0_3 ) );
  INV_X2 \SB1_1_18/INV_5  ( .A(\RI1[1][83] ), .ZN(\SB1_1_18/i0_3 ) );
  INV_X2 \SB1_1_7/INV_5  ( .A(\RI1[1][149] ), .ZN(\SB1_1_7/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_48  ( .A(\RI5[0][48] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[48] ) );
  BUF_X2 \SB4_15/BUF_3  ( .A(\RI3[4][99] ), .Z(\SB4_15/i0[10] ) );
  BUF_X2 \SB4_10/BUF_2  ( .A(\RI3[4][128] ), .Z(\SB4_10/i0_0 ) );
  BUF_X2 \SB4_1/BUF_3  ( .A(\RI3[4][183] ), .Z(\SB4_1/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_168  ( .A(\RI5[1][168] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[168] ) );
  INV_X2 \SB1_3_9/INV_5  ( .A(\RI1[3][137] ), .ZN(\SB1_3_9/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_12  ( .A(\RI5[1][12] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[12] ) );
  INV_X2 \SB1_1_2/INV_5  ( .A(\RI1[1][179] ), .ZN(\SB1_1_2/i0_3 ) );
  INV_X2 \SB1_3_19/INV_5  ( .A(\RI1[3][77] ), .ZN(\SB1_3_19/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_160  ( .A(\RI5[2][160] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[160] ) );
  BUF_X2 \SB2_1_24/BUF_2  ( .A(\RI3[1][44] ), .Z(\SB2_1_24/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_72  ( .A(\RI5[1][72] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[72] ) );
  INV_X2 \SB1_2_24/INV_5  ( .A(\RI1[2][47] ), .ZN(\SB1_2_24/i0_3 ) );
  BUF_X2 \SB4_17/BUF_2  ( .A(\RI3[4][86] ), .Z(\SB4_17/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_36  ( .A(\RI5[1][36] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[36] ) );
  INV_X2 \SB1_3_27/INV_5  ( .A(\RI1[3][29] ), .ZN(\SB1_3_27/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_90  ( .A(\RI5[1][90] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[90] ) );
  INV_X2 \SB1_2_30/INV_5  ( .A(\RI1[2][11] ), .ZN(\SB1_2_30/i0_3 ) );
  BUF_X2 \SB4_13/BUF_3  ( .A(\RI3[4][111] ), .Z(\SB4_13/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_180  ( .A(\RI5[1][180] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[180] ) );
  BUF_X2 \SB2_0_31/BUF_4  ( .A(\RI3[0][4] ), .Z(\SB2_0_31/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_66  ( .A(\RI5[0][66] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[66] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_10  ( .A(\RI5[1][10] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[10] ) );
  INV_X2 \SB1_1_20/INV_5  ( .A(\RI1[1][71] ), .ZN(\SB1_1_20/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_100  ( .A(\RI5[1][100] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[100] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_186  ( .A(\RI5[0][186] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[186] ) );
  BUF_X2 \SB2_3_9/BUF_2  ( .A(\RI3[3][134] ), .Z(\SB2_3_9/i0_0 ) );
  INV_X2 \SB1_1_13/INV_5  ( .A(\RI1[1][113] ), .ZN(\SB1_1_13/i0_3 ) );
  BUF_X2 \SB4_22/BUF_3  ( .A(\RI3[4][57] ), .Z(\SB4_22/i0[10] ) );
  BUF_X2 \SB2_3_27/BUF_3  ( .A(\RI3[3][27] ), .Z(\SB2_3_27/i0[10] ) );
  INV_X1 \SB3_31/INV_5  ( .A(\RI1[4][5] ), .ZN(\SB3_31/i0_3 ) );
  INV_X1 \SB3_6/INV_5  ( .A(\RI1[4][155] ), .ZN(\SB3_6/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_6  ( .A(\RI5[1][6] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[6] ) );
  INV_X1 \SB1_2_14/INV_4  ( .A(\RI1[2][106] ), .ZN(\SB1_2_14/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_156  ( .A(\RI5[2][156] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[156] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_66  ( .A(\RI5[1][66] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[66] ) );
  BUF_X2 \SB4_18/BUF_4  ( .A(\RI3[4][82] ), .Z(\SB4_18/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_114  ( .A(\RI5[0][114] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[114] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_138  ( .A(\RI5[2][138] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[138] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_108  ( .A(\RI5[0][108] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[108] ) );
  INV_X2 \SB1_2_16/INV_5  ( .A(\RI1[2][95] ), .ZN(\SB1_2_16/i0_3 ) );
  INV_X2 \SB1_2_27/INV_5  ( .A(\RI1[2][29] ), .ZN(\SB1_2_27/i0_3 ) );
  INV_X2 \SB1_2_21/INV_5  ( .A(\RI1[2][65] ), .ZN(\SB1_2_21/i0_3 ) );
  BUF_X2 \SB2_3_12/BUF_3  ( .A(\RI3[3][117] ), .Z(\SB2_3_12/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_24  ( .A(\RI5[0][24] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[24] ) );
  BUF_X2 \SB2_3_20/BUF_2  ( .A(\RI3[3][68] ), .Z(\SB2_3_20/i0_0 ) );
  INV_X1 \SB1_2_13/INV_2  ( .A(\RI1[2][110] ), .ZN(\SB1_2_13/i0_0 ) );
  INV_X1 \SB3_8/INV_5  ( .A(\RI1[4][143] ), .ZN(\SB3_8/i0_3 ) );
  INV_X1 \SB3_4/INV_5  ( .A(\RI1[4][167] ), .ZN(\SB3_4/i0_3 ) );
  INV_X1 \SB3_15/INV_5  ( .A(\RI1[4][101] ), .ZN(\SB3_15/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_0  ( .A(\RI5[1][0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[0] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_122  ( .A(\RI5[1][122] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[122] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_180  ( .A(\RI5[0][180] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[180] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_162  ( .A(\RI5[1][162] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[162] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_60  ( .A(\RI5[1][60] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[60] ) );
  BUF_X2 \SB2_3_11/BUF_3  ( .A(\RI3[3][123] ), .Z(\SB2_3_11/i0[10] ) );
  INV_X1 \SB3_5/INV_4  ( .A(\RI1[4][160] ), .ZN(\SB3_5/i0_4 ) );
  INV_X1 \SB1_3_8/INV_4  ( .A(\RI1[3][142] ), .ZN(\SB1_3_8/i0_4 ) );
  INV_X1 \SB1_3_16/INV_4  ( .A(\RI1[3][94] ), .ZN(\SB1_3_16/i0_4 ) );
  INV_X1 \SB1_2_7/INV_4  ( .A(\RI1[2][148] ), .ZN(\SB1_2_7/i0_4 ) );
  BUF_X2 \SB4_5/BUF_3  ( .A(\RI3[4][159] ), .Z(\SB4_5/i0[10] ) );
  INV_X1 \SB1_3_26/INV_4  ( .A(\RI1[3][34] ), .ZN(\SB1_3_26/i0_4 ) );
  INV_X1 \SB3_16/INV_5  ( .A(\RI1[4][95] ), .ZN(\SB3_16/i0_3 ) );
  INV_X1 \SB1_3_25/INV_2  ( .A(\RI1[3][38] ), .ZN(\SB1_3_25/i0_0 ) );
  INV_X1 \SB3_7/INV_5  ( .A(\RI1[4][149] ), .ZN(\SB3_7/i0_3 ) );
  INV_X1 \SB3_25/INV_5  ( .A(\RI1[4][41] ), .ZN(\SB3_25/i0_3 ) );
  BUF_X2 \SB2_2_21/BUF_3  ( .A(\RI3[2][63] ), .Z(\SB2_2_21/i0[10] ) );
  BUF_X1 \SB1_3_23/BUF_5  ( .A(\RI1[3][53] ), .Z(\SB1_3_23/i1_5 ) );
  BUF_X1 \SB1_1_0/BUF_5  ( .A(\RI1[1][191] ), .Z(\SB1_1_0/i1_5 ) );
  INV_X1 \SB1_2_5/INV_2  ( .A(\RI1[2][158] ), .ZN(\SB1_2_5/i0_0 ) );
  INV_X1 \SB2_3_4/INV_2  ( .A(\RI3[3][164] ), .ZN(\SB2_3_4/i1[9] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_45_0  ( .A(Key[168]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[45] ) );
  INV_X1 \SB2_2_2/INV_2  ( .A(\RI3[2][176] ), .ZN(\SB2_2_2/i1[9] ) );
  INV_X1 \SB1_2_20/INV_0  ( .A(\RI1[2][66] ), .ZN(\SB1_2_20/i0[9] ) );
  INV_X1 \SB1_2_26/INV_4  ( .A(\RI1[2][34] ), .ZN(\SB1_2_26/i0_4 ) );
  INV_X1 \SB1_2_3/INV_0  ( .A(\RI1[2][168] ), .ZN(\SB1_2_3/i0[9] ) );
  INV_X1 \SB1_2_12/INV_1  ( .A(\RI1[2][115] ), .ZN(\SB1_2_12/i0[6] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_27_0  ( .A(Key[19]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[27] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_189_0  ( .A(Key[85]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[189] ) );
  INV_X1 \SB2_0_21/INV_2  ( .A(\RI3[0][62] ), .ZN(\SB2_0_21/i1[9] ) );
  INV_X1 \SB1_0_13/INV_0  ( .A(n84), .ZN(\SB1_0_13/i0[9] ) );
  INV_X1 \SB2_2_28/INV_2  ( .A(\RI3[2][20] ), .ZN(\SB2_2_28/i1[9] ) );
  INV_X1 \SB2_2_22/INV_2  ( .A(\RI3[2][56] ), .ZN(\SB2_2_22/i1[9] ) );
  INV_X1 \SB2_2_6/INV_2  ( .A(\RI3[2][152] ), .ZN(\SB2_2_6/i1[9] ) );
  BUF_X1 \SB1_1_24/BUF_5  ( .A(\RI1[1][47] ), .Z(\SB1_1_24/i1_5 ) );
  BUF_X1 \SB1_3_1/BUF_5  ( .A(\RI1[3][185] ), .Z(\SB1_3_1/i1_5 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_84  ( .A(\RI5[0][84] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[84] ) );
  BUF_X2 \SB2_3_21/BUF_3  ( .A(\RI3[3][63] ), .Z(\SB2_3_21/i0[10] ) );
  BUF_X2 \SB4_24/BUF_3  ( .A(\RI3[4][45] ), .Z(\SB4_24/i0[10] ) );
  INV_X1 \SB1_1_3/INV_3  ( .A(\RI1[1][171] ), .ZN(\SB1_1_3/i0[10] ) );
  BUF_X2 \SB2_1_20/BUF_2  ( .A(\RI3[1][68] ), .Z(\SB2_1_20/i0_0 ) );
  INV_X1 \SB3_17/INV_5  ( .A(\RI1[4][89] ), .ZN(\SB3_17/i0_3 ) );
  INV_X1 \SB3_24/INV_5  ( .A(\RI1[4][47] ), .ZN(\SB3_24/i0_3 ) );
  INV_X1 \SB1_2_6/INV_3  ( .A(\RI1[2][153] ), .ZN(\SB1_2_6/i0[10] ) );
  INV_X1 \SB3_20/INV_5  ( .A(\RI1[4][71] ), .ZN(\SB3_20/i0_3 ) );
  INV_X1 \SB2_3_9/INV_2  ( .A(\RI3[3][134] ), .ZN(\SB2_3_9/i1[9] ) );
  INV_X1 \SB2_0_8/INV_2  ( .A(\RI3[0][140] ), .ZN(\SB2_0_8/i1[9] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_89_0  ( .A(Key[73]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[89] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_129_0  ( .A(Key[25]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[129] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_105_0  ( .A(Key[1]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[105] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_62_0  ( .A(Key[6]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[62] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_74_0  ( .A(Key[18]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[74] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_0/BUF_158_0  ( .A(Key[151]), .Z(
        \MC_ARK_ARC_1_0/buf_keyinput[158] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_0/BUF_187_0  ( .A(Key[162]), .Z(
        \MC_ARK_ARC_1_0/buf_keyinput[187] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_137_0  ( .A(Key[121]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[137] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_142_0  ( .A(Key[30]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[142] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_154_0  ( .A(Key[42]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[154] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_173_0  ( .A(Key[157]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[173] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_166_0  ( .A(Key[54]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[166] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_172_0  ( .A(Key[145]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[172] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_112_0  ( .A(Key[109]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[112] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_118_0  ( .A(Key[55]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[118] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_76_0  ( .A(Key[49]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[76] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_69_0  ( .A(Key[144]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[69] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_87_0  ( .A(Key[174]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[87] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_33_0  ( .A(Key[84]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[33] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_184_0  ( .A(Key[37]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[184] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_8_0  ( .A(Key[48]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[8] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_183_0  ( .A(Key[175]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[183] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_176_0  ( .A(Key[24]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[176] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_0/BUF_80_0  ( .A(Key[181]), .Z(
        \MC_ARK_ARC_1_0/buf_keyinput[80] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_152_0  ( .A(Key[0]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[152] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_170_0  ( .A(Key[114]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[170] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_123_0  ( .A(Key[115]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[123] ) );
  CLKBUF_X1 \SB1_0_17/BUF_0  ( .A(n108), .Z(\SB1_0_17/i3[0] ) );
  CLKBUF_X1 \SB1_0_23/BUF_4  ( .A(n140), .Z(\SB1_0_23/i0[7] ) );
  CLKBUF_X1 \SB1_0_20/BUF_0  ( .A(n126), .Z(\SB1_0_20/i3[0] ) );
  CLKBUF_X1 \SB1_0_25/BUF_4  ( .A(n152), .Z(\SB1_0_25/i0[7] ) );
  BUF_X1 \SB1_0_21/BUF_3  ( .A(n129), .Z(\SB1_0_21/i0[8] ) );
  CLKBUF_X1 \SB1_0_8/BUF_4  ( .A(n50), .Z(\SB1_0_8/i0[7] ) );
  CLKBUF_X1 \SB1_0_28/BUF_0  ( .A(n174), .Z(\SB1_0_28/i3[0] ) );
  CLKBUF_X1 \SB1_0_26/BUF_4  ( .A(n158), .Z(\SB1_0_26/i0[7] ) );
  CLKBUF_X1 \SB1_0_26/BUF_0  ( .A(n162), .Z(\SB1_0_26/i3[0] ) );
  CLKBUF_X1 \SB1_0_27/BUF_0  ( .A(n168), .Z(\SB1_0_27/i3[0] ) );
  CLKBUF_X1 \SB1_0_14/BUF_4  ( .A(n86), .Z(\SB1_0_14/i0[7] ) );
  CLKBUF_X1 \SB1_0_31/BUF_4  ( .A(n188), .Z(\SB1_0_31/i0[7] ) );
  CLKBUF_X1 \SB1_0_19/BUF_0  ( .A(n120), .Z(\SB1_0_19/i3[0] ) );
  CLKBUF_X1 \SB1_0_30/BUF_1  ( .A(n185), .Z(\SB1_0_30/i1_7 ) );
  CLKBUF_X1 \SB1_0_5/BUF_4  ( .A(n32), .Z(\SB1_0_5/i0[7] ) );
  CLKBUF_X1 \SB1_0_2/BUF_4  ( .A(n14), .Z(\SB1_0_2/i0[7] ) );
  CLKBUF_X1 \SB1_0_0/BUF_0  ( .A(n6), .Z(\SB1_0_0/i3[0] ) );
  BUF_X1 \SB1_0_20/BUF_2  ( .A(n124), .Z(\SB1_0_20/i1[9] ) );
  CLKBUF_X1 \SB1_0_30/BUF_4  ( .A(n182), .Z(\SB1_0_30/i0[7] ) );
  CLKBUF_X1 \SB1_0_10/BUF_4  ( .A(n62), .Z(\SB1_0_10/i0[7] ) );
  CLKBUF_X1 \SB1_0_29/BUF_4  ( .A(n176), .Z(\SB1_0_29/i0[7] ) );
  CLKBUF_X1 \SB1_0_17/BUF_4  ( .A(n104), .Z(\SB1_0_17/i0[7] ) );
  CLKBUF_X1 \SB1_0_22/BUF_4  ( .A(n134), .Z(\SB1_0_22/i0[7] ) );
  CLKBUF_X1 \SB1_0_14/BUF_0  ( .A(n90), .Z(\SB1_0_14/i3[0] ) );
  BUF_X1 \SB1_0_4/BUF_3  ( .A(n27), .Z(\SB1_0_4/i0[8] ) );
  CLKBUF_X1 \SB1_0_4/BUF_4  ( .A(n26), .Z(\SB1_0_4/i0[7] ) );
  CLKBUF_X1 \SB1_0_16/BUF_0  ( .A(n102), .Z(\SB1_0_16/i3[0] ) );
  BUF_X1 \SB1_0_16/BUF_2  ( .A(n100), .Z(\SB1_0_16/i1[9] ) );
  CLKBUF_X1 \SB1_0_8/BUF_0  ( .A(n54), .Z(\SB1_0_8/i3[0] ) );
  CLKBUF_X1 \SB1_0_12/BUF_0  ( .A(n78), .Z(\SB1_0_12/i3[0] ) );
  CLKBUF_X1 \SB1_0_12/BUF_4  ( .A(n74), .Z(\SB1_0_12/i0[7] ) );
  CLKBUF_X1 \SB1_0_7/BUF_0  ( .A(n48), .Z(\SB1_0_7/i3[0] ) );
  CLKBUF_X1 \SB1_0_9/BUF_0  ( .A(n60), .Z(\SB1_0_9/i3[0] ) );
  CLKBUF_X1 \SB1_0_2/BUF_0  ( .A(n18), .Z(\SB1_0_2/i3[0] ) );
  CLKBUF_X1 \SB1_0_1/BUF_4  ( .A(n8), .Z(\SB1_0_1/i0[7] ) );
  CLKBUF_X1 \SB1_0_6/BUF_4  ( .A(n38), .Z(\SB1_0_6/i0[7] ) );
  CLKBUF_X1 \SB1_0_3/BUF_0  ( .A(n24), .Z(\SB1_0_3/i3[0] ) );
  CLKBUF_X1 \SB1_0_31/BUF_0  ( .A(n192), .Z(\SB1_0_31/i3[0] ) );
  BUF_X1 \SB1_0_31/BUF_3  ( .A(n189), .Z(\SB1_0_31/i0[8] ) );
  CLKBUF_X1 \SB1_0_23/BUF_0  ( .A(n144), .Z(\SB1_0_23/i3[0] ) );
  CLKBUF_X1 \SB1_0_27/BUF_4  ( .A(n164), .Z(\SB1_0_27/i0[7] ) );
  CLKBUF_X1 \SB1_0_19/BUF_4  ( .A(n116), .Z(\SB1_0_19/i0[7] ) );
  CLKBUF_X1 \SB1_0_16/BUF_1  ( .A(n101), .Z(\SB1_0_16/i1_7 ) );
  CLKBUF_X1 \SB1_0_9/BUF_4  ( .A(n56), .Z(\SB1_0_9/i0[7] ) );
  BUF_X1 \SB1_0_26/BUF_3  ( .A(n159), .Z(\SB1_0_26/i0[8] ) );
  CLKBUF_X1 \SB1_0_0/BUF_4  ( .A(n2), .Z(\SB1_0_0/i0[7] ) );
  CLKBUF_X1 \SB1_0_22/BUF_0  ( .A(n138), .Z(\SB1_0_22/i3[0] ) );
  CLKBUF_X1 \SB1_0_15/BUF_1  ( .A(n95), .Z(\SB1_0_15/i1_7 ) );
  CLKBUF_X1 \SB1_0_4/BUF_0  ( .A(n30), .Z(\SB1_0_4/i3[0] ) );
  BUF_X1 \SB1_0_26/BUF_2  ( .A(n160), .Z(\SB1_0_26/i1[9] ) );
  CLKBUF_X1 \SB1_0_15/BUF_0  ( .A(n96), .Z(\SB1_0_15/i3[0] ) );
  CLKBUF_X1 \SB1_0_24/BUF_1  ( .A(n149), .Z(\SB1_0_24/i1_7 ) );
  CLKBUF_X1 \SB1_0_24/BUF_0  ( .A(n150), .Z(\SB1_0_24/i3[0] ) );
  CLKBUF_X1 \SB1_0_21/BUF_4  ( .A(n128), .Z(\SB1_0_21/i0[7] ) );
  CLKBUF_X1 \SB1_0_20/BUF_4  ( .A(n122), .Z(\SB1_0_20/i0[7] ) );
  CLKBUF_X1 \SB1_0_11/BUF_0  ( .A(n72), .Z(\SB1_0_11/i3[0] ) );
  CLKBUF_X1 \SB1_0_13/BUF_4  ( .A(n80), .Z(\SB1_0_13/i0[7] ) );
  CLKBUF_X1 \SB1_0_26/BUF_1  ( .A(n161), .Z(\SB1_0_26/i1_7 ) );
  CLKBUF_X1 \SB1_0_7/BUF_4  ( .A(n44), .Z(\SB1_0_7/i0[7] ) );
  CLKBUF_X1 \SB1_0_15/BUF_4  ( .A(n92), .Z(\SB1_0_15/i0[7] ) );
  CLKBUF_X1 \SB1_0_10/BUF_0  ( .A(n66), .Z(\SB1_0_10/i3[0] ) );
  INV_X1 \SB1_0_14/INV_2  ( .A(n88), .ZN(\SB1_0_14/i0_0 ) );
  CLKBUF_X1 \SB1_0_25/BUF_0  ( .A(n156), .Z(\SB1_0_25/i3[0] ) );
  CLKBUF_X1 \SB1_0_29/BUF_0  ( .A(n180), .Z(\SB1_0_29/i3[0] ) );
  CLKBUF_X1 \SB1_0_30/BUF_0  ( .A(n186), .Z(\SB1_0_30/i3[0] ) );
  BUF_X1 \SB1_0_15/BUF_2  ( .A(n94), .Z(\SB1_0_15/i1[9] ) );
  CLKBUF_X1 \SB1_0_13/BUF_0  ( .A(n84), .Z(\SB1_0_13/i3[0] ) );
  CLKBUF_X1 \SB1_0_3/BUF_4  ( .A(n20), .Z(\SB1_0_3/i0[7] ) );
  CLKBUF_X1 \SB1_0_24/BUF_4  ( .A(n146), .Z(\SB1_0_24/i0[7] ) );
  CLKBUF_X1 \SB1_0_28/BUF_4  ( .A(n170), .Z(\SB1_0_28/i0[7] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_125_0  ( .A(Key[21]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[125] ) );
  CLKBUF_X1 \SB1_1_12/BUF_1  ( .A(\RI1[1][115] ), .Z(\SB1_1_12/i1_7 ) );
  CLKBUF_X1 \SB1_1_2/BUF_4  ( .A(\RI1[1][178] ), .Z(\SB1_1_2/i0[7] ) );
  CLKBUF_X1 \SB1_1_27/BUF_0  ( .A(\RI1[1][24] ), .Z(\SB1_1_27/i3[0] ) );
  CLKBUF_X1 \SB1_1_12/BUF_0  ( .A(\RI1[1][114] ), .Z(\SB1_1_12/i3[0] ) );
  CLKBUF_X1 \SB1_1_23/BUF_0  ( .A(\RI1[1][48] ), .Z(\SB1_1_23/i3[0] ) );
  CLKBUF_X1 \SB1_1_6/BUF_0  ( .A(\RI1[1][150] ), .Z(\SB1_1_6/i3[0] ) );
  INV_X1 \SB1_1_31/INV_4  ( .A(\RI1[1][4] ), .ZN(\SB1_1_31/i0_4 ) );
  INV_X1 \SB1_1_27/INV_0  ( .A(\RI1[1][24] ), .ZN(\SB1_1_27/i0[9] ) );
  INV_X1 \SB1_1_0/INV_0  ( .A(\RI1[1][186] ), .ZN(\SB1_1_0/i0[9] ) );
  CLKBUF_X1 \SB1_1_18/BUF_0  ( .A(\RI1[1][78] ), .Z(\SB1_1_18/i3[0] ) );
  CLKBUF_X1 \SB1_1_14/BUF_0  ( .A(\RI1[1][102] ), .Z(\SB1_1_14/i3[0] ) );
  CLKBUF_X1 \SB1_1_13/BUF_0  ( .A(\RI1[1][108] ), .Z(\SB1_1_13/i3[0] ) );
  CLKBUF_X1 \SB1_1_5/BUF_4  ( .A(\RI1[1][160] ), .Z(\SB1_1_5/i0[7] ) );
  CLKBUF_X1 \SB1_1_3/BUF_0  ( .A(\RI1[1][168] ), .Z(\SB1_1_3/i3[0] ) );
  CLKBUF_X1 \SB1_1_1/BUF_4  ( .A(\RI1[1][184] ), .Z(\SB1_1_1/i0[7] ) );
  CLKBUF_X1 \SB1_1_22/BUF_4  ( .A(\RI1[1][58] ), .Z(\SB1_1_22/i0[7] ) );
  CLKBUF_X1 \SB1_1_5/BUF_0  ( .A(\RI1[1][156] ), .Z(\SB1_1_5/i3[0] ) );
  CLKBUF_X1 \SB1_1_0/BUF_4  ( .A(\RI1[1][190] ), .Z(\SB1_1_0/i0[7] ) );
  BUF_X1 \SB1_1_0/BUF_1  ( .A(\RI1[1][187] ), .Z(\SB1_1_0/i1_7 ) );
  CLKBUF_X1 \SB1_1_9/BUF_4  ( .A(\RI1[1][136] ), .Z(\SB1_1_9/i0[7] ) );
  CLKBUF_X1 \SB1_1_5/BUF_1  ( .A(\RI1[1][157] ), .Z(\SB1_1_5/i1_7 ) );
  CLKBUF_X1 \SB1_1_28/BUF_0  ( .A(\RI1[1][18] ), .Z(\SB1_1_28/i3[0] ) );
  CLKBUF_X1 \SB1_1_0/BUF_0  ( .A(\RI1[1][186] ), .Z(\SB1_1_0/i3[0] ) );
  CLKBUF_X1 \SB1_1_4/BUF_0  ( .A(\RI1[1][162] ), .Z(\SB1_1_4/i3[0] ) );
  CLKBUF_X1 \SB1_1_8/BUF_4  ( .A(\RI1[1][142] ), .Z(\SB1_1_8/i0[7] ) );
  BUF_X1 \SB1_1_20/BUF_3  ( .A(\RI1[1][69] ), .Z(\SB1_1_20/i0[8] ) );
  CLKBUF_X1 \SB1_1_10/BUF_4  ( .A(\RI1[1][130] ), .Z(\SB1_1_10/i0[7] ) );
  CLKBUF_X1 \SB1_1_20/BUF_0  ( .A(\RI1[1][66] ), .Z(\SB1_1_20/i3[0] ) );
  CLKBUF_X1 \SB1_1_20/BUF_4  ( .A(\RI1[1][70] ), .Z(\SB1_1_20/i0[7] ) );
  CLKBUF_X1 \SB1_1_6/BUF_4  ( .A(\RI1[1][154] ), .Z(\SB1_1_6/i0[7] ) );
  CLKBUF_X1 \SB1_1_8/BUF_0  ( .A(\RI1[1][138] ), .Z(\SB1_1_8/i3[0] ) );
  CLKBUF_X1 \SB1_1_15/BUF_4  ( .A(\RI1[1][100] ), .Z(\SB1_1_15/i0[7] ) );
  CLKBUF_X1 \SB1_1_2/BUF_0  ( .A(\RI1[1][174] ), .Z(\SB1_1_2/i3[0] ) );
  CLKBUF_X1 \SB1_1_17/BUF_1  ( .A(\RI1[1][85] ), .Z(\SB1_1_17/i1_7 ) );
  CLKBUF_X1 \SB1_1_17/BUF_0  ( .A(\RI1[1][84] ), .Z(\SB1_1_17/i3[0] ) );
  INV_X1 \SB1_1_26/INV_4  ( .A(\RI1[1][34] ), .ZN(\SB1_1_26/i0_4 ) );
  CLKBUF_X1 \SB1_1_1/BUF_0  ( .A(\RI1[1][180] ), .Z(\SB1_1_1/i3[0] ) );
  CLKBUF_X1 \SB1_1_18/BUF_4  ( .A(\RI1[1][82] ), .Z(\SB1_1_18/i0[7] ) );
  CLKBUF_X1 \SB1_1_22/BUF_0  ( .A(\RI1[1][54] ), .Z(\SB1_1_22/i3[0] ) );
  CLKBUF_X1 \SB1_1_7/BUF_0  ( .A(\RI1[1][144] ), .Z(\SB1_1_7/i3[0] ) );
  CLKBUF_X1 \SB1_1_15/BUF_0  ( .A(\RI1[1][96] ), .Z(\SB1_1_15/i3[0] ) );
  CLKBUF_X1 \SB1_1_30/BUF_0  ( .A(\RI1[1][6] ), .Z(\SB1_1_30/i3[0] ) );
  BUF_X1 \SB1_1_22/BUF_1  ( .A(\RI1[1][55] ), .Z(\SB1_1_22/i1_7 ) );
  CLKBUF_X1 \SB1_1_16/BUF_0  ( .A(\RI1[1][90] ), .Z(\SB1_1_16/i3[0] ) );
  CLKBUF_X1 \SB1_1_3/BUF_4  ( .A(\RI1[1][172] ), .Z(\SB1_1_3/i0[7] ) );
  CLKBUF_X1 \SB1_1_25/BUF_4  ( .A(\RI1[1][40] ), .Z(\SB1_1_25/i0[7] ) );
  CLKBUF_X1 \SB1_1_19/BUF_0  ( .A(\RI1[1][72] ), .Z(\SB1_1_19/i3[0] ) );
  INV_X1 \SB1_1_24/INV_0  ( .A(\RI1[1][42] ), .ZN(\SB1_1_24/i0[9] ) );
  CLKBUF_X1 \SB1_1_24/BUF_1  ( .A(\RI1[1][43] ), .Z(\SB1_1_24/i1_7 ) );
  CLKBUF_X1 \SB1_1_14/BUF_4  ( .A(\RI1[1][106] ), .Z(\SB1_1_14/i0[7] ) );
  INV_X1 \SB1_1_14/INV_2  ( .A(\RI1[1][104] ), .ZN(\SB1_1_14/i0_0 ) );
  INV_X1 \SB1_1_21/INV_4  ( .A(\RI1[1][64] ), .ZN(\SB1_1_21/i0_4 ) );
  CLKBUF_X1 \SB1_1_26/BUF_0  ( .A(\RI1[1][30] ), .Z(\SB1_1_26/i3[0] ) );
  CLKBUF_X1 \SB1_1_31/BUF_4  ( .A(\RI1[1][4] ), .Z(\SB1_1_31/i0[7] ) );
  CLKBUF_X1 \SB1_1_11/BUF_0  ( .A(\RI1[1][120] ), .Z(\SB1_1_11/i3[0] ) );
  CLKBUF_X1 \SB1_1_31/BUF_0  ( .A(\RI1[1][0] ), .Z(\SB1_1_31/i3[0] ) );
  BUF_X1 \SB1_1_3/BUF_1  ( .A(\RI1[1][169] ), .Z(\SB1_1_3/i1_7 ) );
  CLKBUF_X1 \SB1_1_29/BUF_4  ( .A(\RI1[1][16] ), .Z(\SB1_1_29/i0[7] ) );
  CLKBUF_X1 \SB1_1_25/BUF_0  ( .A(\RI1[1][36] ), .Z(\SB1_1_25/i3[0] ) );
  CLKBUF_X1 \SB1_1_26/BUF_4  ( .A(\RI1[1][34] ), .Z(\SB1_1_26/i0[7] ) );
  CLKBUF_X1 \SB1_1_21/BUF_4  ( .A(\RI1[1][64] ), .Z(\SB1_1_21/i0[7] ) );
  CLKBUF_X1 \SB1_1_1/BUF_1  ( .A(\RI1[1][181] ), .Z(\SB1_1_1/i1_7 ) );
  CLKBUF_X1 \SB1_1_9/BUF_0  ( .A(\RI1[1][132] ), .Z(\SB1_1_9/i3[0] ) );
  CLKBUF_X1 \SB1_1_14/BUF_1  ( .A(\RI1[1][103] ), .Z(\SB1_1_14/i1_7 ) );
  CLKBUF_X1 \SB1_1_12/BUF_4  ( .A(\RI1[1][118] ), .Z(\SB1_1_12/i0[7] ) );
  CLKBUF_X1 \SB1_1_21/BUF_0  ( .A(\RI1[1][60] ), .Z(\SB1_1_21/i3[0] ) );
  CLKBUF_X1 \SB1_1_30/BUF_4  ( .A(\RI1[1][10] ), .Z(\SB1_1_30/i0[7] ) );
  CLKBUF_X1 \SB1_1_7/BUF_4  ( .A(\RI1[1][148] ), .Z(\SB1_1_7/i0[7] ) );
  CLKBUF_X1 \SB1_1_10/BUF_0  ( .A(\RI1[1][126] ), .Z(\SB1_1_10/i3[0] ) );
  BUF_X1 \SB1_1_10/BUF_1  ( .A(\RI1[1][127] ), .Z(\SB1_1_10/i1_7 ) );
  INV_X1 \SB1_1_29/INV_0  ( .A(\RI1[1][12] ), .ZN(\SB1_1_29/i0[9] ) );
  INV_X1 \SB1_1_19/INV_0  ( .A(\RI1[1][72] ), .ZN(\SB1_1_19/i0[9] ) );
  CLKBUF_X1 \SB1_1_13/BUF_4  ( .A(\RI1[1][112] ), .Z(\SB1_1_13/i0[7] ) );
  CLKBUF_X1 \SB1_2_22/BUF_0  ( .A(\RI1[2][54] ), .Z(\SB1_2_22/i3[0] ) );
  CLKBUF_X1 \SB1_2_7/BUF_0  ( .A(\RI1[2][144] ), .Z(\SB1_2_7/i3[0] ) );
  CLKBUF_X1 \SB1_2_6/BUF_0  ( .A(\RI1[2][150] ), .Z(\SB1_2_6/i3[0] ) );
  CLKBUF_X1 \SB1_2_4/BUF_4  ( .A(\RI1[2][166] ), .Z(\SB1_2_4/i0[7] ) );
  CLKBUF_X1 \SB1_2_5/BUF_0  ( .A(\RI1[2][156] ), .Z(\SB1_2_5/i3[0] ) );
  INV_X1 \SB1_2_1/INV_4  ( .A(\RI1[2][184] ), .ZN(\SB1_2_1/i0_4 ) );
  CLKBUF_X1 \SB1_2_21/BUF_0  ( .A(\RI1[2][60] ), .Z(\SB1_2_21/i3[0] ) );
  CLKBUF_X1 \SB1_2_25/BUF_0  ( .A(\RI1[2][36] ), .Z(\SB1_2_25/i3[0] ) );
  CLKBUF_X1 \SB1_2_26/BUF_4  ( .A(\RI1[2][34] ), .Z(\SB1_2_26/i0[7] ) );
  CLKBUF_X1 \SB1_2_12/BUF_0  ( .A(\RI1[2][114] ), .Z(\SB1_2_12/i3[0] ) );
  CLKBUF_X1 \SB1_2_16/BUF_4  ( .A(\RI1[2][94] ), .Z(\SB1_2_16/i0[7] ) );
  INV_X1 \SB1_2_15/INV_4  ( .A(\RI1[2][100] ), .ZN(\SB1_2_15/i0_4 ) );
  INV_X1 \SB1_2_29/INV_3  ( .A(\RI1[2][15] ), .ZN(\SB1_2_29/i0[10] ) );
  CLKBUF_X1 \SB1_2_18/BUF_4  ( .A(\RI1[2][82] ), .Z(\SB1_2_18/i0[7] ) );
  INV_X1 \SB1_2_13/INV_4  ( .A(\RI1[2][112] ), .ZN(\SB1_2_13/i0_4 ) );
  CLKBUF_X1 \SB1_2_29/BUF_0  ( .A(\RI1[2][12] ), .Z(\SB1_2_29/i3[0] ) );
  CLKBUF_X1 \SB1_2_26/BUF_0  ( .A(\RI1[2][30] ), .Z(\SB1_2_26/i3[0] ) );
  CLKBUF_X1 \SB1_2_0/BUF_0  ( .A(\RI1[2][186] ), .Z(\SB1_2_0/i3[0] ) );
  CLKBUF_X1 \SB1_2_27/BUF_0  ( .A(\RI1[2][24] ), .Z(\SB1_2_27/i3[0] ) );
  CLKBUF_X1 \SB1_2_9/BUF_4  ( .A(\RI1[2][136] ), .Z(\SB1_2_9/i0[7] ) );
  CLKBUF_X1 \SB1_2_31/BUF_0  ( .A(\RI1[2][0] ), .Z(\SB1_2_31/i3[0] ) );
  CLKBUF_X1 \SB1_2_9/BUF_0  ( .A(\RI1[2][132] ), .Z(\SB1_2_9/i3[0] ) );
  INV_X1 \SB1_2_25/INV_4  ( .A(\RI1[2][40] ), .ZN(\SB1_2_25/i0_4 ) );
  CLKBUF_X1 \SB1_2_13/BUF_0  ( .A(\RI1[2][108] ), .Z(\SB1_2_13/i3[0] ) );
  CLKBUF_X1 \SB1_2_31/BUF_4  ( .A(\RI1[2][4] ), .Z(\SB1_2_31/i0[7] ) );
  CLKBUF_X1 \SB1_2_26/BUF_1  ( .A(\RI1[2][31] ), .Z(\SB1_2_26/i1_7 ) );
  CLKBUF_X1 \SB1_2_2/BUF_0  ( .A(\RI1[2][174] ), .Z(\SB1_2_2/i3[0] ) );
  CLKBUF_X1 \SB1_2_28/BUF_0  ( .A(\RI1[2][18] ), .Z(\SB1_2_28/i3[0] ) );
  CLKBUF_X1 \SB1_2_15/BUF_0  ( .A(\RI1[2][96] ), .Z(\SB1_2_15/i3[0] ) );
  CLKBUF_X1 \SB1_2_8/BUF_4  ( .A(\RI1[2][142] ), .Z(\SB1_2_8/i0[7] ) );
  CLKBUF_X1 \SB1_2_1/BUF_0  ( .A(\RI1[2][180] ), .Z(\SB1_2_1/i3[0] ) );
  INV_X1 \SB1_2_10/INV_4  ( .A(\RI1[2][130] ), .ZN(\SB1_2_10/i0_4 ) );
  CLKBUF_X1 \SB1_2_18/BUF_0  ( .A(\RI1[2][78] ), .Z(\SB1_2_18/i3[0] ) );
  CLKBUF_X1 \SB1_2_4/BUF_0  ( .A(\RI1[2][162] ), .Z(\SB1_2_4/i3[0] ) );
  CLKBUF_X1 \SB1_2_23/BUF_0  ( .A(\RI1[2][48] ), .Z(\SB1_2_23/i3[0] ) );
  CLKBUF_X1 \SB1_2_8/BUF_0  ( .A(\RI1[2][138] ), .Z(\SB1_2_8/i3[0] ) );
  CLKBUF_X1 \SB1_2_14/BUF_4  ( .A(\RI1[2][106] ), .Z(\SB1_2_14/i0[7] ) );
  CLKBUF_X1 \SB1_2_21/BUF_4  ( .A(\RI1[2][64] ), .Z(\SB1_2_21/i0[7] ) );
  CLKBUF_X1 \SB1_2_16/BUF_0  ( .A(\RI1[2][90] ), .Z(\SB1_2_16/i3[0] ) );
  CLKBUF_X1 \SB1_2_30/BUF_0  ( .A(\RI1[2][6] ), .Z(\SB1_2_30/i3[0] ) );
  CLKBUF_X1 \SB1_2_24/BUF_0  ( .A(\RI1[2][42] ), .Z(\SB1_2_24/i3[0] ) );
  INV_X1 \SB1_2_17/INV_0  ( .A(\RI1[2][84] ), .ZN(\SB1_2_17/i0[9] ) );
  CLKBUF_X1 \SB1_2_3/BUF_0  ( .A(\RI1[2][168] ), .Z(\SB1_2_3/i3[0] ) );
  CLKBUF_X1 \SB1_2_19/BUF_0  ( .A(\RI1[2][72] ), .Z(\SB1_2_19/i3[0] ) );
  CLKBUF_X1 \SB1_2_10/BUF_0  ( .A(\RI1[2][126] ), .Z(\SB1_2_10/i3[0] ) );
  INV_X1 \SB1_2_17/INV_4  ( .A(\RI1[2][88] ), .ZN(\SB1_2_17/i0_4 ) );
  CLKBUF_X1 \SB1_2_11/BUF_0  ( .A(\RI1[2][120] ), .Z(\SB1_2_11/i3[0] ) );
  INV_X1 \SB1_2_22/INV_0  ( .A(\RI1[2][54] ), .ZN(\SB1_2_22/i0[9] ) );
  CLKBUF_X1 \SB1_2_17/BUF_0  ( .A(\RI1[2][84] ), .Z(\SB1_2_17/i3[0] ) );
  INV_X1 \SB1_2_24/INV_4  ( .A(\RI1[2][46] ), .ZN(\SB1_2_24/i0_4 ) );
  INV_X1 \SB1_2_3/INV_4  ( .A(\RI1[2][172] ), .ZN(\SB1_2_3/i0_4 ) );
  INV_X1 \SB1_2_30/INV_4  ( .A(\RI1[2][10] ), .ZN(\SB1_2_30/i0_4 ) );
  INV_X1 \SB1_2_22/INV_4  ( .A(\RI1[2][58] ), .ZN(\SB1_2_22/i0_4 ) );
  INV_X1 \SB1_2_7/INV_0  ( .A(\RI1[2][144] ), .ZN(\SB1_2_7/i0[9] ) );
  CLKBUF_X1 \SB1_3_18/BUF_0  ( .A(\RI1[3][78] ), .Z(\SB1_3_18/i3[0] ) );
  CLKBUF_X1 \SB1_3_20/BUF_0  ( .A(\RI1[3][66] ), .Z(\SB1_3_20/i3[0] ) );
  CLKBUF_X1 \SB1_3_15/BUF_4  ( .A(\RI1[3][100] ), .Z(\SB1_3_15/i0[7] ) );
  INV_X1 \SB1_3_7/INV_4  ( .A(\RI1[3][148] ), .ZN(\SB1_3_7/i0_4 ) );
  CLKBUF_X1 \SB1_3_26/BUF_0  ( .A(\RI1[3][30] ), .Z(\SB1_3_26/i3[0] ) );
  CLKBUF_X1 \SB1_3_31/BUF_0  ( .A(\RI1[3][0] ), .Z(\SB1_3_31/i3[0] ) );
  INV_X1 \SB1_3_19/INV_4  ( .A(\RI1[3][76] ), .ZN(\SB1_3_19/i0_4 ) );
  CLKBUF_X1 \SB1_3_6/BUF_0  ( .A(\RI1[3][150] ), .Z(\SB1_3_6/i3[0] ) );
  CLKBUF_X1 \SB1_3_0/BUF_4  ( .A(\RI1[3][190] ), .Z(\SB1_3_0/i0[7] ) );
  CLKBUF_X1 \SB1_3_3/BUF_0  ( .A(\RI1[3][168] ), .Z(\SB1_3_3/i3[0] ) );
  CLKBUF_X1 \SB1_3_16/BUF_0  ( .A(\RI1[3][90] ), .Z(\SB1_3_16/i3[0] ) );
  CLKBUF_X1 \SB1_3_2/BUF_0  ( .A(\RI1[3][174] ), .Z(\SB1_3_2/i3[0] ) );
  INV_X1 \SB1_3_1/INV_4  ( .A(\RI1[3][184] ), .ZN(\SB1_3_1/i0_4 ) );
  CLKBUF_X1 \SB1_3_2/BUF_4  ( .A(\RI1[3][178] ), .Z(\SB1_3_2/i0[7] ) );
  INV_X1 \SB1_3_17/INV_4  ( .A(\RI1[3][88] ), .ZN(\SB1_3_17/i0_4 ) );
  CLKBUF_X1 \SB1_3_12/BUF_0  ( .A(\RI1[3][114] ), .Z(\SB1_3_12/i3[0] ) );
  CLKBUF_X1 \SB1_3_25/BUF_0  ( .A(\RI1[3][36] ), .Z(\SB1_3_25/i3[0] ) );
  CLKBUF_X1 \SB1_3_17/BUF_0  ( .A(\RI1[3][84] ), .Z(\SB1_3_17/i3[0] ) );
  INV_X1 \SB1_3_30/INV_4  ( .A(\RI1[3][10] ), .ZN(\SB1_3_30/i0_4 ) );
  CLKBUF_X1 \SB1_3_9/BUF_0  ( .A(\RI1[3][132] ), .Z(\SB1_3_9/i3[0] ) );
  CLKBUF_X1 \SB1_3_27/BUF_0  ( .A(\RI1[3][24] ), .Z(\SB1_3_27/i3[0] ) );
  CLKBUF_X1 \SB1_3_11/BUF_0  ( .A(\RI1[3][120] ), .Z(\SB1_3_11/i3[0] ) );
  CLKBUF_X1 \SB1_3_24/BUF_0  ( .A(\RI1[3][42] ), .Z(\SB1_3_24/i3[0] ) );
  INV_X1 \SB1_3_23/INV_0  ( .A(\RI1[3][48] ), .ZN(\SB1_3_23/i0[9] ) );
  INV_X1 \SB1_3_12/INV_4  ( .A(\RI1[3][118] ), .ZN(\SB1_3_12/i0_4 ) );
  CLKBUF_X1 \SB1_3_7/BUF_4  ( .A(\RI1[3][148] ), .Z(\SB1_3_7/i0[7] ) );
  CLKBUF_X1 \SB1_3_4/BUF_0  ( .A(\RI1[3][162] ), .Z(\SB1_3_4/i3[0] ) );
  CLKBUF_X1 \SB1_3_23/BUF_0  ( .A(\RI1[3][48] ), .Z(\SB1_3_23/i3[0] ) );
  CLKBUF_X1 \SB1_3_4/BUF_4  ( .A(\RI1[3][166] ), .Z(\SB1_3_4/i0[7] ) );
  CLKBUF_X1 \SB1_3_1/BUF_4  ( .A(\RI1[3][184] ), .Z(\SB1_3_1/i0[7] ) );
  CLKBUF_X1 \SB1_3_22/BUF_0  ( .A(\RI1[3][54] ), .Z(\SB1_3_22/i3[0] ) );
  CLKBUF_X1 \SB1_3_13/BUF_0  ( .A(\RI1[3][108] ), .Z(\SB1_3_13/i3[0] ) );
  CLKBUF_X1 \SB1_3_10/BUF_0  ( .A(\RI1[3][126] ), .Z(\SB1_3_10/i3[0] ) );
  CLKBUF_X1 \SB1_3_8/BUF_0  ( .A(\RI1[3][138] ), .Z(\SB1_3_8/i3[0] ) );
  INV_X1 \SB1_3_22/INV_4  ( .A(\RI1[3][58] ), .ZN(\SB1_3_22/i0_4 ) );
  CLKBUF_X1 \SB1_3_29/BUF_0  ( .A(\RI1[3][12] ), .Z(\SB1_3_29/i3[0] ) );
  INV_X1 \SB1_3_20/INV_0  ( .A(\RI1[3][66] ), .ZN(\SB1_3_20/i0[9] ) );
  CLKBUF_X1 \SB1_3_12/BUF_4  ( .A(\RI1[3][118] ), .Z(\SB1_3_12/i0[7] ) );
  CLKBUF_X1 \SB1_3_29/BUF_4  ( .A(\RI1[3][16] ), .Z(\SB1_3_29/i0[7] ) );
  CLKBUF_X1 \SB1_3_12/BUF_1  ( .A(\RI1[3][115] ), .Z(\SB1_3_12/i1_7 ) );
  INV_X1 \SB1_3_31/INV_4  ( .A(\RI1[3][4] ), .ZN(\SB1_3_31/i0_4 ) );
  CLKBUF_X1 \SB1_3_0/BUF_0  ( .A(\RI1[3][186] ), .Z(\SB1_3_0/i3[0] ) );
  CLKBUF_X1 \SB1_3_17/BUF_4  ( .A(\RI1[3][88] ), .Z(\SB1_3_17/i0[7] ) );
  CLKBUF_X1 \SB1_3_1/BUF_0  ( .A(\RI1[3][180] ), .Z(\SB1_3_1/i3[0] ) );
  CLKBUF_X1 \SB1_3_26/BUF_4  ( .A(\RI1[3][34] ), .Z(\SB1_3_26/i0[7] ) );
  CLKBUF_X1 \SB1_3_30/BUF_0  ( .A(\RI1[3][6] ), .Z(\SB1_3_30/i3[0] ) );
  CLKBUF_X1 \SB1_3_28/BUF_1  ( .A(\RI1[3][19] ), .Z(\SB1_3_28/i1_7 ) );
  CLKBUF_X1 \SB1_3_7/BUF_0  ( .A(\RI1[3][144] ), .Z(\SB1_3_7/i3[0] ) );
  CLKBUF_X1 \SB1_3_28/BUF_0  ( .A(\RI1[3][18] ), .Z(\SB1_3_28/i3[0] ) );
  CLKBUF_X1 \SB1_3_22/BUF_4  ( .A(\RI1[3][58] ), .Z(\SB1_3_22/i0[7] ) );
  INV_X1 \SB1_3_1/INV_0  ( .A(\RI1[3][180] ), .ZN(\SB1_3_1/i0[9] ) );
  CLKBUF_X1 \SB1_3_27/BUF_4  ( .A(\RI1[3][28] ), .Z(\SB1_3_27/i0[7] ) );
  INV_X1 \SB1_3_2/INV_4  ( .A(\RI1[3][178] ), .ZN(\SB1_3_2/i0_4 ) );
  CLKBUF_X1 \SB1_3_24/BUF_4  ( .A(\RI1[3][46] ), .Z(\SB1_3_24/i0[7] ) );
  CLKBUF_X1 \SB1_3_5/BUF_0  ( .A(\RI1[3][156] ), .Z(\SB1_3_5/i3[0] ) );
  CLKBUF_X1 \SB1_3_21/BUF_0  ( .A(\RI1[3][60] ), .Z(\SB1_3_21/i3[0] ) );
  CLKBUF_X1 \SB1_3_9/BUF_4  ( .A(\RI1[3][136] ), .Z(\SB1_3_9/i0[7] ) );
  INV_X1 \SB1_3_28/INV_4  ( .A(\RI1[3][22] ), .ZN(\SB1_3_28/i0_4 ) );
  CLKBUF_X1 \SB1_3_21/BUF_4  ( .A(\RI1[3][64] ), .Z(\SB1_3_21/i0[7] ) );
  INV_X1 \SB1_3_11/INV_4  ( .A(\RI1[3][124] ), .ZN(\SB1_3_11/i0_4 ) );
  INV_X1 \SB1_3_24/INV_4  ( .A(\RI1[3][46] ), .ZN(\SB1_3_24/i0_4 ) );
  CLKBUF_X1 \SB1_3_19/BUF_0  ( .A(\RI1[3][72] ), .Z(\SB1_3_19/i3[0] ) );
  CLKBUF_X1 \SB1_3_19/BUF_4  ( .A(\RI1[3][76] ), .Z(\SB1_3_19/i0[7] ) );
  INV_X1 \SB1_3_14/INV_4  ( .A(\RI1[3][106] ), .ZN(\SB1_3_14/i0_4 ) );
  CLKBUF_X1 \SB1_3_10/BUF_4  ( .A(\RI1[3][130] ), .Z(\SB1_3_10/i0[7] ) );
  CLKBUF_X1 \SB1_3_14/BUF_4  ( .A(\RI1[3][106] ), .Z(\SB1_3_14/i0[7] ) );
  INV_X1 \SB1_3_25/INV_4  ( .A(\RI1[3][40] ), .ZN(\SB1_3_25/i0_4 ) );
  CLKBUF_X1 \SB1_3_15/BUF_0  ( .A(\RI1[3][96] ), .Z(\SB1_3_15/i3[0] ) );
  CLKBUF_X1 \SB1_3_4/BUF_1  ( .A(\RI1[3][163] ), .Z(\SB1_3_4/i1_7 ) );
  INV_X1 \SB1_3_29/INV_4  ( .A(\RI1[3][16] ), .ZN(\SB1_3_29/i0_4 ) );
  CLKBUF_X1 \SB1_3_25/BUF_1  ( .A(\RI1[3][37] ), .Z(\SB1_3_25/i1_7 ) );
  CLKBUF_X1 \SB1_3_14/BUF_0  ( .A(\RI1[3][102] ), .Z(\SB1_3_14/i3[0] ) );
  CLKBUF_X2 \SB2_3_15/BUF_2  ( .A(\RI3[3][98] ), .Z(\SB2_3_15/i0_0 ) );
  CLKBUF_X1 \SB3_3/BUF_0  ( .A(\RI1[4][168] ), .Z(\SB3_3/i3[0] ) );
  CLKBUF_X1 \SB3_31/BUF_0  ( .A(\RI1[4][0] ), .Z(\SB3_31/i3[0] ) );
  CLKBUF_X1 \SB3_30/BUF_0  ( .A(\RI1[4][6] ), .Z(\SB3_30/i3[0] ) );
  CLKBUF_X1 \SB3_28/BUF_0  ( .A(\RI1[4][18] ), .Z(\SB3_28/i3[0] ) );
  CLKBUF_X1 \SB3_0/BUF_0  ( .A(\RI1[4][186] ), .Z(\SB3_0/i3[0] ) );
  INV_X1 \SB3_0/INV_4  ( .A(\RI1[4][190] ), .ZN(\SB3_0/i0_4 ) );
  CLKBUF_X1 \SB3_25/BUF_0  ( .A(\RI1[4][36] ), .Z(\SB3_25/i3[0] ) );
  CLKBUF_X1 \SB3_24/BUF_0  ( .A(\RI1[4][42] ), .Z(\SB3_24/i3[0] ) );
  BUF_X1 \SB3_27/BUF_3  ( .A(\RI1[4][27] ), .Z(\SB3_27/i0[8] ) );
  CLKBUF_X1 \SB3_23/BUF_0  ( .A(\RI1[4][48] ), .Z(\SB3_23/i3[0] ) );
  CLKBUF_X1 \SB3_22/BUF_0  ( .A(\RI1[4][54] ), .Z(\SB3_22/i3[0] ) );
  BUF_X1 \SB3_24/BUF_3  ( .A(\RI1[4][45] ), .Z(\SB3_24/i0[8] ) );
  CLKBUF_X1 \SB3_21/BUF_0  ( .A(\RI1[4][60] ), .Z(\SB3_21/i3[0] ) );
  CLKBUF_X1 \SB3_20/BUF_0  ( .A(\RI1[4][66] ), .Z(\SB3_20/i3[0] ) );
  BUF_X1 \SB3_23/BUF_3  ( .A(\RI1[4][51] ), .Z(\SB3_23/i0[8] ) );
  CLKBUF_X1 \SB3_1/BUF_0  ( .A(\RI1[4][180] ), .Z(\SB3_1/i3[0] ) );
  CLKBUF_X1 \SB3_16/BUF_0  ( .A(\RI1[4][90] ), .Z(\SB3_16/i3[0] ) );
  CLKBUF_X1 \SB3_15/BUF_0  ( .A(\RI1[4][96] ), .Z(\SB3_15/i3[0] ) );
  CLKBUF_X1 \SB3_14/BUF_0  ( .A(\RI1[4][102] ), .Z(\SB3_14/i3[0] ) );
  CLKBUF_X1 \SB3_13/BUF_0  ( .A(\RI1[4][108] ), .Z(\SB3_13/i3[0] ) );
  CLKBUF_X1 \SB3_10/BUF_0  ( .A(\RI1[4][126] ), .Z(\SB3_10/i3[0] ) );
  BUF_X1 \SB3_0/BUF_3  ( .A(\RI1[4][189] ), .Z(\SB3_0/i0[8] ) );
  CLKBUF_X1 \SB3_7/BUF_0  ( .A(\RI1[4][144] ), .Z(\SB3_7/i3[0] ) );
  CLKBUF_X1 \SB3_5/BUF_0  ( .A(\RI1[4][156] ), .Z(\SB3_5/i3[0] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_172_0  ( .A(Key[60]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[172] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_129_0  ( .A(Key[180]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[129] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_165_0  ( .A(Key[61]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[165] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_134_0  ( .A(Key[78]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[134] ) );
  CLKBUF_X1 \SB1_0_3/BUF_1  ( .A(n23), .Z(\SB1_0_3/i1_7 ) );
  CLKBUF_X1 \SB1_0_21/BUF_0  ( .A(n132), .Z(\SB1_0_21/i3[0] ) );
  CLKBUF_X1 \SB1_0_11/BUF_4  ( .A(n68), .Z(\SB1_0_11/i0[7] ) );
  CLKBUF_X1 \SB1_0_18/BUF_0  ( .A(n114), .Z(\SB1_0_18/i3[0] ) );
  CLKBUF_X1 \SB1_0_13/BUF_1  ( .A(n83), .Z(\SB1_0_13/i1_7 ) );
  CLKBUF_X1 \SB1_0_20/BUF_1  ( .A(n125), .Z(\SB1_0_20/i1_7 ) );
  CLKBUF_X1 \SB1_0_6/BUF_1  ( .A(n41), .Z(\SB1_0_6/i1_7 ) );
  BUF_X1 \SB1_0_14/BUF_5  ( .A(n85), .Z(\SB1_0_14/i1_5 ) );
  CLKBUF_X1 \SB1_0_6/BUF_0  ( .A(n42), .Z(\SB1_0_6/i3[0] ) );
  BUF_X1 \SB2_0_20/BUF_1  ( .A(\RI3[0][67] ), .Z(\SB2_0_20/i0[6] ) );
  BUF_X1 \SB2_0_4/BUF_0  ( .A(\RI3[0][162] ), .Z(\SB2_0_4/i0[9] ) );
  CLKBUF_X1 \SB1_1_13/BUF_1  ( .A(\RI1[1][109] ), .Z(\SB1_1_13/i1_7 ) );
  CLKBUF_X1 \SB1_1_17/BUF_4  ( .A(\RI1[1][88] ), .Z(\SB1_1_17/i0[7] ) );
  CLKBUF_X1 \SB1_1_8/BUF_1  ( .A(\RI1[1][139] ), .Z(\SB1_1_8/i1_7 ) );
  CLKBUF_X1 \SB1_1_23/BUF_1  ( .A(\RI1[1][49] ), .Z(\SB1_1_23/i1_7 ) );
  CLKBUF_X1 \SB1_1_25/BUF_1  ( .A(\RI1[1][37] ), .Z(\SB1_1_25/i1_7 ) );
  CLKBUF_X1 \SB1_1_6/BUF_1  ( .A(\RI1[1][151] ), .Z(\SB1_1_6/i1_7 ) );
  CLKBUF_X1 \SB1_1_19/BUF_1  ( .A(\RI1[1][73] ), .Z(\SB1_1_19/i1_7 ) );
  CLKBUF_X1 \SB1_2_5/BUF_1  ( .A(\RI1[2][157] ), .Z(\SB1_2_5/i1_7 ) );
  CLKBUF_X1 \SB1_2_0/BUF_1  ( .A(\RI1[2][187] ), .Z(\SB1_2_0/i1_7 ) );
  CLKBUF_X1 \SB1_2_7/BUF_1  ( .A(\RI1[2][145] ), .Z(\SB1_2_7/i1_7 ) );
  CLKBUF_X1 \SB1_2_23/BUF_1  ( .A(\RI1[2][49] ), .Z(\SB1_2_23/i1_7 ) );
  CLKBUF_X1 \SB1_2_4/BUF_1  ( .A(\RI1[2][163] ), .Z(\SB1_2_4/i1_7 ) );
  CLKBUF_X1 \SB1_2_8/BUF_1  ( .A(\RI1[2][139] ), .Z(\SB1_2_8/i1_7 ) );
  CLKBUF_X1 \SB1_2_23/BUF_4  ( .A(\RI1[2][52] ), .Z(\SB1_2_23/i0[7] ) );
  CLKBUF_X1 \SB1_2_2/BUF_1  ( .A(\RI1[2][175] ), .Z(\SB1_2_2/i1_7 ) );
  CLKBUF_X1 \SB1_2_3/BUF_4  ( .A(\RI1[2][172] ), .Z(\SB1_2_3/i0[7] ) );
  CLKBUF_X1 \SB1_2_27/BUF_1  ( .A(\RI1[2][25] ), .Z(\SB1_2_27/i1_7 ) );
  CLKBUF_X1 \SB1_3_30/BUF_4  ( .A(\RI1[3][10] ), .Z(\SB1_3_30/i0[7] ) );
  CLKBUF_X1 \SB1_3_14/BUF_1  ( .A(\RI1[3][103] ), .Z(\SB1_3_14/i1_7 ) );
  CLKBUF_X1 \SB1_3_15/BUF_1  ( .A(\RI1[3][97] ), .Z(\SB1_3_15/i1_7 ) );
  CLKBUF_X1 \SB1_3_30/BUF_1  ( .A(\RI1[3][7] ), .Z(\SB1_3_30/i1_7 ) );
  CLKBUF_X1 \SB1_3_8/BUF_1  ( .A(\RI1[3][139] ), .Z(\SB1_3_8/i1_7 ) );
  CLKBUF_X1 \SB1_3_19/BUF_1  ( .A(\RI1[3][73] ), .Z(\SB1_3_19/i1_7 ) );
  CLKBUF_X1 \SB1_3_31/BUF_4  ( .A(\RI1[3][4] ), .Z(\SB1_3_31/i0[7] ) );
  CLKBUF_X1 \SB1_3_11/BUF_1  ( .A(\RI1[3][121] ), .Z(\SB1_3_11/i1_7 ) );
  CLKBUF_X1 \SB1_3_6/BUF_1  ( .A(\RI1[3][151] ), .Z(\SB1_3_6/i1_7 ) );
  CLKBUF_X1 \SB1_3_13/BUF_1  ( .A(\RI1[3][109] ), .Z(\SB1_3_13/i1_7 ) );
  BUF_X1 \SB2_3_11/BUF_0  ( .A(\RI3[3][120] ), .Z(\SB2_3_11/i0[9] ) );
  BUF_X2 \SB2_0_21/BUF_3  ( .A(\RI3[0][63] ), .Z(\SB2_0_21/i0[10] ) );
  BUF_X2 \SB2_0_16/BUF_3  ( .A(\RI3[0][93] ), .Z(\SB2_0_16/i0[10] ) );
  BUF_X2 \SB2_0_11/BUF_2  ( .A(\RI3[0][122] ), .Z(\SB2_0_11/i0_0 ) );
  BUF_X2 \SB2_0_6/BUF_2  ( .A(\RI3[0][152] ), .Z(\SB2_0_6/i0_0 ) );
  BUF_X2 \SB2_1_0/BUF_2  ( .A(\RI3[1][188] ), .Z(\SB2_1_0/i0_0 ) );
  BUF_X2 \SB2_0_22/BUF_2  ( .A(\RI3[0][56] ), .Z(\SB2_0_22/i0_0 ) );
  BUF_X2 \SB2_0_0/BUF_2  ( .A(\RI3[0][188] ), .Z(\SB2_0_0/i0_0 ) );
  BUF_X2 \SB2_0_7/BUF_2  ( .A(\RI3[0][146] ), .Z(\SB2_0_7/i0_0 ) );
  BUF_X2 \SB2_0_5/BUF_3  ( .A(\RI3[0][159] ), .Z(\SB2_0_5/i0[10] ) );
  BUF_X2 \SB2_0_27/BUF_3  ( .A(\RI3[0][27] ), .Z(\SB2_0_27/i0[10] ) );
  BUF_X2 \SB2_0_20/BUF_3  ( .A(\RI3[0][69] ), .Z(\SB2_0_20/i0[10] ) );
  BUF_X2 \SB2_0_22/BUF_3  ( .A(\RI3[0][57] ), .Z(\SB2_0_22/i0[10] ) );
  BUF_X2 \SB2_0_19/BUF_2  ( .A(\RI3[0][74] ), .Z(\SB2_0_19/i0_0 ) );
  BUF_X2 \SB2_0_27/BUF_2  ( .A(\RI3[0][26] ), .Z(\SB2_0_27/i0_0 ) );
  BUF_X2 \SB2_0_4/BUF_2  ( .A(\RI3[0][164] ), .Z(\SB2_0_4/i0_0 ) );
  BUF_X2 \SB1_1_28/BUF_2  ( .A(\RI1[1][20] ), .Z(\SB1_1_28/i1[9] ) );
  BUF_X2 \SB2_0_29/BUF_2  ( .A(\RI3[0][14] ), .Z(\SB2_0_29/i0_0 ) );
  BUF_X2 \SB2_0_9/BUF_3  ( .A(\RI3[0][135] ), .Z(\SB2_0_9/i0[10] ) );
  BUF_X2 \SB2_0_12/BUF_2  ( .A(\RI3[0][116] ), .Z(\SB2_0_12/i0_0 ) );
  BUF_X2 \SB2_0_21/BUF_2  ( .A(\RI3[0][62] ), .Z(\SB2_0_21/i0_0 ) );
  BUF_X2 \SB2_0_31/BUF_2  ( .A(\RI3[0][2] ), .Z(\SB2_0_31/i0_0 ) );
  BUF_X2 \SB2_0_13/BUF_3  ( .A(\RI3[0][111] ), .Z(\SB2_0_13/i0[10] ) );
  BUF_X2 \SB2_1_2/BUF_1  ( .A(\RI3[1][175] ), .Z(\SB2_1_2/i0[6] ) );
  BUF_X2 \SB1_1_12/BUF_2  ( .A(\RI1[1][116] ), .Z(\SB1_1_12/i1[9] ) );
  BUF_X2 \SB2_0_24/BUF_3  ( .A(\RI3[0][45] ), .Z(\SB2_0_24/i0[10] ) );
  BUF_X2 \SB2_0_2/BUF_2  ( .A(\RI3[0][176] ), .Z(\SB2_0_2/i0_0 ) );
  BUF_X2 \SB1_1_11/BUF_2  ( .A(\RI1[1][122] ), .Z(\SB1_1_11/i1[9] ) );
  BUF_X2 \SB2_0_26/BUF_3  ( .A(\RI3[0][33] ), .Z(\SB2_0_26/i0[10] ) );
  BUF_X2 \SB2_0_25/BUF_3  ( .A(\RI3[0][39] ), .Z(\SB2_0_25/i0[10] ) );
  BUF_X2 \SB1_1_31/BUF_2  ( .A(\RI1[1][2] ), .Z(\SB1_1_31/i1[9] ) );
  BUF_X2 \SB2_1_27/BUF_1  ( .A(\RI3[1][25] ), .Z(\SB2_1_27/i0[6] ) );
  BUF_X1 \SB1_1_27/BUF_5  ( .A(\RI1[1][29] ), .Z(\SB1_1_27/i1_5 ) );
  BUF_X2 \SB1_2_30/BUF_2  ( .A(\RI1[2][8] ), .Z(\SB1_2_30/i1[9] ) );
  BUF_X1 \SB1_0_13/BUF_5  ( .A(n79), .Z(\SB1_0_13/i1_5 ) );
  BUF_X2 \SB2_0_31/BUF_3  ( .A(\RI3[0][3] ), .Z(\SB2_0_31/i0[10] ) );
  BUF_X1 \SB1_0_31/BUF_5  ( .A(n187), .Z(\SB1_0_31/i1_5 ) );
  BUF_X2 \SB1_2_22/BUF_2  ( .A(\RI1[2][56] ), .Z(\SB1_2_22/i1[9] ) );
  INV_X1 \SB2_0_20/INV_2  ( .A(\RI3[0][68] ), .ZN(\SB2_0_20/i1[9] ) );
  BUF_X2 \SB4_17/BUF_3  ( .A(\RI3[4][87] ), .Z(\SB4_17/i0[10] ) );
  BUF_X2 \SB4_0/BUF_3  ( .A(\RI3[4][189] ), .Z(\SB4_0/i0[10] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_16  ( .A(\RI5[3][16] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[16] ) );
  INV_X1 \SB2_3_21/INV_2  ( .A(\RI3[3][62] ), .ZN(\SB2_3_21/i1[9] ) );
  BUF_X2 \SB4_26/BUF_0  ( .A(\RI3[4][30] ), .Z(\SB4_26/i0[9] ) );
  BUF_X2 \SB4_17/BUF_0  ( .A(\RI3[4][84] ), .Z(\SB4_17/i0[9] ) );
  BUF_X2 \SB4_4/BUF_0  ( .A(\RI3[4][162] ), .Z(\SB4_4/i0[9] ) );
  BUF_X1 \SB1_0_20/BUF_3  ( .A(n123), .Z(\SB1_0_20/i0[8] ) );
  BUF_X1 \SB1_0_21/BUF_5  ( .A(n127), .Z(\SB1_0_21/i1_5 ) );
  INV_X1 \SB1_1_5/INV_0  ( .A(\RI1[1][156] ), .ZN(\SB1_1_5/i0[9] ) );
  INV_X1 \SB1_1_15/INV_0  ( .A(\RI1[1][96] ), .ZN(\SB1_1_15/i0[9] ) );
  INV_X1 \SB1_2_6/INV_0  ( .A(\RI1[2][150] ), .ZN(\SB1_2_6/i0[9] ) );
  INV_X1 \SB1_2_18/INV_0  ( .A(\RI1[2][78] ), .ZN(\SB1_2_18/i0[9] ) );
  INV_X1 \SB1_2_23/INV_0  ( .A(\RI1[2][48] ), .ZN(\SB1_2_23/i0[9] ) );
  INV_X1 \SB1_2_28/INV_0  ( .A(\RI1[2][18] ), .ZN(\SB1_2_28/i0[9] ) );
  INV_X1 \SB1_2_13/INV_0  ( .A(\RI1[2][108] ), .ZN(\SB1_2_13/i0[9] ) );
  INV_X1 \SB1_2_8/INV_0  ( .A(\RI1[2][138] ), .ZN(\SB1_2_8/i0[9] ) );
  BUF_X1 \SB2_2_18/BUF_0  ( .A(\RI3[2][78] ), .Z(\SB2_2_18/i0[9] ) );
  INV_X1 \SB1_3_26/INV_0  ( .A(\RI1[3][30] ), .ZN(\SB1_3_26/i0[9] ) );
  INV_X1 \SB1_3_16/INV_0  ( .A(\RI1[3][90] ), .ZN(\SB1_3_16/i0[9] ) );
  INV_X1 \SB1_3_11/INV_0  ( .A(\RI1[3][120] ), .ZN(\SB1_3_11/i0[9] ) );
  BUF_X1 \SB2_3_29/BUF_0  ( .A(\RI3[3][12] ), .Z(\SB2_3_29/i0[9] ) );
  BUF_X1 \SB3_12/BUF_2  ( .A(\RI1[4][116] ), .Z(\SB3_12/i1[9] ) );
  BUF_X1 \SB3_19/BUF_2  ( .A(\RI1[4][74] ), .Z(\SB3_19/i1[9] ) );
  CLKBUF_X1 U5 ( .A(Key[80]), .Z(n512) );
  CLKBUF_X1 U7 ( .A(Key[97]), .Z(n457) );
  CLKBUF_X1 U10 ( .A(Key[58]), .Z(n482) );
  CLKBUF_X1 U12 ( .A(Key[7]), .Z(n468) );
  CLKBUF_X1 U13 ( .A(Key[35]), .Z(n407) );
  CLKBUF_X1 U14 ( .A(Key[69]), .Z(n449) );
  CLKBUF_X1 U16 ( .A(Key[126]), .Z(n383) );
  CLKBUF_X1 U17 ( .A(Key[140]), .Z(n487) );
  CLKBUF_X1 U18 ( .A(Key[154]), .Z(n489) );
  CLKBUF_X1 U19 ( .A(Key[147]), .Z(n507) );
  CLKBUF_X1 U20 ( .A(Key[125]), .Z(n445) );
  CLKBUF_X1 U21 ( .A(Key[146]), .Z(n476) );
  CLKBUF_X1 U26 ( .A(Key[3]), .Z(n473) );
  CLKBUF_X1 U27 ( .A(Key[129]), .Z(n419) );
  CLKBUF_X1 U28 ( .A(Key[66]), .Z(n428) );
  CLKBUF_X1 U29 ( .A(Key[87]), .Z(n450) );
  CLKBUF_X1 U33 ( .A(Key[86]), .Z(n438) );
  CLKBUF_X1 U35 ( .A(Key[34]), .Z(n464) );
  CLKBUF_X1 U36 ( .A(Key[20]), .Z(n478) );
  CLKBUF_X1 U37 ( .A(Key[170]), .Z(n481) );
  CLKBUF_X1 U38 ( .A(Key[177]), .Z(n484) );
  CLKBUF_X1 U40 ( .A(Key[118]), .Z(n439) );
  CLKBUF_X1 U42 ( .A(Key[62]), .Z(n500) );
  CLKBUF_X1 U43 ( .A(Key[76]), .Z(n458) );
  CLKBUF_X1 U44 ( .A(Key[159]), .Z(n511) );
  CLKBUF_X1 U47 ( .A(Key[134]), .Z(n451) );
  CLKBUF_X1 U48 ( .A(Key[113]), .Z(n396) );
  CLKBUF_X1 U56 ( .A(Key[5]), .Z(n389) );
  CLKBUF_X1 U59 ( .A(Key[33]), .Z(n504) );
  CLKBUF_X1 U60 ( .A(Key[176]), .Z(n421) );
  CLKBUF_X1 U61 ( .A(Key[169]), .Z(n433) );
  CLKBUF_X1 U62 ( .A(Key[190]), .Z(n430) );
  CLKBUF_X1 U64 ( .A(Key[183]), .Z(n508) );
  CLKBUF_X1 U68 ( .A(Key[74]), .Z(n497) );
  CLKBUF_X1 U70 ( .A(Key[96]), .Z(n424) );
  CLKBUF_X1 U71 ( .A(Key[32]), .Z(n460) );
  CLKBUF_X1 U73 ( .A(Key[46]), .Z(n462) );
  CLKBUF_X1 U74 ( .A(Key[165]), .Z(n493) );
  CLKBUF_X1 U75 ( .A(Key[51]), .Z(n496) );
  CLKBUF_X1 U77 ( .A(Key[137]), .Z(n408) );
  CLKBUF_X1 U79 ( .A(Key[166]), .Z(n431) );
  INV_X1 U81 ( .A(\MC_ARK_ARC_1_2/buf_keyinput[112] ), .ZN(n271) );
  CLKBUF_X1 U82 ( .A(Key[123]), .Z(n492) );
  CLKBUF_X1 U83 ( .A(Key[43]), .Z(n384) );
  CLKBUF_X1 U85 ( .A(Key[57]), .Z(n444) );
  INV_X1 U86 ( .A(Key[186]), .ZN(n198) );
  CLKBUF_X1 U87 ( .A(Key[8]), .Z(n499) );
  CLKBUF_X1 U88 ( .A(Key[22]), .Z(n447) );
  CLKBUF_X1 U89 ( .A(Key[15]), .Z(n506) );
  CLKBUF_X1 U91 ( .A(Key[14]), .Z(n379) );
  CLKBUF_X1 U92 ( .A(Key[164]), .Z(n441) );
  CLKBUF_X1 U98 ( .A(Key[98]), .Z(n440) );
  CLKBUF_X1 U101 ( .A(Key[63]), .Z(n505) );
  CLKBUF_X1 U103 ( .A(Key[4]), .Z(n432) );
  XNOR2_X1 U104 ( .A(Key[191]), .B(Plaintext[191]), .ZN(n380) );
  XNOR2_X1 U105 ( .A(Key[119]), .B(Plaintext[119]), .ZN(n381) );
  BUF_X1 U108 ( .A(Key[101]), .Z(n494) );
  BUF_X1 U109 ( .A(Key[23]), .Z(n465) );
  INV_X1 U110 ( .A(Key[138]), .ZN(n244) );
  INV_X1 U114 ( .A(n386), .ZN(n234) );
  INV_X1 U115 ( .A(Key[102]), .ZN(n278) );
  INV_X1 U116 ( .A(n385), .ZN(n216) );
  BUF_X1 U118 ( .A(Key[95]), .Z(n479) );
  BUF_X1 U120 ( .A(Key[149]), .Z(n386) );
  BUF_X1 U124 ( .A(Key[89]), .Z(n390) );
  BUF_X1 U125 ( .A(Key[131]), .Z(n391) );
  BUF_X1 U128 ( .A(Key[59]), .Z(n394) );
  BUF_X1 U129 ( .A(Key[143]), .Z(n395) );
  BUF_X1 U132 ( .A(Key[47]), .Z(n399) );
  BUF_X1 U133 ( .A(Key[41]), .Z(n400) );
  BUF_X1 U134 ( .A(Key[179]), .Z(n401) );
  BUF_X1 U136 ( .A(Key[29]), .Z(n403) );
  BUF_X1 U137 ( .A(Key[65]), .Z(n404) );
  INV_X1 U140 ( .A(\MC_ARK_ARC_1_0/buf_keyinput[11] ), .ZN(n297) );
  INV_X1 U141 ( .A(n454), .ZN(n199) );
  INV_X1 U142 ( .A(n389), .ZN(n369) );
  INV_X1 U145 ( .A(n440), .ZN(n282) );
  INV_X1 U146 ( .A(Key[90]), .ZN(n289) );
  INV_X1 U147 ( .A(Key[187]), .ZN(n197) );
  INV_X1 U148 ( .A(Key[127]), .ZN(n253) );
  INV_X1 U149 ( .A(Key[13]), .ZN(n362) );
  INV_X1 U150 ( .A(Key[151]), .ZN(n232) );
  INV_X1 U154 ( .A(Key[83]), .ZN(n296) );
  INV_X1 U155 ( .A(Key[53]), .ZN(n324) );
  INV_X1 U156 ( .A(Key[155]), .ZN(n228) );
  INV_X1 U157 ( .A(Key[42]), .ZN(n335) );
  INV_X1 U158 ( .A(Key[108]), .ZN(n272) );
  INV_X1 U160 ( .A(Key[72]), .ZN(n306) );
  INV_X1 U161 ( .A(n445), .ZN(n255) );
  INV_X1 U163 ( .A(Key[36]), .ZN(n340) );
  INV_X1 U164 ( .A(Key[120]), .ZN(n260) );
  INV_X1 U166 ( .A(n392), .ZN(n222) );
  INV_X1 U167 ( .A(n387), .ZN(n301) );
  INV_X1 U168 ( .A(Key[117]), .ZN(n263) );
  INV_X1 U173 ( .A(Key[133]), .ZN(n248) );
  INV_X1 U175 ( .A(n422), .ZN(n287) );
  INV_X1 U177 ( .A(\MC_ARK_ARC_1_2/buf_keyinput[143] ), .ZN(n201) );
  INV_X1 U179 ( .A(\MC_ARK_ARC_1_1/buf_keyinput[106] ), .ZN(n327) );
  INV_X1 U180 ( .A(Key[2]), .ZN(n372) );
  INV_X1 U182 ( .A(n421), .ZN(n207) );
  INV_X1 U183 ( .A(Key[158]), .ZN(n225) );
  INV_X1 U184 ( .A(Key[160]), .ZN(n223) );
  INV_X1 U186 ( .A(n432), .ZN(n370) );
  INV_X1 U189 ( .A(n493), .ZN(n218) );
  INV_X1 U191 ( .A(n488), .ZN(n298) );
  INV_X1 U192 ( .A(Key[25]), .ZN(n350) );
  INV_X1 U193 ( .A(Key[1]), .ZN(n373) );
  INV_X1 U194 ( .A(n465), .ZN(n352) );
  INV_X1 U195 ( .A(n394), .ZN(n319) );
  INV_X1 U197 ( .A(n395), .ZN(n240) );
  INV_X1 U198 ( .A(Key[6]), .ZN(n368) );
  INV_X1 U199 ( .A(Key[78]), .ZN(n300) );
  INV_X1 U200 ( .A(Key[0]), .ZN(n374) );
  INV_X1 U202 ( .A(n466), .ZN(n349) );
  INV_X1 U203 ( .A(n480), .ZN(n338) );
  INV_X1 U204 ( .A(n485), .ZN(n231) );
  INV_X1 U207 ( .A(n479), .ZN(n284) );
  INV_X1 U209 ( .A(n400), .ZN(n336) );
  INV_X1 U211 ( .A(n430), .ZN(n194) );
  INV_X1 U212 ( .A(n439), .ZN(n262) );
  INV_X1 U213 ( .A(n437), .ZN(n321) );
  INV_X1 U214 ( .A(n486), .ZN(n310) );
  INV_X1 U215 ( .A(Key[30]), .ZN(n345) );
  INV_X1 U217 ( .A(n477), .ZN(n276) );
  INV_X1 U218 ( .A(n478), .ZN(n355) );
  INV_X1 U219 ( .A(n476), .ZN(n237) );
  INV_X1 U220 ( .A(n438), .ZN(n293) );
  INV_X1 U221 ( .A(Key[144]), .ZN(n239) );
  INV_X1 U222 ( .A(Key[174]), .ZN(n209) );
  INV_X1 U224 ( .A(Key[37]), .ZN(n339) );
  INV_X1 U225 ( .A(Key[55]), .ZN(n322) );
  INV_X1 U226 ( .A(Key[157]), .ZN(n226) );
  INV_X1 U227 ( .A(\MC_ARK_ARC_1_0/buf_keyinput[80] ), .ZN(n202) );
  INV_X1 U228 ( .A(Key[79]), .ZN(n299) );
  INV_X1 U230 ( .A(Key[73]), .ZN(n305) );
  INV_X1 U233 ( .A(n449), .ZN(n309) );
  INV_X1 U234 ( .A(Key[24]), .ZN(n351) );
  INV_X1 U235 ( .A(Key[84]), .ZN(n295) );
  INV_X1 U237 ( .A(\MC_ARK_ARC_1_3/buf_keyinput[172] ), .ZN(n318) );
  INV_X1 U238 ( .A(n393), .ZN(n358) );
  INV_X1 U239 ( .A(\MC_ARK_ARC_1_2/buf_keyinput[177] ), .ZN(n249) );
  INV_X1 U240 ( .A(Key[114]), .ZN(n266) );
  INV_X1 U242 ( .A(Key[54]), .ZN(n323) );
  INV_X1 U243 ( .A(n396), .ZN(n267) );
  INV_X1 U244 ( .A(n399), .ZN(n330) );
  INV_X1 U246 ( .A(Key[49]), .ZN(n328) );
  INV_X1 U248 ( .A(Key[115]), .ZN(n265) );
  INV_X1 U249 ( .A(Key[61]), .ZN(n317) );
  INV_X1 U251 ( .A(n441), .ZN(n219) );
  INV_X1 U252 ( .A(n481), .ZN(n213) );
  INV_X1 U256 ( .A(n431), .ZN(n217) );
  INV_X1 U257 ( .A(n436), .ZN(n205) );
  INV_X1 U258 ( .A(n376), .ZN(n245) );
  INV_X1 U262 ( .A(n377), .ZN(n227) );
  INV_X1 U264 ( .A(n406), .ZN(n193) );
  XNOR2_X1 U265 ( .A(Key[191]), .B(Plaintext[191]), .ZN(n1) );
  XNOR2_X1 U266 ( .A(Key[86]), .B(Plaintext[86]), .ZN(n106) );
  XNOR2_X1 U268 ( .A(Key[75]), .B(Plaintext[75]), .ZN(n117) );
  XNOR2_X1 U271 ( .A(Key[56]), .B(Plaintext[56]), .ZN(n136) );
  INV_X1 U272 ( .A(n443), .ZN(n311) );
  INV_X1 U274 ( .A(n511), .ZN(n224) );
  XNOR2_X1 U275 ( .A(Key[159]), .B(Plaintext[159]), .ZN(n33) );
  XNOR2_X1 U276 ( .A(Key[122]), .B(Plaintext[122]), .ZN(n70) );
  INV_X1 U278 ( .A(n472), .ZN(n337) );
  XNOR2_X1 U279 ( .A(Key[39]), .B(Plaintext[39]), .ZN(n153) );
  XNOR2_X1 U281 ( .A(Key[57]), .B(Plaintext[57]), .ZN(n135) );
  INV_X1 U282 ( .A(n423), .ZN(n288) );
  XNOR2_X1 U284 ( .A(Key[14]), .B(Plaintext[14]), .ZN(n178) );
  INV_X1 U285 ( .A(Key[85]), .ZN(n294) );
  XNOR2_X1 U287 ( .A(Key[51]), .B(Plaintext[51]), .ZN(n141) );
  XNOR2_X1 U288 ( .A(Key[188]), .B(Plaintext[188]), .ZN(n4) );
  XNOR2_X1 U289 ( .A(Key[20]), .B(Plaintext[20]), .ZN(n172) );
  XNOR2_X1 U290 ( .A(Key[17]), .B(Plaintext[17]), .ZN(n175) );
  XNOR2_X1 U291 ( .A(Key[123]), .B(Plaintext[123]), .ZN(n69) );
  INV_X1 U292 ( .A(Key[19]), .ZN(n356) );
  INV_X1 U295 ( .A(n433), .ZN(n214) );
  XNOR2_X1 U299 ( .A(Key[183]), .B(Plaintext[183]), .ZN(n9) );
  INV_X1 U301 ( .A(n504), .ZN(n342) );
  XNOR2_X1 U303 ( .A(Key[15]), .B(Plaintext[15]), .ZN(n177) );
  INV_X1 U306 ( .A(n510), .ZN(n246) );
  XNOR2_X1 U311 ( .A(Key[0]), .B(Plaintext[0]), .ZN(n192) );
  XNOR2_X1 U312 ( .A(Key[1]), .B(Plaintext[1]), .ZN(n191) );
  XNOR2_X1 U313 ( .A(Key[2]), .B(Plaintext[2]), .ZN(n190) );
  XNOR2_X1 U314 ( .A(Key[3]), .B(Plaintext[3]), .ZN(n189) );
  XNOR2_X1 U315 ( .A(Key[4]), .B(Plaintext[4]), .ZN(n188) );
  XNOR2_X1 U316 ( .A(Key[5]), .B(Plaintext[5]), .ZN(n187) );
  XNOR2_X1 U317 ( .A(Key[6]), .B(Plaintext[6]), .ZN(n186) );
  XNOR2_X1 U318 ( .A(Key[7]), .B(Plaintext[7]), .ZN(n185) );
  XNOR2_X1 U319 ( .A(Key[8]), .B(Plaintext[8]), .ZN(n184) );
  XNOR2_X1 U320 ( .A(Key[9]), .B(Plaintext[9]), .ZN(n183) );
  XNOR2_X1 U321 ( .A(Key[10]), .B(Plaintext[10]), .ZN(n182) );
  XNOR2_X1 U322 ( .A(Key[11]), .B(Plaintext[11]), .ZN(n181) );
  XNOR2_X1 U323 ( .A(Key[12]), .B(Plaintext[12]), .ZN(n180) );
  XNOR2_X1 U324 ( .A(Key[13]), .B(Plaintext[13]), .ZN(n179) );
  XNOR2_X1 U325 ( .A(Key[16]), .B(Plaintext[16]), .ZN(n176) );
  XNOR2_X1 U326 ( .A(Key[18]), .B(Plaintext[18]), .ZN(n174) );
  XNOR2_X1 U327 ( .A(Key[19]), .B(Plaintext[19]), .ZN(n173) );
  XNOR2_X1 U328 ( .A(Key[21]), .B(Plaintext[21]), .ZN(n171) );
  XNOR2_X1 U329 ( .A(Key[22]), .B(Plaintext[22]), .ZN(n170) );
  XNOR2_X1 U330 ( .A(Key[23]), .B(Plaintext[23]), .ZN(n169) );
  XNOR2_X1 U331 ( .A(Key[24]), .B(Plaintext[24]), .ZN(n168) );
  XNOR2_X1 U332 ( .A(Key[25]), .B(Plaintext[25]), .ZN(n167) );
  XNOR2_X1 U333 ( .A(Key[26]), .B(Plaintext[26]), .ZN(n166) );
  XNOR2_X1 U334 ( .A(Key[27]), .B(Plaintext[27]), .ZN(n165) );
  XNOR2_X1 U335 ( .A(Key[28]), .B(Plaintext[28]), .ZN(n164) );
  XNOR2_X1 U336 ( .A(Key[29]), .B(Plaintext[29]), .ZN(n163) );
  XNOR2_X1 U337 ( .A(Key[30]), .B(Plaintext[30]), .ZN(n162) );
  XNOR2_X1 U338 ( .A(Key[31]), .B(Plaintext[31]), .ZN(n161) );
  XNOR2_X1 U339 ( .A(Key[32]), .B(Plaintext[32]), .ZN(n160) );
  XNOR2_X1 U340 ( .A(Key[33]), .B(Plaintext[33]), .ZN(n159) );
  XNOR2_X1 U341 ( .A(Key[34]), .B(Plaintext[34]), .ZN(n158) );
  XNOR2_X1 U342 ( .A(Key[35]), .B(Plaintext[35]), .ZN(n157) );
  XNOR2_X1 U343 ( .A(Key[36]), .B(Plaintext[36]), .ZN(n156) );
  XNOR2_X1 U344 ( .A(Key[37]), .B(Plaintext[37]), .ZN(n155) );
  XNOR2_X1 U345 ( .A(Key[38]), .B(Plaintext[38]), .ZN(n154) );
  XNOR2_X1 U346 ( .A(Key[40]), .B(Plaintext[40]), .ZN(n152) );
  XNOR2_X1 U347 ( .A(Key[41]), .B(Plaintext[41]), .ZN(n151) );
  XNOR2_X1 U348 ( .A(Key[42]), .B(Plaintext[42]), .ZN(n150) );
  XNOR2_X1 U349 ( .A(Key[43]), .B(Plaintext[43]), .ZN(n149) );
  XNOR2_X1 U350 ( .A(Key[44]), .B(Plaintext[44]), .ZN(n148) );
  XNOR2_X1 U351 ( .A(Key[45]), .B(Plaintext[45]), .ZN(n147) );
  XNOR2_X1 U352 ( .A(Key[46]), .B(Plaintext[46]), .ZN(n146) );
  XNOR2_X1 U353 ( .A(Key[47]), .B(Plaintext[47]), .ZN(n145) );
  XNOR2_X1 U354 ( .A(Key[48]), .B(Plaintext[48]), .ZN(n144) );
  XNOR2_X1 U355 ( .A(Key[49]), .B(Plaintext[49]), .ZN(n143) );
  XNOR2_X1 U356 ( .A(Key[50]), .B(Plaintext[50]), .ZN(n142) );
  XNOR2_X1 U357 ( .A(Key[52]), .B(Plaintext[52]), .ZN(n140) );
  XNOR2_X1 U358 ( .A(Key[53]), .B(Plaintext[53]), .ZN(n139) );
  XNOR2_X1 U359 ( .A(Key[54]), .B(Plaintext[54]), .ZN(n138) );
  XNOR2_X1 U360 ( .A(Key[55]), .B(Plaintext[55]), .ZN(n137) );
  XNOR2_X1 U361 ( .A(Key[58]), .B(Plaintext[58]), .ZN(n134) );
  XNOR2_X1 U362 ( .A(Key[59]), .B(Plaintext[59]), .ZN(n133) );
  XNOR2_X1 U363 ( .A(Key[60]), .B(Plaintext[60]), .ZN(n132) );
  XNOR2_X1 U364 ( .A(Key[61]), .B(Plaintext[61]), .ZN(n131) );
  XNOR2_X1 U365 ( .A(Key[62]), .B(Plaintext[62]), .ZN(n130) );
  XNOR2_X1 U366 ( .A(Key[63]), .B(Plaintext[63]), .ZN(n129) );
  XNOR2_X1 U367 ( .A(Key[64]), .B(Plaintext[64]), .ZN(n128) );
  XNOR2_X1 U368 ( .A(Key[65]), .B(Plaintext[65]), .ZN(n127) );
  XNOR2_X1 U369 ( .A(Key[66]), .B(Plaintext[66]), .ZN(n126) );
  XNOR2_X1 U370 ( .A(Key[67]), .B(Plaintext[67]), .ZN(n125) );
  XNOR2_X1 U371 ( .A(Key[68]), .B(Plaintext[68]), .ZN(n124) );
  XNOR2_X1 U372 ( .A(Key[69]), .B(Plaintext[69]), .ZN(n123) );
  XNOR2_X1 U373 ( .A(Key[70]), .B(Plaintext[70]), .ZN(n122) );
  XNOR2_X1 U374 ( .A(Key[71]), .B(Plaintext[71]), .ZN(n121) );
  XNOR2_X1 U375 ( .A(Key[72]), .B(Plaintext[72]), .ZN(n120) );
  XNOR2_X1 U376 ( .A(Key[73]), .B(Plaintext[73]), .ZN(n119) );
  XNOR2_X1 U377 ( .A(Key[74]), .B(Plaintext[74]), .ZN(n118) );
  XNOR2_X1 U378 ( .A(Key[76]), .B(Plaintext[76]), .ZN(n116) );
  XNOR2_X1 U379 ( .A(Key[77]), .B(Plaintext[77]), .ZN(n115) );
  XNOR2_X1 U380 ( .A(Key[78]), .B(Plaintext[78]), .ZN(n114) );
  XNOR2_X1 U381 ( .A(Key[79]), .B(Plaintext[79]), .ZN(n113) );
  XNOR2_X1 U382 ( .A(Key[80]), .B(Plaintext[80]), .ZN(n112) );
  XNOR2_X1 U383 ( .A(Key[81]), .B(Plaintext[81]), .ZN(n111) );
  XNOR2_X1 U384 ( .A(Key[82]), .B(Plaintext[82]), .ZN(n110) );
  XNOR2_X1 U385 ( .A(Key[83]), .B(Plaintext[83]), .ZN(n109) );
  XNOR2_X1 U386 ( .A(Key[84]), .B(Plaintext[84]), .ZN(n108) );
  XNOR2_X1 U387 ( .A(Key[85]), .B(Plaintext[85]), .ZN(n107) );
  XNOR2_X1 U388 ( .A(Key[87]), .B(Plaintext[87]), .ZN(n105) );
  XNOR2_X1 U389 ( .A(Key[88]), .B(Plaintext[88]), .ZN(n104) );
  XNOR2_X1 U390 ( .A(Key[89]), .B(Plaintext[89]), .ZN(n103) );
  XNOR2_X1 U391 ( .A(Key[90]), .B(Plaintext[90]), .ZN(n102) );
  XNOR2_X1 U392 ( .A(Key[91]), .B(Plaintext[91]), .ZN(n101) );
  XNOR2_X1 U393 ( .A(Key[92]), .B(Plaintext[92]), .ZN(n100) );
  XNOR2_X1 U394 ( .A(Key[93]), .B(Plaintext[93]), .ZN(n99) );
  XNOR2_X1 U395 ( .A(Key[94]), .B(Plaintext[94]), .ZN(n98) );
  XNOR2_X1 U396 ( .A(Key[95]), .B(Plaintext[95]), .ZN(n97) );
  XNOR2_X1 U397 ( .A(Key[96]), .B(Plaintext[96]), .ZN(n96) );
  XNOR2_X1 U398 ( .A(Key[97]), .B(Plaintext[97]), .ZN(n95) );
  XNOR2_X1 U399 ( .A(Key[98]), .B(Plaintext[98]), .ZN(n94) );
  XNOR2_X1 U400 ( .A(Key[99]), .B(Plaintext[99]), .ZN(n93) );
  XNOR2_X1 U401 ( .A(Key[100]), .B(Plaintext[100]), .ZN(n92) );
  XNOR2_X1 U402 ( .A(Key[101]), .B(Plaintext[101]), .ZN(n91) );
  XNOR2_X1 U403 ( .A(Key[102]), .B(Plaintext[102]), .ZN(n90) );
  XNOR2_X1 U404 ( .A(Key[103]), .B(Plaintext[103]), .ZN(n89) );
  XNOR2_X1 U405 ( .A(Key[104]), .B(Plaintext[104]), .ZN(n88) );
  XNOR2_X1 U406 ( .A(Key[105]), .B(Plaintext[105]), .ZN(n87) );
  XNOR2_X1 U407 ( .A(Key[106]), .B(Plaintext[106]), .ZN(n86) );
  XNOR2_X1 U408 ( .A(Key[107]), .B(Plaintext[107]), .ZN(n85) );
  XNOR2_X1 U409 ( .A(Key[108]), .B(Plaintext[108]), .ZN(n84) );
  XNOR2_X1 U410 ( .A(Key[109]), .B(Plaintext[109]), .ZN(n83) );
  XNOR2_X1 U411 ( .A(Key[110]), .B(Plaintext[110]), .ZN(n82) );
  XNOR2_X1 U412 ( .A(Key[111]), .B(Plaintext[111]), .ZN(n81) );
  XNOR2_X1 U413 ( .A(Key[112]), .B(Plaintext[112]), .ZN(n80) );
  XNOR2_X1 U414 ( .A(Key[113]), .B(Plaintext[113]), .ZN(n79) );
  XNOR2_X1 U415 ( .A(Key[114]), .B(Plaintext[114]), .ZN(n78) );
  XNOR2_X1 U416 ( .A(Key[115]), .B(Plaintext[115]), .ZN(n77) );
  XNOR2_X1 U417 ( .A(Key[116]), .B(Plaintext[116]), .ZN(n76) );
  XNOR2_X1 U418 ( .A(Key[117]), .B(Plaintext[117]), .ZN(n75) );
  XNOR2_X1 U419 ( .A(Key[118]), .B(Plaintext[118]), .ZN(n74) );
  XNOR2_X1 U420 ( .A(Key[119]), .B(Plaintext[119]), .ZN(n73) );
  XNOR2_X1 U421 ( .A(Key[120]), .B(Plaintext[120]), .ZN(n72) );
  XNOR2_X1 U422 ( .A(Key[121]), .B(Plaintext[121]), .ZN(n71) );
  XNOR2_X1 U423 ( .A(Key[124]), .B(Plaintext[124]), .ZN(n68) );
  XNOR2_X1 U424 ( .A(Key[125]), .B(Plaintext[125]), .ZN(n67) );
  XNOR2_X1 U425 ( .A(Key[126]), .B(Plaintext[126]), .ZN(n66) );
  XNOR2_X1 U426 ( .A(Key[127]), .B(Plaintext[127]), .ZN(n65) );
  XNOR2_X1 U427 ( .A(Key[128]), .B(Plaintext[128]), .ZN(n64) );
  XNOR2_X1 U428 ( .A(Key[129]), .B(Plaintext[129]), .ZN(n63) );
  XNOR2_X1 U429 ( .A(Key[130]), .B(Plaintext[130]), .ZN(n62) );
  XNOR2_X1 U430 ( .A(Key[131]), .B(Plaintext[131]), .ZN(n61) );
  XNOR2_X1 U431 ( .A(Key[132]), .B(Plaintext[132]), .ZN(n60) );
  XNOR2_X1 U432 ( .A(Key[133]), .B(Plaintext[133]), .ZN(n59) );
  XNOR2_X1 U433 ( .A(Key[134]), .B(Plaintext[134]), .ZN(n58) );
  XNOR2_X1 U434 ( .A(Key[135]), .B(Plaintext[135]), .ZN(n57) );
  XNOR2_X1 U435 ( .A(Key[136]), .B(Plaintext[136]), .ZN(n56) );
  XNOR2_X1 U436 ( .A(Key[137]), .B(Plaintext[137]), .ZN(n55) );
  XNOR2_X1 U437 ( .A(Key[138]), .B(Plaintext[138]), .ZN(n54) );
  XNOR2_X1 U438 ( .A(Key[139]), .B(Plaintext[139]), .ZN(n53) );
  XNOR2_X1 U439 ( .A(Key[140]), .B(Plaintext[140]), .ZN(n52) );
  XNOR2_X1 U440 ( .A(Key[141]), .B(Plaintext[141]), .ZN(n51) );
  XNOR2_X1 U441 ( .A(Key[142]), .B(Plaintext[142]), .ZN(n50) );
  XNOR2_X1 U442 ( .A(Key[143]), .B(Plaintext[143]), .ZN(n49) );
  XNOR2_X1 U443 ( .A(Key[144]), .B(Plaintext[144]), .ZN(n48) );
  XNOR2_X1 U444 ( .A(Key[145]), .B(Plaintext[145]), .ZN(n47) );
  XNOR2_X1 U445 ( .A(Key[146]), .B(Plaintext[146]), .ZN(n46) );
  XNOR2_X1 U446 ( .A(Key[147]), .B(Plaintext[147]), .ZN(n45) );
  XNOR2_X1 U447 ( .A(Key[148]), .B(Plaintext[148]), .ZN(n44) );
  XNOR2_X1 U448 ( .A(Key[149]), .B(Plaintext[149]), .ZN(n43) );
  XNOR2_X1 U449 ( .A(Key[150]), .B(Plaintext[150]), .ZN(n42) );
  XNOR2_X1 U450 ( .A(Key[151]), .B(Plaintext[151]), .ZN(n41) );
  XNOR2_X1 U451 ( .A(Key[152]), .B(Plaintext[152]), .ZN(n40) );
  XNOR2_X1 U452 ( .A(Key[153]), .B(Plaintext[153]), .ZN(n39) );
  XNOR2_X1 U453 ( .A(Key[154]), .B(Plaintext[154]), .ZN(n38) );
  XNOR2_X1 U454 ( .A(Key[155]), .B(Plaintext[155]), .ZN(n37) );
  XNOR2_X1 U455 ( .A(Key[156]), .B(Plaintext[156]), .ZN(n36) );
  XNOR2_X1 U456 ( .A(Key[157]), .B(Plaintext[157]), .ZN(n35) );
  XNOR2_X1 U457 ( .A(Key[158]), .B(Plaintext[158]), .ZN(n34) );
  XNOR2_X1 U458 ( .A(Key[160]), .B(Plaintext[160]), .ZN(n32) );
  XNOR2_X1 U459 ( .A(Key[161]), .B(Plaintext[161]), .ZN(n31) );
  XNOR2_X1 U460 ( .A(Key[162]), .B(Plaintext[162]), .ZN(n30) );
  XNOR2_X1 U461 ( .A(Key[163]), .B(Plaintext[163]), .ZN(n29) );
  XNOR2_X1 U462 ( .A(Key[164]), .B(Plaintext[164]), .ZN(n28) );
  XNOR2_X1 U463 ( .A(Key[165]), .B(Plaintext[165]), .ZN(n27) );
  XNOR2_X1 U464 ( .A(Key[166]), .B(Plaintext[166]), .ZN(n26) );
  XNOR2_X1 U465 ( .A(Key[167]), .B(Plaintext[167]), .ZN(n25) );
  XNOR2_X1 U466 ( .A(Key[168]), .B(Plaintext[168]), .ZN(n24) );
  XNOR2_X1 U467 ( .A(Key[169]), .B(Plaintext[169]), .ZN(n23) );
  XNOR2_X1 U468 ( .A(Key[170]), .B(Plaintext[170]), .ZN(n22) );
  XNOR2_X1 U469 ( .A(Key[171]), .B(Plaintext[171]), .ZN(n21) );
  XNOR2_X1 U470 ( .A(Key[172]), .B(Plaintext[172]), .ZN(n20) );
  XNOR2_X1 U471 ( .A(Key[173]), .B(Plaintext[173]), .ZN(n19) );
  XNOR2_X1 U472 ( .A(Key[174]), .B(Plaintext[174]), .ZN(n18) );
  XNOR2_X1 U473 ( .A(Key[175]), .B(Plaintext[175]), .ZN(n17) );
  XNOR2_X1 U474 ( .A(Key[176]), .B(Plaintext[176]), .ZN(n16) );
  XNOR2_X1 U475 ( .A(Key[177]), .B(Plaintext[177]), .ZN(n15) );
  XNOR2_X1 U476 ( .A(Key[178]), .B(Plaintext[178]), .ZN(n14) );
  XNOR2_X1 U477 ( .A(Key[179]), .B(Plaintext[179]), .ZN(n13) );
  XNOR2_X1 U478 ( .A(Key[180]), .B(Plaintext[180]), .ZN(n12) );
  XNOR2_X1 U479 ( .A(Key[181]), .B(Plaintext[181]), .ZN(n11) );
  XNOR2_X1 U480 ( .A(Key[182]), .B(Plaintext[182]), .ZN(n10) );
  XNOR2_X1 U481 ( .A(Key[184]), .B(Plaintext[184]), .ZN(n8) );
  XNOR2_X1 U482 ( .A(Key[185]), .B(Plaintext[185]), .ZN(n7) );
  XNOR2_X1 U483 ( .A(Key[186]), .B(Plaintext[186]), .ZN(n6) );
  XNOR2_X1 U484 ( .A(Key[187]), .B(Plaintext[187]), .ZN(n5) );
  XNOR2_X1 U485 ( .A(Key[189]), .B(Plaintext[189]), .ZN(n3) );
  XNOR2_X1 U486 ( .A(Key[190]), .B(Plaintext[190]), .ZN(n2) );
  INV_X1 U487 ( .A(n503), .ZN(n366) );
  INV_X1 U488 ( .A(n501), .ZN(n270) );
  INV_X1 U489 ( .A(n384), .ZN(n334) );
  INV_X1 U490 ( .A(n491), .ZN(n235) );
  INV_X1 U491 ( .A(n489), .ZN(n229) );
  INV_X1 U492 ( .A(n505), .ZN(n315) );
  INV_X1 U493 ( .A(n470), .ZN(n211) );
  INV_X1 U494 ( .A(Key[180]), .ZN(n203) );
  INV_X1 U495 ( .A(n498), .ZN(n196) );
  INV_X1 U496 ( .A(n494), .ZN(n279) );
  INV_X1 U497 ( .A(n378), .ZN(n277) );
  INV_X1 U498 ( .A(n499), .ZN(n367) );
  INV_X1 U499 ( .A(n402), .ZN(n261) );
  INV_X1 U500 ( .A(n448), .ZN(n347) );
  INV_X1 U501 ( .A(n464), .ZN(n341) );
  INV_X1 U503 ( .A(n502), .ZN(n303) );
  INV_X1 U504 ( .A(Key[150]), .ZN(n233) );
  INV_X1 U505 ( .A(n383), .ZN(n254) );
  INV_X1 U506 ( .A(n497), .ZN(n304) );
  INV_X1 U507 ( .A(n461), .ZN(n241) );
  INV_X1 U508 ( .A(n473), .ZN(n371) );
  INV_X1 U509 ( .A(n506), .ZN(n360) );
  INV_X1 U510 ( .A(n463), .ZN(n280) );
  INV_X1 U512 ( .A(n428), .ZN(n312) );
  INV_X1 U513 ( .A(n459), .ZN(n308) );
  INV_X1 U514 ( .A(Key[168]), .ZN(n215) );
  INV_X1 U515 ( .A(n507), .ZN(n236) );
  INV_X1 U517 ( .A(n401), .ZN(n204) );
  INV_X1 U518 ( .A(n424), .ZN(n283) );
  INV_X1 U519 ( .A(n405), .ZN(n210) );
  INV_X1 U520 ( .A(n452), .ZN(n359) );
  INV_X1 U521 ( .A(n500), .ZN(n316) );
  INV_X1 U522 ( .A(n509), .ZN(n269) );
  INV_X1 U524 ( .A(n447), .ZN(n353) );
  INV_X1 U525 ( .A(n446), .ZN(n274) );
  XNOR2_X1 U529 ( .A(\RI4[4][3] ), .B(n274), .ZN(Ciphertext[3]) );
  INV_X1 U547 ( .A(n469), .ZN(n409) );
  INV_X1 U555 ( .A(n468), .ZN(n410) );
  XNOR2_X1 U559 ( .A(\RI4[4][33] ), .B(n256), .ZN(Ciphertext[33]) );
  INV_X1 U560 ( .A(n407), .ZN(n411) );
  XNOR2_X1 U571 ( .A(\RI4[4][45] ), .B(n359), .ZN(Ciphertext[45]) );
  INV_X1 U577 ( .A(n482), .ZN(n412) );
  XNOR2_X1 U578 ( .A(\RI4[4][51] ), .B(n412), .ZN(Ciphertext[51]) );
  INV_X1 U590 ( .A(n474), .ZN(n413) );
  XNOR2_X1 U597 ( .A(\RI4[4][75] ), .B(n341), .ZN(Ciphertext[75]) );
  INV_X1 U598 ( .A(n408), .ZN(n414) );
  XNOR2_X1 U603 ( .A(\RI4[4][81] ), .B(n302), .ZN(Ciphertext[81]) );
  INV_X1 U625 ( .A(n513), .ZN(n415) );
  XNOR2_X1 U627 ( .A(\RI4[4][105] ), .B(n325), .ZN(Ciphertext[105]) );
  INV_X1 U630 ( .A(n512), .ZN(n416) );
  XNOR2_X1 U659 ( .A(\RI4[4][141] ), .B(n268), .ZN(Ciphertext[141]) );
  XNOR2_X1 U674 ( .A(\RI4[4][159] ), .B(n331), .ZN(Ciphertext[159]) );
  INV_X1 U685 ( .A(n471), .ZN(n417) );
  INV_X1 U695 ( .A(n457), .ZN(n418) );
  XNOR2_X1 U699 ( .A(\RI4[4][183] ), .B(n353), .ZN(Ciphertext[183]) );
  XNOR2_X1 U702 ( .A(\RI4[4][187] ), .B(n327), .ZN(Ciphertext[187]) );
  BUF_X2 \SB4_7/BUF_0  ( .A(\RI3[4][144] ), .Z(\SB4_7/i0[9] ) );
  BUF_X2 \SB4_27/BUF_0  ( .A(\RI3[4][24] ), .Z(\SB4_27/i0[9] ) );
  BUF_X2 \SB4_28/BUF_1  ( .A(\RI3[4][19] ), .Z(\SB4_28/i0[6] ) );
  BUF_X1 \SB1_1_11/BUF_1  ( .A(\RI1[1][121] ), .Z(\SB1_1_11/i1_7 ) );
  BUF_X2 \SB2_3_5/BUF_2  ( .A(\RI3[3][158] ), .Z(\SB2_3_5/i0_0 ) );
  BUF_X2 \SB2_0_2/BUF_3  ( .A(\RI3[0][177] ), .Z(\SB2_0_2/i0[10] ) );
  BUF_X2 \SB2_0_26/BUF_2  ( .A(\RI3[0][32] ), .Z(\SB2_0_26/i0_0 ) );
  BUF_X2 \SB4_25/BUF_1  ( .A(\RI3[4][37] ), .Z(\SB4_25/i0[6] ) );
  BUF_X2 \SB2_0_17/BUF_1  ( .A(\RI3[0][85] ), .Z(\SB2_0_17/i0[6] ) );
  BUF_X2 \SB2_0_11/BUF_3  ( .A(\RI3[0][123] ), .Z(\SB2_0_11/i0[10] ) );
  INV_X1 \SB1_2_12/INV_4  ( .A(\RI1[2][118] ), .ZN(\SB1_2_12/i0_4 ) );
  BUF_X2 \SB2_2_8/BUF_1  ( .A(\RI3[2][139] ), .Z(\SB2_2_8/i0[6] ) );
  BUF_X2 \SB2_2_27/BUF_1  ( .A(\RI3[2][25] ), .Z(\SB2_2_27/i0[6] ) );
  BUF_X2 \SB2_1_7/BUF_3  ( .A(\RI3[1][147] ), .Z(\SB2_1_7/i0[10] ) );
  BUF_X2 \SB2_1_24/BUF_1  ( .A(\RI3[1][43] ), .Z(\SB2_1_24/i0[6] ) );
  INV_X1 \SB1_0_20/INV_5  ( .A(n121), .ZN(\SB1_0_20/i0_3 ) );
  BUF_X2 \SB2_1_21/BUF_2  ( .A(\RI3[1][62] ), .Z(\SB2_1_21/i0_0 ) );
  BUF_X2 \SB4_13/BUF_1  ( .A(\RI3[4][109] ), .Z(\SB4_13/i0[6] ) );
  INV_X1 \SB3_9/INV_5  ( .A(\RI1[4][137] ), .ZN(\SB3_9/i0_3 ) );
  INV_X1 \SB2_1_6/INV_2  ( .A(\RI3[1][152] ), .ZN(\SB2_1_6/i1[9] ) );
  INV_X1 \SB3_10/INV_5  ( .A(\RI1[4][131] ), .ZN(\SB3_10/i0_3 ) );
  BUF_X2 \SB2_1_6/BUF_2  ( .A(\RI3[1][152] ), .Z(\SB2_1_6/i0_0 ) );
  BUF_X2 \SB2_0_29/BUF_3  ( .A(\RI3[0][15] ), .Z(\SB2_0_29/i0[10] ) );
  INV_X1 \SB1_3_3/INV_4  ( .A(\RI1[3][172] ), .ZN(\SB1_3_3/i0_4 ) );
  BUF_X2 \SB2_0_15/BUF_3  ( .A(\RI3[0][99] ), .Z(\SB2_0_15/i0[10] ) );
  BUF_X2 \SB4_16/BUF_1  ( .A(\RI3[4][91] ), .Z(\SB4_16/i0[6] ) );
  BUF_X2 \SB3_22/BUF_2  ( .A(\RI1[4][56] ), .Z(\SB3_22/i1[9] ) );
  BUF_X2 \SB2_1_11/BUF_3  ( .A(\RI3[1][123] ), .Z(\SB2_1_11/i0[10] ) );
  BUF_X1 \SB1_3_17/BUF_1  ( .A(\RI1[3][85] ), .Z(\SB1_3_17/i1_7 ) );
  INV_X1 \SB1_3_18/INV_4  ( .A(\RI1[3][82] ), .ZN(\SB1_3_18/i0_4 ) );
  BUF_X2 \SB4_20/BUF_1  ( .A(\RI3[4][67] ), .Z(\SB4_20/i0[6] ) );
  INV_X1 \SB2_3_13/INV_2  ( .A(\RI3[3][110] ), .ZN(\SB2_3_13/i1[9] ) );
  BUF_X2 \SB1_3_6/BUF_3  ( .A(\RI1[3][153] ), .Z(\SB1_3_6/i0[8] ) );
  BUF_X2 \SB2_1_16/BUF_1  ( .A(\RI3[1][91] ), .Z(\SB2_1_16/i0[6] ) );
  BUF_X1 \SB1_2_20/BUF_1  ( .A(\RI1[2][67] ), .Z(\SB1_2_20/i1_7 ) );
  BUF_X2 \SB4_1/BUF_1  ( .A(\RI3[4][181] ), .Z(\SB4_1/i0[6] ) );
  INV_X1 \SB1_0_4/INV_5  ( .A(n25), .ZN(\SB1_0_4/i0_3 ) );
  INV_X1 \SB1_3_4/INV_4  ( .A(\RI1[3][166] ), .ZN(\SB1_3_4/i0_4 ) );
  BUF_X2 \SB2_0_7/BUF_3  ( .A(\RI3[0][147] ), .Z(\SB2_0_7/i0[10] ) );
  BUF_X2 \SB2_2_1/BUF_2  ( .A(\RI3[2][182] ), .Z(\SB2_2_1/i0_0 ) );
  BUF_X2 \SB2_3_2/BUF_2  ( .A(\RI3[3][176] ), .Z(\SB2_3_2/i0_0 ) );
  BUF_X2 \SB2_1_15/BUF_2  ( .A(\RI3[1][98] ), .Z(\SB2_1_15/i0_0 ) );
  INV_X1 \SB2_3_31/INV_2  ( .A(\RI3[3][2] ), .ZN(\SB2_3_31/i1[9] ) );
  INV_X1 \SB2_1_15/INV_2  ( .A(\RI3[1][98] ), .ZN(\SB2_1_15/i1[9] ) );
  BUF_X2 \SB4_8/BUF_0  ( .A(\RI3[4][138] ), .Z(\SB4_8/i0[9] ) );
  BUF_X2 \SB4_22/BUF_1  ( .A(\RI3[4][55] ), .Z(\SB4_22/i0[6] ) );
  BUF_X2 \SB2_1_19/BUF_3  ( .A(\RI3[1][75] ), .Z(\SB2_1_19/i0[10] ) );
  BUF_X2 \SB4_30/BUF_0  ( .A(\RI3[4][6] ), .Z(\SB4_30/i0[9] ) );
  BUF_X1 \SB1_0_0/BUF_1  ( .A(n5), .Z(\SB1_0_0/i1_7 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_76  ( .A(\RI5[2][76] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[76] ) );
  BUF_X2 \SB4_6/BUF_0  ( .A(\RI3[4][150] ), .Z(\SB4_6/i0[9] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_1/BUF_33  ( .A(\RI5[1][33] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[33] ) );
  BUF_X2 \SB2_1_28/BUF_2  ( .A(\RI3[1][20] ), .Z(\SB2_1_28/i0_0 ) );
  BUF_X2 \SB2_2_31/BUF_2  ( .A(\RI3[2][2] ), .Z(\SB2_2_31/i0_0 ) );
  BUF_X2 \SB2_1_12/BUF_3  ( .A(\RI3[1][117] ), .Z(\SB2_1_12/i0[10] ) );
  INV_X1 \SB1_3_0/INV_4  ( .A(\RI1[3][190] ), .ZN(\SB1_3_0/i0_4 ) );
  BUF_X2 \SB3_9/BUF_2  ( .A(\RI1[4][134] ), .Z(\SB3_9/i1[9] ) );
  INV_X1 \SB1_1_26/INV_0  ( .A(\RI1[1][30] ), .ZN(\SB1_1_26/i0[9] ) );
  BUF_X2 \SB2_0_4/BUF_5  ( .A(\RI3[0][167] ), .Z(\SB2_0_4/i0_3 ) );
  BUF_X2 \SB4_3/BUF_0  ( .A(\RI3[4][168] ), .Z(\SB4_3/i0[9] ) );
  BUF_X2 \SB4_3/BUF_1  ( .A(\RI3[4][169] ), .Z(\SB4_3/i0[6] ) );
  INV_X1 \SB1_1_27/INV_4  ( .A(\RI1[1][28] ), .ZN(\SB1_1_27/i0_4 ) );
  BUF_X2 \SB4_27/BUF_1  ( .A(\RI3[4][25] ), .Z(\SB4_27/i0[6] ) );
  BUF_X1 \SB1_2_9/BUF_1  ( .A(\RI1[2][133] ), .Z(\SB1_2_9/i1_7 ) );
  BUF_X2 \SB3_10/BUF_2  ( .A(\RI1[4][128] ), .Z(\SB3_10/i1[9] ) );
  BUF_X2 \SB2_1_21/BUF_1  ( .A(\RI3[1][61] ), .Z(\SB2_1_21/i0[6] ) );
  BUF_X1 \SB1_3_29/BUF_1  ( .A(\RI1[3][13] ), .Z(\SB1_3_29/i1_7 ) );
  BUF_X2 \SB4_21/BUF_0  ( .A(\RI3[4][60] ), .Z(\SB4_21/i0[9] ) );
  BUF_X2 \SB2_3_28/BUF_0  ( .A(\RI3[3][18] ), .Z(\SB2_3_28/i0[9] ) );
  BUF_X2 \SB2_0_18/BUF_3  ( .A(\RI3[0][81] ), .Z(\SB2_0_18/i0[10] ) );
  INV_X1 \SB1_2_6/INV_4  ( .A(\RI1[2][154] ), .ZN(\SB1_2_6/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_28  ( .A(\RI5[1][28] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[28] ) );
  BUF_X2 \SB2_2_21/BUF_2  ( .A(\RI3[2][62] ), .Z(\SB2_2_21/i0_0 ) );
  INV_X1 \SB3_5/INV_5  ( .A(\RI1[4][161] ), .ZN(\SB3_5/i0_3 ) );
  BUF_X1 \SB1_2_29/BUF_1  ( .A(\RI1[2][13] ), .Z(\SB1_2_29/i1_7 ) );
  BUF_X2 \SB2_2_30/BUF_0  ( .A(\RI3[2][6] ), .Z(\SB2_2_30/i0[9] ) );
  BUF_X2 \SB2_0_30/BUF_2  ( .A(\RI3[0][8] ), .Z(\SB2_0_30/i0_0 ) );
  BUF_X2 \SB2_2_4/BUF_2  ( .A(\RI3[2][164] ), .Z(\SB2_2_4/i0_0 ) );
  BUF_X2 \SB2_2_23/BUF_2  ( .A(\RI3[2][50] ), .Z(\SB2_2_23/i0_0 ) );
  BUF_X2 \SB2_1_9/BUF_0  ( .A(\RI3[1][132] ), .Z(\SB2_1_9/i0[9] ) );
  BUF_X2 \SB2_1_4/BUF_1  ( .A(\RI3[1][163] ), .Z(\SB2_1_4/i0[6] ) );
  BUF_X2 \SB2_1_18/BUF_2  ( .A(\RI3[1][80] ), .Z(\SB2_1_18/i0_0 ) );
  BUF_X2 \SB2_1_22/BUF_3  ( .A(\RI3[1][57] ), .Z(\SB2_1_22/i0[10] ) );
  BUF_X2 \SB2_1_25/BUF_2  ( .A(\RI3[1][38] ), .Z(\SB2_1_25/i0_0 ) );
  INV_X1 \SB1_1_16/INV_4  ( .A(\RI1[1][94] ), .ZN(\SB1_1_16/i0_4 ) );
  BUF_X1 \SB1_3_1/BUF_1  ( .A(\RI1[3][181] ), .Z(\SB1_3_1/i1_7 ) );
  INV_X1 \SB1_2_2/INV_4  ( .A(\RI1[2][178] ), .ZN(\SB1_2_2/i0_4 ) );
  BUF_X2 \SB2_0_10/BUF_2  ( .A(\RI3[0][128] ), .Z(\SB2_0_10/i0_0 ) );
  BUF_X2 \SB2_1_27/BUF_2  ( .A(\RI3[1][26] ), .Z(\SB2_1_27/i0_0 ) );
  INV_X1 \SB2_0_10/INV_2  ( .A(\RI3[0][128] ), .ZN(\SB2_0_10/i1[9] ) );
  BUF_X2 \SB2_0_10/BUF_3  ( .A(\RI3[0][129] ), .Z(\SB2_0_10/i0[10] ) );
  BUF_X2 \SB2_0_25/BUF_0  ( .A(\RI3[0][36] ), .Z(\SB2_0_25/i0[9] ) );
  BUF_X2 \SB2_1_11/BUF_2  ( .A(\RI3[1][122] ), .Z(\SB2_1_11/i0_0 ) );
  BUF_X2 \SB4_19/BUF_1  ( .A(\RI3[4][73] ), .Z(\SB4_19/i0[6] ) );
  BUF_X2 \SB4_18/BUF_0  ( .A(\RI3[4][78] ), .Z(\SB4_18/i0[9] ) );
  INV_X1 \SB2_3_7/INV_2  ( .A(\RI3[3][146] ), .ZN(\SB2_3_7/i1[9] ) );
  INV_X1 \SB1_1_13/INV_0  ( .A(\RI1[1][108] ), .ZN(\SB1_1_13/i0[9] ) );
  BUF_X2 \SB2_1_9/BUF_1  ( .A(\RI3[1][133] ), .Z(\SB2_1_9/i0[6] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_82  ( .A(\RI5[0][82] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[82] ) );
  BUF_X1 \SB1_1_9/BUF_1  ( .A(\RI1[1][133] ), .Z(\SB1_1_9/i1_7 ) );
  BUF_X1 \SB1_3_9/BUF_1  ( .A(\RI1[3][133] ), .Z(\SB1_3_9/i1_7 ) );
  BUF_X1 \SB1_3_16/BUF_1  ( .A(\RI1[3][91] ), .Z(\SB1_3_16/i1_7 ) );
  BUF_X2 \SB2_2_16/BUF_2  ( .A(\RI3[2][92] ), .Z(\SB2_2_16/i0_0 ) );
  BUF_X2 \SB2_1_16/BUF_2  ( .A(\RI3[1][92] ), .Z(\SB2_1_16/i0_0 ) );
  BUF_X1 \SB1_2_21/BUF_1  ( .A(\RI1[2][61] ), .Z(\SB1_2_21/i1_7 ) );
  INV_X1 \SB3_26/INV_5  ( .A(\RI1[4][35] ), .ZN(\SB3_26/i0_3 ) );
  BUF_X2 \SB2_0_23/BUF_1  ( .A(\RI3[0][49] ), .Z(\SB2_0_23/i0[6] ) );
  BUF_X2 \SB2_1_23/BUF_2  ( .A(\RI3[1][50] ), .Z(\SB2_1_23/i0_0 ) );
  BUF_X2 \SB4_21/BUF_1  ( .A(\RI3[4][61] ), .Z(\SB4_21/i0[6] ) );
  BUF_X2 \SB2_0_25/BUF_2  ( .A(\RI3[0][38] ), .Z(\SB2_0_25/i0_0 ) );
  INV_X1 \SB1_0_27/INV_5  ( .A(n163), .ZN(\SB1_0_27/i0_3 ) );
  INV_X1 \SB1_0_14/INV_5  ( .A(n85), .ZN(\SB1_0_14/i0_3 ) );
  INV_X1 \SB1_1_9/INV_3  ( .A(\RI1[1][135] ), .ZN(\SB1_1_9/i0[10] ) );
  BUF_X1 \SB1_3_10/BUF_1  ( .A(\RI1[3][127] ), .Z(\SB1_3_10/i1_7 ) );
  BUF_X2 \SB2_3_5/BUF_1  ( .A(\RI3[3][157] ), .Z(\SB2_3_5/i0[6] ) );
  BUF_X2 \SB2_0_10/BUF_4  ( .A(\RI3[0][130] ), .Z(\SB2_0_10/i0_4 ) );
  BUF_X2 \SB2_0_13/BUF_2  ( .A(\RI3[0][110] ), .Z(\SB2_0_13/i0_0 ) );
  INV_X1 \SB1_0_19/INV_5  ( .A(n115), .ZN(\SB1_0_19/i0_3 ) );
  BUF_X2 \SB2_1_10/BUF_2  ( .A(\RI3[1][128] ), .Z(\SB2_1_10/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_172  ( .A(\RI5[2][172] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[172] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_112  ( .A(\RI5[1][112] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[112] ) );
  BUF_X1 \SB1_0_28/BUF_1  ( .A(n173), .Z(\SB1_0_28/i1_7 ) );
  BUF_X2 \SB2_2_30/BUF_1  ( .A(\RI3[2][7] ), .Z(\SB2_2_30/i0[6] ) );
  BUF_X1 \SB1_2_1/BUF_1  ( .A(\RI1[2][181] ), .Z(\SB1_2_1/i1_7 ) );
  INV_X1 \SB3_22/INV_5  ( .A(\RI1[4][59] ), .ZN(\SB3_22/i0_3 ) );
  BUF_X2 \SB4_8/BUF_1  ( .A(\RI3[4][139] ), .Z(\SB4_8/i0[6] ) );
  BUF_X1 \SB1_2_30/BUF_1  ( .A(\RI1[2][7] ), .Z(\SB1_2_30/i1_7 ) );
  BUF_X2 \SB4_25/BUF_0  ( .A(\RI3[4][36] ), .Z(\SB4_25/i0[9] ) );
  BUF_X2 \SB4_31/BUF_1  ( .A(\RI3[4][1] ), .Z(\SB4_31/i0[6] ) );
  BUF_X2 \SB4_4/BUF_1  ( .A(\RI3[4][163] ), .Z(\SB4_4/i0[6] ) );
  BUF_X2 \SB4_6/BUF_1  ( .A(\RI3[4][151] ), .Z(\SB4_6/i0[6] ) );
  BUF_X1 \SB1_2_22/BUF_1  ( .A(\RI1[2][55] ), .Z(\SB1_2_22/i1_7 ) );
  BUF_X2 \SB3_20/BUF_2  ( .A(\RI1[4][68] ), .Z(\SB3_20/i1[9] ) );
  BUF_X2 \SB3_14/BUF_3  ( .A(\RI1[4][105] ), .Z(\SB3_14/i0[8] ) );
  BUF_X1 \SB1_2_18/BUF_1  ( .A(\RI1[2][79] ), .Z(\SB1_2_18/i1_7 ) );
  BUF_X1 \SB1_2_25/BUF_1  ( .A(\RI1[2][37] ), .Z(\SB1_2_25/i1_7 ) );
  INV_X1 \SB1_0_5/INV_2  ( .A(n34), .ZN(\SB1_0_5/i0_0 ) );
  BUF_X2 \SB2_3_0/BUF_2  ( .A(\RI3[3][188] ), .Z(\SB2_3_0/i0_0 ) );
  BUF_X1 \SB1_2_14/BUF_1  ( .A(\RI1[2][103] ), .Z(\SB1_2_14/i1_7 ) );
  BUF_X2 \SB2_3_24/BUF_2  ( .A(\RI3[3][44] ), .Z(\SB2_3_24/i0_0 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_160  ( .A(\RI5[1][160] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[160] ) );
  BUF_X2 \SB2_2_18/BUF_1  ( .A(\RI3[2][79] ), .Z(\SB2_2_18/i0[6] ) );
  BUF_X2 \SB4_10/BUF_0  ( .A(\RI3[4][126] ), .Z(\SB4_10/i0[9] ) );
  BUF_X1 \SB1_1_30/BUF_1  ( .A(\RI1[1][7] ), .Z(\SB1_1_30/i1_7 ) );
  BUF_X2 \SB2_3_14/BUF_0  ( .A(\RI3[3][102] ), .Z(\SB2_3_14/i0[9] ) );
  BUF_X1 \SB1_1_2/BUF_1  ( .A(\RI1[1][175] ), .Z(\SB1_1_2/i1_7 ) );
  BUF_X1 \SB1_3_2/BUF_1  ( .A(\RI1[3][175] ), .Z(\SB1_3_2/i1_7 ) );
  BUF_X2 \SB2_3_27/BUF_2  ( .A(\RI3[3][26] ), .Z(\SB2_3_27/i0_0 ) );
  BUF_X2 \SB2_0_12/BUF_1  ( .A(\RI3[0][115] ), .Z(\SB2_0_12/i0[6] ) );
  BUF_X1 \SB3_6/BUF_0  ( .A(\RI1[4][150] ), .Z(\SB3_6/i3[0] ) );
  INV_X1 \SB1_3_18/INV_0  ( .A(\RI1[3][78] ), .ZN(\SB1_3_18/i0[9] ) );
  BUF_X2 \SB4_30/BUF_1  ( .A(\RI3[4][7] ), .Z(\SB4_30/i0[6] ) );
  BUF_X2 \SB2_3_26/BUF_0  ( .A(\RI3[3][30] ), .Z(\SB2_3_26/i0[9] ) );
  INV_X1 \SB3_2/INV_4  ( .A(\RI1[4][178] ), .ZN(\SB3_2/i0_4 ) );
  BUF_X1 \SB1_2_24/BUF_1  ( .A(\RI1[2][43] ), .Z(\SB1_2_24/i1_7 ) );
  BUF_X2 \SB2_0_29/BUF_0  ( .A(\RI3[0][12] ), .Z(\SB2_0_29/i0[9] ) );
  BUF_X1 \SB1_2_31/BUF_1  ( .A(\RI1[2][1] ), .Z(\SB1_2_31/i1_7 ) );
  INV_X1 \SB1_0_2/INV_5  ( .A(n13), .ZN(\SB1_0_2/i0_3 ) );
  BUF_X2 \SB2_3_12/BUF_2  ( .A(\RI3[3][116] ), .Z(\SB2_3_12/i0_0 ) );
  INV_X1 \SB1_1_8/INV_3  ( .A(\RI1[1][141] ), .ZN(\SB1_1_8/i0[10] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_44_0  ( .A(Key[124]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[44] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_107_0  ( .A(Key[122]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[107] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_0/BUF_40_0  ( .A(Key[93]), .Z(
        \MC_ARK_ARC_1_0/buf_keyinput[40] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_106_0  ( .A(Key[50]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[106] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_179_0  ( .A(Key[163]), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[179] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_94_0  ( .A(Key[79]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[94] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_0/BUF_11_0  ( .A(Key[82]), .Z(
        \MC_ARK_ARC_1_0/buf_keyinput[11] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_0/BUF_95_0  ( .A(Key[94]), .Z(
        \MC_ARK_ARC_1_0/buf_keyinput[95] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_1/BUF_107_0  ( .A(Key[99]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[107] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_143_0  ( .A(Key[182]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[143] ) );
  BUF_X1 \SB1_0_27/BUF_2  ( .A(n166), .Z(\SB1_0_27/i1[9] ) );
  BUF_X1 \SB1_0_11/BUF_3  ( .A(n69), .Z(\SB1_0_11/i0[8] ) );
  CLKBUF_X1 \SB1_0_18/BUF_4  ( .A(n110), .Z(\SB1_0_18/i0[7] ) );
  INV_X1 \SB1_0_6/INV_4  ( .A(n38), .ZN(\SB1_0_6/i0_4 ) );
  BUF_X1 \SB1_0_29/BUF_2  ( .A(n178), .Z(\SB1_0_29/i1[9] ) );
  BUF_X1 \SB1_0_21/BUF_2  ( .A(n130), .Z(\SB1_0_21/i1[9] ) );
  INV_X1 \SB1_0_5/INV_0  ( .A(n36), .ZN(\SB1_0_5/i0[9] ) );
  BUF_X1 \SB1_0_11/BUF_2  ( .A(n70), .Z(\SB1_0_11/i1[9] ) );
  INV_X1 \SB1_0_28/INV_3  ( .A(n171), .ZN(\SB1_0_28/i0[10] ) );
  CLKBUF_X1 \SB1_0_5/BUF_0  ( .A(n36), .Z(\SB1_0_5/i3[0] ) );
  INV_X1 \SB1_0_5/INV_3  ( .A(n33), .ZN(\SB1_0_5/i0[10] ) );
  BUF_X1 \SB1_0_8/BUF_3  ( .A(n51), .Z(\SB1_0_8/i0[8] ) );
  CLKBUF_X1 \SB1_0_16/BUF_4  ( .A(n98), .Z(\SB1_0_16/i0[7] ) );
  BUF_X1 \SB1_0_2/BUF_2  ( .A(n16), .Z(\SB1_0_2/i1[9] ) );
  CLKBUF_X1 \SB1_0_1/BUF_0  ( .A(n12), .Z(\SB1_0_1/i3[0] ) );
  BUF_X1 \SB1_0_4/BUF_2  ( .A(n28), .Z(\SB1_0_4/i1[9] ) );
  BUF_X1 \SB1_0_18/BUF_1  ( .A(n113), .Z(\SB1_0_18/i1_7 ) );
  INV_X1 \SB1_0_1/INV_3  ( .A(n9), .ZN(\SB1_0_1/i0[10] ) );
  BUF_X1 \SB1_0_3/BUF_2  ( .A(n22), .Z(\SB1_0_3/i1[9] ) );
  BUF_X1 \SB1_0_1/BUF_3  ( .A(n9), .Z(\SB1_0_1/i0[8] ) );
  INV_X1 \SB1_0_1/INV_4  ( .A(n8), .ZN(\SB1_0_1/i0_4 ) );
  BUF_X1 \SB1_0_15/BUF_3  ( .A(n93), .Z(\SB1_0_15/i0[8] ) );
  BUF_X1 \SB1_0_8/BUF_2  ( .A(n52), .Z(\SB1_0_8/i1[9] ) );
  BUF_X1 \SB1_0_9/BUF_3  ( .A(n57), .Z(\SB1_0_9/i0[8] ) );
  BUF_X1 \SB2_0_16/BUF_1  ( .A(\RI3[0][91] ), .Z(\SB2_0_16/i0[6] ) );
  BUF_X2 \SB2_0_26/BUF_5  ( .A(\RI3[0][35] ), .Z(\SB2_0_26/i0_3 ) );
  BUF_X1 \SB2_0_22/BUF_1  ( .A(\RI3[0][55] ), .Z(\SB2_0_22/i0[6] ) );
  BUF_X2 \SB2_0_19/BUF_5  ( .A(\RI3[0][77] ), .Z(\SB2_0_19/i0_3 ) );
  BUF_X2 \SB2_0_19/BUF_4  ( .A(\RI3[0][76] ), .Z(\SB2_0_19/i0_4 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_54  ( .A(\RI5[0][54] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[54] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_132  ( .A(\RI5[0][132] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[132] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_121  ( .A(\RI5[0][121] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[121] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_120  ( .A(\RI5[0][120] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[120] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_14  ( .A(\RI5[0][14] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[14] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_31  ( .A(\RI5[0][31] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[31] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_102  ( .A(\RI5[0][102] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[102] ) );
  INV_X1 \SB1_1_18/INV_0  ( .A(\RI1[1][78] ), .ZN(\SB1_1_18/i0[9] ) );
  BUF_X1 \SB1_1_6/BUF_3  ( .A(\RI1[1][153] ), .Z(\SB1_1_6/i0[8] ) );
  CLKBUF_X1 \SB1_1_16/BUF_4  ( .A(\RI1[1][94] ), .Z(\SB1_1_16/i0[7] ) );
  INV_X1 \SB1_1_30/INV_0  ( .A(\RI1[1][6] ), .ZN(\SB1_1_30/i0[9] ) );
  INV_X1 \SB1_1_21/INV_0  ( .A(\RI1[1][60] ), .ZN(\SB1_1_21/i0[9] ) );
  INV_X1 \SB1_1_31/INV_0  ( .A(\RI1[1][0] ), .ZN(\SB1_1_31/i0[9] ) );
  BUF_X1 \SB1_1_23/BUF_3  ( .A(\RI1[1][51] ), .Z(\SB1_1_23/i0[8] ) );
  INV_X1 \SB1_1_11/INV_0  ( .A(\RI1[1][120] ), .ZN(\SB1_1_11/i0[9] ) );
  INV_X1 \SB1_1_8/INV_0  ( .A(\RI1[1][138] ), .ZN(\SB1_1_8/i0[9] ) );
  CLKBUF_X1 \SB1_1_28/BUF_4  ( .A(\RI1[1][22] ), .Z(\SB1_1_28/i0[7] ) );
  INV_X1 \SB1_1_3/INV_0  ( .A(\RI1[1][168] ), .ZN(\SB1_1_3/i0[9] ) );
  INV_X1 \SB1_1_14/INV_0  ( .A(\RI1[1][102] ), .ZN(\SB1_1_14/i0[9] ) );
  BUF_X2 \SB2_1_1/BUF_2  ( .A(\RI3[1][182] ), .Z(\SB2_1_1/i0_0 ) );
  BUF_X1 \SB2_1_11/BUF_0  ( .A(\RI3[1][120] ), .Z(\SB2_1_11/i0[9] ) );
  BUF_X2 \SB2_1_17/BUF_3  ( .A(\RI3[1][87] ), .Z(\SB2_1_17/i0[10] ) );
  BUF_X1 \SB2_1_30/BUF_1  ( .A(\RI3[1][7] ), .Z(\SB2_1_30/i0[6] ) );
  BUF_X1 \SB2_1_12/BUF_0  ( .A(\RI3[1][114] ), .Z(\SB2_1_12/i0[9] ) );
  BUF_X1 \SB2_1_12/BUF_1  ( .A(\RI3[1][115] ), .Z(\SB2_1_12/i0[6] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_30  ( .A(\RI5[1][30] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[30] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_175  ( .A(\RI5[1][175] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[175] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_67  ( .A(\RI5[1][67] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[67] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_169  ( .A(\RI5[1][169] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[169] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_108  ( .A(\RI5[1][108] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[108] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_42  ( .A(\RI5[1][42] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[42] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_184  ( .A(\RI5[1][184] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[184] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_186  ( .A(\RI5[1][186] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[186] ) );
  CLKBUF_X1 \SB1_2_0/BUF_4  ( .A(\RI1[2][190] ), .Z(\SB1_2_0/i0[7] ) );
  INV_X1 \SB1_2_31/INV_1  ( .A(\RI1[2][1] ), .ZN(\SB1_2_31/i0[6] ) );
  CLKBUF_X1 \SB1_2_13/BUF_4  ( .A(\RI1[2][112] ), .Z(\SB1_2_13/i0[7] ) );
  CLKBUF_X1 \SB1_2_7/BUF_4  ( .A(\RI1[2][148] ), .Z(\SB1_2_7/i0[7] ) );
  CLKBUF_X1 \SB1_2_28/BUF_4  ( .A(\RI1[2][22] ), .Z(\SB1_2_28/i0[7] ) );
  CLKBUF_X1 \SB1_2_11/BUF_4  ( .A(\RI1[2][124] ), .Z(\SB1_2_11/i0[7] ) );
  INV_X1 \SB1_2_27/INV_0  ( .A(\RI1[2][24] ), .ZN(\SB1_2_27/i0[9] ) );
  CLKBUF_X1 \SB1_2_12/BUF_4  ( .A(\RI1[2][118] ), .Z(\SB1_2_12/i0[7] ) );
  CLKBUF_X1 \SB1_2_22/BUF_4  ( .A(\RI1[2][58] ), .Z(\SB1_2_22/i0[7] ) );
  CLKBUF_X1 \SB1_2_19/BUF_4  ( .A(\RI1[2][76] ), .Z(\SB1_2_19/i0[7] ) );
  CLKBUF_X1 \SB1_2_25/BUF_4  ( .A(\RI1[2][40] ), .Z(\SB1_2_25/i0[7] ) );
  INV_X1 \SB1_2_24/INV_0  ( .A(\RI1[2][42] ), .ZN(\SB1_2_24/i0[9] ) );
  INV_X1 \SB1_2_30/INV_0  ( .A(\RI1[2][6] ), .ZN(\SB1_2_30/i0[9] ) );
  CLKBUF_X1 \SB1_2_10/BUF_4  ( .A(\RI1[2][130] ), .Z(\SB1_2_10/i0[7] ) );
  BUF_X1 \SB1_2_31/BUF_3  ( .A(\RI1[2][3] ), .Z(\SB1_2_31/i0[8] ) );
  CLKBUF_X1 \SB1_2_24/BUF_4  ( .A(\RI1[2][46] ), .Z(\SB1_2_24/i0[7] ) );
  CLKBUF_X1 \SB1_2_30/BUF_4  ( .A(\RI1[2][10] ), .Z(\SB1_2_30/i0[7] ) );
  INV_X1 \SB1_2_2/INV_0  ( .A(\RI1[2][174] ), .ZN(\SB1_2_2/i0[9] ) );
  INV_X1 \SB1_2_12/INV_0  ( .A(\RI1[2][114] ), .ZN(\SB1_2_12/i0[9] ) );
  BUF_X1 \SB2_2_14/BUF_0  ( .A(\RI3[2][102] ), .Z(\SB2_2_14/i0[9] ) );
  BUF_X1 \SB2_2_25/BUF_0  ( .A(\RI3[2][36] ), .Z(\SB2_2_25/i0[9] ) );
  BUF_X1 \SB2_2_6/BUF_0  ( .A(\RI3[2][150] ), .Z(\SB2_2_6/i0[9] ) );
  BUF_X2 \SB2_2_6/BUF_5  ( .A(\RI3[2][155] ), .Z(\SB2_2_6/i0_3 ) );
  BUF_X1 \SB2_2_9/BUF_0  ( .A(\RI3[2][132] ), .Z(\SB2_2_9/i0[9] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_163  ( .A(\RI5[2][163] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[163] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_144  ( .A(\RI5[2][144] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[144] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_132  ( .A(\RI5[2][132] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[132] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_72  ( .A(\RI5[2][72] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[72] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_0  ( .A(\RI5[2][0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[0] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_168  ( .A(\RI5[2][168] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[168] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_162  ( .A(\RI5[2][162] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[162] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_48  ( .A(\RI5[2][48] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[48] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_79  ( .A(\RI5[2][79] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[79] ) );
  CLKBUF_X1 \SB1_3_16/BUF_4  ( .A(\RI1[3][94] ), .Z(\SB1_3_16/i0[7] ) );
  BUF_X1 \SB1_3_5/BUF_1  ( .A(\RI1[3][157] ), .Z(\SB1_3_5/i1_7 ) );
  BUF_X1 \SB1_3_30/BUF_3  ( .A(\RI1[3][9] ), .Z(\SB1_3_30/i0[8] ) );
  INV_X1 \SB1_3_10/INV_0  ( .A(\RI1[3][126] ), .ZN(\SB1_3_10/i0[9] ) );
  INV_X1 \SB1_3_15/INV_0  ( .A(\RI1[3][96] ), .ZN(\SB1_3_15/i0[9] ) );
  CLKBUF_X1 \SB1_3_3/BUF_4  ( .A(\RI1[3][172] ), .Z(\SB1_3_3/i0[7] ) );
  INV_X1 \SB1_3_30/INV_0  ( .A(\RI1[3][6] ), .ZN(\SB1_3_30/i0[9] ) );
  CLKBUF_X1 \SB1_3_13/BUF_4  ( .A(\RI1[3][112] ), .Z(\SB1_3_13/i0[7] ) );
  CLKBUF_X1 \SB1_3_11/BUF_4  ( .A(\RI1[3][124] ), .Z(\SB1_3_11/i0[7] ) );
  INV_X1 \SB2_3_17/INV_2  ( .A(\RI3[3][86] ), .ZN(\SB2_3_17/i1[9] ) );
  BUF_X1 \SB2_3_7/BUF_0  ( .A(\RI3[3][144] ), .Z(\SB2_3_7/i0[9] ) );
  CLKBUF_X1 \SB3_17/BUF_4  ( .A(\RI1[4][88] ), .Z(\SB3_17/i0[7] ) );
  BUF_X1 \SB3_11/BUF_2  ( .A(\RI1[4][122] ), .Z(\SB3_11/i1[9] ) );
  CLKBUF_X1 \SB3_28/BUF_4  ( .A(\RI1[4][22] ), .Z(\SB3_28/i0[7] ) );
  CLKBUF_X1 \SB3_15/BUF_4  ( .A(\RI1[4][100] ), .Z(\SB3_15/i0[7] ) );
  BUF_X1 \SB3_4/BUF_2  ( .A(\RI1[4][164] ), .Z(\SB3_4/i1[9] ) );
  CLKBUF_X1 \SB3_0/BUF_4  ( .A(\RI1[4][190] ), .Z(\SB3_0/i0[7] ) );
  BUF_X1 \SB3_2/BUF_3  ( .A(\RI1[4][177] ), .Z(\SB3_2/i0[8] ) );
  BUF_X1 \SB3_31/BUF_3  ( .A(\RI1[4][3] ), .Z(\SB3_31/i0[8] ) );
  CLKBUF_X1 \SB3_31/BUF_4  ( .A(\RI1[4][4] ), .Z(\SB3_31/i0[7] ) );
  CLKBUF_X1 \SB3_30/BUF_4  ( .A(\RI1[4][10] ), .Z(\SB3_30/i0[7] ) );
  CLKBUF_X1 \SB3_22/BUF_4  ( .A(\RI1[4][58] ), .Z(\SB3_22/i0[7] ) );
  CLKBUF_X1 \SB3_19/BUF_4  ( .A(\RI1[4][76] ), .Z(\SB3_19/i0[7] ) );
  CLKBUF_X1 \SB3_1/BUF_4  ( .A(\RI1[4][184] ), .Z(\SB3_1/i0[7] ) );
  CLKBUF_X1 \SB3_3/BUF_4  ( .A(\RI1[4][172] ), .Z(\SB3_3/i0[7] ) );
  CLKBUF_X1 \SB3_23/BUF_4  ( .A(\RI1[4][52] ), .Z(\SB3_23/i0[7] ) );
  BUF_X1 \SB4_23/BUF_0  ( .A(\RI3[4][48] ), .Z(\SB4_23/i0[9] ) );
  CLKBUF_X1 U31 ( .A(Key[128]), .Z(n442) );
  CLKBUF_X1 U66 ( .A(Key[88]), .Z(n490) );
  CLKBUF_X1 U65 ( .A(Key[67]), .Z(n443) );
  CLKBUF_X1 U53 ( .A(Key[16]), .Z(n452) );
  BUF_X1 U93 ( .A(Key[171]), .Z(n483) );
  CLKBUF_X1 U122 ( .A(Key[77]), .Z(n387) );
  CLKBUF_X1 U58 ( .A(Key[12]), .Z(n427) );
  BUF_X1 U46 ( .A(Key[148]), .Z(n491) );
  CLKBUF_X1 U50 ( .A(Key[92]), .Z(n422) );
  BUF_X1 \SB1_0_30/BUF_2  ( .A(n184), .Z(\SB1_0_30/i1[9] ) );
  INV_X1 U176 ( .A(n442), .ZN(n252) );
  INV_X1 U151 ( .A(n419), .ZN(n251) );
  BUF_X1 \SB2_0_30/BUF_0  ( .A(\RI3[0][6] ), .Z(\SB2_0_30/i0[9] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_0  ( .A(\RI5[0][0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[0] ) );
  CLKBUF_X1 \SB1_1_4/BUF_4  ( .A(\RI1[1][166] ), .Z(\SB1_1_4/i0[7] ) );
  INV_X1 \SB1_2_4/INV_0  ( .A(\RI1[2][162] ), .ZN(\SB1_2_4/i0[9] ) );
  BUF_X1 \SB2_2_25/BUF_1  ( .A(\RI3[2][37] ), .Z(\SB2_2_25/i0[6] ) );
  BUF_X2 \SB1_1_11/BUF_3  ( .A(\RI1[1][123] ), .Z(\SB1_1_11/i0[8] ) );
  BUF_X2 \SB1_1_4/BUF_2  ( .A(\RI1[1][164] ), .Z(\SB1_1_4/i1[9] ) );
  BUF_X2 \SB2_1_19/BUF_1  ( .A(\RI3[1][73] ), .Z(\SB2_1_19/i0[6] ) );
  BUF_X2 \SB2_0_19/BUF_0  ( .A(\RI3[0][72] ), .Z(\SB2_0_19/i0[9] ) );
  BUF_X2 \SB1_2_24/BUF_3  ( .A(\RI1[2][45] ), .Z(\SB1_2_24/i0[8] ) );
  BUF_X2 \SB2_2_2/BUF_1  ( .A(\RI3[2][175] ), .Z(\SB2_2_2/i0[6] ) );
  BUF_X2 \SB1_2_12/BUF_3  ( .A(\RI1[2][117] ), .Z(\SB1_2_12/i0[8] ) );
  BUF_X1 \SB1_3_0/BUF_1  ( .A(\RI1[3][187] ), .Z(\SB1_3_0/i1_7 ) );
  CLKBUF_X3 \MC_ARK_ARC_1_3/BUF_2  ( .A(\RI5[3][2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[2] ) );
  BUF_X2 \SB1_2_23/BUF_3  ( .A(\RI1[2][51] ), .Z(\SB1_2_23/i0[8] ) );
  BUF_X2 \SB2_0_0/BUF_3  ( .A(\RI3[0][189] ), .Z(\SB2_0_0/i0[10] ) );
  BUF_X2 \SB2_0_24/BUF_1  ( .A(\RI3[0][43] ), .Z(\SB2_0_24/i0[6] ) );
  NAND4_X2 \SB2_0_2/Component_Function_2/N5  ( .A1(
        \SB2_0_2/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_2/Component_Function_2/NAND4_in[0] ), .ZN(\RI5[0][2] ) );
  NAND4_X2 \SB2_1_14/Component_Function_3/N5  ( .A1(
        \SB2_1_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][117] ) );
  INV_X1 U232 ( .A(n483), .ZN(n212) );
  BUF_X1 \SB1_2_25/BUF_3  ( .A(\RI1[2][39] ), .Z(\SB1_2_25/i0[8] ) );
  NAND4_X2 \SB2_3_31/Component_Function_3/N5  ( .A1(
        \SB2_3_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_31/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][15] ) );
  NAND4_X2 \SB2_3_27/Component_Function_2/N5  ( .A1(
        \SB2_3_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_27/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_27/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_27/Component_Function_2/NAND4_in[1] ), .ZN(\RI5[3][44] ) );
  NAND4_X2 \SB2_3_12/Component_Function_3/N5  ( .A1(
        \SB2_3_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_12/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][129] ) );
  NAND4_X2 \SB2_3_13/Component_Function_4/N5  ( .A1(
        \SB2_3_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_13/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_13/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][118] ) );
  NAND4_X2 \SB2_3_16/Component_Function_3/N5  ( .A1(
        \SB2_3_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_16/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][105] ) );
  NAND4_X2 \SB2_3_6/Component_Function_3/N5  ( .A1(
        \SB2_3_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][165] ) );
  NAND4_X2 \SB2_3_17/Component_Function_3/N5  ( .A1(
        \SB2_3_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_17/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][99] ) );
  NAND4_X2 \SB2_3_22/Component_Function_3/N5  ( .A1(
        \SB2_3_22/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_22/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][69] ) );
  BUF_X1 \SB3_7/BUF_2  ( .A(\RI1[4][146] ), .Z(\SB3_7/i1[9] ) );
  BUF_X1 \SB3_15/BUF_2  ( .A(\RI1[4][98] ), .Z(\SB3_15/i1[9] ) );
  BUF_X1 \SB3_17/BUF_2  ( .A(\RI1[4][86] ), .Z(\SB3_17/i1[9] ) );
  BUF_X1 \SB3_22/BUF_3  ( .A(\RI1[4][57] ), .Z(\SB3_22/i0[8] ) );
  BUF_X1 \SB3_8/BUF_3  ( .A(\RI1[4][141] ), .Z(\SB3_8/i0[8] ) );
  BUF_X1 \SB3_11/BUF_3  ( .A(\RI1[4][123] ), .Z(\SB3_11/i0[8] ) );
  BUF_X1 U15 ( .A(\RI1[4][75] ), .Z(\SB3_19/i0[8] ) );
  BUF_X1 U106 ( .A(\RI3[3][91] ), .Z(\SB2_3_16/i0[6] ) );
  CLKBUF_X2 U260 ( .A(\RI1[3][146] ), .Z(\SB1_3_7/i1[9] ) );
  BUF_X2 U261 ( .A(\RI1[3][33] ), .Z(\SB1_3_26/i0[8] ) );
  NAND4_X2 U263 ( .A1(\SB2_2_18/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_18/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_18/Component_Function_3/NAND4_in[2] ), .A4(n1128), .ZN(
        \RI5[2][93] ) );
  BUF_X2 U277 ( .A(\RI3[2][13] ), .Z(\SB2_2_29/i0[6] ) );
  BUF_X2 U280 ( .A(\RI3[2][61] ), .Z(\SB2_2_21/i0[6] ) );
  BUF_X2 U283 ( .A(\RI3[2][109] ), .Z(\SB2_2_13/i0[6] ) );
  BUF_X1 U293 ( .A(\RI3[2][73] ), .Z(\SB2_2_19/i0[6] ) );
  BUF_X2 U302 ( .A(\RI1[2][98] ), .Z(\SB1_2_15/i1[9] ) );
  BUF_X2 U526 ( .A(\RI1[2][14] ), .Z(\SB1_2_29/i1[9] ) );
  BUF_X2 U530 ( .A(\RI3[1][181] ), .Z(\SB2_1_1/i0[6] ) );
  BUF_X2 U534 ( .A(\RI1[1][80] ), .Z(\SB1_1_18/i1[9] ) );
  BUF_X2 U541 ( .A(\RI3[0][92] ), .Z(\SB2_0_16/i0_0 ) );
  BUF_X2 U545 ( .A(\RI3[0][86] ), .Z(\SB2_0_17/i0_0 ) );
  BUF_X2 U548 ( .A(\RI1[2][2] ), .Z(\SB1_2_31/i1[9] ) );
  BUF_X2 U551 ( .A(\RI3[0][19] ), .Z(\SB2_0_28/i0[6] ) );
  BUF_X1 U554 ( .A(\RI1[4][87] ), .Z(\SB3_17/i0[8] ) );
  BUF_X1 U561 ( .A(\RI1[4][113] ), .Z(\SB3_13/i1_5 ) );
  BUF_X1 U562 ( .A(\RI1[4][93] ), .Z(\SB3_16/i0[8] ) );
  BUF_X1 U563 ( .A(\RI1[4][81] ), .Z(\SB3_18/i0[8] ) );
  BUF_X1 U564 ( .A(n107), .Z(\SB1_0_17/i1_7 ) );
  BUF_X1 U565 ( .A(n7), .Z(\SB1_0_1/i1_5 ) );
  NAND4_X2 U569 ( .A1(\SB2_0_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][163] ) );
  NAND4_X2 U572 ( .A1(\SB2_1_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_14/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_14/Component_Function_0/NAND4_in[1] ), .ZN(\RI5[1][132] ) );
  NAND4_X2 U573 ( .A1(\SB2_1_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[1][138] ) );
  NAND4_X2 U575 ( .A1(\SB2_2_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_7/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_2_7/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_7/Component_Function_5/NAND4_in[1] ), .ZN(n816) );
  NAND4_X2 U579 ( .A1(\SB2_2_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[155] ) );
  INV_X2 U580 ( .A(\RI1[3][191] ), .ZN(n809) );
  NAND4_X2 U582 ( .A1(\SB1_3_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_3_7/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_3_7/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][154] ) );
  NAND4_X2 U583 ( .A1(\SB2_3_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][39] ) );
  NAND4_X2 U584 ( .A1(\SB2_3_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_28/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][33] ) );
  NAND4_X2 U585 ( .A1(\SB2_3_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_28/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_28/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_28/Component_Function_4/NAND4_in[1] ), .ZN(\RI5[3][28] ) );
  NAND4_X2 U587 ( .A1(\SB2_3_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_25/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][51] ) );
  NAND4_X2 U588 ( .A1(\SB2_3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_18/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][103] ) );
  NAND4_X2 U589 ( .A1(\SB2_3_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][93] ) );
  NAND4_X2 U591 ( .A1(\SB2_3_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_11/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][135] ) );
  NAND4_X2 U592 ( .A1(\SB2_3_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_12/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[3][134] ) );
  NAND4_X2 U593 ( .A1(\SB2_3_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][123] ) );
  NAND4_X2 U594 ( .A1(\SB2_3_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][169] ) );
  NAND4_X2 U595 ( .A1(\SB2_3_1/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_1/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_1/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_1/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][190] ) );
  NAND4_X2 U596 ( .A1(\SB2_3_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][177] ) );
  NAND4_X2 U599 ( .A1(\SB2_3_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_2/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][189] ) );
  NAND4_X1 U606 ( .A1(\SB2_1_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_0/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_0/Component_Function_5/NAND4_in[0] ), .A4(n947), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[191] ) );
  CLKBUF_X1 U607 ( .A(\RI1[4][161] ), .Z(\SB3_5/i1_5 ) );
  CLKBUF_X1 U611 ( .A(\RI1[3][154] ), .Z(\SB1_3_6/i0[7] ) );
  NAND4_X1 U618 ( .A1(\SB2_1_26/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_26/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[35] ) );
  CLKBUF_X1 U637 ( .A(n145), .Z(\SB1_0_24/i1_5 ) );
  CLKBUF_X1 U643 ( .A(Key[119]), .Z(n402) );
  CLKBUF_X1 U644 ( .A(\MC_ARK_ARC_1_3/buf_datainput[125] ), .Z(n520) );
  NAND4_X1 U646 ( .A1(\SB2_3_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_11/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_11/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_11/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[125] ) );
  BUF_X2 U663 ( .A(\RI1[2][92] ), .Z(\SB1_2_16/i1[9] ) );
  BUF_X2 U673 ( .A(\RI3[4][187] ), .Z(\SB4_0/i0[6] ) );
  CLKBUF_X3 U675 ( .A(\RI1[3][158] ), .Z(\SB1_3_5/i1[9] ) );
  BUF_X2 U676 ( .A(\RI3[4][121] ), .Z(\SB4_11/i0[6] ) );
  BUF_X2 U683 ( .A(\RI3[4][49] ), .Z(\SB4_23/i0[6] ) );
  INV_X2 U688 ( .A(n1), .ZN(\SB1_0_0/i0_3 ) );
  BUF_X2 U690 ( .A(\RI3[0][104] ), .Z(\SB2_0_14/i0_0 ) );
  BUF_X2 U691 ( .A(\RI3[2][39] ), .Z(\SB2_2_25/i0[10] ) );
  BUF_X1 U698 ( .A(n177), .Z(\SB1_0_29/i0[8] ) );
  BUF_X1 U728 ( .A(\RI1[4][135] ), .Z(\SB3_9/i0[8] ) );
  BUF_X1 U730 ( .A(\RI1[4][129] ), .Z(\SB3_10/i0[8] ) );
  NAND4_X1 U734 ( .A1(n1272), .A2(\SB2_3_9/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_3_9/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_9/Component_Function_5/NAND4_in[0] ), .ZN(n784) );
  BUF_X2 U736 ( .A(\RI3[3][56] ), .Z(\SB2_3_22/i0_0 ) );
  BUF_X2 U737 ( .A(\RI3[3][128] ), .Z(\SB2_3_10/i0_0 ) );
  BUF_X1 U743 ( .A(\RI5[2][129] ), .Z(n815) );
  INV_X1 U750 ( .A(\RI1[2][72] ), .ZN(\SB1_2_19/i0[9] ) );
  INV_X1 U751 ( .A(\RI1[2][186] ), .ZN(\SB1_2_0/i0[9] ) );
  INV_X1 U754 ( .A(\RI3[1][104] ), .ZN(\SB2_1_14/i1[9] ) );
  INV_X1 U760 ( .A(\RI3[0][182] ), .ZN(\SB2_0_1/i1[9] ) );
  NAND4_X1 U762 ( .A1(\SB1_0_3/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_3/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_0_3/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_3/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][6] ) );
  BUF_X1 U767 ( .A(n31), .Z(\SB1_0_5/i1_5 ) );
  CLKBUF_X1 U768 ( .A(n89), .Z(\SB1_0_14/i1_7 ) );
  INV_X1 U770 ( .A(n56), .ZN(\SB1_0_9/i0_4 ) );
  INV_X1 U772 ( .A(n110), .ZN(\SB1_0_18/i0_4 ) );
  CLKBUF_X1 U774 ( .A(n157), .Z(\SB1_0_26/i1_5 ) );
  BUF_X1 U775 ( .A(\RI3[0][132] ), .Z(\SB2_0_9/i0[9] ) );
  CLKBUF_X1 U777 ( .A(\RI1[1][76] ), .Z(\SB1_1_19/i0[7] ) );
  CLKBUF_X1 U778 ( .A(\RI1[1][124] ), .Z(\SB1_1_11/i0[7] ) );
  CLKBUF_X1 U779 ( .A(\RI1[1][28] ), .Z(\SB1_1_27/i0[7] ) );
  INV_X1 U781 ( .A(\RI1[1][36] ), .ZN(\SB1_1_25/i0[9] ) );
  INV_X1 U782 ( .A(\RI1[1][126] ), .ZN(\SB1_1_10/i0[9] ) );
  CLKBUF_X1 U783 ( .A(\RI1[1][52] ), .Z(\SB1_1_23/i0[7] ) );
  INV_X1 U784 ( .A(\RI1[1][162] ), .ZN(\SB1_1_4/i0[9] ) );
  CLKBUF_X1 U788 ( .A(\RI1[2][88] ), .Z(\SB1_2_17/i0[7] ) );
  CLKBUF_X1 U789 ( .A(\RI1[2][178] ), .Z(\SB1_2_2/i0[7] ) );
  CLKBUF_X1 U790 ( .A(\RI1[2][184] ), .Z(\SB1_2_1/i0[7] ) );
  CLKBUF_X1 U791 ( .A(\RI1[2][160] ), .Z(\SB1_2_5/i0[7] ) );
  CLKBUF_X1 U792 ( .A(\RI1[2][109] ), .Z(\SB1_2_13/i1_7 ) );
  CLKBUF_X1 U793 ( .A(\RI1[2][16] ), .Z(\SB1_2_29/i0[7] ) );
  CLKBUF_X1 U794 ( .A(\RI1[2][70] ), .Z(\SB1_2_20/i0[7] ) );
  CLKBUF_X1 U795 ( .A(\RI1[2][100] ), .Z(\SB1_2_15/i0[7] ) );
  CLKBUF_X1 U796 ( .A(\RI1[2][28] ), .Z(\SB1_2_27/i0[7] ) );
  CLKBUF_X1 U799 ( .A(\RI1[2][121] ), .Z(\SB1_2_11/i1_7 ) );
  BUF_X1 U800 ( .A(\RI3[2][156] ), .Z(\SB2_2_5/i0[9] ) );
  BUF_X1 U802 ( .A(\RI5[2][129] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[129] ) );
  NAND4_X1 U803 ( .A1(\SB2_2_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_12/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_12/Component_Function_5/NAND4_in[0] ), .ZN(n812) );
  XNOR2_X1 U804 ( .A(\MC_ARK_ARC_1_2/buf_datainput[53] ), .B(n441), .ZN(
        \MC_ARK_ARC_1_2/temp4[17] ) );
  CLKBUF_X1 U805 ( .A(\RI1[3][22] ), .Z(\SB1_3_28/i0[7] ) );
  CLKBUF_X1 U806 ( .A(\RI1[3][70] ), .Z(\SB1_3_20/i0[7] ) );
  CLKBUF_X1 U807 ( .A(\RI1[3][82] ), .Z(\SB1_3_18/i0[7] ) );
  CLKBUF_X1 U808 ( .A(\RI1[3][160] ), .Z(\SB1_3_5/i0[7] ) );
  CLKBUF_X1 U809 ( .A(\RI1[3][40] ), .Z(\SB1_3_25/i0[7] ) );
  INV_X1 U811 ( .A(\RI1[3][102] ), .ZN(\SB1_3_14/i0[9] ) );
  AND2_X1 U813 ( .A1(\RI3[3][12] ), .A2(\RI3[3][13] ), .ZN(n596) );
  INV_X1 U815 ( .A(\RI3[3][152] ), .ZN(\SB2_3_6/i1[9] ) );
  BUF_X1 U817 ( .A(\RI3[3][180] ), .Z(\SB2_3_1/i0[9] ) );
  BUF_X1 U818 ( .A(\RI3[3][66] ), .Z(\SB2_3_20/i0[9] ) );
  CLKBUF_X1 U819 ( .A(Key[150]), .Z(\MC_ARK_ARC_1_3/buf_keyinput[70] ) );
  XNOR2_X1 U820 ( .A(\MC_ARK_ARC_1_3/buf_datainput[47] ), .B(n197), .ZN(
        \MC_ARK_ARC_1_3/temp4[11] ) );
  CLKBUF_X1 U821 ( .A(\RI1[4][166] ), .Z(\SB3_4/i0[7] ) );
  CLKBUF_X1 U823 ( .A(\RI1[4][94] ), .Z(\SB3_16/i0[7] ) );
  CLKBUF_X1 U824 ( .A(\RI1[4][106] ), .Z(\SB3_14/i0[7] ) );
  CLKBUF_X1 U825 ( .A(\RI1[4][118] ), .Z(\SB3_12/i0[7] ) );
  CLKBUF_X1 U826 ( .A(\RI1[4][136] ), .Z(\SB3_9/i0[7] ) );
  CLKBUF_X1 U827 ( .A(\RI1[4][143] ), .Z(\SB3_8/i1_5 ) );
  CLKBUF_X1 U828 ( .A(\RI1[4][154] ), .Z(\SB3_6/i0[7] ) );
  BUF_X1 U829 ( .A(\RI1[4][171] ), .Z(\SB3_3/i0[8] ) );
  CLKBUF_X1 U830 ( .A(\RI1[4][178] ), .Z(\SB3_2/i0[7] ) );
  CLKBUF_X1 U831 ( .A(\RI1[4][35] ), .Z(\SB3_26/i1_5 ) );
  BUF_X1 U832 ( .A(\RI1[4][33] ), .Z(\SB3_26/i0[8] ) );
  CLKBUF_X1 U833 ( .A(\RI1[4][28] ), .Z(\SB3_27/i0[7] ) );
  BUF_X1 U834 ( .A(\RI1[4][99] ), .Z(\SB3_15/i0[8] ) );
  BUF_X1 U835 ( .A(\RI1[4][117] ), .Z(\SB3_12/i0[8] ) );
  CLKBUF_X1 U836 ( .A(\RI1[4][137] ), .Z(\SB3_9/i1_5 ) );
  CLKBUF_X1 U837 ( .A(\RI1[4][148] ), .Z(\SB3_7/i0[7] ) );
  AND4_X1 U842 ( .A1(\SB3_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_4/NAND4_in[3] ), .ZN(n548) );
  AND4_X1 U843 ( .A1(\SB3_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_4/NAND4_in[3] ), .ZN(n549) );
  AND4_X1 U844 ( .A1(\SB3_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_0/NAND4_in[0] ), .A4(n1035), .ZN(n550) );
  AND4_X1 U845 ( .A1(\SB3_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_12/Component_Function_4/NAND4_in[3] ), .ZN(n551) );
  AND4_X1 U846 ( .A1(\SB3_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_28/Component_Function_4/NAND4_in[3] ), .ZN(n552) );
  AND4_X1 U847 ( .A1(\SB3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_15/Component_Function_4/NAND4_in[3] ), .ZN(n553) );
  AND4_X1 U848 ( .A1(\SB3_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_1/Component_Function_1/NAND4_in[3] ), .ZN(n554) );
  AND4_X1 U849 ( .A1(\SB3_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_2/Component_Function_0/NAND4_in[0] ), .A4(n960), .ZN(n555) );
  AND4_X1 U851 ( .A1(\SB3_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_7/Component_Function_0/NAND4_in[0] ), .A4(n1340), .ZN(n556) );
  XNOR2_X1 U854 ( .A(n557), .B(n285), .ZN(Ciphertext[111]) );
  NAND3_X1 U864 ( .A1(\SB2_1_30/i0[9] ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i0[6] ), .ZN(n561) );
  NAND3_X1 U869 ( .A1(\SB1_3_17/i0_0 ), .A2(\SB1_3_17/i0_4 ), .A3(
        \SB1_3_17/i1_5 ), .ZN(\SB1_3_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U870 ( .A1(\SB2_1_7/i0[6] ), .A2(\SB2_1_7/i0_4 ), .A3(\RI3[1][144] ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U872 ( .A1(\SB2_1_29/i0_0 ), .A2(\SB2_1_29/i3[0] ), .ZN(n563) );
  NAND4_X1 U875 ( .A1(\SB3_14/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_5/NAND4_in[0] ), .A4(n565), .ZN(
        \RI3[4][107] ) );
  NAND3_X1 U876 ( .A1(\SB3_14/i1[9] ), .A2(\SB3_14/i0_4 ), .A3(\SB3_14/i0_3 ), 
        .ZN(n565) );
  NAND2_X1 U877 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i3[0] ), .ZN(n566) );
  BUF_X2 U878 ( .A(\RI5[3][113] ), .Z(n797) );
  NAND4_X4 U879 ( .A1(\SB2_2_31/Component_Function_2/NAND4_in[1] ), .A2(n1273), 
        .A3(\SB2_2_31/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_2_31/Component_Function_2/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[20] ) );
  NAND4_X1 U880 ( .A1(\SB4_22/Component_Function_2/NAND4_in[2] ), .A2(n1363), 
        .A3(\SB4_22/Component_Function_2/NAND4_in[1] ), .A4(n567), .ZN(n987)
         );
  NAND4_X2 U882 ( .A1(\SB2_0_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_27/Component_Function_3/NAND4_in[2] ), .A4(n660), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[39] ) );
  NAND4_X1 U884 ( .A1(\SB2_0_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_1/Component_Function_2/NAND4_in[1] ), .A4(n568), .ZN(
        \RI5[0][8] ) );
  NAND4_X1 U886 ( .A1(\SB1_1_8/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_8/Component_Function_3/NAND4_in[0] ), .A4(n569), .ZN(
        \RI3[1][153] ) );
  NAND3_X1 U887 ( .A1(\SB1_1_8/i3[0] ), .A2(\SB1_1_8/i1_5 ), .A3(
        \SB1_1_8/i0[8] ), .ZN(n569) );
  NAND4_X2 U890 ( .A1(\SB2_0_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_11/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[135] ) );
  NAND3_X1 U891 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i0[10] ), .A3(
        \SB2_0_25/i0[6] ), .ZN(\SB2_0_25/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U892 ( .A1(\SB1_0_4/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_0_4/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[0][182] ) );
  XNOR2_X1 U898 ( .A(n573), .B(n227), .ZN(Ciphertext[65]) );
  NAND4_X1 U899 ( .A1(\SB4_21/Component_Function_5/NAND4_in[2] ), .A2(n1041), 
        .A3(\SB4_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_21/Component_Function_5/NAND4_in[0] ), .ZN(n573) );
  NAND4_X1 U900 ( .A1(\SB1_3_21/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_3_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_21/Component_Function_0/NAND4_in[0] ), .A4(n574), .ZN(
        \RI3[3][90] ) );
  NAND3_X1 U901 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[10] ), .A3(
        \SB1_3_21/i0_4 ), .ZN(n574) );
  BUF_X1 U902 ( .A(\RI5[3][131] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[131] ) );
  NAND3_X1 U903 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i0_4 ), .A3(n1964), .ZN(
        \SB4_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U911 ( .A1(\SB2_1_7/i0[9] ), .A2(\SB2_1_7/i0_3 ), .A3(
        \SB2_1_7/i0[8] ), .ZN(\SB2_1_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U912 ( .A1(\SB2_2_27/i0[9] ), .A2(\SB2_2_27/i0[8] ), .A3(
        \SB2_2_27/i0_3 ), .ZN(\SB2_2_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U913 ( .A1(\SB2_1_24/i0[8] ), .A2(\SB2_1_24/i3[0] ), .A3(
        \SB2_1_24/i1_5 ), .ZN(\SB2_1_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U914 ( .A1(\SB2_2_7/i1_5 ), .A2(\SB2_2_7/i3[0] ), .A3(
        \SB2_2_7/i0[8] ), .ZN(\SB2_2_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U915 ( .A1(\SB1_1_31/i0_0 ), .A2(\SB1_1_31/i0_4 ), .A3(
        \SB1_1_31/i1_5 ), .ZN(\SB1_1_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U916 ( .A1(\SB2_1_15/i0[10] ), .A2(\SB2_1_15/i0_0 ), .A3(
        \SB2_1_15/i0[6] ), .ZN(\SB2_1_15/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U918 ( .A(n579), .B(n578), .ZN(\RI1[1][5] ) );
  XNOR2_X1 U919 ( .A(\MC_ARK_ARC_1_0/temp1[5] ), .B(\MC_ARK_ARC_1_0/temp4[5] ), 
        .ZN(n578) );
  XNOR2_X1 U920 ( .A(\MC_ARK_ARC_1_0/temp2[5] ), .B(\MC_ARK_ARC_1_0/temp3[5] ), 
        .ZN(n579) );
  NAND3_X1 U921 ( .A1(\SB2_0_1/i1_5 ), .A2(\SB2_0_1/i3[0] ), .A3(
        \SB2_0_1/i0[8] ), .ZN(n1158) );
  NAND4_X1 U922 ( .A1(\SB1_2_10/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_10/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_10/Component_Function_2/NAND4_in[2] ), .A4(n580), .ZN(
        \RI3[2][146] ) );
  NAND3_X1 U923 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i0_4 ), .A3(
        \SB1_2_10/i1_5 ), .ZN(n580) );
  NAND4_X1 U927 ( .A1(\SB1_0_5/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_0_5/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_5/Component_Function_5/NAND4_in[0] ), .A4(n582), .ZN(
        \RI3[0][161] ) );
  NAND4_X1 U930 ( .A1(\SB3_28/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_5/NAND4_in[0] ), .A4(n583), .ZN(
        \RI3[4][23] ) );
  NAND3_X1 U931 ( .A1(\SB3_28/i0_4 ), .A2(\SB3_28/i0_3 ), .A3(\SB3_28/i1[9] ), 
        .ZN(n583) );
  NAND3_X1 U934 ( .A1(\SB2_2_9/i0_0 ), .A2(\SB2_2_9/i0[10] ), .A3(
        \SB2_2_9/i0[6] ), .ZN(\SB2_2_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U935 ( .A1(\SB2_2_30/i3[0] ), .A2(\SB2_2_30/i1_5 ), .A3(
        \SB2_2_30/i0[8] ), .ZN(\SB2_2_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U936 ( .A1(\SB1_2_0/i0_3 ), .A2(\SB1_2_0/i0_0 ), .A3(\SB1_2_0/i0_4 ), .ZN(\SB1_2_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U937 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i0_4 ), .A3(
        \SB2_3_22/i1[9] ), .ZN(n585) );
  NAND4_X1 U939 ( .A1(\SB1_2_7/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_7/Component_Function_5/NAND4_in[0] ), .A4(n584), .ZN(
        \RI3[2][149] ) );
  NAND3_X1 U940 ( .A1(\SB1_2_7/i0_3 ), .A2(\SB1_2_7/i1[9] ), .A3(
        \SB1_2_7/i0_4 ), .ZN(n584) );
  NAND3_X1 U942 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0_0 ), .A3(
        \SB2_2_19/i0_4 ), .ZN(\SB2_2_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U943 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0_4 ), .A3(
        \SB2_3_19/i1[9] ), .ZN(\SB2_3_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U945 ( .A1(\SB2_3_26/i0_0 ), .A2(\SB2_3_26/i0[10] ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 U947 ( .A1(\SB2_1_5/i0_0 ), .A2(\SB2_1_5/i3[0] ), .ZN(n586) );
  NAND3_X1 U949 ( .A1(\SB1_2_12/i0_0 ), .A2(\SB1_2_12/i0_4 ), .A3(
        \SB1_2_12/i1_5 ), .ZN(\SB1_2_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U950 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0[7] ), .A3(
        \SB1_0_22/i0_0 ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U953 ( .A(\MC_ARK_ARC_1_1/temp5[21] ), .B(n588), .ZN(\RI1[2][21] )
         );
  XNOR2_X1 U954 ( .A(\MC_ARK_ARC_1_1/temp3[21] ), .B(
        \MC_ARK_ARC_1_1/temp4[21] ), .ZN(n588) );
  NAND4_X1 U955 ( .A1(\SB2_2_9/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_9/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_9/Component_Function_2/NAND4_in[1] ), .A4(n589), .ZN(
        \RI5[2][152] ) );
  NAND3_X1 U956 ( .A1(\SB2_2_9/i0_4 ), .A2(\SB2_2_9/i1_5 ), .A3(\SB2_2_9/i0_0 ), .ZN(n589) );
  NAND3_X1 U957 ( .A1(\SB4_5/i0_3 ), .A2(n834), .A3(\SB4_5/i0_0 ), .ZN(
        \SB4_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U958 ( .A1(\SB2_0_14/i0[9] ), .A2(\SB2_0_14/i0_3 ), .A3(
        \SB2_0_14/i0[8] ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U961 ( .A1(\SB1_2_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_3/Component_Function_2/NAND4_in[2] ), .A4(n590), .ZN(
        \RI3[2][188] ) );
  NAND3_X1 U962 ( .A1(\SB1_2_3/i0_0 ), .A2(\SB1_2_3/i0_4 ), .A3(\SB1_2_3/i1_5 ), .ZN(n590) );
  NAND3_X1 U964 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i1_5 ), .A3(\SB4_23/i0_4 ), 
        .ZN(n591) );
  NAND3_X1 U965 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0[10] ), .A3(
        \SB1_3_26/i0[9] ), .ZN(\SB1_3_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U967 ( .A1(\SB2_3_6/i0_0 ), .A2(\SB2_3_6/i1_5 ), .A3(\RI3[3][154] ), 
        .ZN(n592) );
  NAND4_X1 U968 ( .A1(\SB3_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_2/NAND4_in[0] ), .A4(n593), .ZN(
        \RI3[4][50] ) );
  NAND3_X1 U969 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i1_5 ), .A3(\SB3_26/i0_4 ), 
        .ZN(n593) );
  NAND3_X1 U970 ( .A1(n851), .A2(n779), .A3(\SB4_22/i0[8] ), .ZN(
        \SB4_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U971 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i0[10] ), .A3(\SB4_13/i0_4 ), 
        .ZN(\SB4_13/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U976 ( .A1(\SB2_3_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_29/Component_Function_5/NAND4_in[0] ), .A4(n595), .ZN(
        \RI5[3][17] ) );
  NAND2_X1 U977 ( .A1(\SB2_3_29/i0_4 ), .A2(n596), .ZN(n595) );
  NAND3_X1 U978 ( .A1(\SB1_2_8/i0_0 ), .A2(\SB1_2_8/i0_4 ), .A3(\SB1_2_8/i1_5 ), .ZN(\SB1_2_8/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U981 ( .A1(\SB2_2_18/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_18/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_18/Component_Function_4/NAND4_in[1] ), .A4(n598), .ZN(
        \RI5[2][88] ) );
  NAND3_X1 U982 ( .A1(\SB2_2_18/i0_4 ), .A2(\SB2_2_18/i1_5 ), .A3(
        \SB2_2_18/i1[9] ), .ZN(n598) );
  NAND2_X1 U983 ( .A1(\SB2_1_11/i0[6] ), .A2(n599), .ZN(
        \SB2_1_11/Component_Function_5/NAND4_in[3] ) );
  AND2_X1 U984 ( .A1(\RI3[1][124] ), .A2(\RI3[1][120] ), .ZN(n599) );
  NAND3_X1 U985 ( .A1(\SB2_2_23/i0[10] ), .A2(\SB2_2_23/i1_5 ), .A3(
        \SB2_2_23/i1[9] ), .ZN(\SB2_2_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U986 ( .A1(\SB1_1_11/i1[9] ), .A2(\SB1_1_11/i0[10] ), .A3(
        \SB1_1_11/i1_7 ), .ZN(\SB1_1_11/Component_Function_3/NAND4_in[2] ) );
  XNOR2_X1 U987 ( .A(n600), .B(\MC_ARK_ARC_1_2/temp6[15] ), .ZN(\RI1[3][15] )
         );
  XNOR2_X1 U988 ( .A(\MC_ARK_ARC_1_2/temp1[15] ), .B(
        \MC_ARK_ARC_1_2/temp2[15] ), .ZN(n600) );
  NAND4_X1 U989 ( .A1(\SB2_1_11/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_11/Component_Function_4/NAND4_in[1] ), .A4(n601), .ZN(
        \RI5[1][130] ) );
  NAND3_X1 U990 ( .A1(\SB2_1_11/i0_4 ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB2_1_11/i1[9] ), .ZN(n601) );
  NAND3_X1 U992 ( .A1(\SB3_13/i1[9] ), .A2(\SB3_13/i0[10] ), .A3(\SB3_13/i1_7 ), .ZN(\SB3_13/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U996 ( .A1(\SB1_2_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_15/Component_Function_5/NAND4_in[0] ), .A4(n603), .ZN(
        \RI3[2][101] ) );
  NAND4_X1 U998 ( .A1(\SB1_2_10/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_10/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_10/Component_Function_5/NAND4_in[0] ), .A4(n604), .ZN(
        \RI3[2][131] ) );
  NAND3_X1 U999 ( .A1(\SB1_2_10/i0_3 ), .A2(\SB1_2_10/i1[9] ), .A3(
        \SB1_2_10/i0_4 ), .ZN(n604) );
  XNOR2_X1 U1000 ( .A(n605), .B(n374), .ZN(Ciphertext[125]) );
  NAND4_X1 U1001 ( .A1(\SB4_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_11/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_11/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_11/Component_Function_5/NAND4_in[0] ), .ZN(n605) );
  NAND3_X1 U1004 ( .A1(\SB2_0_18/i0_3 ), .A2(\SB2_0_18/i0_4 ), .A3(
        \SB2_0_18/i1[9] ), .ZN(\SB2_0_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1005 ( .A1(\SB2_1_11/i0_4 ), .A2(\SB2_1_11/i0_3 ), .A3(
        \SB2_1_11/i0_0 ), .ZN(\SB2_1_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1006 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0[9] ), .A3(
        \SB1_0_21/i0[8] ), .ZN(\SB1_0_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1007 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0_0 ), .A3(
        \SB1_0_21/i0_4 ), .ZN(\SB1_0_21/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U1008 ( .A(\RI1[1][65] ), .ZN(\SB1_1_21/i0_3 ) );
  XNOR2_X1 U1009 ( .A(\MC_ARK_ARC_1_0/temp6[65] ), .B(
        \MC_ARK_ARC_1_0/temp5[65] ), .ZN(\RI1[1][65] ) );
  NAND3_X1 U1010 ( .A1(\SB2_0_2/i0_0 ), .A2(\SB2_0_2/i0[7] ), .A3(
        \SB2_0_2/i0_3 ), .ZN(\SB2_0_2/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U1012 ( .A1(\SB2_1_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_5/NAND4_in[1] ), .A3(n927), .A4(
        \SB2_1_11/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[125] ) );
  NAND3_X1 U1013 ( .A1(n2149), .A2(\SB1_1_4/i0_0 ), .A3(\SB1_1_4/i0_4 ), .ZN(
        \SB1_1_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1014 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i1[9] ), .A3(\SB4_2/i0[6] ), 
        .ZN(\SB4_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1017 ( .A1(\SB2_2_11/i0_3 ), .A2(\SB2_2_11/i1[9] ), .A3(
        \SB2_2_11/i0[6] ), .ZN(\SB2_2_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1020 ( .A1(\SB1_3_18/i0[10] ), .A2(\SB1_3_18/i1[9] ), .A3(
        \SB1_3_18/i1_5 ), .ZN(\SB1_3_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1021 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i3[0] ), .A3(\SB4_31/i1_7 ), 
        .ZN(\SB4_31/Component_Function_4/NAND4_in[1] ) );
  NAND4_X1 U1022 ( .A1(\SB1_1_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_12/Component_Function_2/NAND4_in[2] ), .A4(n609), .ZN(
        \RI3[1][134] ) );
  NAND3_X1 U1023 ( .A1(\SB1_1_12/i0_0 ), .A2(\SB1_1_12/i0_4 ), .A3(
        \SB1_1_12/i1_5 ), .ZN(n609) );
  NAND3_X1 U1026 ( .A1(\SB2_0_2/i0_3 ), .A2(\SB2_0_2/i0[9] ), .A3(
        \SB2_0_2/i0[10] ), .ZN(\SB2_0_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1030 ( .A1(\SB2_1_24/i0_4 ), .A2(\SB2_1_24/i0[9] ), .A3(
        \SB2_1_24/i0[6] ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1031 ( .A1(\SB2_1_8/i0_4 ), .A2(\SB2_1_8/i0_3 ), .A3(
        \SB2_1_8/i0_0 ), .ZN(\SB2_1_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1033 ( .A1(\SB2_1_21/i0_3 ), .A2(\SB2_1_21/i0[9] ), .A3(
        \SB2_1_21/i0[8] ), .ZN(n611) );
  NAND3_X1 U1037 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i1_5 ), .A3(
        \SB2_1_3/i0_0 ), .ZN(n613) );
  NAND3_X1 U1038 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0[9] ), .A3(
        \SB2_1_25/i0[10] ), .ZN(\SB2_1_25/Component_Function_4/NAND4_in[2] )
         );
  AND2_X1 U1041 ( .A1(\RI3[1][139] ), .A2(\RI3[1][142] ), .ZN(n718) );
  XNOR2_X1 U1042 ( .A(n615), .B(n344), .ZN(Ciphertext[6]) );
  NAND3_X1 U1044 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i0_0 ), .A3(
        \SB2_3_19/i0[6] ), .ZN(\SB2_3_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1045 ( .A1(\SB2_2_14/i0[9] ), .A2(\SB2_2_14/i0_3 ), .A3(
        \SB2_2_14/i0[8] ), .ZN(\SB2_2_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1047 ( .A1(\SB1_2_29/i0_0 ), .A2(\SB1_2_29/i0_4 ), .A3(
        \SB1_2_29/i0_3 ), .ZN(\SB1_2_29/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U1049 ( .A(\MC_ARK_ARC_1_3/temp6[86] ), .B(n616), .ZN(\RI1[4][86] )
         );
  XNOR2_X1 U1050 ( .A(\MC_ARK_ARC_1_3/temp2[86] ), .B(
        \MC_ARK_ARC_1_3/temp1[86] ), .ZN(n616) );
  NAND4_X2 U1052 ( .A1(\SB2_2_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_13/Component_Function_5/NAND4_in[1] ), .A4(n617), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[113] ) );
  NAND2_X1 U1053 ( .A1(\SB2_2_13/i0_0 ), .A2(\SB2_2_13/i3[0] ), .ZN(n617) );
  NAND3_X1 U1054 ( .A1(\SB1_2_12/i1[9] ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i1_7 ), .ZN(\SB1_2_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1055 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i0_0 ), .A3(
        \SB2_1_21/i0[6] ), .ZN(\SB2_1_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1057 ( .A1(\SB2_3_19/i0_4 ), .A2(\RI3[3][72] ), .A3(
        \SB2_3_19/i0[6] ), .ZN(\SB2_3_19/Component_Function_5/NAND4_in[3] ) );
  NAND4_X1 U1060 ( .A1(\SB1_3_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_31/Component_Function_4/NAND4_in[3] ), .A4(n618), .ZN(
        \RI3[3][10] ) );
  NAND3_X1 U1061 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[9] ), .A3(
        \SB1_3_31/i0[10] ), .ZN(n618) );
  NAND4_X1 U1062 ( .A1(\SB2_3_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_30/Component_Function_5/NAND4_in[0] ), .A4(n619), .ZN(
        \RI5[3][11] ) );
  NAND3_X1 U1063 ( .A1(\SB2_3_30/i0_4 ), .A2(\RI3[3][6] ), .A3(
        \SB2_3_30/i0[6] ), .ZN(n619) );
  NAND3_X1 U1065 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0_4 ), .A3(
        \SB2_1_25/i1[9] ), .ZN(n1422) );
  NAND4_X1 U1066 ( .A1(\SB4_31/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_31/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_31/Component_Function_4/NAND4_in[1] ), .A4(n620), .ZN(n1466) );
  NAND3_X1 U1068 ( .A1(\SB2_0_27/i0_0 ), .A2(\SB2_0_27/i3[0] ), .A3(
        \SB2_0_27/i1_7 ), .ZN(\SB2_0_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1070 ( .A1(\SB1_3_22/i0_0 ), .A2(\SB1_3_22/i0_4 ), .A3(
        \SB1_3_22/i1_5 ), .ZN(\SB1_3_22/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U1071 ( .A1(\SB1_3_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_3_25/Component_Function_4/NAND4_in[1] ), .A4(n621), .ZN(
        \RI3[3][46] ) );
  NAND3_X1 U1072 ( .A1(\SB1_3_25/i0[10] ), .A2(n804), .A3(\SB1_3_25/i0[9] ), 
        .ZN(n621) );
  NAND3_X1 U1076 ( .A1(\SB2_1_3/i0_0 ), .A2(\SB2_1_3/i3[0] ), .A3(
        \SB2_1_3/i1_7 ), .ZN(\SB2_1_3/Component_Function_4/NAND4_in[1] ) );
  NAND4_X1 U1077 ( .A1(\SB1_2_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_8/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_8/Component_Function_5/NAND4_in[0] ), .A4(n623), .ZN(
        \RI3[2][143] ) );
  NAND3_X1 U1078 ( .A1(\SB1_2_8/i0_4 ), .A2(\SB1_2_8/i0[9] ), .A3(
        \SB1_2_8/i0[6] ), .ZN(n623) );
  NAND3_X1 U1079 ( .A1(\SB2_2_8/i0_0 ), .A2(\SB2_2_8/i0[7] ), .A3(
        \SB2_2_8/i0_3 ), .ZN(\SB2_2_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1080 ( .A1(\SB1_3_30/i0[9] ), .A2(\SB1_3_30/i1_5 ), .A3(
        \SB1_3_30/i0[6] ), .ZN(\SB1_3_30/Component_Function_1/NAND4_in[2] ) );
  NAND4_X1 U1084 ( .A1(\SB1_2_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_13/Component_Function_2/NAND4_in[2] ), .A4(n625), .ZN(
        \RI3[2][128] ) );
  NAND3_X1 U1085 ( .A1(\SB1_2_13/i0_0 ), .A2(\SB1_2_13/i0_4 ), .A3(
        \SB1_2_13/i1_5 ), .ZN(n625) );
  NAND3_X1 U1086 ( .A1(\SB4_2/i0_4 ), .A2(n785), .A3(\SB4_2/i0[6] ), .ZN(
        \SB4_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1089 ( .A1(\SB2_1_8/i0_0 ), .A2(\SB2_1_8/i3[0] ), .A3(
        \SB2_1_8/i1_7 ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[1] ) );
  XNOR2_X1 U1090 ( .A(n627), .B(n321), .ZN(Ciphertext[133]) );
  NAND4_X1 U1091 ( .A1(\SB4_9/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_9/Component_Function_1/NAND4_in[0] ), .A3(
        \SB4_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_9/Component_Function_1/NAND4_in[3] ), .ZN(n627) );
  NAND3_X1 U1092 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i0[9] ), .A3(
        \SB2_1_28/i0[6] ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1093 ( .A1(\SB1_2_1/i1[9] ), .A2(\SB1_2_1/i0[10] ), .A3(
        \SB1_2_1/i1_7 ), .ZN(\SB1_2_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1094 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i0_4 ), .A3(\SB4_7/i0_0 ), 
        .ZN(\SB4_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1095 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i0_4 ), .A3(\SB4_7/i0[10] ), 
        .ZN(\SB4_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1096 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i1[9] ), .A3(
        \SB2_2_18/i0[6] ), .ZN(\SB2_2_18/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U1100 ( .A(\RI1[3][185] ), .ZN(\SB1_3_1/i0_3 ) );
  XNOR2_X1 U1101 ( .A(\MC_ARK_ARC_1_2/temp6[185] ), .B(
        \MC_ARK_ARC_1_2/temp5[185] ), .ZN(\RI1[3][185] ) );
  NAND3_X1 U1102 ( .A1(\SB2_1_4/i0_4 ), .A2(\SB2_1_4/i0[9] ), .A3(
        \SB2_1_4/i0[6] ), .ZN(\SB2_1_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1103 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0[10] ), .A3(
        \SB1_0_22/i0_4 ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1110 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[10] ), .A3(
        \SB1_3_21/i0[9] ), .ZN(\SB1_3_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1111 ( .A1(\SB4_2/i0_0 ), .A2(n785), .A3(\SB4_2/i0[8] ), .ZN(
        \SB4_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1112 ( .A1(\SB2_3_23/i0[9] ), .A2(\SB2_3_23/i0_3 ), .A3(
        \SB2_3_23/i0[8] ), .ZN(\SB2_3_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1113 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0[7] ), .ZN(\SB2_2_0/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U1114 ( .A1(\SB3_21/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_21/Component_Function_1/NAND4_in[0] ), .A3(
        \SB3_21/Component_Function_1/NAND4_in[1] ), .A4(n631), .ZN(
        \RI3[4][85] ) );
  NAND3_X1 U1115 ( .A1(\SB3_21/i1_7 ), .A2(\SB3_21/i0_4 ), .A3(\SB3_21/i0[8] ), 
        .ZN(n631) );
  NAND3_X1 U1116 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0_4 ), .ZN(\SB2_2_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1117 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i1_5 ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1120 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i1[9] ), .A3(
        \SB1_1_3/i0_4 ), .ZN(\SB1_1_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1121 ( .A1(\SB2_0_14/i0_4 ), .A2(\SB2_0_14/i0_3 ), .A3(
        \SB2_0_14/i1[9] ), .ZN(\SB2_0_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1122 ( .A1(\SB2_3_31/i0_3 ), .A2(n1651), .A3(\SB2_3_31/i1[9] ), 
        .ZN(\SB2_3_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1124 ( .A1(\SB2_2_17/i0[9] ), .A2(\SB2_2_17/i0_3 ), .A3(
        \SB2_2_17/i0[8] ), .ZN(n633) );
  NAND3_X1 U1127 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0[9] ), .A3(\SB4_12/i0[8] ), .ZN(\SB4_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1128 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i1_5 ), .A3(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U1129 ( .A1(\SB1_2_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_23/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_23/Component_Function_2/NAND4_in[2] ), .A4(n634), .ZN(
        \RI3[2][68] ) );
  NAND3_X1 U1130 ( .A1(\SB1_2_23/i0_0 ), .A2(\SB1_2_23/i0_4 ), .A3(
        \SB1_2_23/i1_5 ), .ZN(n634) );
  NAND3_X1 U1131 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0_0 ), .A3(
        \SB2_2_4/i0_4 ), .ZN(\SB2_2_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1132 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i0_4 ), .A3(
        \SB1_3_5/i0_0 ), .ZN(\SB1_3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1134 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i1[9] ), .A3(n554), .ZN(
        n635) );
  XNOR2_X1 U1135 ( .A(n636), .B(n312), .ZN(Ciphertext[107]) );
  NAND4_X1 U1136 ( .A1(\SB4_14/Component_Function_5/NAND4_in[2] ), .A2(n637), 
        .A3(\SB4_14/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_14/Component_Function_5/NAND4_in[0] ), .ZN(n636) );
  NAND3_X1 U1137 ( .A1(\SB2_3_18/i0_0 ), .A2(\SB2_3_18/i0_4 ), .A3(
        \SB2_3_18/i0_3 ), .ZN(\SB2_3_18/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U1138 ( .A(\MC_ARK_ARC_1_3/temp5[147] ), .B(
        \MC_ARK_ARC_1_3/temp6[147] ), .ZN(\RI1[4][147] ) );
  XNOR2_X1 U1139 ( .A(\MC_ARK_ARC_1_3/temp2[147] ), .B(
        \MC_ARK_ARC_1_3/temp1[147] ), .ZN(\MC_ARK_ARC_1_3/temp5[147] ) );
  NAND3_X1 U1140 ( .A1(\SB4_14/i0[10] ), .A2(\SB4_14/i0_0 ), .A3(n806), .ZN(
        n637) );
  NAND3_X1 U1141 ( .A1(\SB4_5/i0[8] ), .A2(\SB4_5/i1_5 ), .A3(\SB4_5/i3[0] ), 
        .ZN(\SB4_5/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U1142 ( .A1(\SB3_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_7/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_7/Component_Function_3/NAND4_in[3] ), .A4(n638), .ZN(
        \RI3[4][159] ) );
  NAND3_X1 U1143 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i1[9] ), .A3(\SB3_7/i1_7 ), 
        .ZN(n638) );
  NAND3_X1 U1144 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i0_4 ), .A3(
        \SB1_1_3/i0[10] ), .ZN(\SB1_1_3/Component_Function_0/NAND4_in[2] ) );
  XNOR2_X1 U1145 ( .A(n640), .B(n639), .ZN(\RI1[2][29] ) );
  XNOR2_X1 U1146 ( .A(\MC_ARK_ARC_1_1/temp4[29] ), .B(
        \MC_ARK_ARC_1_1/temp2[29] ), .ZN(n639) );
  XNOR2_X1 U1147 ( .A(\MC_ARK_ARC_1_1/temp1[29] ), .B(
        \MC_ARK_ARC_1_1/temp3[29] ), .ZN(n640) );
  XNOR2_X1 U1148 ( .A(n642), .B(n641), .ZN(\RI1[1][77] ) );
  XNOR2_X1 U1149 ( .A(\MC_ARK_ARC_1_0/temp2[77] ), .B(
        \MC_ARK_ARC_1_0/temp4[77] ), .ZN(n641) );
  XNOR2_X1 U1150 ( .A(\MC_ARK_ARC_1_0/temp1[77] ), .B(
        \MC_ARK_ARC_1_0/temp3[77] ), .ZN(n642) );
  NAND3_X1 U1151 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0_4 ), .A3(
        \SB1_0_10/i1[9] ), .ZN(\SB1_0_10/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U1154 ( .A(n644), .B(n296), .ZN(Ciphertext[178]) );
  NAND4_X1 U1155 ( .A1(\SB4_2/Component_Function_4/NAND4_in[2] ), .A2(n758), 
        .A3(\SB4_2/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_2/Component_Function_4/NAND4_in[1] ), .ZN(n644) );
  XNOR2_X1 U1156 ( .A(n645), .B(n646), .ZN(\RI1[4][178] ) );
  XNOR2_X1 U1157 ( .A(\MC_ARK_ARC_1_3/temp1[178] ), .B(
        \MC_ARK_ARC_1_3/temp4[178] ), .ZN(n645) );
  XNOR2_X1 U1158 ( .A(\MC_ARK_ARC_1_3/temp3[178] ), .B(
        \MC_ARK_ARC_1_3/temp2[178] ), .ZN(n646) );
  NAND4_X1 U1159 ( .A1(\SB3_2/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_2/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_2/Component_Function_4/NAND4_in[2] ), .A4(n647), .ZN(
        \RI3[4][184] ) );
  NAND3_X1 U1160 ( .A1(\SB3_2/i0_4 ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i1_5 ), 
        .ZN(n647) );
  XNOR2_X1 U1164 ( .A(n650), .B(n349), .ZN(Ciphertext[19]) );
  NAND4_X1 U1165 ( .A1(n1278), .A2(\SB4_28/Component_Function_1/NAND4_in[2] ), 
        .A3(\SB4_28/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_28/Component_Function_1/NAND4_in[0] ), .ZN(n650) );
  NAND4_X1 U1168 ( .A1(\SB3_1/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_1/Component_Function_0/NAND4_in[0] ), .A4(n652), .ZN(\RI3[4][18] ) );
  NAND3_X1 U1169 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i0[7] ), .A3(\SB3_1/i0_0 ), 
        .ZN(n652) );
  XNOR2_X1 U1171 ( .A(\MC_ARK_ARC_1_0/temp3[11] ), .B(
        \MC_ARK_ARC_1_0/temp4[11] ), .ZN(n653) );
  XNOR2_X1 U1172 ( .A(\MC_ARK_ARC_1_0/temp2[11] ), .B(
        \MC_ARK_ARC_1_0/temp1[11] ), .ZN(n654) );
  NAND4_X1 U1173 ( .A1(\SB2_1_5/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_5/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_5/Component_Function_4/NAND4_in[1] ), .A4(n655), .ZN(
        \RI5[1][166] ) );
  NAND3_X1 U1174 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0[9] ), .A3(
        \SB2_1_5/i0[10] ), .ZN(n655) );
  NAND4_X1 U1175 ( .A1(\SB2_0_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_29/Component_Function_2/NAND4_in[1] ), .A4(n656), .ZN(
        \RI5[0][32] ) );
  NAND3_X1 U1176 ( .A1(\SB2_0_29/i0_0 ), .A2(\SB2_0_29/i1_5 ), .A3(
        \SB2_0_29/i0_4 ), .ZN(n656) );
  NAND4_X1 U1177 ( .A1(n963), .A2(\SB1_1_17/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB1_1_17/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_1_17/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[1][104] ) );
  NAND3_X1 U1178 ( .A1(\SB1_0_30/i0[9] ), .A2(\SB1_0_30/i0[10] ), .A3(
        \SB1_0_30/i0_3 ), .ZN(\SB1_0_30/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U1179 ( .A(n657), .B(n330), .ZN(Ciphertext[118]) );
  NAND4_X1 U1180 ( .A1(\SB4_12/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_12/Component_Function_4/NAND4_in[3] ), .A3(
        \SB4_12/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_12/Component_Function_4/NAND4_in[1] ), .ZN(n657) );
  NAND3_X1 U1182 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i0_4 ), .A3(
        \SB2_0_6/i0_0 ), .ZN(\SB2_0_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1183 ( .A1(\SB2_2_24/i0_4 ), .A2(\SB2_2_24/i0_3 ), .A3(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U1185 ( .A(\MC_ARK_ARC_1_2/temp1[155] ), .B(
        \MC_ARK_ARC_1_2/temp4[155] ), .ZN(n658) );
  NAND3_X1 U1187 ( .A1(\SB1_2_14/i0_4 ), .A2(\SB1_2_14/i0_0 ), .A3(
        \SB1_2_14/i1_5 ), .ZN(n937) );
  NAND4_X2 U1189 ( .A1(\SB2_2_29/Component_Function_5/NAND4_in[3] ), .A2(n1193), .A3(\SB2_2_29/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[17] ) );
  NAND3_X1 U1190 ( .A1(\SB2_0_27/i3[0] ), .A2(\SB2_0_27/i1_5 ), .A3(
        \SB2_0_27/i0[8] ), .ZN(n660) );
  NAND3_X1 U1192 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i1_5 ), .A3(
        \SB4_30/i1[9] ), .ZN(n661) );
  NAND3_X1 U1193 ( .A1(\SB1_2_0/i1[9] ), .A2(\SB1_2_0/i0_4 ), .A3(
        \SB1_2_0/i1_5 ), .ZN(\SB1_2_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1194 ( .A1(\SB2_2_31/i0_0 ), .A2(\SB2_2_31/i0_4 ), .A3(
        \SB2_2_31/i1_5 ), .ZN(\SB2_2_31/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U1195 ( .A1(\SB3_0/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_0/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_0/Component_Function_3/NAND4_in[2] ), .A4(n662), .ZN(\RI3[4][9] )
         );
  NAND3_X1 U1196 ( .A1(\SB3_0/i3[0] ), .A2(\SB3_0/i1_5 ), .A3(\SB3_0/i0[8] ), 
        .ZN(n662) );
  NAND3_X1 U1198 ( .A1(\SB3_24/i3[0] ), .A2(\SB3_24/i1_5 ), .A3(\SB3_24/i0[8] ), .ZN(n663) );
  XNOR2_X1 U1199 ( .A(\MC_ARK_ARC_1_3/buf_datainput[144] ), .B(\RI5[3][108] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[42] ) );
  NAND4_X2 U1200 ( .A1(\SB2_3_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_18/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_18/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][108] ) );
  NAND3_X1 U1201 ( .A1(\SB2_2_15/i0[10] ), .A2(\SB2_2_15/i1_5 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U1202 ( .A1(\SB2_2_17/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_17/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_17/Component_Function_4/NAND4_in[1] ), .A4(n664), .ZN(
        \RI5[2][94] ) );
  NAND3_X1 U1203 ( .A1(\SB2_2_17/i0_4 ), .A2(\SB2_2_17/i1_5 ), .A3(
        \SB2_2_17/i1[9] ), .ZN(n664) );
  XNOR2_X1 U1205 ( .A(n666), .B(n355), .ZN(Ciphertext[73]) );
  NAND4_X1 U1206 ( .A1(\SB4_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_19/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_19/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_19/Component_Function_1/NAND4_in[2] ), .ZN(n666) );
  NAND4_X1 U1207 ( .A1(\SB1_3_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_7/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_7/Component_Function_2/NAND4_in[2] ), .A4(n667), .ZN(
        \RI3[3][164] ) );
  NAND2_X1 U1210 ( .A1(\SB2_2_11/i0_0 ), .A2(\SB2_2_11/i3[0] ), .ZN(n668) );
  NAND3_X1 U1211 ( .A1(\SB2_1_0/i0_0 ), .A2(\SB2_1_0/i0[10] ), .A3(
        \SB2_1_0/i0[6] ), .ZN(\SB2_1_0/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1212 ( .A1(\SB2_3_31/i0[6] ), .A2(\SB2_3_31/i0_0 ), .A3(
        \SB2_3_31/i0[10] ), .ZN(\SB2_3_31/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U1214 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i1[9] ), .A3(\SB4_5/i1_7 ), 
        .ZN(\SB4_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1216 ( .A1(\SB2_3_18/i0[8] ), .A2(\SB2_3_18/i1_5 ), .A3(
        \SB2_3_18/i3[0] ), .ZN(\SB2_3_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1217 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i1_5 ), .A3(\SB4_16/i0_4 ), 
        .ZN(\SB4_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1218 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0[8] ), .ZN(\SB2_2_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1219 ( .A1(\SB1_3_7/i1[9] ), .A2(\SB1_3_7/i0_3 ), .A3(
        \SB1_3_7/i0_4 ), .ZN(n978) );
  NAND3_X1 U1220 ( .A1(\SB2_1_19/i0_3 ), .A2(\SB2_1_19/i1[9] ), .A3(
        \SB2_1_19/i0[6] ), .ZN(\SB2_1_19/Component_Function_3/NAND4_in[0] ) );
  INV_X1 U1222 ( .A(\RI1[4][16] ), .ZN(\SB3_29/i0_4 ) );
  XNOR2_X1 U1223 ( .A(\MC_ARK_ARC_1_3/temp5[16] ), .B(
        \MC_ARK_ARC_1_3/temp6[16] ), .ZN(\RI1[4][16] ) );
  NAND3_X1 U1225 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i0_0 ), .A3(
        \SB2_2_17/i0[7] ), .ZN(\SB2_2_17/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U1226 ( .A(n669), .B(n337), .ZN(Ciphertext[62]) );
  NAND4_X1 U1227 ( .A1(n681), .A2(\SB4_21/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB4_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB4_21/Component_Function_2/NAND4_in[1] ), .ZN(n669) );
  NAND3_X1 U1228 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i3[0] ), .A3(\SB4_13/i1_7 ), 
        .ZN(\SB4_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1229 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB2_1_13/i0_4 ), .A3(
        \SB2_1_13/i0_0 ), .ZN(\SB2_1_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1230 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0_0 ), .A3(
        \SB1_3_10/i0_4 ), .ZN(\SB1_3_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1231 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i0_0 ), .A3(
        \SB1_1_8/i0_4 ), .ZN(\SB1_1_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1232 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i0_3 ), .A3(\SB3_26/i0[7] ), 
        .ZN(n1352) );
  NAND3_X1 U1233 ( .A1(\SB2_1_6/i0[8] ), .A2(\SB2_1_6/i1_5 ), .A3(
        \SB2_1_6/i3[0] ), .ZN(\SB2_1_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1234 ( .A1(\SB2_0_11/i0[10] ), .A2(\SB2_0_11/i0_0 ), .A3(
        \SB2_0_11/i0[6] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U1235 ( .A(\MC_ARK_ARC_1_2/temp5[75] ), .B(n670), .ZN(\RI1[3][75] )
         );
  XNOR2_X1 U1236 ( .A(\MC_ARK_ARC_1_2/temp3[75] ), .B(
        \MC_ARK_ARC_1_2/temp4[75] ), .ZN(n670) );
  NAND3_X1 U1237 ( .A1(\SB4_14/i0[9] ), .A2(\SB4_14/i1_5 ), .A3(n806), .ZN(
        \SB4_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1238 ( .A1(\SB2_2_14/i0_4 ), .A2(\SB2_2_14/i1_5 ), .A3(
        \SB2_2_14/i0_0 ), .ZN(\SB2_2_14/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U1239 ( .A1(n1332), .A2(\SB4_21/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB4_21/Component_Function_1/NAND4_in[0] ), .A4(n671), .ZN(n966)
         );
  NAND3_X1 U1240 ( .A1(\SB4_21/i0[9] ), .A2(\SB4_21/i1_5 ), .A3(\SB4_21/i0[6] ), .ZN(n671) );
  NAND3_X1 U1241 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0[9] ), .A3(
        \SB1_1_23/i0[10] ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[2] )
         );
  XNOR2_X1 U1242 ( .A(n672), .B(n368), .ZN(Ciphertext[71]) );
  NAND4_X1 U1243 ( .A1(\SB4_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_20/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_20/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_20/Component_Function_5/NAND4_in[3] ), .ZN(n672) );
  NAND3_X1 U1253 ( .A1(\SB1_3_29/i0_0 ), .A2(\SB1_3_29/i0_4 ), .A3(
        \SB1_3_29/i1_5 ), .ZN(\SB1_3_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1256 ( .A1(\SB4_21/i0_4 ), .A2(\SB4_21/i1_5 ), .A3(\SB4_21/i1[9] ), 
        .ZN(n679) );
  NAND3_X1 U1258 ( .A1(n2114), .A2(\SB2_3_16/i0_3 ), .A3(\SB2_3_16/i0[8] ), 
        .ZN(n680) );
  NAND3_X1 U1259 ( .A1(\SB2_3_20/i0_3 ), .A2(\SB2_3_20/i0[9] ), .A3(
        \SB2_3_20/i0[8] ), .ZN(\SB2_3_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1260 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0_0 ), .A3(
        \SB2_2_28/i0[7] ), .ZN(\SB2_2_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1261 ( .A1(\SB4_21/i0_0 ), .A2(\SB4_21/i0_4 ), .A3(\SB4_21/i1_5 ), 
        .ZN(n681) );
  NAND3_X1 U1263 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i1[9] ), .A3(
        \SB2_0_27/i0[6] ), .ZN(\SB2_0_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1265 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i0[10] ), .A3(
        \SB1_3_5/i0[9] ), .ZN(n682) );
  XNOR2_X1 U1266 ( .A(n684), .B(n683), .ZN(\RI1[2][58] ) );
  XNOR2_X1 U1267 ( .A(\MC_ARK_ARC_1_1/temp1[58] ), .B(
        \MC_ARK_ARC_1_1/temp4[58] ), .ZN(n683) );
  XNOR2_X1 U1268 ( .A(\MC_ARK_ARC_1_1/temp3[58] ), .B(
        \MC_ARK_ARC_1_1/temp2[58] ), .ZN(n684) );
  XNOR2_X1 U1269 ( .A(n686), .B(n685), .ZN(\RI1[3][89] ) );
  XNOR2_X1 U1270 ( .A(\MC_ARK_ARC_1_2/temp4[89] ), .B(
        \MC_ARK_ARC_1_2/temp3[89] ), .ZN(n685) );
  XNOR2_X1 U1271 ( .A(\MC_ARK_ARC_1_2/temp2[89] ), .B(
        \MC_ARK_ARC_1_2/temp1[89] ), .ZN(n686) );
  AND2_X1 U1272 ( .A1(\RI3[2][78] ), .A2(\RI3[2][82] ), .ZN(n728) );
  NAND3_X1 U1275 ( .A1(\SB1_2_22/i0[8] ), .A2(\SB1_2_22/i0_4 ), .A3(
        \SB1_2_22/i1_7 ), .ZN(\SB1_2_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1276 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i3[0] ), .A3(\SB4_23/i1_7 ), 
        .ZN(\SB4_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1278 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0_0 ), .A3(
        \SB1_0_22/i0_4 ), .ZN(\SB1_0_22/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U1279 ( .A(n689), .B(n688), .ZN(\RI1[4][167] ) );
  XNOR2_X1 U1280 ( .A(\MC_ARK_ARC_1_3/temp4[167] ), .B(
        \MC_ARK_ARC_1_3/temp2[167] ), .ZN(n688) );
  XNOR2_X1 U1281 ( .A(\MC_ARK_ARC_1_3/temp1[167] ), .B(
        \MC_ARK_ARC_1_3/temp3[167] ), .ZN(n689) );
  NAND3_X1 U1283 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0[7] ), .A3(
        \SB1_0_0/i0_0 ), .ZN(\SB1_0_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1284 ( .A1(\SB2_2_30/i0[9] ), .A2(\SB2_2_30/i0_4 ), .A3(
        \SB2_2_30/i0[6] ), .ZN(\SB2_2_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1285 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i1[9] ), .A3(
        \SB2_3_27/i0_4 ), .ZN(n690) );
  NAND3_X1 U1286 ( .A1(\SB4_9/i0_0 ), .A2(\SB4_9/i1_5 ), .A3(\RI3[4][136] ), 
        .ZN(\SB4_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1288 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i1_5 ), .A3(
        \SB4_10/i1[9] ), .ZN(n691) );
  XNOR2_X1 U1292 ( .A(n693), .B(n357), .ZN(Ciphertext[155]) );
  NAND4_X1 U1293 ( .A1(\SB4_6/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_6/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_6/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_6/Component_Function_5/NAND4_in[0] ), .ZN(n693) );
  NAND3_X1 U1296 ( .A1(\SB4_7/i0_0 ), .A2(\SB4_7/i3[0] ), .A3(\SB4_7/i1_7 ), 
        .ZN(\SB4_7/Component_Function_4/NAND4_in[1] ) );
  NAND4_X1 U1299 ( .A1(\SB4_1/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_1/Component_Function_2/NAND4_in[3] ), .A3(
        \SB4_1/Component_Function_2/NAND4_in[1] ), .A4(n695), .ZN(n1333) );
  NAND3_X1 U1300 ( .A1(\SB4_1/i0[10] ), .A2(\SB4_1/i1_5 ), .A3(\SB4_1/i1[9] ), 
        .ZN(n695) );
  INV_X2 U1301 ( .A(\RI1[3][53] ), .ZN(\SB1_3_23/i0_3 ) );
  XNOR2_X1 U1302 ( .A(\MC_ARK_ARC_1_2/temp6[53] ), .B(
        \MC_ARK_ARC_1_2/temp5[53] ), .ZN(\RI1[3][53] ) );
  NAND3_X1 U1303 ( .A1(\SB2_2_29/i0_4 ), .A2(\SB2_2_29/i0_3 ), .A3(
        \SB2_2_29/i1[9] ), .ZN(n1193) );
  NAND3_X1 U1304 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i0_4 ), .A3(
        \SB2_2_13/i1[9] ), .ZN(\SB2_2_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1305 ( .A1(\SB2_1_3/i0[9] ), .A2(\SB2_1_3/i0_3 ), .A3(
        \SB2_1_3/i0[8] ), .ZN(\SB2_1_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1306 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0_4 ), .A3(
        \SB2_2_22/i0_0 ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1307 ( .A1(\SB2_0_14/i0[6] ), .A2(\SB2_0_14/i0_3 ), .A3(
        \SB2_0_14/i0[10] ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[1] )
         );
  XNOR2_X1 U1309 ( .A(n696), .B(n697), .ZN(\RI1[2][107] ) );
  XNOR2_X1 U1310 ( .A(\MC_ARK_ARC_1_1/temp4[107] ), .B(
        \MC_ARK_ARC_1_1/temp2[107] ), .ZN(n696) );
  XNOR2_X1 U1311 ( .A(\MC_ARK_ARC_1_1/temp3[107] ), .B(
        \MC_ARK_ARC_1_1/temp1[107] ), .ZN(n697) );
  NAND3_X1 U1312 ( .A1(\SB1_3_25/i0_0 ), .A2(\SB1_3_25/i0[6] ), .A3(
        \SB1_3_25/i0[10] ), .ZN(\SB1_3_25/Component_Function_5/NAND4_in[1] )
         );
  NAND4_X1 U1315 ( .A1(\SB3_3/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_3/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_3/Component_Function_0/NAND4_in[1] ), .A4(n699), .ZN(\RI3[4][6] )
         );
  NAND3_X1 U1316 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i0_3 ), .A3(\SB3_3/i0_4 ), 
        .ZN(n699) );
  NAND3_X1 U1317 ( .A1(\SB2_1_8/i0_3 ), .A2(\SB2_1_8/i0[9] ), .A3(
        \SB2_1_8/i0[10] ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U1318 ( .A1(\SB2_0_25/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_25/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_25/Component_Function_4/NAND4_in[1] ), .A4(n700), .ZN(
        \RI5[0][46] ) );
  NAND3_X1 U1319 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0[9] ), .A3(
        \SB2_0_25/i0[10] ), .ZN(n700) );
  NAND3_X1 U1320 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i1[9] ), .A3(
        \SB1_3_12/i0[6] ), .ZN(\SB1_3_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1322 ( .A1(\RI3[0][10] ), .A2(\SB2_0_30/i1_5 ), .A3(
        \SB2_0_30/i0_0 ), .ZN(n701) );
  NAND3_X1 U1325 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0[9] ), .A3(
        \SB1_1_14/i0[8] ), .ZN(\SB1_1_14/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U1326 ( .A(n703), .B(n238), .ZN(Ciphertext[132]) );
  NAND4_X1 U1327 ( .A1(\SB4_9/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_9/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_9/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_9/Component_Function_0/NAND4_in[1] ), .ZN(n703) );
  NAND4_X1 U1328 ( .A1(\SB1_2_1/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_1/Component_Function_2/NAND4_in[2] ), .A4(n704), .ZN(
        \RI3[2][8] ) );
  NAND3_X1 U1329 ( .A1(\SB1_2_1/i0_0 ), .A2(\SB1_2_1/i0_4 ), .A3(
        \SB1_2_1/i1_5 ), .ZN(n704) );
  NAND3_X1 U1330 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0[10] ), .A3(\SB3_2/i0[9] ), 
        .ZN(\SB3_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1331 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0_0 ), .A3(
        \SB1_3_21/i0_4 ), .ZN(\SB1_3_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1332 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i0_0 ), .A3(
        \SB2_0_27/i0[6] ), .ZN(\SB2_0_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1333 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i1_5 ), .A3(
        \SB4_20/i1[9] ), .ZN(\SB4_20/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U1334 ( .A1(\SB4_15/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_15/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_15/Component_Function_1/NAND4_in[0] ), .A4(n705), .ZN(n1303) );
  NAND3_X1 U1335 ( .A1(\SB4_15/i0[9] ), .A2(\SB4_15/i1_5 ), .A3(\SB4_15/i0[6] ), .ZN(n705) );
  NAND3_X1 U1336 ( .A1(\SB3_20/i0_0 ), .A2(\SB3_20/i0[7] ), .A3(n864), .ZN(
        \SB3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1338 ( .A1(\SB4_22/i1_5 ), .A2(\SB4_22/i0_4 ), .A3(\SB4_22/i1[9] ), 
        .ZN(n706) );
  NAND4_X1 U1339 ( .A1(\SB4_20/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_20/Component_Function_1/NAND4_in[0] ), .A4(n707), .ZN(n1253) );
  NAND3_X1 U1340 ( .A1(\SB4_20/i0[9] ), .A2(\SB4_20/i1_5 ), .A3(\SB4_20/i0[6] ), .ZN(n707) );
  NAND3_X1 U1341 ( .A1(\SB2_1_18/i0[10] ), .A2(\SB2_1_18/i1[9] ), .A3(
        \SB2_1_18/i1_7 ), .ZN(\SB2_1_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1342 ( .A1(\SB4_2/i0_0 ), .A2(n556), .A3(\SB4_2/i1_7 ), .ZN(
        \SB4_2/Component_Function_4/NAND4_in[1] ) );
  NAND4_X1 U1343 ( .A1(\SB1_2_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_2/NAND4_in[2] ), .A4(n708), .ZN(
        \RI3[2][26] ) );
  NAND3_X1 U1344 ( .A1(\SB1_2_30/i0_0 ), .A2(\SB1_2_30/i0_4 ), .A3(
        \SB1_2_30/i1_5 ), .ZN(n708) );
  NAND3_X1 U1346 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0_0 ), .A3(
        \SB2_2_7/i0_4 ), .ZN(\SB2_2_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1347 ( .A1(\SB1_1_3/i1[9] ), .A2(\SB1_1_3/i0_4 ), .A3(
        \SB1_1_3/i1_5 ), .ZN(\SB1_1_3/Component_Function_4/NAND4_in[3] ) );
  NAND4_X1 U1348 ( .A1(\SB2_1_19/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_19/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_19/Component_Function_3/NAND4_in[2] ), .A4(n709), .ZN(
        \RI5[1][87] ) );
  NAND3_X1 U1350 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i0[9] ), .A3(
        \SB2_3_21/i0[8] ), .ZN(\SB2_3_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1351 ( .A1(\SB3_31/i1[9] ), .A2(\SB3_31/i0[10] ), .A3(
        \SB3_31/i1_7 ), .ZN(\SB3_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1354 ( .A1(\SB2_1_18/i0_4 ), .A2(\SB2_1_18/i1_7 ), .A3(
        \SB2_1_18/i0[8] ), .ZN(\SB2_1_18/Component_Function_1/NAND4_in[3] ) );
  XNOR2_X1 U1355 ( .A(n711), .B(n249), .ZN(Ciphertext[89]) );
  NAND4_X1 U1356 ( .A1(\SB4_17/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_17/Component_Function_5/NAND4_in[1] ), .A3(n772), .A4(
        \SB4_17/Component_Function_5/NAND4_in[0] ), .ZN(n711) );
  NAND4_X1 U1359 ( .A1(\SB2_1_16/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_16/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_16/Component_Function_1/NAND4_in[0] ), .A4(n713), .ZN(
        \RI5[1][115] ) );
  NAND3_X1 U1360 ( .A1(\SB2_1_16/i0_4 ), .A2(\SB2_1_16/i1_7 ), .A3(
        \SB2_1_16/i0[8] ), .ZN(n713) );
  NAND4_X2 U1367 ( .A1(\SB2_2_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_19/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[77] ) );
  NAND2_X1 U1370 ( .A1(\RI3[1][138] ), .A2(n718), .ZN(
        \SB2_1_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1371 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0[10] ), .A3(
        \SB1_1_13/i0_4 ), .ZN(\SB1_1_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1372 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0_4 ), .A3(
        \SB2_2_19/i1[9] ), .ZN(\SB2_2_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1373 ( .A1(\SB2_1_16/i0[10] ), .A2(\SB2_1_16/i1_5 ), .A3(
        \SB2_1_16/i1[9] ), .ZN(\SB2_1_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1376 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0[10] ), .A3(
        \SB1_0_12/i0[9] ), .ZN(\SB1_0_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1378 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i0[10] ), .A3(
        \SB2_1_12/i0[6] ), .ZN(\SB2_1_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1379 ( .A1(\SB2_1_3/i0_0 ), .A2(\SB2_1_3/i0[10] ), .A3(
        \SB2_1_3/i0[6] ), .ZN(\SB2_1_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1380 ( .A1(\SB2_0_11/i0_4 ), .A2(\RI3[0][120] ), .A3(
        \SB2_0_11/i0[6] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1381 ( .A1(\SB3_2/i0_4 ), .A2(\SB3_2/i0_3 ), .A3(\SB3_2/i0_0 ), 
        .ZN(\SB3_2/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U1382 ( .A1(\SB2_1_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_8/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_8/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_1_8/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[143] ) );
  NAND3_X1 U1383 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0_0 ), .A3(
        \SB2_2_30/i0_4 ), .ZN(\SB2_2_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1384 ( .A1(\SB2_1_20/i0_3 ), .A2(\SB2_1_20/i1[9] ), .A3(
        \SB2_1_20/i0[6] ), .ZN(\SB2_1_20/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U1386 ( .A1(\SB3_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_7/Component_Function_0/NAND4_in[0] ), .A4(n1340), .ZN(n785) );
  XNOR2_X1 U1387 ( .A(n720), .B(n343), .ZN(Ciphertext[157]) );
  NAND4_X1 U1388 ( .A1(\SB4_5/Component_Function_1/NAND4_in[1] ), .A2(n1202), 
        .A3(\SB4_5/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_5/Component_Function_1/NAND4_in[2] ), .ZN(n720) );
  XNOR2_X1 U1389 ( .A(\MC_ARK_ARC_1_1/temp2[59] ), .B(
        \MC_ARK_ARC_1_1/temp1[59] ), .ZN(n721) );
  NAND4_X1 U1390 ( .A1(\SB4_17/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_17/Component_Function_2/NAND4_in[1] ), .A3(n1309), .A4(n722), 
        .ZN(n1306) );
  NAND3_X1 U1391 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i1_5 ), .A3(
        \SB4_17/i1[9] ), .ZN(n722) );
  NAND3_X1 U1392 ( .A1(\SB3_8/i0[10] ), .A2(\SB3_8/i0_3 ), .A3(\SB3_8/i0_4 ), 
        .ZN(\SB3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1393 ( .A1(n1623), .A2(\SB2_3_19/i0_3 ), .A3(\SB2_3_19/i0[10] ), 
        .ZN(\SB2_3_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1394 ( .A1(\SB2_1_12/i0_4 ), .A2(\SB2_1_12/i1_7 ), .A3(
        \SB2_1_12/i0[8] ), .ZN(\SB2_1_12/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 U1395 ( .A1(\SB4_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB4_8/Component_Function_2/NAND4_in[0] ), .A4(n723), .ZN(n1184) );
  NAND3_X1 U1396 ( .A1(\SB4_8/i0_0 ), .A2(n1638), .A3(\SB4_8/i1_5 ), .ZN(n723)
         );
  NAND4_X1 U1397 ( .A1(\SB2_1_3/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_3/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_3/Component_Function_1/NAND4_in[0] ), .A4(n724), .ZN(
        \RI5[1][1] ) );
  NAND3_X1 U1398 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i1_7 ), .A3(
        \SB2_1_3/i0[8] ), .ZN(n724) );
  NAND3_X1 U1401 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i3[0] ), .A3(\SB4_8/i1_7 ), 
        .ZN(\SB4_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1402 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0_0 ), .A3(\SB3_19/i0_4 ), 
        .ZN(\SB3_19/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U1403 ( .A(n726), .B(n318), .ZN(Ciphertext[161]) );
  NAND4_X1 U1404 ( .A1(\SB4_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_5/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_5/Component_Function_5/NAND4_in[3] ), .ZN(n726) );
  NAND4_X2 U1405 ( .A1(\SB2_2_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_18/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_18/Component_Function_5/NAND4_in[0] ), .A4(n727), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[83] ) );
  NAND2_X1 U1406 ( .A1(\SB2_2_18/i0[6] ), .A2(n728), .ZN(n727) );
  NAND3_X1 U1407 ( .A1(n851), .A2(\SB4_22/i0[7] ), .A3(\SB4_22/i0_0 ), .ZN(
        \SB4_22/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U1408 ( .A1(\SB4_3/Component_Function_1/NAND4_in[1] ), .A2(n1298), 
        .A3(\SB4_3/Component_Function_1/NAND4_in[0] ), .A4(n729), .ZN(n1094)
         );
  NAND3_X1 U1409 ( .A1(\SB4_3/i0[9] ), .A2(\SB4_3/i1_5 ), .A3(\SB4_3/i0[6] ), 
        .ZN(n729) );
  NAND3_X1 U1410 ( .A1(n1663), .A2(\SB4_9/i1[9] ), .A3(\RI3[4][136] ), .ZN(
        \SB4_9/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U1411 ( .A1(\SB4_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_20/Component_Function_3/NAND4_in[3] ), .A4(n730), .ZN(n970) );
  NAND3_X1 U1412 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i1[9] ), .A3(
        \SB4_20/i1_7 ), .ZN(n730) );
  NAND3_X1 U1413 ( .A1(\SB1_2_30/i1[9] ), .A2(\SB1_2_30/i0[10] ), .A3(
        \SB1_2_30/i1_7 ), .ZN(\SB1_2_30/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U1414 ( .A1(\SB2_2_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_0/NAND4_in[0] ), .A4(n731), .ZN(
        \RI5[2][144] ) );
  NAND3_X1 U1415 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0_0 ), .A3(
        \SB2_2_12/i0[7] ), .ZN(n731) );
  XNOR2_X1 U1416 ( .A(n732), .B(n291), .ZN(Ciphertext[165]) );
  NAND3_X1 U1418 ( .A1(\SB4_9/i0_3 ), .A2(\SB4_9/i1[9] ), .A3(\SB4_9/i0[6] ), 
        .ZN(\SB4_9/Component_Function_3/NAND4_in[0] ) );
  XNOR2_X1 U1419 ( .A(\MC_ARK_ARC_1_0/temp5[119] ), .B(n733), .ZN(
        \RI1[1][119] ) );
  XNOR2_X1 U1420 ( .A(\MC_ARK_ARC_1_0/temp3[119] ), .B(
        \MC_ARK_ARC_1_0/temp4[119] ), .ZN(n733) );
  NAND3_X1 U1422 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i0[10] ), .A3(
        \SB1_3_17/i0[9] ), .ZN(n734) );
  XNOR2_X1 U1423 ( .A(n735), .B(n300), .ZN(Ciphertext[191]) );
  NAND4_X1 U1424 ( .A1(\SB4_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_0/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_0/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_0/Component_Function_5/NAND4_in[0] ), .ZN(n735) );
  XNOR2_X1 U1426 ( .A(\MC_ARK_ARC_1_0/temp4[185] ), .B(
        \MC_ARK_ARC_1_0/temp3[185] ), .ZN(n736) );
  XNOR2_X1 U1433 ( .A(n740), .B(n293), .ZN(Ciphertext[55]) );
  NAND4_X1 U1434 ( .A1(\SB4_22/Component_Function_1/NAND4_in[1] ), .A2(n1036), 
        .A3(\SB4_22/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_22/Component_Function_1/NAND4_in[3] ), .ZN(n740) );
  NAND3_X1 U1435 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i3[0] ), .A3(\SB4_14/i1_7 ), 
        .ZN(\SB4_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1436 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i3[0] ), .A3(\SB4_1/i1_7 ), 
        .ZN(n741) );
  NAND3_X1 U1437 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i3[0] ), .A3(\SB4_12/i1_7 ), 
        .ZN(\SB4_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1438 ( .A1(\SB1_0_3/i0_3 ), .A2(\SB1_0_3/i0[9] ), .A3(
        \SB1_0_3/i0[10] ), .ZN(\SB1_0_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1439 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i0_4 ), .A3(
        \SB1_3_1/i1_5 ), .ZN(\SB1_3_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1443 ( .A1(\SB2_1_10/i0[9] ), .A2(\SB2_1_10/i0_3 ), .A3(
        \SB2_1_10/i0[8] ), .ZN(n743) );
  NAND3_X1 U1445 ( .A1(\SB4_26/i0_0 ), .A2(\SB4_26/i3[0] ), .A3(\SB4_26/i1_7 ), 
        .ZN(n744) );
  XNOR2_X1 U1446 ( .A(n745), .B(n313), .ZN(Ciphertext[148]) );
  NAND4_X1 U1447 ( .A1(\SB4_7/Component_Function_4/NAND4_in[2] ), .A2(n1062), 
        .A3(\SB4_7/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_7/Component_Function_4/NAND4_in[1] ), .ZN(n745) );
  NAND3_X1 U1450 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i3[0] ), .A3(\SB4_6/i1_7 ), 
        .ZN(n747) );
  NAND3_X1 U1451 ( .A1(\SB4_0/i0_0 ), .A2(\SB4_0/i3[0] ), .A3(\SB4_0/i1_7 ), 
        .ZN(\SB4_0/Component_Function_4/NAND4_in[1] ) );
  XNOR2_X1 U1456 ( .A(n750), .B(n197), .ZN(Ciphertext[138]) );
  NAND4_X1 U1457 ( .A1(\SB4_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_8/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_8/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_8/Component_Function_0/NAND4_in[1] ), .ZN(n750) );
  NAND2_X1 U1459 ( .A1(\SB2_0_2/i0_0 ), .A2(\SB2_0_2/i3[0] ), .ZN(n751) );
  XNOR2_X1 U1462 ( .A(\MC_ARK_ARC_1_1/temp5[186] ), .B(
        \MC_ARK_ARC_1_1/temp6[186] ), .ZN(\RI1[2][186] ) );
  NAND3_X1 U1464 ( .A1(\SB3_2/i0_4 ), .A2(\SB3_2/i1_7 ), .A3(\SB3_2/i0[8] ), 
        .ZN(\SB3_2/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U1465 ( .A1(\SB2_2_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_28/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_28/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_28/Component_Function_5/NAND4_in[0] ), .ZN(n800) );
  XNOR2_X1 U1466 ( .A(n754), .B(n755), .ZN(\RI1[3][23] ) );
  XNOR2_X1 U1467 ( .A(\MC_ARK_ARC_1_2/temp1[23] ), .B(
        \MC_ARK_ARC_1_2/temp4[23] ), .ZN(n754) );
  XNOR2_X1 U1468 ( .A(\MC_ARK_ARC_1_2/temp3[23] ), .B(
        \MC_ARK_ARC_1_2/temp2[23] ), .ZN(n755) );
  NAND3_X1 U1469 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[10] ), .A3(
        \SB1_1_20/i0_4 ), .ZN(\SB1_1_20/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U1470 ( .A1(\SB1_2_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_5/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_2_5/Component_Function_5/NAND4_in[0] ), .A4(n756), .ZN(
        \RI3[2][161] ) );
  NAND3_X1 U1471 ( .A1(\SB1_2_5/i0_4 ), .A2(\SB1_2_5/i0[6] ), .A3(
        \SB1_2_5/i0[9] ), .ZN(n756) );
  NAND4_X1 U1472 ( .A1(\SB1_1_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_2/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_2/Component_Function_1/NAND4_in[0] ), .A4(n757), .ZN(
        \RI3[1][7] ) );
  NAND3_X1 U1473 ( .A1(\SB1_1_2/i1_7 ), .A2(\SB1_1_2/i0_4 ), .A3(
        \SB1_1_2/i0[8] ), .ZN(n757) );
  NAND3_X1 U1474 ( .A1(\SB4_2/i0_4 ), .A2(\SB4_2/i1[9] ), .A3(\SB4_2/i1_5 ), 
        .ZN(n758) );
  NAND3_X1 U1479 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i1[9] ), .A3(\SB4_0/i1_7 ), 
        .ZN(n761) );
  NAND4_X1 U1480 ( .A1(\SB1_3_20/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_20/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_20/Component_Function_2/NAND4_in[2] ), .A4(n762), .ZN(
        \RI3[3][86] ) );
  XNOR2_X1 U1482 ( .A(n763), .B(n246), .ZN(Ciphertext[158]) );
  NAND4_X1 U1483 ( .A1(\SB4_5/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_5/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_5/Component_Function_2/NAND4_in[0] ), .A4(
        \SB4_5/Component_Function_2/NAND4_in[3] ), .ZN(n763) );
  NAND3_X1 U1484 ( .A1(\SB1_2_29/i0_0 ), .A2(\SB1_2_29/i1_5 ), .A3(
        \SB1_2_29/i0_4 ), .ZN(\SB1_2_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1485 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i0_3 ), .A3(
        \SB2_0_4/i0[9] ), .ZN(\SB2_0_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1486 ( .A1(\SB1_1_2/i0_4 ), .A2(\SB1_1_2/i0[9] ), .A3(
        \SB1_1_2/i0[6] ), .ZN(\SB1_1_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1487 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i1_7 ), .A3(
        \SB2_1_28/i0[8] ), .ZN(\SB2_1_28/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 U1488 ( .A1(\SB1_1_7/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_7/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_7/Component_Function_4/NAND4_in[3] ), .A4(n764), .ZN(
        \RI3[1][154] ) );
  NAND3_X1 U1489 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i0[10] ), .A3(
        \SB1_1_7/i0[9] ), .ZN(n764) );
  XNOR2_X1 U1490 ( .A(n765), .B(n289), .ZN(Ciphertext[83]) );
  NAND3_X1 U1492 ( .A1(\SB1_1_11/i0_4 ), .A2(\SB1_1_11/i0[8] ), .A3(
        \SB1_1_11/i1_7 ), .ZN(\SB1_1_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1493 ( .A1(\SB1_0_30/i1_7 ), .A2(\SB1_0_30/i0[8] ), .A3(
        \SB1_0_30/i0_3 ), .ZN(\SB1_0_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1496 ( .A1(\SB2_2_10/i0[10] ), .A2(\SB2_2_10/i1_5 ), .A3(
        \SB2_2_10/i1[9] ), .ZN(\SB2_2_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1497 ( .A1(n1663), .A2(\RI3[4][136] ), .A3(\SB4_9/i0_0 ), .ZN(
        \SB4_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1498 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0_0 ), .A3(
        \SB1_2_26/i0_4 ), .ZN(\SB1_2_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1505 ( .A1(\SB4_14/i0_0 ), .A2(n799), .A3(\SB4_14/i1_5 ), .ZN(n769) );
  NAND4_X2 U1508 ( .A1(\SB2_3_29/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_29/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_29/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[32] ) );
  XNOR2_X1 U1509 ( .A(\MC_ARK_ARC_1_1/temp6[72] ), .B(
        \MC_ARK_ARC_1_1/temp5[72] ), .ZN(\RI1[2][72] ) );
  NAND3_X1 U1510 ( .A1(\SB2_0_21/i1_5 ), .A2(\SB2_0_21/i3[0] ), .A3(
        \SB2_0_21/i0[8] ), .ZN(\SB2_0_21/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U1512 ( .A1(\SB2_3_24/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_24/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_3_24/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_3_24/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[62] ) );
  NAND3_X1 U1514 ( .A1(\SB2_1_16/i3[0] ), .A2(\SB2_1_16/i1_5 ), .A3(
        \SB2_1_16/i0[8] ), .ZN(n771) );
  NAND3_X1 U1515 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i1[9] ), .A3(\SB4_17/i0_4 ), 
        .ZN(n772) );
  NAND3_X1 U1516 ( .A1(\SB4_29/i0_0 ), .A2(n790), .A3(\SB4_29/i0[8] ), .ZN(
        n773) );
  NAND3_X1 U1517 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i3[0] ), .A3(\SB4_28/i1_7 ), 
        .ZN(\SB4_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1518 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i1[9] ), .A3(
        \SB2_2_2/i0[6] ), .ZN(\SB2_2_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1519 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i1[9] ), .A3(
        \SB2_2_1/i0[6] ), .ZN(\SB2_2_1/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U1520 ( .A1(\SB2_1_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_1_12/Component_Function_2/NAND4_in[1] ), .A4(n774), .ZN(
        \RI5[1][134] ) );
  NAND3_X1 U1521 ( .A1(\SB2_1_12/i0_3 ), .A2(\SB2_1_12/i0[9] ), .A3(
        \SB2_1_12/i0[8] ), .ZN(n774) );
  NAND3_X1 U1522 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i1[9] ), .A3(
        \SB2_0_16/i0[6] ), .ZN(\SB2_0_16/Component_Function_3/NAND4_in[0] ) );
  XNOR2_X1 U1525 ( .A(n777), .B(n776), .ZN(\RI1[4][35] ) );
  XNOR2_X1 U1526 ( .A(\MC_ARK_ARC_1_3/temp2[35] ), .B(
        \MC_ARK_ARC_1_3/temp4[35] ), .ZN(n776) );
  XNOR2_X1 U1527 ( .A(\MC_ARK_ARC_1_3/temp1[35] ), .B(
        \MC_ARK_ARC_1_3/temp3[35] ), .ZN(n777) );
  XNOR2_X1 U1528 ( .A(\MC_ARK_ARC_1_1/temp4[11] ), .B(n778), .ZN(
        \MC_ARK_ARC_1_1/temp6[11] ) );
  XNOR2_X1 U1529 ( .A(\MC_ARK_ARC_1_1/buf_datainput[77] ), .B(n808), .ZN(n778)
         );
  INV_X1 U1531 ( .A(\RI3[0][50] ), .ZN(\SB2_0_23/i1[9] ) );
  BUF_X1 U1534 ( .A(\RI3[4][18] ), .Z(\SB4_28/i0[9] ) );
  NAND4_X2 U1535 ( .A1(\SB3_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_28/Component_Function_4/NAND4_in[3] ), .ZN(n780) );
  NAND4_X1 U1537 ( .A1(n1225), .A2(\SB2_2_23/Component_Function_5/NAND4_in[3] ), .A3(\SB2_2_23/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_23/Component_Function_5/NAND4_in[0] ), .ZN(n782) );
  NAND4_X1 U1538 ( .A1(n1225), .A2(\SB2_2_23/Component_Function_5/NAND4_in[3] ), .A3(\SB2_2_23/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[53] ) );
  NAND4_X2 U1540 ( .A1(\SB2_1_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][93] ) );
  NAND4_X1 U1543 ( .A1(\SB2_0_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_22/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_22/Component_Function_5/NAND4_in[0] ), .ZN(n787) );
  NAND4_X1 U1544 ( .A1(\SB2_0_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_22/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_22/Component_Function_5/NAND4_in[0] ), .ZN(n788) );
  INV_X1 U1545 ( .A(\RI1[1][89] ), .ZN(n789) );
  NAND4_X1 U1546 ( .A1(\SB2_0_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_22/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_22/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[59] ) );
  INV_X1 U1547 ( .A(\RI1[1][89] ), .ZN(\SB1_1_17/i0_3 ) );
  BUF_X1 U1548 ( .A(\RI1[4][183] ), .Z(\SB3_1/i0[8] ) );
  NAND4_X1 U1551 ( .A1(\SB2_2_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_22/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_22/Component_Function_5/NAND4_in[0] ), .ZN(n793) );
  CLKBUF_X1 U1553 ( .A(\RI1[4][149] ), .Z(\SB3_7/i1_5 ) );
  BUF_X1 U1554 ( .A(\RI3[3][42] ), .Z(\SB2_3_24/i0[9] ) );
  NAND4_X1 U1557 ( .A1(n1230), .A2(\SB2_0_1/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_1/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[185] ) );
  XNOR2_X1 U1559 ( .A(\MC_ARK_ARC_1_3/temp5[147] ), .B(
        \MC_ARK_ARC_1_3/temp6[147] ), .ZN(n798) );
  NAND4_X2 U1560 ( .A1(\SB3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_15/Component_Function_4/NAND4_in[2] ), .A3(
        \SB3_15/Component_Function_4/NAND4_in[1] ), .A4(
        \SB3_15/Component_Function_4/NAND4_in[3] ), .ZN(n799) );
  NAND4_X1 U1561 ( .A1(\SB2_2_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_28/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_28/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[23] ) );
  NAND4_X1 U1563 ( .A1(\SB2_2_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_2/Component_Function_5/NAND4_in[3] ), .A4(n1028), .ZN(n803) );
  INV_X1 U1564 ( .A(\RI1[3][41] ), .ZN(n804) );
  INV_X1 U1566 ( .A(\RI1[3][41] ), .ZN(\SB1_3_25/i0_3 ) );
  NAND4_X1 U1568 ( .A1(\SB3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_1/NAND4_in[3] ), .ZN(n806) );
  INV_X1 U1569 ( .A(\RI3[4][86] ), .ZN(\SB4_17/i1[9] ) );
  BUF_X1 U1570 ( .A(\RI1[4][80] ), .Z(\SB3_18/i1[9] ) );
  NAND4_X1 U1573 ( .A1(\SB3_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_1/NAND4_in[3] ), .ZN(n810) );
  NAND4_X1 U1576 ( .A1(\SB2_1_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_18/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_18/Component_Function_5/NAND4_in[0] ), .ZN(n813) );
  INV_X1 U1577 ( .A(\RI1[2][17] ), .ZN(n814) );
  NAND4_X1 U1578 ( .A1(\SB2_1_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_18/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[83] ) );
  INV_X1 U1579 ( .A(\RI1[2][17] ), .ZN(\SB1_2_29/i0_3 ) );
  NAND4_X1 U1580 ( .A1(\SB2_2_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_7/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_7/Component_Function_5/NAND4_in[0] ), .ZN(n817) );
  NAND4_X1 U1581 ( .A1(\SB2_3_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_0/NAND4_in[3] ), .ZN(n818) );
  NAND4_X1 U1582 ( .A1(\SB2_3_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][138] ) );
  INV_X1 U1583 ( .A(\RI1[4][29] ), .ZN(n819) );
  AND4_X1 U1586 ( .A1(\SB3_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_4/NAND4_in[3] ), .ZN(n821) );
  NAND4_X1 U1587 ( .A1(\SB2_2_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_1/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_1/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_1/Component_Function_5/NAND4_in[0] ), .ZN(n822) );
  NAND4_X1 U1588 ( .A1(\SB2_2_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_1/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_1/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_1/Component_Function_5/NAND4_in[0] ), .ZN(n823) );
  NAND4_X1 U1589 ( .A1(\SB2_2_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_1/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_1/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[185] ) );
  NAND4_X1 U1590 ( .A1(\SB2_2_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_6/Component_Function_5/NAND4_in[0] ), .ZN(n824) );
  INV_X1 U1591 ( .A(\RI1[4][76] ), .ZN(\SB3_19/i0_4 ) );
  INV_X1 U1593 ( .A(\RI1[1][131] ), .ZN(n826) );
  INV_X1 U1595 ( .A(\RI1[1][131] ), .ZN(\SB1_1_10/i0_3 ) );
  NAND4_X1 U1596 ( .A1(\SB2_2_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_3/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_3/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[173] ) );
  BUF_X1 U1597 ( .A(\RI3[4][119] ), .Z(n828) );
  BUF_X1 U1598 ( .A(\RI3[4][119] ), .Z(\SB4_12/i0_3 ) );
  NAND4_X1 U1599 ( .A1(\SB2_2_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_0/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_0/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_0/Component_Function_5/NAND4_in[0] ), .ZN(n829) );
  NAND4_X1 U1600 ( .A1(\SB2_2_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_0/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_0/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_0/Component_Function_5/NAND4_in[0] ), .ZN(n830) );
  INV_X1 U1601 ( .A(\RI1[3][125] ), .ZN(n831) );
  NAND4_X1 U1602 ( .A1(\SB2_2_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_0/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_0/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[191] ) );
  INV_X1 U1603 ( .A(\RI1[3][125] ), .ZN(\SB1_3_11/i0_3 ) );
  INV_X1 U1605 ( .A(\RI1[4][155] ), .ZN(n833) );
  NAND4_X2 U1606 ( .A1(\SB3_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_4/NAND4_in[3] ), .ZN(n834) );
  INV_X1 U1607 ( .A(\RI1[4][131] ), .ZN(n835) );
  AND4_X1 U1608 ( .A1(\SB3_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_4/NAND4_in[3] ), .A4(n1114), .ZN(n836) );
  BUF_X2 U1612 ( .A(\RI5[3][185] ), .Z(n839) );
  INV_X1 U1614 ( .A(\RI1[4][125] ), .ZN(n840) );
  INV_X1 U1618 ( .A(\RI1[4][65] ), .ZN(n843) );
  NAND4_X2 U1619 ( .A1(\SB3_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_4/NAND4_in[3] ), .ZN(n844) );
  CLKBUF_X1 U1620 ( .A(\RI1[4][11] ), .Z(\SB3_30/i1_5 ) );
  INV_X1 U1621 ( .A(\RI1[4][41] ), .ZN(n845) );
  NAND4_X2 U1622 ( .A1(\SB2_2_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_25/Component_Function_5/NAND4_in[3] ), .ZN(n846) );
  NAND4_X1 U1623 ( .A1(\SB2_2_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_25/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[41] ) );
  INV_X1 U1624 ( .A(\RI1[4][53] ), .ZN(n847) );
  NAND4_X1 U1631 ( .A1(\SB2_1_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_1_14/Component_Function_5/NAND4_in[3] ), .ZN(n852) );
  NAND4_X1 U1632 ( .A1(\SB2_1_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_1_14/Component_Function_5/NAND4_in[3] ), .ZN(n853) );
  NAND4_X1 U1633 ( .A1(\SB2_1_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_1_14/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[107] ) );
  BUF_X1 U1634 ( .A(\RI3[4][65] ), .Z(n854) );
  BUF_X1 U1635 ( .A(\RI3[4][65] ), .Z(\SB4_21/i0_3 ) );
  INV_X1 U1638 ( .A(\RI1[4][185] ), .ZN(n856) );
  BUF_X1 U1639 ( .A(\RI3[4][185] ), .Z(n857) );
  BUF_X1 U1640 ( .A(\RI3[4][185] ), .Z(\SB4_1/i0_3 ) );
  BUF_X1 U1641 ( .A(\RI3[4][155] ), .Z(n858) );
  BUF_X1 U1642 ( .A(\RI3[4][155] ), .Z(\SB4_6/i0_3 ) );
  BUF_X1 U1643 ( .A(\RI3[4][173] ), .Z(n859) );
  BUF_X1 U1644 ( .A(\RI3[4][173] ), .Z(\SB4_3/i0_3 ) );
  INV_X1 U1646 ( .A(\RI1[4][107] ), .ZN(n860) );
  BUF_X1 U1647 ( .A(\RI1[1][137] ), .Z(\SB1_1_9/i1_5 ) );
  INV_X1 U1648 ( .A(\RI1[4][17] ), .ZN(n861) );
  INV_X1 U1649 ( .A(n85), .ZN(n862) );
  INV_X1 U1650 ( .A(\RI3[4][56] ), .ZN(\SB4_22/i1[9] ) );
  BUF_X1 U1651 ( .A(\RI3[4][143] ), .Z(n863) );
  BUF_X1 U1652 ( .A(\RI3[4][143] ), .Z(\SB4_8/i0_3 ) );
  INV_X1 U1654 ( .A(\RI1[4][191] ), .ZN(\SB3_0/i0_3 ) );
  CLKBUF_X1 U1655 ( .A(\RI1[4][191] ), .Z(\SB3_0/i1_5 ) );
  INV_X1 U1656 ( .A(\RI1[4][71] ), .ZN(n864) );
  INV_X1 U1657 ( .A(\RI1[4][23] ), .ZN(n865) );
  BUF_X1 U1658 ( .A(\RI3[4][23] ), .Z(n866) );
  BUF_X1 U1659 ( .A(\RI3[4][23] ), .Z(\SB4_28/i0_3 ) );
  INV_X1 U1660 ( .A(\RI1[4][89] ), .ZN(n867) );
  BUF_X1 U1661 ( .A(\RI3[4][89] ), .Z(n868) );
  BUF_X1 U1662 ( .A(\RI3[4][89] ), .Z(\SB4_17/i0_3 ) );
  INV_X1 U1663 ( .A(\RI1[4][83] ), .ZN(n869) );
  BUF_X1 U1664 ( .A(\RI3[4][83] ), .Z(n870) );
  BUF_X1 U1665 ( .A(\RI3[4][83] ), .Z(\SB4_18/i0_3 ) );
  BUF_X1 U1666 ( .A(\RI3[4][101] ), .Z(n871) );
  BUF_X1 U1667 ( .A(\RI3[4][101] ), .Z(\SB4_15/i0_3 ) );
  INV_X1 U1668 ( .A(\RI1[4][47] ), .ZN(n872) );
  INV_X1 U1669 ( .A(n115), .ZN(n873) );
  NAND4_X1 U1670 ( .A1(\SB2_0_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_16/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_16/Component_Function_5/NAND4_in[0] ), .ZN(n874) );
  NAND4_X1 U1672 ( .A1(\SB2_0_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_16/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[95] ) );
  INV_X1 U1673 ( .A(\RI1[4][95] ), .ZN(n876) );
  BUF_X1 U1675 ( .A(\RI3[4][149] ), .Z(\SB4_7/i0_3 ) );
  INV_X1 U1676 ( .A(\RI3[4][62] ), .ZN(\SB4_21/i1[9] ) );
  NAND3_X1 U1679 ( .A1(\SB1_2_25/i0_0 ), .A2(\SB1_2_25/i0_4 ), .A3(
        \SB1_2_25/i1_5 ), .ZN(n976) );
  NAND3_X1 U1680 ( .A1(\SB2_0_4/i0_4 ), .A2(\SB2_0_4/i0_0 ), .A3(
        \SB2_0_4/i0_3 ), .ZN(\SB2_0_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1681 ( .A1(\SB2_0_19/i0_4 ), .A2(\SB2_0_19/i0_3 ), .A3(
        \SB2_0_19/i1[9] ), .ZN(\SB2_0_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1682 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i1_5 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(\SB2_1_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1683 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i0_4 ), .A3(
        \SB2_2_13/i0_0 ), .ZN(\SB2_2_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1684 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0[9] ), .A3(
        \SB2_2_12/i0[10] ), .ZN(\SB2_2_12/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1685 ( .A1(n871), .A2(\SB4_15/i0_4 ), .A3(\SB4_15/i1[9] ), .ZN(
        \SB4_15/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1689 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i0_4 ), .A3(
        \SB1_1_2/i1_5 ), .ZN(\SB1_1_2/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U1690 ( .A1(\SB1_3_21/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_21/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_3_21/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_3_21/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_20/i0_4 ) );
  NAND3_X1 U1691 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0_4 ), .A3(
        \SB2_2_12/i0_0 ), .ZN(\SB2_2_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1692 ( .A1(\SB2_0_26/i0_3 ), .A2(\RI3[0][30] ), .A3(
        \SB2_0_26/i0[8] ), .ZN(\SB2_0_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1694 ( .A1(\SB2_3_22/i0[8] ), .A2(\SB2_3_22/i1_5 ), .A3(
        \SB2_3_22/i3[0] ), .ZN(\SB2_3_22/Component_Function_3/NAND4_in[3] ) );
  XNOR2_X1 U1695 ( .A(\MC_ARK_ARC_1_2/temp5[62] ), .B(n880), .ZN(\RI1[3][62] )
         );
  XNOR2_X1 U1696 ( .A(\MC_ARK_ARC_1_2/temp3[62] ), .B(
        \MC_ARK_ARC_1_2/temp4[62] ), .ZN(n880) );
  NAND3_X1 U1697 ( .A1(\SB2_2_5/i0_4 ), .A2(\SB2_2_5/i1_5 ), .A3(
        \SB2_2_5/i0_0 ), .ZN(\SB2_2_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1698 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0[9] ), .A3(\SB3_0/i0[10] ), 
        .ZN(\SB3_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1699 ( .A1(\SB3_26/i0[10] ), .A2(\SB3_26/i1_7 ), .A3(
        \SB3_26/i1[9] ), .ZN(\SB3_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1700 ( .A1(\SB2_0_22/i0_4 ), .A2(\SB2_0_22/i0[9] ), .A3(
        \SB2_0_22/i0[6] ), .ZN(\SB2_0_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1701 ( .A1(\SB2_0_30/i0_0 ), .A2(\SB2_0_30/i0[7] ), .A3(
        \SB2_0_30/i0_3 ), .ZN(\SB2_0_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1702 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0_4 ), .A3(\SB3_0/i1[9] ), 
        .ZN(\SB3_0/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U1706 ( .A1(\SB1_2_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_18/Component_Function_5/NAND4_in[0] ), .A4(n882), .ZN(
        \RI3[2][83] ) );
  NAND3_X1 U1707 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i1[9] ), .A3(
        \SB1_2_18/i0_4 ), .ZN(n882) );
  NAND3_X1 U1708 ( .A1(\SB1_3_7/i0_3 ), .A2(\SB1_3_7/i0_0 ), .A3(
        \SB1_3_7/i0_4 ), .ZN(\SB1_3_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1709 ( .A1(\SB2_2_27/i0_4 ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1710 ( .A1(\SB2_3_5/i0[10] ), .A2(\SB2_3_5/i0_0 ), .A3(
        \SB2_3_5/i0[6] ), .ZN(\SB2_3_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1713 ( .A1(\SB2_0_1/i0[9] ), .A2(\SB2_0_1/i0_4 ), .A3(
        \SB2_0_1/i0[6] ), .ZN(\SB2_0_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1715 ( .A1(\SB4_26/i0_4 ), .A2(\SB4_26/i1_7 ), .A3(\SB4_26/i0[8] ), 
        .ZN(\SB4_26/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U1716 ( .A(\RI1[4][29] ), .ZN(\SB3_27/i0_3 ) );
  NAND4_X1 U1717 ( .A1(\SB1_2_21/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_21/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_21/Component_Function_2/NAND4_in[2] ), .A4(n883), .ZN(
        \RI3[2][80] ) );
  NAND4_X2 U1719 ( .A1(\SB2_3_4/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_4/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[182] ) );
  NAND4_X1 U1720 ( .A1(\SB1_2_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_2/NAND4_in[2] ), .A4(n884), .ZN(
        \RI3[2][38] ) );
  NAND3_X1 U1721 ( .A1(\SB1_2_28/i0_0 ), .A2(\SB1_2_28/i0_4 ), .A3(
        \SB1_2_28/i1_5 ), .ZN(n884) );
  NAND3_X1 U1723 ( .A1(\SB2_1_19/i0[10] ), .A2(\SB2_1_19/i0_0 ), .A3(
        \SB2_1_19/i0[6] ), .ZN(\SB2_1_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1724 ( .A1(\SB2_1_25/i0_4 ), .A2(\SB2_1_25/i0[9] ), .A3(
        \SB2_1_25/i0[6] ), .ZN(\SB2_1_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1725 ( .A1(\SB2_2_29/i0[9] ), .A2(\SB2_2_29/i0_4 ), .A3(
        \SB2_2_29/i0[6] ), .ZN(\SB2_2_29/Component_Function_5/NAND4_in[3] ) );
  NAND4_X4 U1727 ( .A1(\SB2_0_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_18/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[83] ) );
  NAND3_X1 U1729 ( .A1(\SB1_3_15/i0_0 ), .A2(\SB1_3_15/i0_4 ), .A3(
        \SB1_3_15/i1_5 ), .ZN(n1212) );
  NAND3_X1 U1730 ( .A1(\SB2_2_6/i0[8] ), .A2(\SB2_2_6/i3[0] ), .A3(
        \SB2_2_6/i1_5 ), .ZN(\SB2_2_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1731 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i1_7 ), .ZN(\SB1_3_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1733 ( .A1(\SB2_0_20/i0_0 ), .A2(\SB2_0_20/i0_4 ), .A3(
        \SB2_0_20/i1_5 ), .ZN(n885) );
  NAND4_X1 U1734 ( .A1(\SB1_1_3/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_3/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_3/Component_Function_2/NAND4_in[2] ), .A4(n886), .ZN(
        \RI3[1][188] ) );
  NAND3_X1 U1735 ( .A1(\SB1_1_3/i0_0 ), .A2(\SB1_1_3/i0_4 ), .A3(
        \SB1_1_3/i1_5 ), .ZN(n886) );
  NAND3_X1 U1736 ( .A1(\SB2_1_10/i0_4 ), .A2(\RI3[1][126] ), .A3(
        \SB2_1_10/i0[6] ), .ZN(\SB2_1_10/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U1737 ( .A1(\SB1_3_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_3_9/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_3_9/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_8/i0_4 ) );
  NAND3_X1 U1738 ( .A1(\SB4_30/i0_4 ), .A2(\SB4_30/i1[9] ), .A3(\SB4_30/i1_5 ), 
        .ZN(\SB4_30/Component_Function_4/NAND4_in[3] ) );
  XNOR2_X1 U1739 ( .A(n888), .B(n887), .ZN(\RI1[3][129] ) );
  XNOR2_X1 U1740 ( .A(\MC_ARK_ARC_1_2/temp4[129] ), .B(
        \MC_ARK_ARC_1_2/temp1[129] ), .ZN(n887) );
  XNOR2_X1 U1741 ( .A(\MC_ARK_ARC_1_2/temp3[129] ), .B(
        \MC_ARK_ARC_1_2/temp2[129] ), .ZN(n888) );
  INV_X2 U1742 ( .A(\RI1[1][101] ), .ZN(\SB1_1_15/i0_3 ) );
  XNOR2_X1 U1743 ( .A(\MC_ARK_ARC_1_0/temp6[101] ), .B(
        \MC_ARK_ARC_1_0/temp5[101] ), .ZN(\RI1[1][101] ) );
  XNOR2_X1 U1744 ( .A(n890), .B(n889), .ZN(\RI1[3][29] ) );
  XNOR2_X1 U1745 ( .A(\MC_ARK_ARC_1_2/temp1[29] ), .B(
        \MC_ARK_ARC_1_2/temp4[29] ), .ZN(n889) );
  XNOR2_X1 U1746 ( .A(\MC_ARK_ARC_1_2/temp3[29] ), .B(
        \MC_ARK_ARC_1_2/temp2[29] ), .ZN(n890) );
  NAND4_X1 U1748 ( .A1(\SB1_3_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_25/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_25/Component_Function_1/NAND4_in[0] ), .A4(n891), .ZN(
        \RI3[3][61] ) );
  NAND3_X1 U1749 ( .A1(\SB1_3_25/i1_7 ), .A2(\SB1_3_25/i0_4 ), .A3(
        \SB1_3_25/i0[8] ), .ZN(n891) );
  NAND3_X1 U1751 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0_4 ), .A3(
        \SB2_1_10/i0_0 ), .ZN(\SB2_1_10/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U1752 ( .A(n893), .B(n892), .ZN(\RI1[3][125] ) );
  XNOR2_X1 U1753 ( .A(\MC_ARK_ARC_1_2/temp3[125] ), .B(
        \MC_ARK_ARC_1_2/temp4[125] ), .ZN(n892) );
  XNOR2_X1 U1754 ( .A(\MC_ARK_ARC_1_2/temp1[125] ), .B(
        \MC_ARK_ARC_1_2/temp2[125] ), .ZN(n893) );
  NAND3_X1 U1755 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i0[10] ), .A3(
        \SB1_2_5/i0[9] ), .ZN(\SB1_2_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1757 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0[9] ), .A3(
        \SB1_1_10/i0[10] ), .ZN(\SB1_1_10/Component_Function_4/NAND4_in[2] )
         );
  NAND4_X1 U1758 ( .A1(\SB2_1_9/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_9/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_9/Component_Function_2/NAND4_in[1] ), .A4(n894), .ZN(
        \RI5[1][152] ) );
  NAND3_X1 U1761 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i0_4 ), .ZN(\SB1_2_3/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U1762 ( .A1(n1438), .A2(n1235), .A3(
        \SB2_0_20/Component_Function_5/NAND4_in[1] ), .A4(n1263), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[71] ) );
  NAND3_X1 U1763 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0[10] ), .A3(
        \SB1_1_9/i0[9] ), .ZN(\SB1_1_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1764 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0[8] ), .A3(
        \SB1_2_12/i1_7 ), .ZN(\SB1_2_12/Component_Function_1/NAND4_in[1] ) );
  NAND4_X1 U1765 ( .A1(\SB2_2_11/Component_Function_2/NAND4_in[0] ), .A2(n1210), .A3(\SB2_2_11/Component_Function_2/NAND4_in[1] ), .A4(n895), .ZN(
        \RI5[2][140] ) );
  NAND3_X1 U1766 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i1_5 ), .A3(
        \SB2_2_11/i0_0 ), .ZN(n895) );
  NAND4_X1 U1767 ( .A1(\SB1_2_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_2/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_2_2/Component_Function_1/NAND4_in[0] ), .A4(n896), .ZN(
        \RI3[2][7] ) );
  NAND3_X1 U1768 ( .A1(\SB1_2_2/i0[9] ), .A2(\SB1_2_2/i1_5 ), .A3(
        \SB1_2_2/i0[6] ), .ZN(n896) );
  NAND4_X2 U1769 ( .A1(\SB2_1_7/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_7/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_7/Component_Function_0/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[174] ) );
  NAND3_X1 U1770 ( .A1(\SB2_0_10/i0_0 ), .A2(\SB2_0_10/i0[10] ), .A3(
        \SB2_0_10/i0[6] ), .ZN(\SB2_0_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1773 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0[10] ), .A3(
        \SB1_1_15/i0[9] ), .ZN(\SB1_1_15/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U1778 ( .A1(\SB2_2_25/i0[6] ), .A2(n899), .ZN(
        \SB2_2_25/Component_Function_5/NAND4_in[3] ) );
  AND2_X1 U1779 ( .A1(\RI3[2][40] ), .A2(\RI3[2][36] ), .ZN(n899) );
  NAND3_X1 U1781 ( .A1(\SB1_2_12/i3[0] ), .A2(\SB1_2_12/i1_5 ), .A3(
        \SB1_2_12/i0[8] ), .ZN(\SB1_2_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1782 ( .A1(\SB2_2_8/i0_3 ), .A2(\SB2_2_8/i0[6] ), .A3(
        \SB2_2_8/i1[9] ), .ZN(\SB2_2_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1783 ( .A1(\SB3_3/i0_3 ), .A2(\SB3_3/i1[9] ), .A3(\SB3_3/i0_4 ), 
        .ZN(n900) );
  NAND4_X1 U1784 ( .A1(\SB3_3/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_3/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_3/Component_Function_5/NAND4_in[0] ), .A4(n900), .ZN(
        \RI3[4][173] ) );
  NAND3_X1 U1785 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i1[9] ), .A3(
        \RI3[3][64] ), .ZN(\SB2_3_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1787 ( .A1(\SB1_3_21/i1[9] ), .A2(\SB1_3_21/i0_3 ), .A3(
        \SB1_3_21/i0_4 ), .ZN(\SB1_3_21/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U1788 ( .A1(\SB3_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_20/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_20/Component_Function_5/NAND4_in[0] ), .A4(n902), .ZN(
        \RI3[4][71] ) );
  NAND3_X1 U1789 ( .A1(\SB3_20/i1[9] ), .A2(\SB3_20/i0_4 ), .A3(\SB3_20/i0_3 ), 
        .ZN(n902) );
  NAND4_X1 U1790 ( .A1(\SB1_2_9/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_9/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_9/Component_Function_2/NAND4_in[2] ), .A4(n903), .ZN(
        \RI3[2][152] ) );
  NAND4_X1 U1793 ( .A1(\SB4_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_24/Component_Function_1/NAND4_in[0] ), .A4(n904), .ZN(n908) );
  NAND3_X1 U1794 ( .A1(\SB4_24/i0[9] ), .A2(\SB4_24/i1_5 ), .A3(\SB4_24/i0[6] ), .ZN(n904) );
  NAND2_X1 U1797 ( .A1(\SB2_1_3/i0_0 ), .A2(\SB2_1_3/i3[0] ), .ZN(n906) );
  AND2_X1 U1798 ( .A1(\RI3[2][136] ), .A2(\RI3[2][132] ), .ZN(n907) );
  NAND2_X1 U1801 ( .A1(\SB2_2_9/i0[6] ), .A2(n907), .ZN(
        \SB2_2_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1802 ( .A1(\SB1_3_11/i0_0 ), .A2(\SB1_3_11/i0_4 ), .A3(
        \SB1_3_11/i1_5 ), .ZN(\SB1_3_11/Component_Function_2/NAND4_in[3] ) );
  XNOR2_X1 U1803 ( .A(n908), .B(n372), .ZN(Ciphertext[43]) );
  NAND3_X1 U1804 ( .A1(n1664), .A2(\SB1_0_8/i0[10] ), .A3(\SB1_0_8/i0[9] ), 
        .ZN(\SB1_0_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1806 ( .A1(\SB2_3_28/i0[10] ), .A2(\SB2_3_28/i0_0 ), .A3(
        \SB2_3_28/i0[6] ), .ZN(\SB2_3_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1807 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i1_5 ), .A3(
        \SB2_1_29/i1[9] ), .ZN(\SB2_1_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1808 ( .A1(n848), .A2(\SB4_23/i1[9] ), .A3(\SB4_23/i0[6] ), .ZN(
        \SB4_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1809 ( .A1(\SB2_1_25/i0[10] ), .A2(\SB2_1_25/i0_0 ), .A3(
        \SB2_1_25/i0[6] ), .ZN(\SB2_1_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1810 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i0_0 ), .A3(
        \SB1_0_26/i0_4 ), .ZN(\SB1_0_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1811 ( .A1(\SB2_2_9/i0_4 ), .A2(\SB2_2_9/i0_0 ), .A3(
        \SB2_2_9/i0_3 ), .ZN(\SB2_2_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1814 ( .A1(\SB1_0_24/i0_3 ), .A2(\SB1_0_24/i0[9] ), .A3(
        \SB1_0_24/i0[10] ), .ZN(\SB1_0_24/Component_Function_4/NAND4_in[2] )
         );
  NAND4_X1 U1819 ( .A1(\SB2_1_20/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_20/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_20/Component_Function_4/NAND4_in[1] ), .A4(n912), .ZN(
        \RI5[1][76] ) );
  NAND3_X1 U1820 ( .A1(\SB2_1_20/i0_4 ), .A2(\SB2_1_20/i1_5 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(n912) );
  XNOR2_X1 U1825 ( .A(n914), .B(n282), .ZN(Ciphertext[139]) );
  NAND3_X1 U1828 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0_0 ), .A3(
        \SB2_1_17/i0_4 ), .ZN(n915) );
  NAND3_X1 U1832 ( .A1(\SB2_0_0/i0_4 ), .A2(\SB2_0_0/i1_5 ), .A3(
        \SB2_0_0/i0_0 ), .ZN(n917) );
  NAND3_X1 U1835 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0_0 ), .A3(
        \SB1_0_18/i0_4 ), .ZN(\SB1_0_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1836 ( .A1(\SB3_11/i0[6] ), .A2(\SB3_11/i1_5 ), .A3(\SB3_11/i0[9] ), .ZN(\SB3_11/Component_Function_1/NAND4_in[2] ) );
  XNOR2_X1 U1837 ( .A(n919), .B(\MC_ARK_ARC_1_3/temp6[121] ), .ZN(
        \RI1[4][121] ) );
  XNOR2_X1 U1838 ( .A(\MC_ARK_ARC_1_3/temp1[121] ), .B(
        \MC_ARK_ARC_1_3/temp2[121] ), .ZN(n919) );
  NAND4_X1 U1839 ( .A1(\SB2_0_18/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_18/Component_Function_3/NAND4_in[0] ), .A4(n920), .ZN(
        \RI5[0][93] ) );
  NAND3_X1 U1840 ( .A1(\SB2_0_18/i3[0] ), .A2(\SB2_0_18/i1_5 ), .A3(
        \SB2_0_18/i0[8] ), .ZN(n920) );
  NAND3_X1 U1842 ( .A1(\SB2_0_1/i0[6] ), .A2(\SB2_0_1/i0[10] ), .A3(
        \SB2_0_1/i0_0 ), .ZN(\SB2_0_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1843 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i0[10] ), .A3(
        \SB1_1_26/i0[9] ), .ZN(\SB1_1_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1844 ( .A1(\SB1_2_24/i0_0 ), .A2(\SB1_2_24/i0_4 ), .A3(
        \SB1_2_24/i1_5 ), .ZN(n981) );
  XNOR2_X1 U1847 ( .A(\MC_ARK_ARC_1_0/temp2[27] ), .B(
        \MC_ARK_ARC_1_0/temp1[27] ), .ZN(n922) );
  NAND3_X1 U1849 ( .A1(\SB1_2_25/i1[9] ), .A2(\SB1_2_25/i0_3 ), .A3(
        \SB1_2_25/i0_4 ), .ZN(n1266) );
  XNOR2_X1 U1854 ( .A(n925), .B(n924), .ZN(\RI1[1][191] ) );
  XNOR2_X1 U1855 ( .A(\MC_ARK_ARC_1_0/temp4[191] ), .B(
        \MC_ARK_ARC_1_0/temp1[191] ), .ZN(n924) );
  XNOR2_X1 U1856 ( .A(\MC_ARK_ARC_1_0/temp2[191] ), .B(
        \MC_ARK_ARC_1_0/temp3[191] ), .ZN(n925) );
  NAND4_X1 U1857 ( .A1(\SB1_1_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_6/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_6/Component_Function_2/NAND4_in[2] ), .A4(n926), .ZN(
        \RI3[1][170] ) );
  NAND3_X1 U1858 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i1_5 ), .A3(
        \SB1_1_6/i0_4 ), .ZN(n926) );
  NAND3_X1 U1859 ( .A1(\SB2_1_7/i0[10] ), .A2(\SB2_1_7/i0_0 ), .A3(
        \RI3[1][145] ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U1861 ( .A1(\SB2_0_20/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_20/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[81] ) );
  NAND3_X1 U1862 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i0_4 ), .A3(
        \SB2_1_31/i1[9] ), .ZN(\SB2_1_31/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U1863 ( .A1(\SB2_1_11/i0_0 ), .A2(\SB2_1_11/i3[0] ), .ZN(n927) );
  NAND4_X1 U1864 ( .A1(\SB3_16/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_4/NAND4_in[0] ), .A4(n928), .ZN(
        \RI3[4][100] ) );
  NAND3_X1 U1865 ( .A1(\SB3_16/i0[9] ), .A2(\SB3_16/i0_3 ), .A3(
        \SB3_16/i0[10] ), .ZN(n928) );
  NAND3_X1 U1867 ( .A1(\SB4_15/i0_4 ), .A2(\SB4_15/i0[9] ), .A3(\SB4_15/i0[6] ), .ZN(n929) );
  NAND3_X1 U1872 ( .A1(\SB1_2_29/i0[8] ), .A2(\SB1_2_29/i0_4 ), .A3(
        \SB1_2_29/i1_7 ), .ZN(\SB1_2_29/Component_Function_1/NAND4_in[3] ) );
  XNOR2_X1 U1873 ( .A(\MC_ARK_ARC_1_3/temp5[76] ), .B(
        \MC_ARK_ARC_1_3/temp6[76] ), .ZN(\RI1[4][76] ) );
  OR3_X1 U1876 ( .A1(\RI1[1][3] ), .A2(\RI1[1][2] ), .A3(\RI1[1][1] ), .ZN(
        \SB1_1_31/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U1877 ( .A(n934), .B(n329), .ZN(Ciphertext[77]) );
  NAND4_X1 U1878 ( .A1(\SB4_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_19/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_19/Component_Function_5/NAND4_in[0] ), .ZN(n934) );
  NAND3_X1 U1882 ( .A1(\SB1_0_19/i0[6] ), .A2(\SB1_0_19/i0[9] ), .A3(
        \SB1_0_19/i0_4 ), .ZN(\SB1_0_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1883 ( .A1(\SB1_2_17/i0_0 ), .A2(\SB1_2_17/i0_4 ), .A3(
        \SB1_2_17/i1_5 ), .ZN(\SB1_2_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1884 ( .A1(\SB2_2_9/i0[10] ), .A2(\SB2_2_9/i1_5 ), .A3(
        \SB2_2_9/i1[9] ), .ZN(\SB2_2_9/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U1885 ( .A1(\SB1_1_21/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_21/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_1_21/Component_Function_1/NAND4_in[0] ), .A4(n936), .ZN(
        \RI3[1][85] ) );
  NAND3_X1 U1886 ( .A1(\SB1_1_21/i0[9] ), .A2(\SB1_1_21/i1_5 ), .A3(
        \SB1_1_21/i0[6] ), .ZN(n936) );
  NAND3_X1 U1887 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i0_0 ), .A3(
        \SB2_0_27/i0[7] ), .ZN(\SB2_0_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1888 ( .A1(\SB2_2_10/i3[0] ), .A2(\SB2_2_10/i1_5 ), .A3(
        \SB2_2_10/i0[8] ), .ZN(n1214) );
  NAND4_X1 U1889 ( .A1(\SB1_2_14/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_14/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_14/Component_Function_2/NAND4_in[2] ), .A4(n937), .ZN(
        \RI3[2][122] ) );
  NAND3_X1 U1891 ( .A1(\SB2_0_3/i0_0 ), .A2(\SB2_0_3/i1_5 ), .A3(
        \SB2_0_3/i0_4 ), .ZN(n938) );
  NAND4_X1 U1892 ( .A1(\SB1_0_18/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_18/Component_Function_0/NAND4_in[0] ), .A4(n939), .ZN(
        \RI3[0][108] ) );
  NAND3_X1 U1893 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0[10] ), .A3(
        \SB1_0_18/i0_4 ), .ZN(n939) );
  NAND3_X1 U1895 ( .A1(\SB2_2_31/i0_0 ), .A2(\SB2_2_31/i0[10] ), .A3(
        \SB2_2_31/i0[6] ), .ZN(\SB2_2_31/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U1898 ( .A1(\SB1_2_1/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_2_1/Component_Function_5/NAND4_in[3] ), .A4(n940), .ZN(
        \RI3[2][185] ) );
  NAND3_X1 U1899 ( .A1(\SB1_2_1/i0_3 ), .A2(\SB1_2_1/i1[9] ), .A3(
        \SB1_2_1/i0_4 ), .ZN(n940) );
  NAND3_X1 U1900 ( .A1(\SB1_3_12/i0_0 ), .A2(\SB1_3_12/i0_4 ), .A3(
        \SB1_3_12/i1_5 ), .ZN(\SB1_3_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1902 ( .A1(\SB1_2_6/i0_0 ), .A2(\SB1_2_6/i0_4 ), .A3(
        \SB1_2_6/i1_5 ), .ZN(n967) );
  NAND3_X1 U1903 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i0[9] ), .A3(
        \SB1_1_17/i0[10] ), .ZN(\SB1_1_17/Component_Function_4/NAND4_in[2] )
         );
  NAND4_X1 U1904 ( .A1(\SB1_1_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_15/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_15/Component_Function_0/NAND4_in[0] ), .A4(n941), .ZN(
        \RI3[1][126] ) );
  NAND3_X1 U1905 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0[10] ), .A3(
        \SB1_1_15/i0_4 ), .ZN(n941) );
  INV_X1 U1907 ( .A(\RI3[2][158] ), .ZN(\SB2_2_5/i1[9] ) );
  NAND4_X1 U1908 ( .A1(\SB1_2_8/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_8/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_2_8/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_2_8/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[2][158] ) );
  NAND3_X1 U1909 ( .A1(\SB2_1_11/i0[9] ), .A2(\SB2_1_11/i0_3 ), .A3(
        \SB2_1_11/i0[10] ), .ZN(\SB2_1_11/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1910 ( .A1(n866), .A2(\SB4_28/i0_4 ), .A3(\SB4_28/i1[9] ), .ZN(
        \SB4_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1911 ( .A1(\SB2_3_28/i0_3 ), .A2(\SB2_3_28/i0_4 ), .A3(
        \SB2_3_28/i1[9] ), .ZN(\SB2_3_28/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U1912 ( .A1(\SB1_2_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_0/Component_Function_2/NAND4_in[2] ), .A4(n942), .ZN(
        \RI3[2][14] ) );
  NAND3_X1 U1913 ( .A1(\SB1_2_0/i0_0 ), .A2(\SB1_2_0/i0_4 ), .A3(
        \SB1_2_0/i1_5 ), .ZN(n942) );
  NAND3_X1 U1914 ( .A1(\SB1_0_31/i0[9] ), .A2(\SB1_0_31/i0_3 ), .A3(
        \SB1_0_31/i0[10] ), .ZN(\SB1_0_31/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1917 ( .A1(\SB1_0_27/i0[10] ), .A2(\SB1_0_27/i0_3 ), .A3(
        \SB1_0_27/i0[6] ), .ZN(\SB1_0_27/Component_Function_2/NAND4_in[1] ) );
  XNOR2_X1 U1918 ( .A(n945), .B(n944), .ZN(\RI1[1][89] ) );
  XNOR2_X1 U1919 ( .A(\MC_ARK_ARC_1_0/temp1[89] ), .B(
        \MC_ARK_ARC_1_0/temp4[89] ), .ZN(n944) );
  XNOR2_X1 U1920 ( .A(\MC_ARK_ARC_1_0/temp3[89] ), .B(
        \MC_ARK_ARC_1_0/temp2[89] ), .ZN(n945) );
  NAND3_X1 U1921 ( .A1(\SB2_1_8/i0_4 ), .A2(\SB2_1_8/i0_3 ), .A3(
        \SB2_1_8/i1[9] ), .ZN(\SB2_1_8/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U1922 ( .A1(\SB2_2_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_24/Component_Function_0/NAND4_in[0] ), .A4(n946), .ZN(
        \RI5[2][72] ) );
  NAND3_X1 U1923 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0_0 ), .A3(
        \SB2_2_24/i0[7] ), .ZN(n946) );
  NAND2_X1 U1924 ( .A1(\SB2_1_0/i0[6] ), .A2(n948), .ZN(n947) );
  AND2_X1 U1925 ( .A1(\RI3[1][186] ), .A2(\RI3[1][190] ), .ZN(n948) );
  NAND3_X1 U1926 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0[10] ), .A3(
        \SB1_1_6/i0_4 ), .ZN(\SB1_1_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1927 ( .A1(\SB2_1_0/i0_3 ), .A2(\SB2_1_0/i1[9] ), .A3(
        \SB2_1_0/i0[6] ), .ZN(\SB2_1_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1928 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0_4 ), .A3(
        \SB2_1_25/i0_0 ), .ZN(\SB2_1_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1929 ( .A1(\SB1_3_19/i0_0 ), .A2(\SB1_3_19/i0_4 ), .A3(
        \SB1_3_19/i1_5 ), .ZN(\SB1_3_19/Component_Function_2/NAND4_in[3] ) );
  XNOR2_X1 U1930 ( .A(\MC_ARK_ARC_1_1/temp6[63] ), .B(n949), .ZN(\RI1[2][63] )
         );
  XNOR2_X1 U1931 ( .A(\MC_ARK_ARC_1_1/temp2[63] ), .B(
        \MC_ARK_ARC_1_1/temp1[63] ), .ZN(n949) );
  NAND3_X1 U1933 ( .A1(\SB2_1_23/i0[10] ), .A2(\SB2_1_23/i0_0 ), .A3(
        \SB2_1_23/i0[6] ), .ZN(\SB2_1_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1934 ( .A1(\SB1_1_25/i0_3 ), .A2(\SB1_1_25/i0_0 ), .A3(
        \SB1_1_25/i0_4 ), .ZN(\SB1_1_25/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U1935 ( .A(\RI1[2][119] ), .ZN(\SB1_2_12/i0_3 ) );
  XNOR2_X1 U1936 ( .A(\MC_ARK_ARC_1_1/temp5[119] ), .B(
        \MC_ARK_ARC_1_1/temp6[119] ), .ZN(\RI1[2][119] ) );
  NAND2_X1 U1937 ( .A1(\SB2_0_30/i0_0 ), .A2(\SB2_0_30/i3[0] ), .ZN(n950) );
  NAND3_X1 U1939 ( .A1(\SB4_24/i0[6] ), .A2(\SB4_24/i0[8] ), .A3(
        \SB4_24/i0[7] ), .ZN(n951) );
  NAND3_X1 U1940 ( .A1(\SB1_1_25/i0_3 ), .A2(\SB1_1_25/i0[9] ), .A3(
        \SB1_1_25/i0[8] ), .ZN(\SB1_1_25/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U1941 ( .A1(\SB3_1/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_5/NAND4_in[0] ), .A4(n952), .ZN(
        \RI3[4][185] ) );
  NAND3_X1 U1942 ( .A1(\SB3_1/i1[9] ), .A2(\SB3_1/i0_3 ), .A3(\SB3_1/i0_4 ), 
        .ZN(n952) );
  NAND3_X1 U1945 ( .A1(n857), .A2(\SB4_1/i0[10] ), .A3(\SB4_1/i0[9] ), .ZN(
        \SB4_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1947 ( .A1(\SB1_2_17/i0_3 ), .A2(\SB1_2_17/i0[9] ), .A3(
        \SB1_2_17/i0[10] ), .ZN(\SB1_2_17/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1948 ( .A1(\SB2_1_18/i0_4 ), .A2(\SB2_1_18/i0[9] ), .A3(
        \SB2_1_18/i0[6] ), .ZN(\SB2_1_18/Component_Function_5/NAND4_in[3] ) );
  XNOR2_X1 U1949 ( .A(n954), .B(n955), .ZN(\RI1[2][17] ) );
  XNOR2_X1 U1950 ( .A(\MC_ARK_ARC_1_1/temp2[17] ), .B(
        \MC_ARK_ARC_1_1/temp4[17] ), .ZN(n954) );
  XNOR2_X1 U1951 ( .A(\MC_ARK_ARC_1_1/temp3[17] ), .B(
        \MC_ARK_ARC_1_1/temp1[17] ), .ZN(n955) );
  NAND3_X1 U1952 ( .A1(\SB1_2_13/i1_7 ), .A2(\SB1_2_13/i0_4 ), .A3(
        \SB1_2_13/i0[8] ), .ZN(\SB1_2_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1953 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i1_5 ), .A3(
        \SB1_1_29/i0_4 ), .ZN(\SB1_1_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1954 ( .A1(n1649), .A2(\SB1_2_19/i0_0 ), .A3(\SB1_2_19/i0_4 ), 
        .ZN(\SB1_2_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1955 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i0_4 ), .A3(
        \SB2_3_24/i1[9] ), .ZN(\SB2_3_24/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1956 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i0_3 ), .A3(
        \SB2_1_3/i0_0 ), .ZN(\SB2_1_3/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U1957 ( .A1(\SB2_2_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_10/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_10/Component_Function_1/NAND4_in[0] ), .A4(n956), .ZN(
        \RI5[2][151] ) );
  NAND3_X1 U1958 ( .A1(\SB2_2_10/i0_4 ), .A2(\SB2_2_10/i1_7 ), .A3(
        \SB2_2_10/i0[8] ), .ZN(n956) );
  NAND4_X1 U1959 ( .A1(\SB1_1_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_30/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_30/Component_Function_1/NAND4_in[0] ), .A4(n957), .ZN(
        \RI3[1][31] ) );
  NAND3_X1 U1960 ( .A1(\SB1_1_30/i1_7 ), .A2(\SB1_1_30/i0_4 ), .A3(
        \SB1_1_30/i0[8] ), .ZN(n957) );
  NAND3_X1 U1961 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0_4 ), .A3(
        \SB2_1_9/i0_0 ), .ZN(\SB2_1_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1962 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i0[9] ), .A3(
        \SB1_1_19/i0[10] ), .ZN(\SB1_1_19/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1963 ( .A1(\SB1_0_14/i0[7] ), .A2(\SB1_0_14/i0_0 ), .A3(n862), 
        .ZN(\SB1_0_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1964 ( .A1(\SB2_2_20/i0_0 ), .A2(\SB2_2_20/i0[10] ), .A3(
        \SB2_2_20/i0[6] ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1965 ( .A1(\SB2_1_0/i0_4 ), .A2(\SB2_1_0/i0_3 ), .A3(
        \SB2_1_0/i1[9] ), .ZN(\SB2_1_0/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U1968 ( .A(n958), .B(n363), .ZN(Ciphertext[17]) );
  NAND4_X1 U1969 ( .A1(\SB4_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_29/Component_Function_5/NAND4_in[1] ), .A3(n1002), .A4(
        \SB4_29/Component_Function_5/NAND4_in[0] ), .ZN(n958) );
  NAND3_X1 U1970 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0_0 ), .A3(
        \SB2_2_14/i0[7] ), .ZN(\SB2_2_14/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U1971 ( .A1(\SB2_1_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_6/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_6/Component_Function_2/NAND4_in[1] ), .A4(n959), .ZN(
        \RI5[1][170] ) );
  NAND3_X1 U1972 ( .A1(\SB2_1_6/i0_0 ), .A2(\SB2_1_6/i1_5 ), .A3(\RI3[1][154] ), .ZN(n959) );
  NAND3_X1 U1973 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0[7] ), .A3(\SB3_2/i0_0 ), 
        .ZN(n960) );
  NAND3_X1 U1974 ( .A1(\SB2_2_1/i3[0] ), .A2(\SB2_2_1/i1_5 ), .A3(
        \SB2_2_1/i0[8] ), .ZN(n961) );
  NAND3_X1 U1975 ( .A1(\SB2_1_12/i0_4 ), .A2(\SB2_1_12/i0[9] ), .A3(
        \SB2_1_12/i0[6] ), .ZN(\SB2_1_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1976 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0[9] ), .A3(
        \SB1_1_13/i0[10] ), .ZN(\SB1_1_13/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1977 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i0[10] ), .A3(
        \SB1_1_3/i0[9] ), .ZN(\SB1_1_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1978 ( .A1(\SB1_2_22/i0_0 ), .A2(\SB1_2_22/i0_4 ), .A3(
        \SB1_2_22/i1_5 ), .ZN(\SB1_2_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1979 ( .A1(\SB2_1_14/i0[10] ), .A2(\SB2_1_14/i1_5 ), .A3(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1983 ( .A1(\SB1_1_17/i0_4 ), .A2(\SB1_1_17/i0_0 ), .A3(
        \SB1_1_17/i1_5 ), .ZN(n963) );
  NAND4_X1 U1984 ( .A1(\SB1_1_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_1_12/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_1_12/Component_Function_0/NAND4_in[1] ), .A4(n964), .ZN(
        \RI3[1][144] ) );
  NAND3_X1 U1985 ( .A1(\SB1_1_12/i0_3 ), .A2(\SB1_1_12/i0[10] ), .A3(
        \SB1_1_12/i0_4 ), .ZN(n964) );
  NAND3_X1 U1986 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i0[10] ), .A3(
        \SB2_0_27/i0[9] ), .ZN(n965) );
  NAND3_X1 U1987 ( .A1(\SB1_2_21/i1[9] ), .A2(\SB1_2_21/i0[10] ), .A3(
        \SB1_2_21/i1_7 ), .ZN(\SB1_2_21/Component_Function_3/NAND4_in[2] ) );
  XNOR2_X1 U1988 ( .A(n966), .B(n252), .ZN(Ciphertext[61]) );
  NAND3_X1 U1989 ( .A1(\SB2_1_29/i0[8] ), .A2(\SB2_1_29/i3[0] ), .A3(
        \SB2_1_29/i1_5 ), .ZN(n1252) );
  NAND3_X1 U1990 ( .A1(\SB1_1_31/i0_3 ), .A2(\SB1_1_31/i0[9] ), .A3(
        \SB1_1_31/i0[8] ), .ZN(\SB1_1_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1991 ( .A1(\SB2_1_29/i0[9] ), .A2(\SB2_1_29/i0_3 ), .A3(
        \SB2_1_29/i0[8] ), .ZN(\SB2_1_29/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U1992 ( .A1(\SB1_2_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_6/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_6/Component_Function_2/NAND4_in[2] ), .A4(n967), .ZN(
        \RI3[2][170] ) );
  XNOR2_X1 U1998 ( .A(n970), .B(n413), .ZN(Ciphertext[69]) );
  NAND3_X1 U1999 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0_0 ), .A3(n548), .ZN(
        \SB4_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2002 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i0_4 ), .A3(
        \SB2_0_27/i1[9] ), .ZN(\SB2_0_27/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2005 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0_4 ), .A3(
        \SB2_1_4/i0_0 ), .ZN(\SB2_1_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2006 ( .A1(\SB2_3_18/i0[10] ), .A2(\SB2_3_18/i0_0 ), .A3(
        \SB2_3_18/i0[6] ), .ZN(\SB2_3_18/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U2007 ( .A(\RI1[1][77] ), .ZN(\SB1_1_19/i0_3 ) );
  NAND4_X2 U2008 ( .A1(\SB2_1_19/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_19/Component_Function_2/NAND4_in[1] ), .A3(n1134), .A4(
        \SB2_1_19/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[92] ) );
  NAND4_X1 U2009 ( .A1(\SB2_2_11/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_11/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_11/Component_Function_4/NAND4_in[1] ), .A4(n972), .ZN(
        \RI5[2][130] ) );
  NAND3_X1 U2010 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i1_5 ), .A3(
        \SB2_2_11/i1[9] ), .ZN(n972) );
  NAND4_X1 U2011 ( .A1(\SB1_2_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_19/Component_Function_5/NAND4_in[0] ), .A4(n973), .ZN(
        \RI3[2][77] ) );
  NAND3_X1 U2012 ( .A1(\SB1_2_19/i0_3 ), .A2(\SB1_2_19/i1[9] ), .A3(
        \SB1_2_19/i0_4 ), .ZN(n973) );
  NAND3_X1 U2013 ( .A1(n814), .A2(\SB1_2_29/i1_7 ), .A3(\SB1_2_29/i0[8] ), 
        .ZN(\SB1_2_29/Component_Function_1/NAND4_in[1] ) );
  XNOR2_X1 U2014 ( .A(n975), .B(n974), .ZN(\RI1[3][149] ) );
  XNOR2_X1 U2015 ( .A(\MC_ARK_ARC_1_2/temp1[149] ), .B(
        \MC_ARK_ARC_1_2/temp4[149] ), .ZN(n974) );
  XNOR2_X1 U2016 ( .A(\MC_ARK_ARC_1_2/temp2[149] ), .B(
        \MC_ARK_ARC_1_2/temp3[149] ), .ZN(n975) );
  NAND3_X1 U2017 ( .A1(n857), .A2(\SB4_1/i1[9] ), .A3(\SB4_1/i0[6] ), .ZN(
        \SB4_1/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U2018 ( .A1(\SB1_2_25/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_25/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_25/Component_Function_2/NAND4_in[2] ), .A4(n976), .ZN(
        \RI3[2][56] ) );
  NAND4_X1 U2019 ( .A1(\SB1_2_19/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_19/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_19/Component_Function_4/NAND4_in[3] ), .A4(n977), .ZN(
        \RI3[2][82] ) );
  NAND3_X1 U2020 ( .A1(\SB1_2_19/i0_3 ), .A2(\SB1_2_19/i0[9] ), .A3(
        \SB1_2_19/i0[10] ), .ZN(n977) );
  NAND4_X1 U2021 ( .A1(\SB1_3_7/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_7/Component_Function_5/NAND4_in[0] ), .A4(n978), .ZN(
        \RI3[3][149] ) );
  NAND3_X1 U2022 ( .A1(n859), .A2(\SB4_3/i0_4 ), .A3(\SB4_3/i1[9] ), .ZN(
        \SB4_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2025 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i0[10] ), .A3(
        \SB1_2_14/i0_4 ), .ZN(\SB1_2_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2026 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i0[9] ), .A3(
        \SB1_1_21/i0[8] ), .ZN(\SB1_1_21/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U2027 ( .A1(\SB3_23/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_23/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_23/Component_Function_5/NAND4_in[0] ), .A4(n980), .ZN(
        \RI3[4][53] ) );
  NAND3_X1 U2028 ( .A1(\SB3_23/i1[9] ), .A2(\SB3_23/i0_3 ), .A3(\SB3_23/i0_4 ), 
        .ZN(n980) );
  NAND3_X1 U2029 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0[9] ), .A3(
        \SB2_1_17/i0[8] ), .ZN(\SB2_1_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2030 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i0_0 ), .A3(
        \SB1_1_19/i0_4 ), .ZN(\SB1_1_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2031 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i0_3 ), .A3(
        \SB2_2_11/i1[9] ), .ZN(\SB2_2_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2032 ( .A1(\SB2_0_15/i0_0 ), .A2(\SB2_0_15/i0[7] ), .A3(
        \SB2_0_15/i0_3 ), .ZN(\SB2_0_15/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U2033 ( .A1(\SB1_2_24/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_24/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_24/Component_Function_2/NAND4_in[2] ), .A4(n981), .ZN(
        \RI3[2][62] ) );
  NAND4_X2 U2034 ( .A1(\SB2_0_4/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_0_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_0_4/Component_Function_2/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[182] ) );
  NAND3_X1 U2035 ( .A1(\SB2_1_16/i0_4 ), .A2(\RI3[1][90] ), .A3(
        \SB2_1_16/i0[6] ), .ZN(\SB2_1_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2036 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i1_7 ), .A3(
        \SB2_1_2/i0[8] ), .ZN(\SB2_1_2/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U2037 ( .A1(\SB2_0_15/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_15/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_15/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[111] ) );
  XNOR2_X1 U2041 ( .A(\MC_ARK_ARC_1_1/temp1[89] ), .B(
        \MC_ARK_ARC_1_1/temp3[89] ), .ZN(n984) );
  NAND4_X1 U2044 ( .A1(\SB2_2_18/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_18/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_18/Component_Function_1/NAND4_in[0] ), .A4(n986), .ZN(
        \RI5[2][103] ) );
  NAND3_X1 U2045 ( .A1(\SB2_2_18/i0[9] ), .A2(\SB2_2_18/i1_5 ), .A3(
        \SB2_2_18/i0[6] ), .ZN(n986) );
  NAND3_X1 U2046 ( .A1(\SB2_1_17/i0_0 ), .A2(\SB2_1_17/i0[10] ), .A3(
        \SB2_1_17/i0[6] ), .ZN(\SB2_1_17/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U2047 ( .A(n987), .B(n195), .ZN(Ciphertext[56]) );
  NAND3_X1 U2048 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0_4 ), .A3(
        \SB2_1_10/i1[9] ), .ZN(n988) );
  NAND3_X1 U2054 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0_0 ), .A3(\SB4_28/i0[7] ), 
        .ZN(\SB4_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2055 ( .A1(\SB3_28/i0[7] ), .A2(\SB3_28/i0_0 ), .A3(\SB3_28/i0_3 ), 
        .ZN(\SB3_28/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U2056 ( .A(n991), .B(\MC_ARK_ARC_1_2/temp5[59] ), .ZN(\RI1[3][59] )
         );
  XNOR2_X1 U2057 ( .A(\MC_ARK_ARC_1_2/temp4[59] ), .B(
        \MC_ARK_ARC_1_2/temp3[59] ), .ZN(n991) );
  XNOR2_X1 U2058 ( .A(\MC_ARK_ARC_1_2/temp3[14] ), .B(
        \MC_ARK_ARC_1_2/temp4[14] ), .ZN(n992) );
  NAND3_X1 U2059 ( .A1(n2106), .A2(\SB4_31/i1[9] ), .A3(\SB4_31/i0[6] ), .ZN(
        \SB4_31/Component_Function_3/NAND4_in[0] ) );
  NAND4_X4 U2060 ( .A1(n1276), .A2(\SB2_3_5/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_3_5/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[161] ) );
  NAND4_X1 U2062 ( .A1(\SB2_2_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_14/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_14/Component_Function_1/NAND4_in[0] ), .A4(n993), .ZN(
        \RI5[2][127] ) );
  NAND3_X1 U2063 ( .A1(\SB2_2_14/i0_4 ), .A2(\SB2_2_14/i1_7 ), .A3(
        \SB2_2_14/i0[8] ), .ZN(n993) );
  NAND4_X2 U2064 ( .A1(\SB1_3_16/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_16/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_3_16/Component_Function_4/NAND4_in[2] ), .ZN(\SB2_3_15/i0_4 ) );
  NAND3_X1 U2066 ( .A1(\SB4_13/i0_4 ), .A2(\SB4_13/i1[9] ), .A3(\SB4_13/i1_5 ), 
        .ZN(\SB4_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2067 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0_4 ), .A3(
        \SB2_3_15/i1[9] ), .ZN(n1280) );
  NAND3_X1 U2068 ( .A1(\SB4_14/i0_3 ), .A2(n799), .A3(\SB4_14/i1[9] ), .ZN(
        \SB4_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2069 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i0[10] ), .A3(
        \SB1_1_21/i0_4 ), .ZN(\SB1_1_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2071 ( .A1(\SB2_1_13/i0_4 ), .A2(\SB2_1_13/i0_3 ), .A3(
        \SB2_1_13/i1[9] ), .ZN(\SB2_1_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2072 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0_4 ), .A3(
        \SB2_2_7/i1[9] ), .ZN(\SB2_2_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2073 ( .A1(\SB3_31/i1[9] ), .A2(\SB3_31/i0_3 ), .A3(\SB3_31/i0_4 ), 
        .ZN(\SB3_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2074 ( .A1(\SB1_3_25/i0_0 ), .A2(\SB1_3_25/i0_4 ), .A3(
        \SB1_3_25/i1_5 ), .ZN(n1191) );
  NAND3_X1 U2077 ( .A1(\SB3_4/i0[9] ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0[10] ), 
        .ZN(\SB3_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2078 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0_4 ), .A3(
        \SB2_2_16/i1[9] ), .ZN(n996) );
  NAND3_X1 U2079 ( .A1(\SB2_3_9/i0_4 ), .A2(n546), .A3(\SB2_3_9/i0[6] ), .ZN(
        \SB2_3_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2081 ( .A1(\SB4_3/i0_4 ), .A2(\SB4_3/i1[9] ), .A3(\SB4_3/i1_5 ), 
        .ZN(\SB4_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2082 ( .A1(\SB1_2_20/i0_0 ), .A2(\SB1_2_20/i0_4 ), .A3(
        \SB1_2_20/i1_5 ), .ZN(\SB1_2_20/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U2084 ( .A1(\SB1_1_15/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_1_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_5/NAND4_in[0] ), .A4(n997), .ZN(
        \RI3[1][101] ) );
  NAND3_X1 U2085 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i1[9] ), .A3(
        \SB1_1_15/i0_4 ), .ZN(n997) );
  XNOR2_X1 U2086 ( .A(n999), .B(n998), .ZN(\RI1[4][5] ) );
  XNOR2_X1 U2087 ( .A(\MC_ARK_ARC_1_3/temp4[5] ), .B(\MC_ARK_ARC_1_3/temp1[5] ), .ZN(n998) );
  XNOR2_X1 U2088 ( .A(\MC_ARK_ARC_1_3/temp3[5] ), .B(\MC_ARK_ARC_1_3/temp2[5] ), .ZN(n999) );
  NAND4_X1 U2089 ( .A1(\SB2_3_20/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_3_20/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_5/NAND4_in[0] ), .A4(n1000), .ZN(
        \RI5[3][71] ) );
  NAND3_X1 U2090 ( .A1(\SB2_3_20/i0_3 ), .A2(\SB2_3_20/i0_4 ), .A3(
        \SB2_3_20/i1[9] ), .ZN(n1000) );
  NAND4_X1 U2091 ( .A1(\SB2_3_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_5/NAND4_in[0] ), .A4(n1001), .ZN(
        \RI5[3][23] ) );
  NAND3_X1 U2092 ( .A1(\SB2_3_28/i0[9] ), .A2(\SB2_3_28/i0_4 ), .A3(
        \RI3[3][19] ), .ZN(n1001) );
  NAND3_X1 U2093 ( .A1(n2131), .A2(n790), .A3(n791), .ZN(n1002) );
  XNOR2_X1 U2094 ( .A(n1003), .B(n239), .ZN(Ciphertext[173]) );
  NAND3_X1 U2096 ( .A1(n780), .A2(\SB4_27/i1[9] ), .A3(\SB4_27/i1_5 ), .ZN(
        \SB4_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2099 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i0_0 ), .A3(
        \SB1_2_24/i0[6] ), .ZN(\SB1_2_24/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2100 ( .A1(\SB1_3_6/i0_0 ), .A2(\SB1_3_6/i0_4 ), .A3(
        \SB1_3_6/i1_5 ), .ZN(\SB1_3_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2101 ( .A1(\SB2_2_15/i0_4 ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(\SB2_2_15/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2102 ( .A1(n873), .A2(\SB1_0_19/i0[9] ), .A3(\SB1_0_19/i0[10] ), 
        .ZN(\SB1_0_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2103 ( .A1(\SB1_2_10/i0_3 ), .A2(\SB1_2_10/i0[10] ), .A3(
        \SB1_2_10/i0[9] ), .ZN(\SB1_2_10/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U2104 ( .A1(\SB2_2_9/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_9/Component_Function_5/NAND4_in[1] ), .A3(n1005), .A4(
        \SB2_2_9/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[137] ) );
  NAND2_X1 U2105 ( .A1(\SB2_2_9/i0_0 ), .A2(\SB2_2_9/i3[0] ), .ZN(n1005) );
  NAND3_X1 U2107 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0[7] ), .A3(
        \SB1_1_9/i0_0 ), .ZN(\SB1_1_9/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U2108 ( .A1(\SB1_3_9/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_9/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_9/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_3_9/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[3][152] ) );
  XNOR2_X1 U2109 ( .A(n1007), .B(n1006), .ZN(\RI1[4][83] ) );
  XNOR2_X1 U2110 ( .A(\MC_ARK_ARC_1_3/temp2[83] ), .B(
        \MC_ARK_ARC_1_3/temp4[83] ), .ZN(n1006) );
  XNOR2_X1 U2111 ( .A(\MC_ARK_ARC_1_3/temp3[83] ), .B(
        \MC_ARK_ARC_1_3/temp1[83] ), .ZN(n1007) );
  NAND3_X1 U2112 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i0[9] ), .A3(
        \SB1_3_25/i0[8] ), .ZN(\SB1_3_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2114 ( .A1(\SB1_3_23/i0[8] ), .A2(\SB1_3_23/i0[9] ), .A3(
        \SB1_3_23/i0_0 ), .ZN(\SB1_3_23/Component_Function_4/NAND4_in[0] ) );
  XNOR2_X1 U2115 ( .A(\MC_ARK_ARC_1_2/temp5[50] ), .B(n1008), .ZN(\RI1[3][50] ) );
  XNOR2_X1 U2116 ( .A(\MC_ARK_ARC_1_2/temp3[50] ), .B(
        \MC_ARK_ARC_1_2/temp4[50] ), .ZN(n1008) );
  NAND3_X1 U2117 ( .A1(\SB2_1_16/i0[9] ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0[8] ), .ZN(n1009) );
  NAND3_X1 U2118 ( .A1(\SB3_4/i0_4 ), .A2(\SB3_4/i1[9] ), .A3(\SB3_4/i0_3 ), 
        .ZN(\SB3_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2120 ( .A1(\SB1_0_24/i0_3 ), .A2(\SB1_0_24/i0[9] ), .A3(
        \SB1_0_24/i0[8] ), .ZN(\SB1_0_24/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2122 ( .A(n1011), .B(n1010), .ZN(\RI1[2][143] ) );
  XNOR2_X1 U2123 ( .A(\MC_ARK_ARC_1_1/temp4[143] ), .B(
        \MC_ARK_ARC_1_1/temp2[143] ), .ZN(n1010) );
  XNOR2_X1 U2124 ( .A(\MC_ARK_ARC_1_1/temp1[143] ), .B(
        \MC_ARK_ARC_1_1/temp3[143] ), .ZN(n1011) );
  NAND4_X1 U2125 ( .A1(\SB1_3_12/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_12/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_3_12/Component_Function_3/NAND4_in[0] ), .A4(n1012), .ZN(
        \RI3[3][129] ) );
  NAND3_X1 U2126 ( .A1(\SB1_3_12/i3[0] ), .A2(\SB1_3_12/i1_5 ), .A3(
        \SB1_3_12/i0[8] ), .ZN(n1012) );
  NAND3_X1 U2130 ( .A1(\SB2_2_23/i1_5 ), .A2(\SB2_2_23/i3[0] ), .A3(
        \SB2_2_23/i0[8] ), .ZN(n1014) );
  NAND4_X1 U2131 ( .A1(\SB2_1_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_0/NAND4_in[0] ), .A4(n1015), .ZN(
        \RI5[1][66] ) );
  NAND3_X1 U2132 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0_0 ), .A3(
        \SB2_1_25/i0[7] ), .ZN(n1015) );
  XNOR2_X1 U2133 ( .A(n1017), .B(n1016), .ZN(\RI1[2][179] ) );
  XNOR2_X1 U2134 ( .A(\MC_ARK_ARC_1_1/temp1[179] ), .B(
        \MC_ARK_ARC_1_1/temp4[179] ), .ZN(n1016) );
  XNOR2_X1 U2135 ( .A(\MC_ARK_ARC_1_1/temp2[179] ), .B(
        \MC_ARK_ARC_1_1/temp3[179] ), .ZN(n1017) );
  NAND3_X1 U2139 ( .A1(\SB2_1_20/i0_4 ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(\SB2_1_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2140 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i0_0 ), .A3(
        \SB2_1_24/i0[6] ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2141 ( .A1(\SB1_2_4/i0_0 ), .A2(\SB1_2_4/i0_4 ), .A3(
        \SB1_2_4/i1_5 ), .ZN(\SB1_2_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2142 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i0_0 ), .A3(
        \SB1_0_13/i0_4 ), .ZN(\SB1_0_13/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2143 ( .A(n1020), .B(\MC_ARK_ARC_1_1/temp5[110] ), .ZN(
        \RI1[2][110] ) );
  XNOR2_X1 U2144 ( .A(\MC_ARK_ARC_1_1/temp3[110] ), .B(
        \MC_ARK_ARC_1_1/temp4[110] ), .ZN(n1020) );
  NAND4_X2 U2149 ( .A1(\SB2_0_3/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_3/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_3/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[183] ) );
  NAND3_X1 U2150 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i1[9] ), .A3(
        \SB2_1_26/i0[6] ), .ZN(\SB2_1_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2151 ( .A1(\SB1_1_5/i0_3 ), .A2(\SB1_1_5/i0[9] ), .A3(
        \SB1_1_5/i0[8] ), .ZN(\SB1_1_5/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2155 ( .A(n1025), .B(n1024), .ZN(\RI1[3][173] ) );
  XNOR2_X1 U2156 ( .A(\MC_ARK_ARC_1_2/temp4[173] ), .B(
        \MC_ARK_ARC_1_2/temp1[173] ), .ZN(n1024) );
  XNOR2_X1 U2157 ( .A(\MC_ARK_ARC_1_2/temp3[173] ), .B(
        \MC_ARK_ARC_1_2/temp2[173] ), .ZN(n1025) );
  NAND3_X1 U2158 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i1[9] ), .A3(\SB4_30/i0[6] ), .ZN(\SB4_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2161 ( .A1(\SB2_1_7/i0[10] ), .A2(\SB2_1_7/i1[9] ), .A3(
        \SB2_1_7/i1_7 ), .ZN(\SB2_1_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2163 ( .A1(\SB2_1_29/i0_4 ), .A2(\SB2_1_29/i0_0 ), .A3(
        \SB2_1_29/i0_3 ), .ZN(n1026) );
  NAND2_X1 U2166 ( .A1(\SB2_2_2/i0_0 ), .A2(\SB2_2_2/i3[0] ), .ZN(n1028) );
  NAND3_X1 U2169 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i0_0 ), .A3(\SB4_30/i0[7] ), 
        .ZN(\SB4_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2170 ( .A1(\SB1_1_5/i0_3 ), .A2(\SB1_1_5/i0[10] ), .A3(
        \SB1_1_5/i0[9] ), .ZN(\SB1_1_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2171 ( .A1(\SB4_28/i0_4 ), .A2(\SB4_28/i1[9] ), .A3(\SB4_28/i1_5 ), 
        .ZN(\SB4_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2172 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i0_4 ), .A3(
        \SB1_0_19/i1[9] ), .ZN(\SB1_0_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2173 ( .A1(\SB2_1_29/i0_3 ), .A2(\SB2_1_29/i0_0 ), .A3(
        \SB2_1_29/i0[7] ), .ZN(\SB2_1_29/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U2174 ( .A(n1030), .B(n304), .ZN(Ciphertext[163]) );
  NAND3_X1 U2176 ( .A1(\SB1_3_13/i0_0 ), .A2(\SB1_3_13/i0_4 ), .A3(
        \SB1_3_13/i1_5 ), .ZN(\SB1_3_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2177 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i0_4 ), .A3(
        \SB1_3_21/i1_5 ), .ZN(\SB1_3_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2179 ( .A1(\SB2_2_5/i0[10] ), .A2(\SB2_2_5/i0_0 ), .A3(
        \SB2_2_5/i0[6] ), .ZN(\SB2_2_5/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U2180 ( .A1(\SB2_2_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_8/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_8/Component_Function_4/NAND4_in[1] ), .A4(n1031), .ZN(
        \RI5[2][148] ) );
  NAND3_X1 U2181 ( .A1(\SB2_2_8/i0_4 ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i1[9] ), .ZN(n1031) );
  NAND3_X1 U2186 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0_4 ), .A3(
        \SB2_1_22/i0_0 ), .ZN(n1032) );
  NAND3_X1 U2187 ( .A1(\SB2_0_30/i0[10] ), .A2(\SB2_0_30/i1_5 ), .A3(
        \SB2_0_30/i1[9] ), .ZN(\SB2_0_30/Component_Function_2/NAND4_in[0] ) );
  XNOR2_X1 U2189 ( .A(n1033), .B(n338), .ZN(Ciphertext[103]) );
  NAND4_X1 U2190 ( .A1(\SB4_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_14/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_14/Component_Function_1/NAND4_in[0] ), .A4(n1255), .ZN(n1033) );
  NAND3_X1 U2191 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i0[10] ), .A3(
        \SB1_1_7/i0_4 ), .ZN(\SB1_1_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2192 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i0_4 ), .A3(
        \SB1_3_27/i1_5 ), .ZN(n1063) );
  NAND3_X1 U2193 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i0_0 ), .A3(
        \SB2_3_11/i0[6] ), .ZN(\SB2_3_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2194 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i0_4 ), .A3(
        \SB1_3_23/i1_5 ), .ZN(\SB1_3_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2195 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0_4 ), .A3(
        \SB2_1_24/i0_0 ), .ZN(\SB2_1_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2196 ( .A1(n1667), .A2(\SB4_4/i1[9] ), .A3(\SB4_4/i0_4 ), .ZN(
        \SB4_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2199 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i0_0 ), .A3(\SB4_6/i0[7] ), 
        .ZN(\SB4_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2201 ( .A1(n819), .A2(\SB3_27/i0_0 ), .A3(\SB3_27/i0[7] ), .ZN(
        n1035) );
  NAND3_X1 U2205 ( .A1(\SB2_2_9/i0_3 ), .A2(\SB2_2_9/i0[9] ), .A3(
        \SB2_2_9/i0[10] ), .ZN(\SB2_2_9/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U2206 ( .A(n1038), .B(\MC_ARK_ARC_1_0/temp6[117] ), .ZN(
        \RI1[1][117] ) );
  XNOR2_X1 U2207 ( .A(\MC_ARK_ARC_1_0/temp2[117] ), .B(
        \MC_ARK_ARC_1_0/temp1[117] ), .ZN(n1038) );
  NAND3_X1 U2208 ( .A1(\SB2_0_15/i0_0 ), .A2(\SB2_0_15/i0_4 ), .A3(
        \SB2_0_15/i0_3 ), .ZN(\SB2_0_15/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2211 ( .A(n1040), .B(n271), .ZN(Ciphertext[72]) );
  NAND4_X1 U2212 ( .A1(\SB4_19/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_19/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_19/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_19/Component_Function_0/NAND4_in[1] ), .ZN(n1040) );
  NAND3_X1 U2214 ( .A1(\SB2_3_15/i0[8] ), .A2(\SB2_3_15/i1_5 ), .A3(
        \SB2_3_15/i3[0] ), .ZN(\SB2_3_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2215 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i1_7 ), .ZN(\SB1_3_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2216 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0[9] ), .A3(
        \SB1_1_16/i0[8] ), .ZN(\SB1_1_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2217 ( .A1(\SB2_2_5/i3[0] ), .A2(\SB2_2_5/i1_5 ), .A3(
        \SB2_2_5/i0[8] ), .ZN(\SB2_2_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2218 ( .A1(\SB4_21/i0[9] ), .A2(\SB4_21/i0_4 ), .A3(\SB4_21/i0[6] ), .ZN(n1041) );
  NAND3_X1 U2219 ( .A1(\SB4_25/i0_4 ), .A2(\SB4_25/i1[9] ), .A3(\SB4_25/i0_3 ), 
        .ZN(\SB4_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2220 ( .A1(\SB2_3_6/i3[0] ), .A2(\SB2_3_6/i1_5 ), .A3(
        \SB2_3_6/i0[8] ), .ZN(\SB2_3_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2223 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i0[10] ), .A3(
        \SB4_25/i0[9] ), .ZN(\SB4_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2224 ( .A1(\SB1_2_25/i0_3 ), .A2(\SB1_2_25/i0[9] ), .A3(
        \SB1_2_25/i0[8] ), .ZN(\SB1_2_25/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U2225 ( .A1(\SB2_0_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_15/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_15/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[101] ) );
  NAND3_X1 U2227 ( .A1(\SB1_2_0/i0_3 ), .A2(\SB1_2_0/i0_4 ), .A3(
        \SB1_2_0/i0[10] ), .ZN(\SB1_2_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2228 ( .A1(\SB2_1_23/i0_3 ), .A2(\RI3[1][48] ), .A3(
        \SB2_1_23/i0[8] ), .ZN(n1283) );
  AND2_X1 U2229 ( .A1(\RI3[2][28] ), .A2(\RI3[2][24] ), .ZN(n1043) );
  NAND2_X1 U2230 ( .A1(\SB2_2_27/i0[6] ), .A2(n1043), .ZN(
        \SB2_2_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2231 ( .A1(\SB2_2_10/i0_4 ), .A2(\SB2_2_10/i0_3 ), .A3(
        \SB2_2_10/i1[9] ), .ZN(\SB2_2_10/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U2232 ( .A1(\SB2_2_27/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_27/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_27/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_27/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[29] ) );
  NAND4_X1 U2233 ( .A1(\SB1_2_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_24/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_2_24/Component_Function_4/NAND4_in[1] ), .A4(n1044), .ZN(
        \RI3[2][52] ) );
  NAND3_X1 U2234 ( .A1(\SB1_2_24/i0_3 ), .A2(\SB1_2_24/i0[10] ), .A3(
        \SB1_2_24/i0[9] ), .ZN(n1044) );
  NAND3_X1 U2236 ( .A1(\SB2_1_14/i0_0 ), .A2(\SB2_1_14/i0[10] ), .A3(
        \SB2_1_14/i0[6] ), .ZN(\SB2_1_14/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2237 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0_0 ), .A3(
        \SB2_1_20/i0[6] ), .ZN(\SB2_1_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2238 ( .A1(\SB1_2_1/i0_3 ), .A2(\SB1_2_1/i0[10] ), .A3(
        \SB1_2_1/i0[9] ), .ZN(\SB1_2_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2239 ( .A1(\SB2_1_8/i0[9] ), .A2(\SB2_1_8/i0_3 ), .A3(
        \SB2_1_8/i0[8] ), .ZN(\SB2_1_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2240 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0_4 ), .A3(
        \SB2_0_21/i1[9] ), .ZN(\SB2_0_21/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U2241 ( .A1(\SB1_3_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_3_19/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_3_19/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_18/i0_4 ) );
  NAND3_X1 U2242 ( .A1(\SB2_3_1/i3[0] ), .A2(\SB2_3_1/i1_5 ), .A3(
        \SB2_3_1/i0[8] ), .ZN(\SB2_3_1/Component_Function_3/NAND4_in[3] ) );
  XNOR2_X1 U2243 ( .A(n1045), .B(n241), .ZN(Ciphertext[63]) );
  NAND3_X1 U2245 ( .A1(\SB2_3_13/i3[0] ), .A2(\SB2_3_13/i1_5 ), .A3(
        \SB2_3_13/i0[8] ), .ZN(\SB2_3_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2246 ( .A1(\SB2_1_20/i3[0] ), .A2(\SB2_1_20/i1_5 ), .A3(
        \SB2_1_20/i0[8] ), .ZN(n1046) );
  NAND3_X1 U2248 ( .A1(\SB2_1_8/i3[0] ), .A2(\SB2_1_8/i1_5 ), .A3(
        \SB2_1_8/i0[8] ), .ZN(n1047) );
  NAND3_X1 U2249 ( .A1(\SB2_2_11/i3[0] ), .A2(\SB2_2_11/i1_5 ), .A3(
        \SB2_2_11/i0[8] ), .ZN(n1048) );
  NAND3_X1 U2250 ( .A1(\SB1_2_29/i1[9] ), .A2(\SB1_2_29/i0[10] ), .A3(
        \SB1_2_29/i1_7 ), .ZN(\SB1_2_29/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U2251 ( .A1(\SB1_1_28/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_28/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_28/Component_Function_4/NAND4_in[3] ), .A4(n1049), .ZN(
        \RI3[1][28] ) );
  NAND3_X1 U2252 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i0[10] ), .A3(
        \SB1_1_28/i0[9] ), .ZN(n1049) );
  NAND4_X1 U2253 ( .A1(\SB2_0_21/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_21/Component_Function_2/NAND4_in[0] ), .A4(n1050), .ZN(
        \RI5[0][80] ) );
  NAND3_X1 U2254 ( .A1(\SB2_0_21/i0_4 ), .A2(\SB2_0_21/i0_0 ), .A3(
        \SB2_0_21/i1_5 ), .ZN(n1050) );
  NAND4_X1 U2256 ( .A1(\SB1_1_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_2/NAND4_in[2] ), .A4(n1051), .ZN(
        \RI3[1][128] ) );
  NAND3_X1 U2257 ( .A1(\SB1_1_13/i0_0 ), .A2(\SB1_1_13/i0_4 ), .A3(
        \SB1_1_13/i1_5 ), .ZN(n1051) );
  NAND3_X1 U2258 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i1_5 ), .A3(
        \SB2_1_3/i1[9] ), .ZN(n1052) );
  NAND4_X1 U2261 ( .A1(\SB1_1_14/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_14/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_14/Component_Function_5/NAND4_in[0] ), .A4(n1054), .ZN(
        \RI3[1][107] ) );
  NAND3_X1 U2262 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i0_4 ), .ZN(n1054) );
  XNOR2_X1 U2264 ( .A(\MC_ARK_ARC_1_1/temp5[39] ), .B(n1055), .ZN(\RI1[2][39] ) );
  XNOR2_X1 U2265 ( .A(\MC_ARK_ARC_1_1/temp3[39] ), .B(
        \MC_ARK_ARC_1_1/temp4[39] ), .ZN(n1055) );
  NAND3_X1 U2266 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0[9] ), .A3(
        \SB1_1_30/i0[10] ), .ZN(\SB1_1_30/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2267 ( .A1(\SB1_1_23/i1_7 ), .A2(\SB1_1_23/i0[10] ), .A3(
        \SB1_1_23/i1[9] ), .ZN(\SB1_1_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2270 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i0[10] ), .A3(
        \SB1_1_28/i0_4 ), .ZN(\SB1_1_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2271 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i0[10] ), .A3(
        \SB1_2_4/i0_4 ), .ZN(\SB1_2_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2272 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0[6] ), .A3(
        \SB2_0_4/i1[9] ), .ZN(n1056) );
  NAND3_X1 U2273 ( .A1(\SB1_3_0/i0_0 ), .A2(\SB1_3_0/i0_4 ), .A3(
        \SB1_3_0/i1_5 ), .ZN(\SB1_3_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2274 ( .A1(\SB2_1_19/i0[10] ), .A2(\SB2_1_19/i1_5 ), .A3(
        \SB2_1_19/i1[9] ), .ZN(\SB2_1_19/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U2275 ( .A1(\SB1_2_11/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_11/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_11/Component_Function_2/NAND4_in[2] ), .A4(n1057), .ZN(
        \RI3[2][140] ) );
  NAND3_X1 U2276 ( .A1(\SB1_2_11/i0_0 ), .A2(\SB1_2_11/i0_4 ), .A3(
        \SB1_2_11/i1_5 ), .ZN(n1057) );
  NAND4_X1 U2277 ( .A1(\SB2_2_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_27/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_27/Component_Function_4/NAND4_in[1] ), .A4(n1058), .ZN(
        \RI5[2][34] ) );
  NAND3_X1 U2278 ( .A1(\SB2_2_27/i0_4 ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB2_2_27/i1[9] ), .ZN(n1058) );
  NAND3_X1 U2279 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0_0 ), .A3(
        \SB2_0_16/i0[7] ), .ZN(\SB2_0_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2280 ( .A1(\SB2_0_31/i0_3 ), .A2(\SB2_0_31/i0_0 ), .A3(
        \SB2_0_31/i0[7] ), .ZN(\SB2_0_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2281 ( .A1(\SB1_1_11/i0[9] ), .A2(\SB1_1_11/i1_5 ), .A3(
        \SB1_1_11/i0[6] ), .ZN(\SB1_1_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2282 ( .A1(\SB2_0_21/i0[10] ), .A2(\SB2_0_21/i0_0 ), .A3(
        \SB2_0_21/i0[6] ), .ZN(\SB2_0_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2283 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i1[9] ), .A3(\SB4_25/i0[6] ), .ZN(\SB4_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2284 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i0_0 ), .A3(
        \SB4_15/i0[6] ), .ZN(n1059) );
  NAND4_X1 U2285 ( .A1(\SB1_3_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_9/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_9/Component_Function_3/NAND4_in[2] ), .A4(n1060), .ZN(
        \RI3[3][147] ) );
  NAND3_X1 U2286 ( .A1(\SB1_3_9/i3[0] ), .A2(\SB1_3_9/i1_5 ), .A3(
        \SB1_3_9/i0[8] ), .ZN(n1060) );
  NAND3_X1 U2287 ( .A1(\SB2_3_28/i0[8] ), .A2(\SB2_3_28/i3[0] ), .A3(
        \SB2_3_28/i1_5 ), .ZN(\SB2_3_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2289 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i0_0 ), .A3(
        \SB2_1_31/i0[7] ), .ZN(\SB2_1_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2291 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[8] ), .A3(
        \SB2_2_22/i0[9] ), .ZN(\SB2_2_22/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2292 ( .A(\MC_ARK_ARC_1_0/temp5[149] ), .B(n1061), .ZN(
        \RI1[1][149] ) );
  XNOR2_X1 U2293 ( .A(\MC_ARK_ARC_1_0/temp3[149] ), .B(
        \MC_ARK_ARC_1_0/temp4[149] ), .ZN(n1061) );
  NAND3_X1 U2295 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i1[9] ), .A3(\SB4_7/i1_5 ), 
        .ZN(n1062) );
  NAND3_X1 U2296 ( .A1(n2136), .A2(\SB1_0_6/i0[7] ), .A3(\SB1_0_6/i0_0 ), .ZN(
        \SB1_0_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2297 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0_4 ), .A3(
        \SB2_2_1/i1[9] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2298 ( .A1(\SB2_2_31/i0_4 ), .A2(\SB2_2_31/i1_7 ), .A3(
        \SB2_2_31/i0[8] ), .ZN(\SB2_2_31/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 U2299 ( .A1(\SB1_3_27/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_27/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_27/Component_Function_2/NAND4_in[2] ), .A4(n1063), .ZN(
        \RI3[3][44] ) );
  NAND3_X1 U2300 ( .A1(n2149), .A2(\SB1_1_4/i0[8] ), .A3(\SB1_1_4/i1_7 ), .ZN(
        \SB1_1_4/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2301 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0[9] ), .A3(
        \SB2_2_12/i0[8] ), .ZN(\SB2_2_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2302 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i1[9] ), .A3(
        \SB2_0_4/i1_7 ), .ZN(n1064) );
  NAND3_X1 U2303 ( .A1(\SB2_2_24/i1_5 ), .A2(\SB2_2_24/i3[0] ), .A3(
        \SB2_2_24/i0[8] ), .ZN(n1065) );
  XNOR2_X1 U2304 ( .A(n1066), .B(n1067), .ZN(\RI1[2][83] ) );
  XNOR2_X1 U2305 ( .A(\MC_ARK_ARC_1_1/temp3[83] ), .B(
        \MC_ARK_ARC_1_1/temp4[83] ), .ZN(n1066) );
  XNOR2_X1 U2306 ( .A(\MC_ARK_ARC_1_1/temp1[83] ), .B(
        \MC_ARK_ARC_1_1/temp2[83] ), .ZN(n1067) );
  NAND3_X1 U2311 ( .A1(\SB4_24/i0_0 ), .A2(\SB4_24/i3[0] ), .A3(\SB4_24/i1_7 ), 
        .ZN(\SB4_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2314 ( .A1(\SB3_27/i0_0 ), .A2(\SB3_27/i1_5 ), .A3(\SB3_27/i0_4 ), 
        .ZN(\SB3_27/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U2315 ( .A1(\SB1_2_26/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_26/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_26/Component_Function_0/NAND4_in[1] ), .A4(n1071), .ZN(
        \RI3[2][60] ) );
  NAND3_X1 U2316 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0[10] ), .A3(
        \SB1_2_26/i0_4 ), .ZN(n1071) );
  NAND3_X1 U2317 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i1[9] ), .A3(
        \SB1_2_16/i0_4 ), .ZN(n1087) );
  NAND3_X1 U2318 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i0[9] ), .A3(
        \SB2_0_27/i0[8] ), .ZN(\SB2_0_27/Component_Function_2/NAND4_in[2] ) );
  AND2_X1 U2319 ( .A1(\RI3[2][160] ), .A2(\RI3[2][156] ), .ZN(n1113) );
  NAND3_X1 U2320 ( .A1(\SB2_2_17/i0_4 ), .A2(\SB2_2_17/i1_5 ), .A3(
        \SB2_2_17/i0_0 ), .ZN(\SB2_2_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2321 ( .A1(\SB2_2_20/i0_4 ), .A2(\SB2_2_20/i0[9] ), .A3(
        \SB2_2_20/i0[6] ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2322 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0_4 ), .A3(
        \SB2_2_16/i0_0 ), .ZN(\SB2_2_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2323 ( .A1(\SB2_2_3/i0[10] ), .A2(\SB2_2_3/i0_0 ), .A3(
        \SB2_2_3/i0[6] ), .ZN(\SB2_2_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2324 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0[9] ), .A3(
        \SB1_2_21/i0[10] ), .ZN(\SB1_2_21/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2325 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i0[9] ), .ZN(\SB1_2_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2327 ( .A1(\RI3[2][178] ), .A2(\SB2_2_2/i1_5 ), .A3(\SB2_2_2/i0_0 ), .ZN(n1072) );
  NAND4_X1 U2328 ( .A1(\SB1_3_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_24/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_3_24/Component_Function_5/NAND4_in[3] ), .A4(n1073), .ZN(
        \RI3[3][47] ) );
  NAND3_X1 U2329 ( .A1(\SB1_3_24/i0_3 ), .A2(\SB1_3_24/i1[9] ), .A3(
        \SB1_3_24/i0_4 ), .ZN(n1073) );
  NAND3_X1 U2330 ( .A1(\SB1_2_10/i0_3 ), .A2(\SB1_2_10/i0[9] ), .A3(
        \SB1_2_10/i0[8] ), .ZN(\SB1_2_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2331 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0[9] ), .A3(
        \SB1_2_21/i0[8] ), .ZN(\SB1_2_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2333 ( .A1(\SB2_3_17/i0_4 ), .A2(\RI3[3][84] ), .A3(
        \SB2_3_17/i0[6] ), .ZN(n1074) );
  NAND4_X1 U2334 ( .A1(\SB1_1_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_24/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_24/Component_Function_1/NAND4_in[0] ), .A4(n1075), .ZN(
        \RI3[1][67] ) );
  NAND3_X1 U2335 ( .A1(\SB1_1_24/i1_7 ), .A2(\SB1_1_24/i0_4 ), .A3(
        \SB1_1_24/i0[8] ), .ZN(n1075) );
  NAND4_X1 U2336 ( .A1(\SB1_3_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_5/NAND4_in[0] ), .A4(n1076), .ZN(
        \RI3[3][155] ) );
  NAND3_X1 U2337 ( .A1(\SB1_3_6/i0_4 ), .A2(\SB1_3_6/i0[6] ), .A3(
        \SB1_3_6/i0[9] ), .ZN(n1076) );
  NAND3_X1 U2338 ( .A1(\SB2_2_10/i0_3 ), .A2(\SB2_2_10/i1[9] ), .A3(
        \SB2_2_10/i0[6] ), .ZN(\SB2_2_10/Component_Function_3/NAND4_in[0] ) );
  XNOR2_X1 U2339 ( .A(n1077), .B(\MC_ARK_ARC_1_2/temp6[81] ), .ZN(\RI1[3][81] ) );
  XNOR2_X1 U2340 ( .A(\MC_ARK_ARC_1_2/temp1[81] ), .B(
        \MC_ARK_ARC_1_2/temp2[81] ), .ZN(n1077) );
  NAND3_X1 U2343 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[9] ), .A3(
        \SB2_2_16/i0[10] ), .ZN(\SB2_2_16/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2344 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i0[10] ), .A3(
        \SB1_2_18/i0[9] ), .ZN(\SB1_2_18/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U2345 ( .A1(\SB2_1_14/i0[6] ), .A2(n1079), .ZN(
        \SB2_1_14/Component_Function_5/NAND4_in[3] ) );
  AND2_X1 U2346 ( .A1(\RI3[1][106] ), .A2(\RI3[1][102] ), .ZN(n1079) );
  NAND3_X1 U2347 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0_0 ), .A3(
        \SB2_0_21/i0[7] ), .ZN(\SB2_0_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2348 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i0_3 ), .A3(
        \SB1_3_24/i0[9] ), .ZN(\SB1_3_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2350 ( .A1(\SB1_2_30/i0[9] ), .A2(\SB1_2_30/i0_3 ), .A3(
        \SB1_2_30/i0[10] ), .ZN(\SB1_2_30/Component_Function_4/NAND4_in[2] )
         );
  INV_X1 U2351 ( .A(\RI3[1][86] ), .ZN(\SB2_1_17/i1[9] ) );
  NAND4_X1 U2352 ( .A1(\SB2_1_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_2/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_2/Component_Function_2/NAND4_in[1] ), .A4(n1080), .ZN(
        \RI5[1][2] ) );
  NAND3_X1 U2353 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i0_0 ), .A3(
        \SB2_1_2/i1_5 ), .ZN(n1080) );
  NAND4_X1 U2354 ( .A1(\SB1_0_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_31/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_0_31/Component_Function_2/NAND4_in[0] ), .A4(n1081), .ZN(
        \RI3[0][20] ) );
  NAND3_X1 U2355 ( .A1(\SB1_0_31/i0_0 ), .A2(\SB1_0_31/i0_4 ), .A3(
        \SB1_0_31/i1_5 ), .ZN(n1081) );
  NAND4_X1 U2358 ( .A1(\SB1_3_1/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_1/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_1/Component_Function_5/NAND4_in[0] ), .A4(n1083), .ZN(
        \RI3[3][185] ) );
  NAND3_X1 U2359 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i1[9] ), .A3(
        \SB1_3_1/i0_4 ), .ZN(n1083) );
  NAND3_X1 U2360 ( .A1(\SB4_21/i0_0 ), .A2(\SB4_21/i1_7 ), .A3(\SB4_21/i3[0] ), 
        .ZN(\SB4_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2361 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0_0 ), .A3(\SB4_15/i0[7] ), 
        .ZN(\SB4_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2362 ( .A1(\SB1_0_1/i0_3 ), .A2(\SB1_0_1/i0_4 ), .A3(
        \SB1_0_1/i1[9] ), .ZN(\SB1_0_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2365 ( .A1(\SB2_0_26/i3[0] ), .A2(\SB2_0_26/i0[8] ), .A3(
        \SB2_0_26/i1_5 ), .ZN(\SB2_0_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2366 ( .A1(\SB1_0_31/i0_3 ), .A2(\SB1_0_31/i0[10] ), .A3(
        \SB1_0_31/i0_4 ), .ZN(\SB1_0_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2367 ( .A1(\SB1_3_15/i0[9] ), .A2(\SB1_3_15/i0_3 ), .A3(
        \SB1_3_15/i0[10] ), .ZN(\SB1_3_15/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2368 ( .A1(\SB2_0_9/i0[8] ), .A2(\SB2_0_9/i1_5 ), .A3(
        \SB2_0_9/i3[0] ), .ZN(\SB2_0_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2369 ( .A1(\SB2_3_16/i0[10] ), .A2(\SB2_3_16/i0_0 ), .A3(
        \SB2_3_16/i0[6] ), .ZN(\SB2_3_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2370 ( .A1(\SB2_0_18/i0_3 ), .A2(\SB2_0_18/i0[9] ), .A3(
        \SB2_0_18/i0[10] ), .ZN(\SB2_0_18/Component_Function_4/NAND4_in[2] )
         );
  XNOR2_X1 U2372 ( .A(n1086), .B(n1085), .ZN(\RI1[2][53] ) );
  XNOR2_X1 U2373 ( .A(\MC_ARK_ARC_1_1/temp2[53] ), .B(
        \MC_ARK_ARC_1_1/temp4[53] ), .ZN(n1085) );
  XNOR2_X1 U2374 ( .A(\MC_ARK_ARC_1_1/temp3[53] ), .B(
        \MC_ARK_ARC_1_1/temp1[53] ), .ZN(n1086) );
  NAND3_X1 U2375 ( .A1(\SB1_1_8/i1_7 ), .A2(\SB1_1_8/i0_4 ), .A3(
        \SB1_1_8/i0[8] ), .ZN(\SB1_1_8/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 U2376 ( .A1(\SB1_2_16/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_16/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_16/Component_Function_5/NAND4_in[0] ), .A4(n1087), .ZN(
        \RI3[2][95] ) );
  NAND3_X1 U2377 ( .A1(\SB1_3_18/i0_4 ), .A2(\SB1_3_18/i0[9] ), .A3(
        \SB1_3_18/i0[6] ), .ZN(\SB1_3_18/Component_Function_5/NAND4_in[3] ) );
  NAND4_X1 U2378 ( .A1(\SB4_25/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_25/Component_Function_4/NAND4_in[1] ), .A4(n1088), .ZN(n1449) );
  NAND3_X1 U2379 ( .A1(\SB4_25/i0_4 ), .A2(\SB4_25/i1[9] ), .A3(\SB4_25/i1_5 ), 
        .ZN(n1088) );
  NAND3_X1 U2381 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0[10] ), .A3(
        \SB2_2_28/i0[9] ), .ZN(n1089) );
  NAND4_X1 U2383 ( .A1(\SB2_0_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_6/Component_Function_4/NAND4_in[1] ), .A4(n1090), .ZN(
        \RI5[0][160] ) );
  NAND3_X1 U2384 ( .A1(\SB2_0_6/i0_4 ), .A2(\SB2_0_6/i1_5 ), .A3(
        \SB2_0_6/i1[9] ), .ZN(n1090) );
  NAND3_X1 U2385 ( .A1(\SB1_1_31/i0_3 ), .A2(\SB1_1_31/i0[10] ), .A3(
        \SB1_1_31/i0_4 ), .ZN(\SB1_1_31/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U2387 ( .A1(\SB2_1_29/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_29/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_29/Component_Function_2/NAND4_in[1] ), .A4(n1092), .ZN(
        \RI5[1][32] ) );
  NAND3_X1 U2388 ( .A1(\SB2_1_29/i0_4 ), .A2(\SB2_1_29/i1_5 ), .A3(
        \SB2_1_29/i0_0 ), .ZN(n1092) );
  NAND3_X1 U2389 ( .A1(\SB1_3_10/i0_0 ), .A2(\SB1_3_10/i1_5 ), .A3(
        \SB1_3_10/i0_4 ), .ZN(\SB1_3_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2390 ( .A1(\SB2_2_0/i0[10] ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0[6] ), .ZN(\SB2_2_0/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2391 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i0_0 ), .A3(
        \SB2_2_12/i0[6] ), .ZN(\SB2_2_12/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U2392 ( .A(\RI3[3][38] ), .ZN(\SB2_3_25/i1[9] ) );
  NAND3_X1 U2393 ( .A1(\SB2_2_2/i0_3 ), .A2(\RI3[2][174] ), .A3(
        \SB2_2_2/i0[8] ), .ZN(\SB2_2_2/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U2394 ( .A(\RI1[2][53] ), .ZN(\SB1_2_23/i0_3 ) );
  NAND3_X1 U2395 ( .A1(\SB2_0_25/i0[8] ), .A2(\SB2_0_25/i1_5 ), .A3(
        \SB2_0_25/i3[0] ), .ZN(\SB2_0_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2396 ( .A1(\SB1_0_27/i0[10] ), .A2(\SB1_0_27/i1_7 ), .A3(
        \SB1_0_27/i1[9] ), .ZN(\SB1_0_27/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U2400 ( .A1(\SB1_3_28/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_28/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_3_28/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_28/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[3][38] ) );
  NAND3_X1 U2401 ( .A1(\SB4_4/i0_3 ), .A2(\SB4_4/i1[9] ), .A3(\SB4_4/i0[6] ), 
        .ZN(\SB4_4/Component_Function_3/NAND4_in[0] ) );
  XNOR2_X1 U2402 ( .A(n1094), .B(n264), .ZN(Ciphertext[169]) );
  NAND3_X1 U2403 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i0_4 ), .A3(
        \SB1_2_3/i1[9] ), .ZN(n1453) );
  NAND4_X1 U2404 ( .A1(\SB4_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_11/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_11/Component_Function_0/NAND4_in[0] ), .A4(n1095), .ZN(n1154) );
  NAND3_X1 U2405 ( .A1(\SB4_11/i0[6] ), .A2(\SB4_11/i0[8] ), .A3(n551), .ZN(
        n1095) );
  NAND3_X1 U2406 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i0[10] ), .A3(
        \SB1_1_1/i0[9] ), .ZN(\SB1_1_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2407 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0[9] ), .A3(
        \SB2_0_4/i0[8] ), .ZN(\SB2_0_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2409 ( .A1(n1667), .A2(\SB4_4/i0_4 ), .A3(\SB4_4/i0_0 ), .ZN(
        \SB4_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2410 ( .A1(\SB1_2_20/i1[9] ), .A2(\SB1_2_20/i0[10] ), .A3(
        \SB1_2_20/i1_7 ), .ZN(\SB1_2_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2411 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[9] ), .A3(
        \SB2_0_5/i0[10] ), .ZN(\SB2_0_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2413 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[9] ), .A3(
        \SB1_3_23/i0[10] ), .ZN(n1096) );
  NAND4_X2 U2414 ( .A1(\SB1_3_29/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_29/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_29/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_28/i0_4 ) );
  XNOR2_X1 U2418 ( .A(n1100), .B(n1099), .ZN(\RI1[1][17] ) );
  XNOR2_X1 U2419 ( .A(\MC_ARK_ARC_1_0/temp2[17] ), .B(
        \MC_ARK_ARC_1_0/temp4[17] ), .ZN(n1099) );
  XNOR2_X1 U2420 ( .A(\MC_ARK_ARC_1_0/temp1[17] ), .B(
        \MC_ARK_ARC_1_0/temp3[17] ), .ZN(n1100) );
  NAND3_X1 U2423 ( .A1(\SB1_1_29/i0_3 ), .A2(\SB1_1_29/i0[9] ), .A3(
        \SB1_1_29/i0[10] ), .ZN(\SB1_1_29/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2424 ( .A1(\SB1_1_19/i1_7 ), .A2(\SB1_1_19/i0[10] ), .A3(
        \SB1_1_19/i1[9] ), .ZN(\SB1_1_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2425 ( .A1(\SB4_7/i0[6] ), .A2(\SB4_7/i1_5 ), .A3(\SB4_7/i0[9] ), 
        .ZN(n1101) );
  NAND4_X1 U2426 ( .A1(\SB1_3_23/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_23/Component_Function_5/NAND4_in[0] ), .A4(n1102), .ZN(
        \RI3[3][53] ) );
  NAND3_X1 U2427 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i1[9] ), .A3(
        \SB1_3_23/i0_4 ), .ZN(n1102) );
  NAND3_X1 U2430 ( .A1(\SB1_2_27/i0_3 ), .A2(\SB1_2_27/i0[9] ), .A3(
        \SB1_2_27/i0[8] ), .ZN(\SB1_2_27/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U2433 ( .A(\RI1[3][107] ), .ZN(\SB1_3_14/i0_3 ) );
  XNOR2_X1 U2434 ( .A(\MC_ARK_ARC_1_2/temp5[107] ), .B(
        \MC_ARK_ARC_1_2/temp6[107] ), .ZN(\RI1[3][107] ) );
  NAND4_X1 U2436 ( .A1(\SB1_2_25/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_25/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_25/Component_Function_4/NAND4_in[3] ), .A4(n1104), .ZN(
        \RI3[2][46] ) );
  NAND3_X1 U2437 ( .A1(\SB1_2_25/i0_3 ), .A2(\SB1_2_25/i0[9] ), .A3(
        \SB1_2_25/i0[10] ), .ZN(n1104) );
  NAND3_X1 U2438 ( .A1(\SB4_21/i0[6] ), .A2(\SB4_21/i0[8] ), .A3(
        \SB4_21/i0[7] ), .ZN(n1105) );
  NAND4_X1 U2441 ( .A1(\SB4_4/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_4/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_4/Component_Function_0/NAND4_in[0] ), .A4(n1107), .ZN(n1446) );
  NAND3_X1 U2442 ( .A1(\SB4_4/i0[6] ), .A2(\SB4_4/i0[8] ), .A3(\SB4_4/i0[7] ), 
        .ZN(n1107) );
  NAND3_X1 U2444 ( .A1(\SB4_31/i0[6] ), .A2(\SB4_31/i0[8] ), .A3(
        \SB4_31/i0[7] ), .ZN(n1108) );
  NAND3_X1 U2446 ( .A1(\SB2_2_29/i0[10] ), .A2(\SB2_2_29/i1_7 ), .A3(
        \SB2_2_29/i1[9] ), .ZN(n1109) );
  NAND3_X1 U2447 ( .A1(\SB2_3_16/i3[0] ), .A2(\SB2_3_16/i1_5 ), .A3(
        \SB2_3_16/i0[8] ), .ZN(\SB2_3_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2448 ( .A1(\SB2_3_4/i3[0] ), .A2(\SB2_3_4/i1_5 ), .A3(
        \SB2_3_4/i0[8] ), .ZN(\SB2_3_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2449 ( .A1(\SB1_3_6/i1_7 ), .A2(\SB1_3_6/i0[10] ), .A3(
        \SB1_3_6/i1[9] ), .ZN(\SB1_3_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2451 ( .A1(\SB2_3_31/i0[8] ), .A2(\SB2_3_31/i1_5 ), .A3(
        \SB2_3_31/i3[0] ), .ZN(\SB2_3_31/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U2452 ( .A1(\SB2_0_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_25/Component_Function_0/NAND4_in[0] ), .A4(n1110), .ZN(
        \RI5[0][66] ) );
  NAND3_X1 U2453 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0[7] ), .A3(
        \SB2_0_25/i0_0 ), .ZN(n1110) );
  NAND3_X1 U2456 ( .A1(\SB2_2_26/i0_4 ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i1[9] ), .ZN(\SB2_2_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2457 ( .A1(\SB2_1_13/i0_0 ), .A2(\SB2_1_13/i0[10] ), .A3(
        \SB2_1_13/i0[6] ), .ZN(\SB2_1_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2458 ( .A1(\SB1_2_20/i0_3 ), .A2(\SB1_2_20/i0_0 ), .A3(
        \SB1_2_20/i0_4 ), .ZN(\SB1_2_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2459 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0_0 ), .A3(
        \SB2_2_28/i0_4 ), .ZN(\SB2_2_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2460 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0_0 ), .A3(
        \SB2_1_5/i0_4 ), .ZN(\SB2_1_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2461 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0_0 ), .A3(
        \SB1_1_15/i0_4 ), .ZN(\SB1_1_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2462 ( .A1(\SB2_2_21/i0_4 ), .A2(\RI3[2][60] ), .A3(
        \SB2_2_21/i0[6] ), .ZN(\SB2_2_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2463 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i0[9] ), .A3(
        \SB1_2_31/i0[10] ), .ZN(\SB1_2_31/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2466 ( .A1(\SB2_2_0/i0[10] ), .A2(\SB2_2_0/i1_5 ), .A3(
        \SB2_2_0/i1[9] ), .ZN(\SB2_2_0/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U2467 ( .A1(\SB2_2_5/i0[6] ), .A2(n1113), .ZN(
        \SB2_2_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2470 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0[9] ), .A3(
        \SB1_1_13/i0[8] ), .ZN(\SB1_1_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2471 ( .A1(\SB1_2_30/i0_3 ), .A2(\SB1_2_30/i0[9] ), .A3(
        \SB1_2_30/i0[8] ), .ZN(\SB1_2_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2472 ( .A1(\SB2_2_8/i0_0 ), .A2(\SB2_2_8/i0[10] ), .A3(
        \SB2_2_8/i0[6] ), .ZN(\SB2_2_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2473 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB2_3_23/i0[10] ), .A3(
        \SB2_3_23/i0[6] ), .ZN(\SB2_3_23/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U2475 ( .A(n1117), .B(n1116), .ZN(\RI1[1][59] ) );
  XNOR2_X1 U2476 ( .A(\MC_ARK_ARC_1_0/temp1[59] ), .B(
        \MC_ARK_ARC_1_0/temp4[59] ), .ZN(n1116) );
  XNOR2_X1 U2477 ( .A(\MC_ARK_ARC_1_0/temp3[59] ), .B(
        \MC_ARK_ARC_1_0/temp2[59] ), .ZN(n1117) );
  NAND3_X1 U2478 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0[10] ), .A3(
        \SB1_0_5/i0_4 ), .ZN(\SB1_0_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2479 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0_4 ), .A3(
        \SB1_0_0/i1[9] ), .ZN(\SB1_0_0/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U2481 ( .A1(\SB1_2_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_5/NAND4_in[0] ), .A4(n1118), .ZN(
        \RI3[2][155] ) );
  NAND4_X1 U2483 ( .A1(\SB1_2_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_24/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_24/Component_Function_5/NAND4_in[0] ), .A4(n1119), .ZN(
        \RI3[2][47] ) );
  NAND3_X1 U2484 ( .A1(\SB1_2_24/i0_3 ), .A2(\SB1_2_24/i1[9] ), .A3(
        \SB1_2_24/i0_4 ), .ZN(n1119) );
  NAND3_X1 U2485 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i0[9] ), .A3(
        \SB1_2_31/i0[8] ), .ZN(n1247) );
  NAND3_X1 U2486 ( .A1(n2136), .A2(\SB1_0_6/i0[10] ), .A3(\SB1_0_6/i0_4 ), 
        .ZN(\SB1_0_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2487 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i1[9] ), .A3(
        \SB1_2_31/i0[6] ), .ZN(\SB1_2_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2488 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0[9] ), .A3(
        \SB1_2_13/i0[10] ), .ZN(\SB1_2_13/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2489 ( .A1(\SB2_0_6/i1_5 ), .A2(\SB2_0_6/i3[0] ), .A3(
        \SB2_0_6/i0[8] ), .ZN(\SB2_0_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2490 ( .A1(\SB2_3_9/i0[10] ), .A2(\SB2_3_9/i0_0 ), .A3(
        \SB2_3_9/i0[6] ), .ZN(\SB2_3_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2493 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0_0 ), .A3(
        \SB1_1_14/i0_4 ), .ZN(\SB1_1_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2496 ( .A1(\SB2_3_1/i0_4 ), .A2(\SB2_3_1/i0[9] ), .A3(
        \RI3[3][181] ), .ZN(\SB2_3_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2498 ( .A1(\SB2_0_8/i1_5 ), .A2(\SB2_0_8/i3[0] ), .A3(
        \SB2_0_8/i0[8] ), .ZN(n1121) );
  NAND4_X2 U2501 ( .A1(\SB1_3_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_4/NAND4_in[1] ), .A3(n1250), .A4(
        \SB1_3_14/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_13/i0_4 ) );
  NAND3_X1 U2502 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0_0 ), .A3(
        \SB1_0_10/i0_4 ), .ZN(\SB1_0_10/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U2503 ( .A1(\SB1_3_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_4/NAND4_in[3] ), .A4(n1123), .ZN(
        \RI3[3][184] ) );
  NAND4_X1 U2505 ( .A1(\SB1_1_12/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_12/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_12/Component_Function_4/NAND4_in[3] ), .A4(n1124), .ZN(
        \RI3[1][124] ) );
  NAND3_X1 U2506 ( .A1(\SB1_1_12/i0_3 ), .A2(\SB1_1_12/i0[10] ), .A3(
        \SB1_1_12/i0[9] ), .ZN(n1124) );
  NAND3_X1 U2508 ( .A1(\SB1_2_27/i0_3 ), .A2(\SB1_2_27/i0_0 ), .A3(
        \SB1_2_27/i0_4 ), .ZN(\SB1_2_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2509 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i0_0 ), .A3(
        \SB2_2_1/i0[6] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U2510 ( .A1(\SB2_1_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_26/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_26/Component_Function_3/NAND4_in[2] ), .A4(n1125), .ZN(
        \RI5[1][45] ) );
  NAND3_X1 U2511 ( .A1(\SB2_1_26/i3[0] ), .A2(\SB2_1_26/i1_5 ), .A3(
        \SB2_1_26/i0[8] ), .ZN(n1125) );
  NAND3_X1 U2512 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i0[9] ), .A3(
        \SB1_2_2/i0[10] ), .ZN(\SB1_2_2/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U2513 ( .A(n1127), .B(n1126), .ZN(\RI1[3][123] ) );
  XNOR2_X1 U2514 ( .A(\MC_ARK_ARC_1_2/temp1[123] ), .B(
        \MC_ARK_ARC_1_2/temp4[123] ), .ZN(n1126) );
  XNOR2_X1 U2515 ( .A(\MC_ARK_ARC_1_2/temp3[123] ), .B(
        \MC_ARK_ARC_1_2/temp2[123] ), .ZN(n1127) );
  NAND3_X1 U2516 ( .A1(\SB2_2_18/i3[0] ), .A2(\SB2_2_18/i1_5 ), .A3(
        \SB2_2_18/i0[8] ), .ZN(n1128) );
  NAND4_X1 U2517 ( .A1(\SB2_1_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_14/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_14/Component_Function_2/NAND4_in[1] ), .A4(n1129), .ZN(
        \RI5[1][122] ) );
  NAND3_X1 U2518 ( .A1(\SB2_1_14/i0_4 ), .A2(\SB2_1_14/i1_5 ), .A3(
        \SB2_1_14/i0_0 ), .ZN(n1129) );
  NAND4_X1 U2519 ( .A1(\SB1_3_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_30/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_30/Component_Function_2/NAND4_in[2] ), .A4(n1130), .ZN(
        \RI3[3][26] ) );
  NAND3_X1 U2520 ( .A1(\SB1_3_30/i0_0 ), .A2(\SB1_3_30/i0_4 ), .A3(
        \SB1_3_30/i1_5 ), .ZN(n1130) );
  XNOR2_X1 U2521 ( .A(n1131), .B(n1132), .ZN(\RI1[1][113] ) );
  XNOR2_X1 U2522 ( .A(\MC_ARK_ARC_1_0/temp1[113] ), .B(
        \MC_ARK_ARC_1_0/temp4[113] ), .ZN(n1131) );
  XNOR2_X1 U2523 ( .A(\MC_ARK_ARC_1_0/temp3[113] ), .B(
        \MC_ARK_ARC_1_0/temp2[113] ), .ZN(n1132) );
  NAND3_X1 U2524 ( .A1(\SB2_1_30/i3[0] ), .A2(\SB2_1_30/i1_5 ), .A3(
        \SB2_1_30/i0[8] ), .ZN(\SB2_1_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2526 ( .A1(\SB2_1_19/i0_4 ), .A2(\SB2_1_19/i1_5 ), .A3(
        \SB2_1_19/i0_0 ), .ZN(n1134) );
  NAND3_X1 U2527 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0_0 ), .A3(
        \SB1_0_20/i0_4 ), .ZN(\SB1_0_20/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U2528 ( .A1(\SB1_2_14/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_14/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_14/Component_Function_4/NAND4_in[3] ), .A4(n1135), .ZN(
        \RI3[2][112] ) );
  NAND3_X1 U2529 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i0[9] ), .A3(
        \SB1_2_14/i0[10] ), .ZN(n1135) );
  NAND4_X1 U2530 ( .A1(\SB1_0_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_4/NAND4_in[2] ), .A4(n1136), .ZN(
        \RI3[0][58] ) );
  NAND3_X1 U2531 ( .A1(\SB1_0_23/i1_5 ), .A2(\SB1_0_23/i1[9] ), .A3(
        \SB1_0_23/i0_4 ), .ZN(n1136) );
  NAND3_X1 U2532 ( .A1(\SB2_2_6/i0_4 ), .A2(\SB2_2_6/i0_3 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2533 ( .A1(\SB2_1_19/i0_4 ), .A2(\SB2_1_19/i0[9] ), .A3(
        \SB2_1_19/i0[6] ), .ZN(\SB2_1_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2534 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i0_4 ), .A3(
        \SB2_0_27/i0_0 ), .ZN(\SB2_0_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2535 ( .A1(\SB1_0_27/i0_3 ), .A2(\SB1_0_27/i1[9] ), .A3(
        \SB1_0_27/i0_4 ), .ZN(\SB1_0_27/Component_Function_5/NAND4_in[2] ) );
  NAND4_X4 U2536 ( .A1(\SB2_0_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_24/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_24/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_24/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[47] ) );
  NAND3_X1 U2537 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i0[9] ), .A3(
        \SB1_1_26/i0[8] ), .ZN(\SB1_1_26/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2538 ( .A(n1138), .B(n1137), .ZN(\RI1[3][41] ) );
  XNOR2_X1 U2539 ( .A(\MC_ARK_ARC_1_2/temp4[41] ), .B(
        \MC_ARK_ARC_1_2/temp1[41] ), .ZN(n1137) );
  XNOR2_X1 U2540 ( .A(\MC_ARK_ARC_1_2/temp3[41] ), .B(
        \MC_ARK_ARC_1_2/temp2[41] ), .ZN(n1138) );
  INV_X2 U2542 ( .A(\RI1[2][89] ), .ZN(\SB1_2_17/i0_3 ) );
  NAND3_X1 U2546 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i0[9] ), .A3(
        \SB1_1_1/i0[8] ), .ZN(\SB1_1_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2547 ( .A1(\SB2_1_9/i0_4 ), .A2(\SB2_1_9/i0[9] ), .A3(
        \SB2_1_9/i0[6] ), .ZN(\SB2_1_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2550 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0[9] ), .A3(
        \SB2_1_18/i0[8] ), .ZN(\SB2_1_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2551 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[9] ), .A3(
        \SB2_2_23/i0[8] ), .ZN(\SB2_2_23/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U2552 ( .A(\RI1[2][23] ), .ZN(\SB1_2_28/i0_3 ) );
  XNOR2_X1 U2553 ( .A(\MC_ARK_ARC_1_1/temp5[23] ), .B(
        \MC_ARK_ARC_1_1/temp6[23] ), .ZN(\RI1[2][23] ) );
  NAND3_X1 U2554 ( .A1(\SB1_2_25/i0_3 ), .A2(\SB1_2_25/i0_0 ), .A3(
        \SB1_2_25/i0_4 ), .ZN(\SB1_2_25/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2555 ( .A(n1140), .B(n254), .ZN(Ciphertext[143]) );
  NAND4_X1 U2556 ( .A1(\SB4_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_8/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_8/Component_Function_5/NAND4_in[0] ), .ZN(n1140) );
  NAND3_X1 U2557 ( .A1(\SB2_0_26/i0_0 ), .A2(\SB2_0_26/i0[6] ), .A3(
        \SB2_0_26/i0[10] ), .ZN(n1141) );
  NAND3_X1 U2558 ( .A1(\SB2_2_22/i0_4 ), .A2(\SB2_2_22/i1_7 ), .A3(
        \SB2_2_22/i0[8] ), .ZN(\SB2_2_22/Component_Function_1/NAND4_in[3] ) );
  XNOR2_X1 U2562 ( .A(n1145), .B(n1144), .ZN(\RI1[1][189] ) );
  XNOR2_X1 U2563 ( .A(\MC_ARK_ARC_1_0/temp2[189] ), .B(
        \MC_ARK_ARC_1_0/temp4[189] ), .ZN(n1144) );
  XNOR2_X1 U2564 ( .A(\MC_ARK_ARC_1_0/temp1[189] ), .B(
        \MC_ARK_ARC_1_0/temp3[189] ), .ZN(n1145) );
  NAND3_X1 U2565 ( .A1(n834), .A2(\SB4_5/i1[9] ), .A3(\SB4_5/i1_5 ), .ZN(n1146) );
  NAND3_X1 U2566 ( .A1(\SB2_3_9/i3[0] ), .A2(\SB2_3_9/i0[8] ), .A3(
        \SB2_3_9/i1_5 ), .ZN(\SB2_3_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2569 ( .A1(\SB2_0_22/i1_5 ), .A2(\SB2_0_22/i3[0] ), .A3(
        \SB2_0_22/i0[8] ), .ZN(\SB2_0_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2570 ( .A1(\SB1_1_31/i1[9] ), .A2(\SB1_1_31/i0[10] ), .A3(
        \SB1_1_31/i1_7 ), .ZN(\SB1_1_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2571 ( .A1(\SB1_1_0/i3[0] ), .A2(\SB1_1_0/i1_5 ), .A3(
        \SB1_1_0/i0[8] ), .ZN(\SB1_1_0/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U2572 ( .A1(\SB2_0_28/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_28/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_28/Component_Function_3/NAND4_in[0] ), .A4(n1148), .ZN(
        \RI5[0][33] ) );
  NAND3_X1 U2573 ( .A1(\SB2_0_28/i3[0] ), .A2(\SB2_0_28/i1_5 ), .A3(
        \SB2_0_28/i0[8] ), .ZN(n1148) );
  NAND3_X1 U2574 ( .A1(\SB2_2_22/i3[0] ), .A2(\SB2_2_22/i1_5 ), .A3(
        \SB2_2_22/i0[8] ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2577 ( .A1(\SB1_0_30/i0_3 ), .A2(\SB1_0_30/i0_0 ), .A3(
        \SB1_0_30/i0_4 ), .ZN(\SB1_0_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2578 ( .A1(\SB4_18/i0_4 ), .A2(\SB4_18/i0[8] ), .A3(\SB4_18/i1_7 ), 
        .ZN(\SB4_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2581 ( .A1(n871), .A2(\SB4_15/i1[9] ), .A3(\SB4_15/i0[6] ), .ZN(
        \SB4_15/Component_Function_3/NAND4_in[0] ) );
  XNOR2_X1 U2582 ( .A(n1151), .B(n204), .ZN(Ciphertext[82]) );
  NAND4_X1 U2583 ( .A1(\SB4_18/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_18/Component_Function_4/NAND4_in[0] ), .A3(n1285), .A4(
        \SB4_18/Component_Function_4/NAND4_in[1] ), .ZN(n1151) );
  NAND4_X1 U2584 ( .A1(\SB1_0_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_24/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_24/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][47] ) );
  XNOR2_X1 U2587 ( .A(n1153), .B(n253), .ZN(Ciphertext[102]) );
  NAND4_X1 U2588 ( .A1(\SB4_14/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_14/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_14/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_14/Component_Function_0/NAND4_in[1] ), .ZN(n1153) );
  XNOR2_X1 U2589 ( .A(n1154), .B(n317), .ZN(Ciphertext[120]) );
  NAND3_X1 U2591 ( .A1(\SB2_3_8/i0_4 ), .A2(\SB2_3_8/i0_3 ), .A3(
        \SB2_3_8/i1[9] ), .ZN(\SB2_3_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2592 ( .A1(\SB1_3_4/i0_0 ), .A2(\SB1_3_4/i0_4 ), .A3(
        \SB1_3_4/i1_5 ), .ZN(\SB1_3_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2593 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i0_0 ), .A3(
        \SB1_1_24/i0_4 ), .ZN(\SB1_1_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2594 ( .A1(\RI3[0][190] ), .A2(\RI3[0][186] ), .A3(\RI3[0][187] ), 
        .ZN(n1155) );
  NAND4_X1 U2596 ( .A1(\SB1_0_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_26/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_0_26/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[0][50] ) );
  NAND3_X1 U2598 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0_4 ), .A3(
        \SB1_0_18/i1[9] ), .ZN(n1156) );
  NAND3_X1 U2599 ( .A1(\SB1_2_9/i1[9] ), .A2(\SB1_2_9/i0[10] ), .A3(
        \SB1_2_9/i1_7 ), .ZN(\SB1_2_9/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U2600 ( .A1(\SB1_2_27/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_27/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_27/Component_Function_2/NAND4_in[2] ), .A4(n1157), .ZN(
        \RI3[2][44] ) );
  NAND4_X1 U2602 ( .A1(\SB2_0_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_1/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_1/Component_Function_3/NAND4_in[2] ), .A4(n1158), .ZN(
        \RI5[0][3] ) );
  NAND4_X1 U2604 ( .A1(\SB1_1_26/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_1_26/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_26/Component_Function_5/NAND4_in[0] ), .A4(n1159), .ZN(
        \RI3[1][35] ) );
  NAND3_X1 U2605 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i1[9] ), .A3(
        \SB1_1_26/i0_4 ), .ZN(n1159) );
  XNOR2_X1 U2606 ( .A(n1160), .B(n411), .ZN(Ciphertext[34]) );
  NAND3_X1 U2607 ( .A1(\SB2_2_6/i0[9] ), .A2(\SB2_2_6/i0_3 ), .A3(
        \SB2_2_6/i0[8] ), .ZN(n1161) );
  NAND2_X1 U2608 ( .A1(\SB2_0_24/i0[6] ), .A2(n1162), .ZN(
        \SB2_0_24/Component_Function_5/NAND4_in[3] ) );
  AND2_X1 U2609 ( .A1(\RI3[0][42] ), .A2(\RI3[0][46] ), .ZN(n1162) );
  NAND4_X1 U2612 ( .A1(\SB1_1_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_24/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_1_24/Component_Function_5/NAND4_in[3] ), .A4(n1164), .ZN(
        \RI3[1][47] ) );
  NAND3_X1 U2613 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i1[9] ), .A3(
        \SB1_1_24/i0_4 ), .ZN(n1164) );
  NAND3_X1 U2614 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i0[9] ), .A3(
        \SB1_1_3/i0[8] ), .ZN(\SB1_1_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2615 ( .A1(\SB1_1_2/i0_3 ), .A2(\SB1_1_2/i0[9] ), .A3(
        \SB1_1_2/i0[8] ), .ZN(\SB1_1_2/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2616 ( .A(\MC_ARK_ARC_1_2/temp5[56] ), .B(n1165), .ZN(\RI1[3][56] ) );
  XNOR2_X1 U2617 ( .A(\MC_ARK_ARC_1_2/temp3[56] ), .B(
        \MC_ARK_ARC_1_2/temp4[56] ), .ZN(n1165) );
  NAND3_X1 U2618 ( .A1(\SB2_3_0/i0_4 ), .A2(\SB2_3_0/i0_3 ), .A3(
        \SB2_3_0/i1[9] ), .ZN(n1166) );
  NAND3_X1 U2620 ( .A1(\SB1_1_18/i0_3 ), .A2(\SB1_1_18/i0_0 ), .A3(
        \SB1_1_18/i0_4 ), .ZN(\SB1_1_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2621 ( .A1(\SB1_1_29/i0_3 ), .A2(\SB1_1_29/i0[9] ), .A3(
        \SB1_1_29/i0[8] ), .ZN(\SB1_1_29/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U2622 ( .A1(\SB2_3_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_31/Component_Function_5/NAND4_in[0] ), .A4(n1167), .ZN(
        \RI5[3][5] ) );
  NAND3_X1 U2623 ( .A1(n1652), .A2(\RI3[3][0] ), .A3(\RI3[3][1] ), .ZN(n1167)
         );
  NAND3_X1 U2624 ( .A1(n1671), .A2(\SB4_26/i1[9] ), .A3(\SB4_26/i0[6] ), .ZN(
        \SB4_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2625 ( .A1(\SB1_3_20/i0_3 ), .A2(\SB1_3_20/i0_0 ), .A3(
        \SB1_3_20/i0_4 ), .ZN(\SB1_3_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2626 ( .A1(\SB2_2_17/i0_4 ), .A2(\SB2_2_17/i0_3 ), .A3(
        \SB2_2_17/i1[9] ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2627 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0[7] ), .A3(\SB4_2/i0_0 ), 
        .ZN(\SB4_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2628 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i0_4 ), 
        .ZN(\SB4_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2629 ( .A1(\SB1_2_11/i0_3 ), .A2(\SB1_2_11/i0_0 ), .A3(
        \SB1_2_11/i0_4 ), .ZN(\SB1_2_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2630 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i0_0 ), .A3(
        \SB1_1_26/i0_4 ), .ZN(\SB1_1_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2636 ( .A1(\SB2_3_27/i3[0] ), .A2(n1630), .A3(\SB2_3_27/i0[8] ), 
        .ZN(\SB2_3_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2637 ( .A1(\SB2_2_8/i3[0] ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i0[8] ), .ZN(n1169) );
  NAND3_X1 U2638 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i0_4 ), .A3(
        \SB1_1_19/i1_5 ), .ZN(\SB1_1_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2639 ( .A1(n848), .A2(\SB4_23/i0[8] ), .A3(\SB4_23/i1_7 ), .ZN(
        \SB4_23/Component_Function_1/NAND4_in[1] ) );
  XNOR2_X1 U2640 ( .A(n1170), .B(n1171), .ZN(\RI1[3][191] ) );
  XNOR2_X1 U2641 ( .A(\MC_ARK_ARC_1_2/temp4[191] ), .B(
        \MC_ARK_ARC_1_2/temp1[191] ), .ZN(n1170) );
  XNOR2_X1 U2642 ( .A(\MC_ARK_ARC_1_2/temp2[191] ), .B(
        \MC_ARK_ARC_1_2/temp3[191] ), .ZN(n1171) );
  NAND3_X1 U2643 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0_4 ), .A3(
        \SB2_1_22/i1[9] ), .ZN(n1172) );
  NAND3_X1 U2644 ( .A1(\SB2_2_8/i0[10] ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i1[9] ), .ZN(\SB2_2_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2648 ( .A1(\SB2_0_7/i3[0] ), .A2(\SB2_0_7/i1_5 ), .A3(
        \SB2_0_7/i0[8] ), .ZN(n1174) );
  NAND3_X1 U2650 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i0_0 ), .A3(
        \SB1_2_3/i0_4 ), .ZN(\SB1_2_3/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U2651 ( .A1(\SB2_2_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_20/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_20/Component_Function_2/NAND4_in[1] ), .A4(n1175), .ZN(
        \RI5[2][86] ) );
  NAND3_X1 U2652 ( .A1(\SB2_2_20/i0_4 ), .A2(\SB2_2_20/i0_0 ), .A3(
        \SB2_2_20/i1_5 ), .ZN(n1175) );
  NAND4_X1 U2657 ( .A1(\SB3_6/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_6/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_6/Component_Function_0/NAND4_in[1] ), .A4(n1178), .ZN(
        \RI3[4][180] ) );
  NAND3_X1 U2658 ( .A1(\SB3_6/i0[7] ), .A2(\SB3_6/i0_0 ), .A3(n833), .ZN(n1178) );
  AND2_X1 U2659 ( .A1(\RI3[2][142] ), .A2(\RI3[2][138] ), .ZN(n1205) );
  NAND4_X2 U2660 ( .A1(\SB2_3_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_20/Component_Function_1/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[91] ) );
  NAND3_X1 U2661 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0_0 ), .A3(
        \SB1_0_28/i0_4 ), .ZN(\SB1_0_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2662 ( .A1(\SB1_2_22/i0_3 ), .A2(\SB1_2_22/i0[9] ), .A3(
        \SB1_2_22/i0[8] ), .ZN(\SB1_2_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2665 ( .A1(\SB2_2_1/i0_4 ), .A2(\RI3[2][180] ), .A3(
        \SB2_2_1/i0[6] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[3] ) );
  NAND4_X4 U2666 ( .A1(\SB2_0_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_12/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[119] ) );
  NAND3_X1 U2667 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0[10] ), .A3(
        \SB1_0_5/i0[9] ), .ZN(\SB1_0_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2668 ( .A1(\SB2_1_11/i0[9] ), .A2(\SB2_1_11/i0_3 ), .A3(
        \SB2_1_11/i0[8] ), .ZN(\SB2_1_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2669 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i0_4 ), .A3(
        \SB1_1_23/i1_5 ), .ZN(\SB1_1_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2670 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0_0 ), .A3(
        \SB1_1_13/i0_4 ), .ZN(\SB1_1_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2671 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i0_0 ), .A3(
        \SB1_1_3/i0_4 ), .ZN(\SB1_1_3/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U2672 ( .A1(\SB2_1_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_2/Component_Function_5/NAND4_in[0] ), .A4(n1180), .ZN(
        \RI5[1][179] ) );
  NAND3_X1 U2673 ( .A1(\SB2_1_2/i0_4 ), .A2(\RI3[1][174] ), .A3(
        \SB2_1_2/i0[6] ), .ZN(n1180) );
  NAND4_X1 U2674 ( .A1(\SB1_1_20/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_1_20/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[1][86] ) );
  NAND3_X1 U2675 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0_0 ), .A3(
        \SB1_1_30/i0_4 ), .ZN(\SB1_1_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2678 ( .A1(\SB1_1_21/i1[9] ), .A2(\SB1_1_21/i0[10] ), .A3(
        \SB1_1_21/i1_7 ), .ZN(\SB1_1_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2681 ( .A1(\SB4_7/i0[6] ), .A2(\SB4_7/i0_0 ), .A3(\SB4_7/i0[10] ), 
        .ZN(n1182) );
  NAND3_X1 U2682 ( .A1(\SB2_2_14/i0[8] ), .A2(\SB2_2_14/i1_5 ), .A3(
        \SB2_2_14/i3[0] ), .ZN(\SB2_2_14/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U2684 ( .A1(\SB2_2_30/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_30/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_2_30/Component_Function_1/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[31] ) );
  NAND3_X1 U2685 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i0_0 ), .A3(\SB4_3/i0[7] ), 
        .ZN(\SB4_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2686 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0[9] ), .A3(
        \SB1_0_22/i0[8] ), .ZN(\SB1_0_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2687 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i0_0 ), .A3(
        \SB2_0_4/i0[6] ), .ZN(\SB2_0_4/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U2690 ( .A(n1184), .B(n366), .ZN(Ciphertext[140]) );
  NAND3_X1 U2691 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i0[9] ), .ZN(\SB1_2_12/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U2693 ( .A1(\SB4_27/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_27/Component_Function_1/NAND4_in[0] ), .A4(n1185), .ZN(n1339) );
  NAND3_X1 U2694 ( .A1(n780), .A2(\SB4_27/i1_7 ), .A3(\SB4_27/i0[8] ), .ZN(
        n1185) );
  NAND3_X1 U2695 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i0[10] ), .A3(
        \SB1_1_26/i0_4 ), .ZN(\SB1_1_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2696 ( .A1(\SB1_2_7/i0_3 ), .A2(\SB1_2_7/i0_0 ), .A3(
        \SB1_2_7/i0_4 ), .ZN(\SB1_2_7/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U2700 ( .A1(\SB4_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_3/Component_Function_0/NAND4_in[0] ), .A4(n1187), .ZN(n1338) );
  NAND3_X1 U2701 ( .A1(\SB4_3/i0[6] ), .A2(\SB4_3/i0[8] ), .A3(\SB4_3/i0[7] ), 
        .ZN(n1187) );
  NAND3_X1 U2702 ( .A1(\SB2_3_27/i0[9] ), .A2(\SB2_3_27/i0_3 ), .A3(
        \SB2_3_27/i0[8] ), .ZN(\SB2_3_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2703 ( .A1(\SB2_3_6/i0[9] ), .A2(\SB2_3_6/i0_3 ), .A3(
        \SB2_3_6/i0[8] ), .ZN(\SB2_3_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2704 ( .A1(\SB1_3_28/i0_0 ), .A2(\SB1_3_28/i0_4 ), .A3(
        \SB1_3_28/i1_5 ), .ZN(\SB1_3_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2705 ( .A1(\SB2_1_19/i0_4 ), .A2(\SB2_1_19/i0_3 ), .A3(
        \SB2_1_19/i1[9] ), .ZN(\SB2_1_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2706 ( .A1(\SB2_2_25/i3[0] ), .A2(\SB2_2_25/i1_5 ), .A3(
        \SB2_2_25/i0[8] ), .ZN(\SB2_2_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2707 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i0_0 ), .A3(\SB4_0/i0[7] ), 
        .ZN(\SB4_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2708 ( .A1(\SB4_8/i0_3 ), .A2(\SB4_8/i0_0 ), .A3(n1512), .ZN(
        \SB4_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2709 ( .A1(\SB4_22/i0_0 ), .A2(n779), .A3(\SB4_22/i0[8] ), .ZN(
        \SB4_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2710 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i0_0 ), .A3(
        \SB1_1_7/i0_4 ), .ZN(\SB1_1_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2711 ( .A1(\SB3_11/i1[9] ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i0_3 ), 
        .ZN(\SB3_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2713 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i1[9] ), .A3(\SB4_3/i0[6] ), 
        .ZN(\SB4_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2714 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0[9] ), .A3(
        \SB2_2_4/i0[8] ), .ZN(\SB2_2_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2715 ( .A1(\SB1_3_9/i0_0 ), .A2(\SB1_3_9/i1_5 ), .A3(
        \SB1_3_9/i0_4 ), .ZN(\SB1_3_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2716 ( .A1(\SB2_2_1/i0[9] ), .A2(\SB2_2_1/i0_3 ), .A3(
        \SB2_2_1/i0[8] ), .ZN(\SB2_2_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2717 ( .A1(\SB2_2_25/i1[9] ), .A2(\SB2_2_25/i0_3 ), .A3(
        \SB2_2_25/i0_4 ), .ZN(\SB2_2_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2718 ( .A1(\SB1_2_15/i0_3 ), .A2(\SB1_2_15/i0[10] ), .A3(
        \SB1_2_15/i0[9] ), .ZN(\SB1_2_15/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U2720 ( .A1(\SB4_11/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_11/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_11/Component_Function_1/NAND4_in[0] ), .A4(n1188), .ZN(n1190) );
  NAND3_X1 U2721 ( .A1(n805), .A2(\SB4_11/i1_7 ), .A3(\SB4_11/i0[8] ), .ZN(
        n1188) );
  NAND2_X1 U2722 ( .A1(\SB2_2_26/i0_0 ), .A2(\SB2_2_26/i3[0] ), .ZN(n1189) );
  NAND3_X1 U2723 ( .A1(n851), .A2(\SB4_22/i0[8] ), .A3(\SB4_22/i1_7 ), .ZN(
        \SB4_22/Component_Function_1/NAND4_in[1] ) );
  XNOR2_X1 U2724 ( .A(n1190), .B(n219), .ZN(Ciphertext[121]) );
  NAND3_X1 U2725 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0[7] ), .A3(
        \SB1_0_12/i0_0 ), .ZN(\SB1_0_12/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U2726 ( .A1(\SB1_3_25/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_25/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_25/Component_Function_2/NAND4_in[2] ), .A4(n1191), .ZN(
        \RI3[3][56] ) );
  NAND3_X1 U2730 ( .A1(\SB1_1_14/i3[0] ), .A2(\SB1_1_14/i1_5 ), .A3(
        \SB1_1_14/i0[8] ), .ZN(\SB1_1_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2731 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i0[9] ), .A3(
        \SB4_14/i0[10] ), .ZN(\SB4_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2732 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0_0 ), .A3(
        \SB1_0_12/i0_4 ), .ZN(\SB1_0_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2733 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0_0 ), .A3(
        \SB1_0_15/i0_4 ), .ZN(\SB1_0_15/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2736 ( .A(n1197), .B(n1196), .ZN(\RI1[1][74] ) );
  XNOR2_X1 U2737 ( .A(\MC_ARK_ARC_1_0/temp1[74] ), .B(
        \MC_ARK_ARC_1_0/temp2[74] ), .ZN(n1196) );
  XNOR2_X1 U2738 ( .A(\MC_ARK_ARC_1_0/temp3[74] ), .B(
        \MC_ARK_ARC_1_0/temp4[74] ), .ZN(n1197) );
  NAND3_X1 U2739 ( .A1(\SB1_2_15/i0_3 ), .A2(\SB1_2_15/i0_0 ), .A3(
        \SB1_2_15/i0_4 ), .ZN(\SB1_2_15/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U2740 ( .A1(\SB2_0_11/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_0_11/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_11/Component_Function_4/NAND4_in[1] ), .A4(n1198), .ZN(
        \RI5[0][130] ) );
  NAND3_X1 U2741 ( .A1(\SB2_0_11/i0_4 ), .A2(\SB2_0_11/i1[9] ), .A3(
        \SB2_0_11/i1_5 ), .ZN(n1198) );
  NAND4_X1 U2742 ( .A1(\SB2_2_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_14/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_14/Component_Function_4/NAND4_in[1] ), .A4(n1199), .ZN(
        \RI5[2][112] ) );
  NAND3_X1 U2745 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0[9] ), .A3(
        \SB1_1_16/i0[10] ), .ZN(\SB1_1_16/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2746 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i0[8] ), .A3(\SB4_6/i1_7 ), 
        .ZN(\SB4_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2747 ( .A1(\SB1_2_6/i0_3 ), .A2(\SB1_2_6/i0[9] ), .A3(
        \SB1_2_6/i0[8] ), .ZN(\SB1_2_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2748 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0_4 ), .A3(
        \SB1_0_6/i1[9] ), .ZN(n1318) );
  NAND4_X1 U2749 ( .A1(\SB3_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_23/Component_Function_4/NAND4_in[3] ), .A3(
        \SB3_23/Component_Function_4/NAND4_in[1] ), .A4(n1200), .ZN(
        \RI3[4][58] ) );
  NAND3_X1 U2753 ( .A1(n834), .A2(\SB4_5/i1_7 ), .A3(\SB4_5/i0[8] ), .ZN(n1202) );
  NAND3_X1 U2754 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i1[9] ), .A3(
        \SB1_1_9/i1_7 ), .ZN(\SB1_1_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2755 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0_0 ), .A3(
        \SB1_0_2/i0_4 ), .ZN(\SB1_0_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2756 ( .A1(\SB1_2_6/i0_3 ), .A2(\SB1_2_6/i0_0 ), .A3(
        \SB1_2_6/i0_4 ), .ZN(\SB1_2_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2758 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0[10] ), .A3(
        \SB2_0_21/i0[9] ), .ZN(n1203) );
  NAND4_X1 U2759 ( .A1(\SB1_0_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_29/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][17] ) );
  NAND3_X1 U2760 ( .A1(\SB1_2_24/i0_3 ), .A2(\SB1_2_24/i0[9] ), .A3(
        \SB1_2_24/i0[8] ), .ZN(\SB1_2_24/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2764 ( .A(\MC_ARK_ARC_1_3/temp5[179] ), .B(n1204), .ZN(
        \RI1[4][179] ) );
  XNOR2_X1 U2765 ( .A(\MC_ARK_ARC_1_3/temp3[179] ), .B(
        \MC_ARK_ARC_1_3/temp4[179] ), .ZN(n1204) );
  NAND2_X1 U2766 ( .A1(\SB2_2_8/i0[6] ), .A2(n1205), .ZN(
        \SB2_2_8/Component_Function_5/NAND4_in[3] ) );
  NAND4_X1 U2767 ( .A1(\SB2_2_10/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_10/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_10/Component_Function_2/NAND4_in[1] ), .A4(n1206), .ZN(
        \RI5[2][146] ) );
  NAND3_X1 U2768 ( .A1(\SB2_2_10/i0_4 ), .A2(\SB2_2_10/i1_5 ), .A3(
        \SB2_2_10/i0_0 ), .ZN(n1206) );
  XNOR2_X1 U2769 ( .A(n1208), .B(n1207), .ZN(\RI1[1][83] ) );
  XNOR2_X1 U2770 ( .A(\MC_ARK_ARC_1_0/temp1[83] ), .B(
        \MC_ARK_ARC_1_0/temp4[83] ), .ZN(n1207) );
  XNOR2_X1 U2771 ( .A(\MC_ARK_ARC_1_0/temp2[83] ), .B(
        \MC_ARK_ARC_1_0/temp3[83] ), .ZN(n1208) );
  NAND3_X1 U2773 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i0_3 ), .A3(
        \SB2_1_1/i1[9] ), .ZN(n1209) );
  NAND3_X1 U2774 ( .A1(\SB3_11/i0[7] ), .A2(\SB3_11/i0_0 ), .A3(n840), .ZN(
        \SB3_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2775 ( .A1(\SB2_3_12/i0_3 ), .A2(\SB2_3_12/i0[9] ), .A3(
        \SB2_3_12/i0[8] ), .ZN(\SB2_3_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2777 ( .A1(\SB2_3_12/i0_4 ), .A2(\SB2_3_12/i0_3 ), .A3(
        \SB2_3_12/i1[9] ), .ZN(n1211) );
  NAND3_X1 U2778 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i1[9] ), .A3(\SB4_16/i0[6] ), .ZN(\SB4_16/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U2779 ( .A1(\SB1_3_15/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_15/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_15/Component_Function_2/NAND4_in[2] ), .A4(n1212), .ZN(
        \RI3[3][116] ) );
  NAND3_X1 U2780 ( .A1(\SB1_3_14/i0_3 ), .A2(\SB1_3_14/i0_0 ), .A3(
        \SB1_3_14/i0_4 ), .ZN(\SB1_3_14/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2782 ( .A(n1213), .B(n266), .ZN(Ciphertext[59]) );
  NAND4_X1 U2783 ( .A1(\SB4_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_22/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_22/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_22/Component_Function_5/NAND4_in[0] ), .ZN(n1213) );
  NAND3_X1 U2784 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i1[9] ), .A3(n806), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2785 ( .A1(\SB1_3_29/i0_3 ), .A2(\SB1_3_29/i0[10] ), .A3(
        \SB1_3_29/i0[9] ), .ZN(\SB1_3_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2787 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i1[9] ), .A3(\SB4_20/i0[6] ), .ZN(\SB4_20/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U2788 ( .A1(\SB2_2_0/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_0/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_0/Component_Function_2/NAND4_in[1] ), .A4(n1215), .ZN(
        \RI5[2][14] ) );
  NAND3_X1 U2789 ( .A1(\SB2_2_0/i0_4 ), .A2(\SB2_2_0/i1_5 ), .A3(
        \SB2_2_0/i0_0 ), .ZN(n1215) );
  XNOR2_X1 U2792 ( .A(n1217), .B(n247), .ZN(Ciphertext[7]) );
  NAND4_X1 U2793 ( .A1(\SB4_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_30/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_30/Component_Function_1/NAND4_in[2] ), .ZN(n1217) );
  NAND3_X1 U2796 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i0[9] ), .A3(\SB3_5/i0[10] ), 
        .ZN(\SB3_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2797 ( .A1(\SB4_10/i0_4 ), .A2(\SB4_10/i1[9] ), .A3(\SB4_10/i1_5 ), 
        .ZN(\SB4_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2798 ( .A1(\SB4_15/i0_4 ), .A2(\SB4_15/i1[9] ), .A3(\SB4_15/i1_5 ), 
        .ZN(\SB4_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2800 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i0[7] ), .A3(\SB3_5/i0_0 ), 
        .ZN(n1277) );
  NAND3_X1 U2802 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i0_0 ), .A3(
        \SB1_2_2/i0_4 ), .ZN(\SB1_2_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2803 ( .A1(\SB2_2_0/i0[8] ), .A2(\SB2_2_0/i1_5 ), .A3(
        \SB2_2_0/i3[0] ), .ZN(\SB2_2_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2804 ( .A1(\SB1_2_23/i0_3 ), .A2(\SB1_2_23/i0[9] ), .A3(
        \SB1_2_23/i0[10] ), .ZN(\SB1_2_23/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2805 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i1[9] ), .A3(
        \SB1_0_22/i0_4 ), .ZN(\SB1_0_22/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U2806 ( .A(n1219), .B(n305), .ZN(Ciphertext[12]) );
  NAND4_X1 U2807 ( .A1(\SB4_29/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_29/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_29/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_29/Component_Function_0/NAND4_in[1] ), .ZN(n1219) );
  NAND3_X1 U2808 ( .A1(\SB2_2_8/i0_4 ), .A2(\SB2_2_8/i1[9] ), .A3(
        \SB2_2_8/i0_3 ), .ZN(\SB2_2_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2809 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i1[9] ), .A3(\SB4_11/i0[6] ), .ZN(\SB4_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2810 ( .A1(\SB2_2_31/i0_4 ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i1[9] ), .ZN(\SB2_2_31/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U2811 ( .A(\RI3[2][182] ), .ZN(\SB2_2_1/i1[9] ) );
  NAND4_X1 U2812 ( .A1(\SB4_4/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_4/Component_Function_4/NAND4_in[3] ), .A3(
        \SB4_4/Component_Function_4/NAND4_in[0] ), .A4(n1220), .ZN(n1310) );
  NAND3_X1 U2813 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i3[0] ), .A3(\SB4_4/i1_7 ), 
        .ZN(n1220) );
  NAND3_X1 U2814 ( .A1(n1657), .A2(\SB1_2_9/i0_0 ), .A3(\SB1_2_9/i0_4 ), .ZN(
        \SB1_2_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2815 ( .A1(\SB1_2_28/i0_3 ), .A2(\SB1_2_28/i0_0 ), .A3(
        \SB1_2_28/i0_4 ), .ZN(\SB1_2_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2816 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i0_0 ), .A3(
        \SB1_1_21/i0_4 ), .ZN(\SB1_1_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2817 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i0_3 ), .A3(\SB3_3/i0[9] ), 
        .ZN(\SB3_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2818 ( .A1(\SB3_7/i0_0 ), .A2(\SB3_7/i1_5 ), .A3(\SB3_7/i0_4 ), 
        .ZN(\SB3_7/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2819 ( .A1(\SB4_2/i0_4 ), .A2(\SB4_2/i1_7 ), .A3(\SB4_2/i0[8] ), 
        .ZN(n1221) );
  NAND3_X1 U2820 ( .A1(\SB2_1_26/i0_4 ), .A2(\RI3[1][30] ), .A3(
        \SB2_1_26/i0[6] ), .ZN(\SB2_1_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2821 ( .A1(\SB4_19/i0_4 ), .A2(\SB4_19/i1[9] ), .A3(\SB4_19/i1_5 ), 
        .ZN(\SB4_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2823 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i0[9] ), .A3(
        \SB2_2_13/i0[10] ), .ZN(\SB2_2_13/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2824 ( .A1(\SB1_2_20/i0_3 ), .A2(\SB1_2_20/i0[9] ), .A3(
        \SB1_2_20/i0[10] ), .ZN(\SB1_2_20/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2827 ( .A1(\SB1_2_31/i0[10] ), .A2(\SB1_2_31/i1_7 ), .A3(
        \SB1_2_31/i1[9] ), .ZN(\SB1_2_31/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U2828 ( .A1(\SB2_2_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_15/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_15/Component_Function_4/NAND4_in[1] ), .A4(n1223), .ZN(
        \RI5[2][106] ) );
  NAND3_X1 U2829 ( .A1(\SB2_2_15/i0_4 ), .A2(\SB2_2_15/i1_5 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(n1223) );
  NAND3_X1 U2832 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i0_0 ), .A3(
        \SB1_2_4/i0_4 ), .ZN(\SB1_2_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2833 ( .A1(\SB2_2_23/i0_4 ), .A2(\SB2_2_23/i0_3 ), .A3(
        \SB2_2_23/i1[9] ), .ZN(n1225) );
  NAND3_X1 U2836 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i0_0 ), .A3(
        \SB2_2_22/i0[6] ), .ZN(\SB2_2_22/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2838 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i1_7 ), .A3(
        \SB1_2_24/i1[9] ), .ZN(\SB1_2_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2839 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i0[9] ), .A3(
        \SB1_1_24/i0[8] ), .ZN(\SB1_1_24/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U2840 ( .A1(\SB1_2_19/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_19/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_19/Component_Function_2/NAND4_in[2] ), .A4(n1227), .ZN(
        \RI3[2][92] ) );
  NAND3_X1 U2841 ( .A1(\SB1_2_19/i0_0 ), .A2(\SB1_2_19/i0_4 ), .A3(
        \SB1_2_19/i1_5 ), .ZN(n1227) );
  NAND3_X1 U2842 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0_0 ), .A3(
        \SB1_0_0/i0_4 ), .ZN(\SB1_0_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2846 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i0_0 ), .A3(\SB4_1/i0_4 ), 
        .ZN(\SB4_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2851 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0_4 ), .A3(
        \SB1_0_14/i1[9] ), .ZN(\SB1_0_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2854 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0_0 ), .A3(
        \SB1_0_14/i0_4 ), .ZN(\SB1_0_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2855 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0[10] ), .A3(
        \SB1_1_9/i0_4 ), .ZN(\SB1_1_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2856 ( .A1(\SB2_0_1/i0_3 ), .A2(\SB2_0_1/i0_4 ), .A3(
        \SB2_0_1/i1[9] ), .ZN(n1230) );
  NAND3_X1 U2857 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0_0 ), .A3(
        \SB1_0_9/i0_4 ), .ZN(\SB1_0_9/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2858 ( .A(\MC_ARK_ARC_1_1/temp5[159] ), .B(n1231), .ZN(
        \RI1[2][159] ) );
  XNOR2_X1 U2859 ( .A(\MC_ARK_ARC_1_1/temp3[159] ), .B(
        \MC_ARK_ARC_1_1/temp4[159] ), .ZN(n1231) );
  NAND3_X1 U2860 ( .A1(\SB2_1_22/i1_5 ), .A2(\SB2_1_22/i3[0] ), .A3(
        \SB2_1_22/i0[8] ), .ZN(n1232) );
  NAND3_X1 U2861 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0[9] ), .A3(
        \SB1_1_0/i0[10] ), .ZN(\SB1_1_0/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U2862 ( .A(n1233), .B(n373), .ZN(Ciphertext[84]) );
  NAND4_X1 U2863 ( .A1(\SB4_17/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_17/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_17/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_17/Component_Function_0/NAND4_in[1] ), .ZN(n1233) );
  NAND3_X1 U2864 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i0_4 ), .A3(
        \SB2_1_11/i1[9] ), .ZN(\SB2_1_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2865 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i1[9] ), .A3(
        \SB1_1_22/i0_4 ), .ZN(n1366) );
  NAND3_X1 U2866 ( .A1(\SB1_3_14/i0_3 ), .A2(\SB1_3_14/i0[10] ), .A3(
        \SB1_3_14/i0[9] ), .ZN(n1250) );
  NAND4_X1 U2867 ( .A1(\SB2_3_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_5/NAND4_in[0] ), .A4(n1234), .ZN(
        \RI5[3][113] ) );
  NAND3_X1 U2868 ( .A1(\SB2_3_13/i0_4 ), .A2(\RI3[3][108] ), .A3(\RI3[3][109] ), .ZN(n1234) );
  INV_X2 U2869 ( .A(\RI1[1][155] ), .ZN(\SB1_1_6/i0_3 ) );
  XNOR2_X1 U2870 ( .A(\MC_ARK_ARC_1_0/temp5[155] ), .B(
        \MC_ARK_ARC_1_0/temp6[155] ), .ZN(\RI1[1][155] ) );
  NAND3_X1 U2871 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0[9] ), .A3(
        \SB1_2_26/i0[8] ), .ZN(\SB1_2_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2873 ( .A1(\SB2_0_31/i0[10] ), .A2(\SB2_0_31/i0_0 ), .A3(
        \SB2_0_31/i0[6] ), .ZN(\SB2_0_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 U2874 ( .A1(\SB2_0_20/i0_0 ), .A2(\SB2_0_20/i3[0] ), .ZN(n1235) );
  NAND3_X1 U2875 ( .A1(\SB2_1_15/i0[9] ), .A2(\SB2_1_15/i0_3 ), .A3(
        \SB2_1_15/i0[8] ), .ZN(n1236) );
  XNOR2_X1 U2880 ( .A(\MC_ARK_ARC_1_1/temp1[35] ), .B(
        \MC_ARK_ARC_1_1/temp3[35] ), .ZN(n1239) );
  XNOR2_X1 U2881 ( .A(n1241), .B(n1240), .ZN(\RI1[2][65] ) );
  XNOR2_X1 U2882 ( .A(\MC_ARK_ARC_1_1/temp4[65] ), .B(
        \MC_ARK_ARC_1_1/temp2[65] ), .ZN(n1240) );
  XNOR2_X1 U2883 ( .A(\MC_ARK_ARC_1_1/temp1[65] ), .B(
        \MC_ARK_ARC_1_1/temp3[65] ), .ZN(n1241) );
  NAND3_X1 U2884 ( .A1(\SB1_1_27/i0_3 ), .A2(\SB1_1_27/i0[10] ), .A3(
        \SB1_1_27/i0[9] ), .ZN(\SB1_1_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2885 ( .A1(\RI3[3][94] ), .A2(\SB2_3_16/i0_3 ), .A3(
        \SB2_3_16/i1[9] ), .ZN(n1242) );
  XNOR2_X1 U2887 ( .A(\MC_ARK_ARC_1_2/temp5[20] ), .B(n1244), .ZN(\RI1[3][20] ) );
  XNOR2_X1 U2888 ( .A(\MC_ARK_ARC_1_2/temp3[20] ), .B(
        \MC_ARK_ARC_1_2/temp4[20] ), .ZN(n1244) );
  NAND4_X1 U2889 ( .A1(\SB2_2_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_8/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_8/Component_Function_2/NAND4_in[1] ), .A4(n1245), .ZN(
        \RI5[2][158] ) );
  NAND3_X1 U2890 ( .A1(\SB2_2_8/i0_4 ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i0_0 ), .ZN(n1245) );
  NAND2_X1 U2892 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB2_3_23/i3[0] ), .ZN(n1246) );
  NAND4_X1 U2893 ( .A1(\SB1_2_31/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_2_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_31/Component_Function_2/NAND4_in[1] ), .A4(n1247), .ZN(
        \RI3[2][20] ) );
  XNOR2_X1 U2894 ( .A(n1248), .B(n1315), .ZN(\RI1[4][59] ) );
  XNOR2_X1 U2895 ( .A(\MC_ARK_ARC_1_3/temp1[59] ), .B(
        \MC_ARK_ARC_1_3/temp4[59] ), .ZN(n1248) );
  NAND3_X1 U2897 ( .A1(\SB2_2_28/i0_0 ), .A2(\SB2_2_28/i0_4 ), .A3(
        \SB2_2_28/i1_5 ), .ZN(\SB2_2_28/Component_Function_2/NAND4_in[3] ) );
  INV_X2 U2898 ( .A(\RI1[3][95] ), .ZN(\SB1_3_16/i0_3 ) );
  XNOR2_X1 U2899 ( .A(\MC_ARK_ARC_1_2/temp6[95] ), .B(
        \MC_ARK_ARC_1_2/temp5[95] ), .ZN(\RI1[3][95] ) );
  NAND3_X1 U2902 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0[9] ), .A3(
        \SB1_0_15/i0[10] ), .ZN(\SB1_0_15/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2903 ( .A1(\SB1_1_27/i0_3 ), .A2(\SB1_1_27/i0_0 ), .A3(
        \SB1_1_27/i0_4 ), .ZN(\SB1_1_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2904 ( .A1(\SB1_2_29/i0_3 ), .A2(\SB1_2_29/i0[10] ), .A3(
        \SB1_2_29/i0[9] ), .ZN(\SB1_2_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2905 ( .A1(\SB1_3_20/i1_7 ), .A2(\SB1_3_20/i0[10] ), .A3(
        \SB1_3_20/i1[9] ), .ZN(\SB1_3_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2906 ( .A1(\SB2_2_27/i0[8] ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB2_2_27/i3[0] ), .ZN(\SB2_2_27/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U2907 ( .A1(\SB2_0_4/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[167] ) );
  NAND3_X1 U2908 ( .A1(\SB1_2_15/i0_3 ), .A2(\SB1_2_15/i0[7] ), .A3(
        \SB1_2_15/i0_0 ), .ZN(\SB1_2_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2909 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i0[9] ), .A3(
        \SB1_0_26/i0[8] ), .ZN(\SB1_0_26/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2913 ( .A(n1253), .B(n213), .ZN(Ciphertext[67]) );
  NAND3_X1 U2914 ( .A1(n858), .A2(\SB4_6/i1[9] ), .A3(\SB4_6/i0[6] ), .ZN(
        \SB4_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2915 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i0_0 ), .A3(
        \SB2_3_21/i0[6] ), .ZN(\SB2_3_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2916 ( .A1(n828), .A2(\SB4_12/i1[9] ), .A3(\SB4_12/i0[6] ), .ZN(
        \SB4_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2917 ( .A1(n863), .A2(\SB4_8/i1[9] ), .A3(\SB4_8/i0[6] ), .ZN(
        \SB4_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2918 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0_0 ), .A3(
        \SB1_2_21/i0_4 ), .ZN(\SB1_2_21/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2919 ( .A(n1254), .B(n298), .ZN(Ciphertext[68]) );
  NAND4_X1 U2920 ( .A1(\SB4_20/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_20/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_20/Component_Function_2/NAND4_in[3] ), .A4(
        \SB4_20/Component_Function_2/NAND4_in[0] ), .ZN(n1254) );
  NAND3_X1 U2921 ( .A1(\SB2_0_26/i0_4 ), .A2(\SB2_0_26/i0_3 ), .A3(
        \SB2_0_26/i1[9] ), .ZN(\SB2_0_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2922 ( .A1(\SB4_25/i0_4 ), .A2(\SB4_25/i1_7 ), .A3(\SB4_25/i0[8] ), 
        .ZN(\SB4_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2923 ( .A1(\SB3_21/i0[9] ), .A2(\SB3_21/i0[10] ), .A3(
        \SB3_21/i0_3 ), .ZN(\SB3_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2924 ( .A1(n799), .A2(\SB4_14/i1_7 ), .A3(\SB4_14/i0[8] ), .ZN(
        n1255) );
  NAND3_X1 U2927 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0[9] ), .A3(
        \SB1_0_12/i0[8] ), .ZN(\SB1_0_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2928 ( .A1(\SB1_2_1/i0_3 ), .A2(\SB1_2_1/i0_0 ), .A3(
        \SB1_2_1/i0_4 ), .ZN(\SB1_2_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2929 ( .A1(\SB2_2_8/i0[9] ), .A2(\SB2_2_8/i0_3 ), .A3(
        \SB2_2_8/i0[8] ), .ZN(\SB2_2_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2930 ( .A1(\SB2_2_25/i0[9] ), .A2(\SB2_2_25/i0_3 ), .A3(
        \SB2_2_25/i0[8] ), .ZN(\SB2_2_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2931 ( .A1(\SB2_2_5/i0[9] ), .A2(\SB2_2_5/i0_3 ), .A3(
        \SB2_2_5/i0[8] ), .ZN(\SB2_2_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2932 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i0_3 ), .A3(
        \SB2_1_28/i1[9] ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2933 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0_0 ), .A3(
        \SB1_1_6/i0_4 ), .ZN(\SB1_1_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2936 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0[9] ), .A3(
        \SB2_0_16/i0[8] ), .ZN(\SB2_0_16/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U2937 ( .A1(\SB2_2_20/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_20/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_20/Component_Function_4/NAND4_in[1] ), .A4(n1257), .ZN(
        \RI5[2][76] ) );
  NAND3_X1 U2938 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0[10] ), .A3(
        \SB2_2_20/i0[9] ), .ZN(n1257) );
  NAND4_X1 U2941 ( .A1(\SB3_21/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_21/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_5/NAND4_in[0] ), .A4(n1259), .ZN(
        \RI3[4][65] ) );
  NAND3_X1 U2942 ( .A1(\SB3_21/i1[9] ), .A2(\SB3_21/i0_3 ), .A3(\SB3_21/i0_4 ), 
        .ZN(n1259) );
  NAND3_X1 U2944 ( .A1(\SB2_2_2/i1_5 ), .A2(\SB2_2_2/i3[0] ), .A3(
        \SB2_2_2/i0[8] ), .ZN(n1260) );
  NAND3_X1 U2945 ( .A1(\SB2_1_7/i0_4 ), .A2(\SB2_1_7/i1_7 ), .A3(
        \SB2_1_7/i0[8] ), .ZN(\SB2_1_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2947 ( .A1(\SB2_1_0/i3[0] ), .A2(\SB2_1_0/i1_5 ), .A3(
        \SB2_1_0/i0[8] ), .ZN(n1261) );
  NAND3_X1 U2948 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i1[9] ), .A3(\SB4_28/i0[6] ), .ZN(\SB4_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2949 ( .A1(\SB1_1_2/i1_7 ), .A2(\SB1_1_2/i0[10] ), .A3(
        \SB1_1_2/i1[9] ), .ZN(\SB1_1_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2950 ( .A1(\SB3_25/i0[9] ), .A2(\SB3_25/i0_3 ), .A3(
        \SB3_25/i0[10] ), .ZN(\SB3_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2951 ( .A1(\SB4_5/i0_3 ), .A2(\SB4_5/i0[10] ), .A3(\SB4_5/i0[9] ), 
        .ZN(\SB4_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2952 ( .A1(\SB1_0_4/i0_3 ), .A2(\SB1_0_4/i0_4 ), .A3(
        \SB1_0_4/i1[9] ), .ZN(\SB1_0_4/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U2953 ( .A1(\SB1_2_14/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_14/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_14/Component_Function_5/NAND4_in[0] ), .A4(n1262), .ZN(
        \RI3[2][107] ) );
  NAND3_X1 U2954 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i1[9] ), .A3(
        \SB1_2_14/i0_4 ), .ZN(n1262) );
  NAND3_X1 U2955 ( .A1(\SB1_0_9/i0[10] ), .A2(\SB1_0_9/i1_7 ), .A3(
        \SB1_0_9/i1[9] ), .ZN(\SB1_0_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2956 ( .A1(\SB2_0_11/i0_4 ), .A2(\SB2_0_11/i0_0 ), .A3(
        \SB2_0_11/i0_3 ), .ZN(\SB2_0_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2957 ( .A1(\SB4_5/i0_3 ), .A2(\SB4_5/i1[9] ), .A3(n810), .ZN(
        \SB4_5/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U2959 ( .A1(\SB2_2_6/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_6/Component_Function_4/NAND4_in[1] ), .A4(n1264), .ZN(
        \RI5[2][160] ) );
  NAND3_X1 U2960 ( .A1(\SB2_2_6/i0_4 ), .A2(\SB2_2_6/i1_5 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(n1264) );
  NAND4_X1 U2962 ( .A1(\SB1_1_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_3/NAND4_in[2] ), .A4(n1265), .ZN(
        \RI3[1][81] ) );
  NAND3_X1 U2963 ( .A1(\SB1_1_20/i3[0] ), .A2(\SB1_1_20/i1_5 ), .A3(
        \SB1_1_20/i0[8] ), .ZN(n1265) );
  NAND4_X1 U2964 ( .A1(\SB1_2_25/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_25/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_25/Component_Function_5/NAND4_in[0] ), .A4(n1266), .ZN(
        \RI3[2][41] ) );
  NAND4_X1 U2965 ( .A1(\SB1_0_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_25/Component_Function_0/NAND4_in[0] ), .A4(n1267), .ZN(
        \RI3[0][66] ) );
  NAND3_X1 U2967 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0_4 ), .A3(\SB4_15/i0_0 ), 
        .ZN(\SB4_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2969 ( .A1(\SB2_1_1/i0[9] ), .A2(\SB2_1_1/i0_3 ), .A3(
        \SB2_1_1/i0[8] ), .ZN(n1268) );
  NAND3_X1 U2970 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i0[10] ), .A3(
        \SB1_2_16/i0[9] ), .ZN(\SB1_2_16/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2971 ( .A1(\SB1_1_3/i1[9] ), .A2(\SB1_1_3/i0[10] ), .A3(
        \SB1_1_3/i1_7 ), .ZN(\SB1_1_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2972 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[9] ), .A3(
        \SB1_1_22/i0[10] ), .ZN(\SB1_1_22/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2973 ( .A1(\SB2_1_3/i1_5 ), .A2(\SB2_1_3/i3[0] ), .A3(
        \SB2_1_3/i0[8] ), .ZN(\SB2_1_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2974 ( .A1(\SB1_1_5/i0_3 ), .A2(\SB1_1_5/i0_0 ), .A3(
        \SB1_1_5/i0_4 ), .ZN(\SB1_1_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2975 ( .A1(\SB2_0_4/i0_4 ), .A2(\SB2_0_4/i0[9] ), .A3(
        \SB2_0_4/i0[6] ), .ZN(\SB2_0_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2976 ( .A1(\SB2_0_20/i0_0 ), .A2(\SB2_0_20/i0[7] ), .A3(
        \SB2_0_20/i0_3 ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U2977 ( .A(n1269), .B(n1314), .ZN(\RI1[2][189] ) );
  XNOR2_X1 U2978 ( .A(\MC_ARK_ARC_1_1/temp2[189] ), .B(
        \MC_ARK_ARC_1_1/temp3[189] ), .ZN(n1269) );
  NAND3_X1 U2979 ( .A1(\SB2_1_11/i3[0] ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB2_1_11/i0[8] ), .ZN(\SB2_1_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2980 ( .A1(\SB2_1_1/i3[0] ), .A2(\SB2_1_1/i1_5 ), .A3(
        \SB2_1_1/i0[8] ), .ZN(\SB2_1_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2981 ( .A1(\SB1_2_0/i1_7 ), .A2(\SB1_2_0/i0[10] ), .A3(
        \SB1_2_0/i1[9] ), .ZN(\SB1_2_0/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U2987 ( .A1(\SB1_0_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_1/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_1/Component_Function_1/NAND4_in[0] ), .A4(n1270), .ZN(
        \RI3[0][13] ) );
  NAND4_X4 U2989 ( .A1(\SB2_0_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_19/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[77] ) );
  XNOR2_X1 U2990 ( .A(\MC_ARK_ARC_1_2/temp5[131] ), .B(n1271), .ZN(
        \RI1[3][131] ) );
  XNOR2_X1 U2991 ( .A(\MC_ARK_ARC_1_2/temp3[131] ), .B(
        \MC_ARK_ARC_1_2/temp4[131] ), .ZN(n1271) );
  NAND3_X1 U2992 ( .A1(\SB2_3_9/i0_4 ), .A2(\SB2_3_9/i0_3 ), .A3(
        \SB2_3_9/i1[9] ), .ZN(n1272) );
  NAND3_X1 U2993 ( .A1(\SB4_21/i0_3 ), .A2(\SB4_21/i1[9] ), .A3(\SB4_21/i0[6] ), .ZN(\SB4_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2994 ( .A1(\SB1_1_18/i0_3 ), .A2(\SB1_1_18/i0[9] ), .A3(
        \SB1_1_18/i0[8] ), .ZN(\SB1_1_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2995 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i0_0 ), .A3(
        \SB2_1_9/i0[6] ), .ZN(\SB2_1_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2996 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i0_0 ), .A3(\SB4_16/i0_4 ), 
        .ZN(\SB4_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2997 ( .A1(\SB1_1_11/i0_3 ), .A2(\SB1_1_11/i0_0 ), .A3(
        \SB1_1_11/i0_4 ), .ZN(\SB1_1_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2998 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i0_0 ), .A3(
        \SB1_2_16/i0_4 ), .ZN(\SB1_2_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2999 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0[9] ), .A3(
        \SB1_2_26/i0[10] ), .ZN(\SB1_2_26/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3000 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i0[8] ), .ZN(n1273) );
  NAND3_X1 U3001 ( .A1(\SB1_2_28/i0_3 ), .A2(\SB1_2_28/i0[10] ), .A3(
        \SB1_2_28/i0[9] ), .ZN(\SB1_2_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3002 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i1[9] ), .A3(\SB4_0/i0[6] ), 
        .ZN(\SB4_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3003 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i0_0 ), .A3(
        \SB1_0_19/i0_4 ), .ZN(\SB1_0_19/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U3004 ( .A1(\SB2_1_20/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_20/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_20/Component_Function_2/NAND4_in[1] ), .A4(n1274), .ZN(
        \RI5[1][86] ) );
  NAND3_X1 U3005 ( .A1(\SB2_1_20/i0_4 ), .A2(\SB2_1_20/i1_5 ), .A3(
        \SB2_1_20/i0_0 ), .ZN(n1274) );
  NAND3_X1 U3006 ( .A1(n1672), .A2(\SB4_0/i0[9] ), .A3(\SB4_0/i0[10] ), .ZN(
        \SB4_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3007 ( .A1(n1672), .A2(\SB4_0/i0_4 ), .A3(\SB4_0/i1[9] ), .ZN(
        \SB4_0/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U3008 ( .A1(\SB4_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_0/Component_Function_1/NAND4_in[0] ), .A3(
        \SB4_0/Component_Function_1/NAND4_in[3] ), .A4(n1275), .ZN(
        \RI4[4][187] ) );
  NAND3_X1 U3009 ( .A1(\SB4_0/i0[9] ), .A2(\SB4_0/i0[6] ), .A3(\SB4_0/i1_5 ), 
        .ZN(n1275) );
  NAND3_X1 U3011 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i0_0 ), .A3(
        \SB1_2_18/i0_4 ), .ZN(\SB1_2_18/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U3012 ( .A1(\SB3_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_0/NAND4_in[0] ), .A4(n1277), .ZN(
        \RI3[4][186] ) );
  NAND4_X2 U3013 ( .A1(\SB1_3_27/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_27/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_3_27/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_26/i0_4 ) );
  NAND3_X1 U3014 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i0[9] ), .A3(
        \SB1_3_5/i0[8] ), .ZN(\SB1_3_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3015 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i0[7] ), .A3(\SB4_1/i0_0 ), 
        .ZN(\SB4_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3016 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0_0 ), .A3(
        \SB1_0_8/i0_4 ), .ZN(\SB1_0_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3018 ( .A1(\SB4_28/i0_4 ), .A2(\SB4_28/i1_7 ), .A3(\SB4_28/i0[8] ), 
        .ZN(n1278) );
  NAND3_X1 U3019 ( .A1(\SB1_2_15/i1_7 ), .A2(\SB1_2_15/i0[10] ), .A3(
        \SB1_2_15/i1[9] ), .ZN(\SB1_2_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3020 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0_0 ), .A3(
        \SB1_1_23/i0_4 ), .ZN(\SB1_1_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3021 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i0_0 ), .A3(
        \SB1_2_8/i0_4 ), .ZN(\SB1_2_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3023 ( .A1(\SB2_2_10/i0_3 ), .A2(\SB2_2_10/i0[9] ), .A3(
        \SB2_2_10/i0[8] ), .ZN(\SB2_2_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3024 ( .A1(\SB2_2_9/i0_3 ), .A2(\SB2_2_9/i0[9] ), .A3(
        \SB2_2_9/i0[8] ), .ZN(\SB2_2_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3026 ( .A1(\SB2_1_0/i0[9] ), .A2(\SB2_1_0/i0_3 ), .A3(
        \SB2_1_0/i0[8] ), .ZN(\SB2_1_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3027 ( .A1(\SB4_29/i0_3 ), .A2(\SB4_29/i1[9] ), .A3(n791), .ZN(
        \SB4_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3028 ( .A1(\SB2_2_7/i0_4 ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0[6] ), .ZN(\SB2_2_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3029 ( .A1(n1668), .A2(\SB4_30/i0_4 ), .A3(\SB4_30/i0_0 ), .ZN(
        \SB4_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3030 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i0_0 ), .A3(n799), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3031 ( .A1(\SB1_2_11/i1_7 ), .A2(\SB1_2_11/i0[10] ), .A3(
        \SB1_2_11/i1[9] ), .ZN(\SB1_2_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3032 ( .A1(\SB1_1_2/i0_3 ), .A2(\SB1_1_2/i0_0 ), .A3(
        \SB1_1_2/i0_4 ), .ZN(\SB1_1_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3033 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0_0 ), .A3(
        \SB1_2_12/i0_4 ), .ZN(\SB1_2_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3034 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i0[9] ), .A3(
        \SB1_2_8/i0[10] ), .ZN(\SB1_2_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3035 ( .A1(\SB1_2_6/i0_3 ), .A2(\SB1_2_6/i0[10] ), .A3(
        \SB1_2_6/i0[9] ), .ZN(\SB1_2_6/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U3036 ( .A1(\SB2_3_15/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_3_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_15/Component_Function_5/NAND4_in[0] ), .A4(n1280), .ZN(
        \RI5[3][101] ) );
  NAND4_X1 U3037 ( .A1(\SB4_20/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_20/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_20/Component_Function_0/NAND4_in[0] ), .A4(n1281), .ZN(n1401) );
  NAND3_X1 U3038 ( .A1(\SB4_20/i0[6] ), .A2(\SB4_20/i0[8] ), .A3(n548), .ZN(
        n1281) );
  NAND3_X1 U3039 ( .A1(\SB2_2_31/i3[0] ), .A2(\SB2_2_31/i1_5 ), .A3(
        \SB2_2_31/i0[8] ), .ZN(\SB2_2_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3041 ( .A1(\SB2_0_16/i0[8] ), .A2(\SB2_0_16/i1_5 ), .A3(
        \SB2_0_16/i3[0] ), .ZN(\SB2_0_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3042 ( .A1(\SB2_1_9/i0[8] ), .A2(\SB2_1_9/i1_5 ), .A3(
        \SB2_1_9/i3[0] ), .ZN(\SB2_1_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3044 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i0[9] ), .A3(
        \SB1_2_2/i0[8] ), .ZN(\SB1_2_2/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3045 ( .A(\MC_ARK_ARC_1_2/temp5[69] ), .B(n1282), .ZN(\RI1[3][69] ) );
  XNOR2_X1 U3046 ( .A(\MC_ARK_ARC_1_2/temp3[69] ), .B(
        \MC_ARK_ARC_1_2/temp4[69] ), .ZN(n1282) );
  NAND3_X1 U3047 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i1[9] ), .A3(\SB4_24/i0[6] ), .ZN(\SB4_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3050 ( .A1(n2135), .A2(\SB4_24/i0[9] ), .A3(\SB4_24/i0[10] ), .ZN(
        \SB4_24/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U3051 ( .A1(\SB2_1_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_23/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_23/Component_Function_2/NAND4_in[3] ), .A4(n1283), .ZN(
        \RI5[1][68] ) );
  NAND3_X1 U3052 ( .A1(\SB4_18/i0_4 ), .A2(n2113), .A3(\SB4_18/i1_5 ), .ZN(
        n1285) );
  NAND4_X1 U3053 ( .A1(\SB1_2_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_26/Component_Function_2/NAND4_in[2] ), .A4(n1286), .ZN(
        \RI3[2][50] ) );
  NAND3_X1 U3054 ( .A1(\SB1_2_26/i0_0 ), .A2(\SB1_2_26/i1_5 ), .A3(
        \SB1_2_26/i0_4 ), .ZN(n1286) );
  XNOR2_X1 U3057 ( .A(n1288), .B(n265), .ZN(Ciphertext[18]) );
  NAND4_X1 U3058 ( .A1(\SB4_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_28/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_28/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_28/Component_Function_0/NAND4_in[1] ), .ZN(n1288) );
  XNOR2_X1 U3059 ( .A(n1289), .B(n409), .ZN(Ciphertext[21]) );
  NAND3_X1 U3061 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0[9] ), .A3(
        \SB1_1_30/i0[8] ), .ZN(\SB1_1_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3062 ( .A1(n1672), .A2(\SB4_0/i0[8] ), .A3(\SB4_0/i1_7 ), .ZN(
        \SB4_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3063 ( .A1(\SB1_1_2/i0_3 ), .A2(\SB1_1_2/i0_4 ), .A3(
        \SB1_1_2/i1[9] ), .ZN(n1394) );
  NAND3_X1 U3064 ( .A1(n2135), .A2(\SB4_24/i0_4 ), .A3(\SB4_24/i0_0 ), .ZN(
        \SB4_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3065 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0_0 ), .A3(\SB4_24/i0[7] ), 
        .ZN(\SB4_24/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U3066 ( .A1(\SB1_2_4/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_2_4/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[2][182] ) );
  NAND3_X1 U3068 ( .A1(\SB2_0_17/i0_4 ), .A2(\RI3[0][84] ), .A3(
        \SB2_0_17/i0[6] ), .ZN(n1290) );
  NAND3_X1 U3070 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0_0 ), .A3(
        \SB1_1_22/i0_4 ), .ZN(\SB1_1_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3071 ( .A1(\SB4_29/i0_3 ), .A2(n2131), .A3(\SB4_29/i1[9] ), .ZN(
        \SB4_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3072 ( .A1(\SB4_29/i0_3 ), .A2(n790), .A3(\SB4_29/i0[10] ), .ZN(
        \SB4_29/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U3073 ( .A(n1291), .B(n1292), .ZN(\RI1[3][122] ) );
  XNOR2_X1 U3074 ( .A(\MC_ARK_ARC_1_2/temp3[122] ), .B(
        \MC_ARK_ARC_1_2/temp1[122] ), .ZN(n1291) );
  XNOR2_X1 U3075 ( .A(\MC_ARK_ARC_1_2/temp2[122] ), .B(
        \MC_ARK_ARC_1_2/temp4[122] ), .ZN(n1292) );
  NAND4_X1 U3076 ( .A1(\SB3_20/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_20/Component_Function_2/NAND4_in[3] ), .A4(
        \SB3_20/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[4][86] ) );
  NAND3_X1 U3079 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0_0 ), .A3(
        \SB1_1_0/i0_4 ), .ZN(\SB1_1_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3080 ( .A1(\SB2_1_21/i0[8] ), .A2(\SB2_1_21/i1_5 ), .A3(
        \SB2_1_21/i3[0] ), .ZN(\SB2_1_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3085 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0_4 ), .A3(\SB3_2/i0[10] ), 
        .ZN(\SB3_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3086 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0_4 ), .A3(
        \SB1_0_15/i1[9] ), .ZN(n1308) );
  NAND3_X1 U3088 ( .A1(\SB1_0_3/i0_3 ), .A2(\SB1_0_3/i0_4 ), .A3(
        \SB1_0_3/i1[9] ), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3089 ( .A1(\SB2_0_20/i0_0 ), .A2(\SB2_0_20/i0_4 ), .A3(
        \SB2_0_20/i0_3 ), .ZN(\SB2_0_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3091 ( .A1(n790), .A2(\SB4_29/i1_5 ), .A3(n791), .ZN(n1296) );
  NAND3_X1 U3092 ( .A1(\SB2_1_28/i3[0] ), .A2(\SB2_1_28/i1_5 ), .A3(
        \SB2_1_28/i0[8] ), .ZN(\SB2_1_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3093 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i0_0 ), .A3(
        \SB1_0_17/i0_4 ), .ZN(\SB1_0_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3095 ( .A1(\SB4_31/i0_4 ), .A2(\SB4_31/i1_7 ), .A3(\SB4_31/i0[8] ), 
        .ZN(n1297) );
  NAND3_X1 U3096 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i0[9] ), .A3(
        \SB1_2_4/i0[10] ), .ZN(\SB1_2_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3097 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB2_3_30/i1[9] ), .ZN(\SB2_3_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3099 ( .A1(n2100), .A2(\SB4_23/i0_4 ), .A3(\SB4_23/i0_0 ), .ZN(
        \SB4_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3101 ( .A1(\SB4_26/i0_3 ), .A2(\SB4_26/i0_0 ), .A3(\SB4_26/i0_4 ), 
        .ZN(\SB4_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3102 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0_0 ), .A3(
        \SB1_1_20/i0_4 ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3103 ( .A1(\SB4_3/i0_4 ), .A2(\SB4_3/i1_7 ), .A3(\SB4_3/i0[8] ), 
        .ZN(n1298) );
  NAND3_X1 U3104 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i0_4 ), .ZN(\SB1_2_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3105 ( .A1(\SB4_16/i0_4 ), .A2(\SB4_16/i1_7 ), .A3(\SB4_16/i0[8] ), 
        .ZN(n1299) );
  NAND4_X1 U3106 ( .A1(\SB2_2_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_26/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_26/Component_Function_3/NAND4_in[2] ), .A4(n1300), .ZN(
        \RI5[2][45] ) );
  NAND3_X1 U3107 ( .A1(\SB2_2_26/i3[0] ), .A2(\SB2_2_26/i1_5 ), .A3(
        \SB2_2_26/i0[8] ), .ZN(n1300) );
  NAND3_X1 U3108 ( .A1(\SB2_2_15/i0[8] ), .A2(\SB2_2_15/i1_5 ), .A3(
        \SB2_2_15/i3[0] ), .ZN(\SB2_2_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3110 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0[9] ), .A3(
        \SB1_1_23/i0[8] ), .ZN(\SB1_1_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3112 ( .A1(n2100), .A2(\SB4_23/i0_4 ), .A3(\SB4_23/i0[10] ), .ZN(
        \SB4_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3113 ( .A1(\SB2_0_3/i0[8] ), .A2(\SB2_0_3/i1_5 ), .A3(
        \SB2_0_3/i3[0] ), .ZN(\SB2_0_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3118 ( .A1(\SB2_2_21/i0[8] ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB2_2_21/i3[0] ), .ZN(\SB2_2_21/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U3119 ( .A(\RI3[1][179] ), .ZN(\SB2_1_2/i1_5 ) );
  NAND4_X1 U3120 ( .A1(\SB1_1_2/Component_Function_5/NAND4_in[1] ), .A2(n1394), 
        .A3(\SB1_1_2/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_1_2/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[1][179] ) );
  NAND3_X1 U3121 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0[9] ), .A3(
        \SB2_2_24/i0[10] ), .ZN(\SB2_2_24/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3122 ( .A1(\SB1_2_23/i0[10] ), .A2(\SB1_2_23/i1_7 ), .A3(
        \SB1_2_23/i1[9] ), .ZN(\SB1_2_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3123 ( .A1(\SB4_10/i0_3 ), .A2(\SB4_10/i1[9] ), .A3(\SB4_10/i0[6] ), .ZN(\SB4_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3124 ( .A1(\SB4_10/i0_4 ), .A2(\SB4_10/i0_3 ), .A3(\SB4_10/i1[9] ), 
        .ZN(\SB4_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3125 ( .A1(\SB4_10/i0_3 ), .A2(\SB4_10/i0[9] ), .A3(
        \SB4_10/i0[10] ), .ZN(\SB4_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3127 ( .A1(\SB3_22/i0_3 ), .A2(\SB3_22/i0_4 ), .A3(\SB3_22/i1[9] ), 
        .ZN(\SB3_22/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3128 ( .A(n1303), .B(n196), .ZN(Ciphertext[97]) );
  NAND3_X1 U3129 ( .A1(n859), .A2(\SB4_3/i0_4 ), .A3(\SB4_3/i0_0 ), .ZN(
        \SB4_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3131 ( .A1(n854), .A2(\SB4_21/i0_4 ), .A3(\SB4_21/i0_0 ), .ZN(
        \SB4_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3132 ( .A1(\RI3[4][136] ), .A2(\SB4_9/i1_7 ), .A3(\SB4_9/i0[8] ), 
        .ZN(\SB4_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3133 ( .A1(\SB2_2_22/i0_4 ), .A2(\SB2_2_22/i0[9] ), .A3(
        \SB2_2_22/i0[6] ), .ZN(\SB2_2_22/Component_Function_5/NAND4_in[3] ) );
  NAND4_X1 U3134 ( .A1(\SB1_2_31/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_31/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_2_31/Component_Function_3/NAND4_in[2] ), .A4(n1304), .ZN(
        \RI3[2][15] ) );
  NAND3_X1 U3135 ( .A1(\SB1_2_31/i3[0] ), .A2(\SB1_2_31/i1_5 ), .A3(
        \SB1_2_31/i0[8] ), .ZN(n1304) );
  NAND3_X1 U3136 ( .A1(\SB1_1_29/i0_3 ), .A2(\SB1_1_29/i0_0 ), .A3(
        \SB1_1_29/i0_4 ), .ZN(\SB1_1_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3137 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0_0 ), .A3(
        \SB1_1_10/i0_4 ), .ZN(\SB1_1_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3138 ( .A1(\SB2_1_27/i0[8] ), .A2(\SB2_1_27/i1_5 ), .A3(
        \SB2_1_27/i3[0] ), .ZN(\SB2_1_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3141 ( .A1(\SB1_0_27/i0_3 ), .A2(\SB1_0_27/i0[9] ), .A3(
        \SB1_0_27/i0[8] ), .ZN(\SB1_0_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3142 ( .A1(\SB1_2_23/i0_3 ), .A2(\SB1_2_23/i0_0 ), .A3(
        \SB1_2_23/i0_4 ), .ZN(\SB1_2_23/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U3143 ( .A(n1306), .B(n360), .ZN(Ciphertext[86]) );
  NAND3_X1 U3144 ( .A1(\SB2_1_23/i0_4 ), .A2(\SB2_1_23/i0_3 ), .A3(
        \SB2_1_23/i1[9] ), .ZN(n1307) );
  NAND4_X1 U3145 ( .A1(\SB1_0_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_0_15/Component_Function_5/NAND4_in[0] ), .A4(n1308), .ZN(
        \RI3[0][101] ) );
  NAND3_X1 U3146 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0[9] ), .A3(
        \SB1_1_14/i0[10] ), .ZN(\SB1_1_14/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3147 ( .A1(\SB4_17/i0_0 ), .A2(\SB4_17/i1_5 ), .A3(\SB4_17/i0_4 ), 
        .ZN(n1309) );
  NAND3_X1 U3149 ( .A1(n851), .A2(\SB4_22/i1[9] ), .A3(\SB4_22/i0_4 ), .ZN(
        \SB4_22/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3150 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i1_7 ), .A3(n550), .ZN(
        \SB4_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3151 ( .A1(\SB1_0_31/i0_3 ), .A2(\SB1_0_31/i0[9] ), .A3(
        \SB1_0_31/i0[8] ), .ZN(\SB1_0_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3152 ( .A1(\SB2_0_11/i0_4 ), .A2(\SB2_0_11/i0_3 ), .A3(
        \SB2_0_11/i1[9] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3153 ( .A1(\SB1_1_25/i0_3 ), .A2(\SB1_1_25/i0[10] ), .A3(
        \SB1_1_25/i0[9] ), .ZN(\SB1_1_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3154 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i0_0 ), .A3(
        \SB1_2_31/i0_4 ), .ZN(\SB1_2_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3155 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i0_0 ), .A3(
        \SB1_1_17/i0_4 ), .ZN(\SB1_1_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3156 ( .A1(\SB2_2_12/i0[8] ), .A2(\SB2_2_12/i3[0] ), .A3(
        \SB2_2_12/i1_5 ), .ZN(\SB2_2_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3157 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[9] ), .A3(
        \SB2_2_29/i0[8] ), .ZN(\SB2_2_29/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3158 ( .A(n1310), .B(n193), .ZN(Ciphertext[166]) );
  NAND3_X1 U3159 ( .A1(\SB2_1_15/i3[0] ), .A2(\SB2_1_15/i1_5 ), .A3(
        \SB2_1_15/i0[8] ), .ZN(\SB2_1_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3162 ( .A1(\SB2_2_17/i3[0] ), .A2(\SB2_2_17/i1_5 ), .A3(
        \SB2_2_17/i0[8] ), .ZN(n1311) );
  NAND3_X1 U3164 ( .A1(\SB4_15/i0_4 ), .A2(\SB4_15/i1_5 ), .A3(\SB4_15/i0_0 ), 
        .ZN(n1312) );
  NAND3_X1 U3165 ( .A1(n854), .A2(\SB4_21/i0_4 ), .A3(\SB4_21/i1[9] ), .ZN(
        \SB4_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3166 ( .A1(\SB1_1_12/i0_3 ), .A2(\SB1_1_12/i0_0 ), .A3(
        \SB1_1_12/i0_4 ), .ZN(\SB1_1_12/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U3167 ( .A(n1313), .B(n306), .ZN(Ciphertext[53]) );
  NAND4_X1 U3168 ( .A1(\SB4_23/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_23/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_23/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_23/Component_Function_5/NAND4_in[0] ), .ZN(n1313) );
  NAND3_X1 U3169 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i0_4 ), .A3(
        \SB1_0_26/i1[9] ), .ZN(n1336) );
  XNOR2_X1 U3170 ( .A(\MC_ARK_ARC_1_1/temp1[189] ), .B(
        \MC_ARK_ARC_1_1/temp4[189] ), .ZN(n1314) );
  NAND3_X1 U3171 ( .A1(\SB1_1_25/i1_7 ), .A2(\SB1_1_25/i0[10] ), .A3(
        \SB1_1_25/i1[9] ), .ZN(\SB1_1_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3172 ( .A1(\SB2_1_23/i3[0] ), .A2(\SB2_1_23/i1_5 ), .A3(
        \SB2_1_23/i0[8] ), .ZN(\SB2_1_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3173 ( .A1(\SB4_12/i0_3 ), .A2(\SB4_12/i0_0 ), .A3(\SB4_12/i0_4 ), 
        .ZN(\SB4_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3174 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i0_0 ), .A3(
        \SB1_1_1/i0_4 ), .ZN(\SB1_1_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3175 ( .A1(\SB2_1_31/i0[8] ), .A2(\SB2_1_31/i1_5 ), .A3(
        \SB2_1_31/i3[0] ), .ZN(\SB2_1_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3176 ( .A1(\SB2_1_7/i0[8] ), .A2(\SB2_1_7/i1_5 ), .A3(
        \SB2_1_7/i3[0] ), .ZN(\SB2_1_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3177 ( .A1(\SB4_6/i0_4 ), .A2(\SB4_6/i1_7 ), .A3(\SB4_6/i0[8] ), 
        .ZN(\SB4_6/Component_Function_1/NAND4_in[3] ) );
  XNOR2_X1 U3178 ( .A(\MC_ARK_ARC_1_3/temp2[59] ), .B(
        \MC_ARK_ARC_1_3/temp3[59] ), .ZN(n1315) );
  OR3_X1 U3181 ( .A1(\RI1[3][156] ), .A2(\RI1[3][157] ), .A3(\RI1[3][160] ), 
        .ZN(\SB1_3_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3182 ( .A1(\SB1_1_31/i0_3 ), .A2(\SB1_1_31/i0_0 ), .A3(
        \SB1_1_31/i0_4 ), .ZN(\SB1_1_31/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U3183 ( .A1(\SB1_1_9/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_9/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_1_9/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[1][137] ) );
  NAND4_X1 U3184 ( .A1(\SB3_9/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_9/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_5/NAND4_in[0] ), .A4(n1316), .ZN(
        \RI3[4][137] ) );
  NAND3_X1 U3185 ( .A1(\SB3_9/i0_3 ), .A2(\SB3_9/i0_4 ), .A3(\SB3_9/i1[9] ), 
        .ZN(n1316) );
  NAND4_X1 U3187 ( .A1(\SB1_0_6/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_6/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_0_6/Component_Function_5/NAND4_in[1] ), .A4(n1318), .ZN(
        \RI3[0][155] ) );
  NAND4_X1 U3188 ( .A1(\SB4_13/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_13/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_13/Component_Function_0/NAND4_in[0] ), .A4(n1319), .ZN(n1441) );
  NAND3_X1 U3189 ( .A1(\SB4_13/i0[6] ), .A2(\SB4_13/i0[8] ), .A3(
        \SB4_13/i0[7] ), .ZN(n1319) );
  NAND3_X1 U3190 ( .A1(n1638), .A2(\SB4_8/i1_7 ), .A3(\SB4_8/i0[8] ), .ZN(
        n1320) );
  NAND3_X1 U3191 ( .A1(\SB3_9/i0_3 ), .A2(\SB3_9/i0[9] ), .A3(\SB3_9/i0[10] ), 
        .ZN(\SB3_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3192 ( .A1(\SB2_1_21/i0_4 ), .A2(\RI3[1][60] ), .A3(
        \SB2_1_21/i0[6] ), .ZN(\SB2_1_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3193 ( .A1(\SB4_8/i0_3 ), .A2(\SB4_8/i0_0 ), .A3(n1638), .ZN(
        \SB4_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3194 ( .A1(n1672), .A2(\SB4_0/i0_0 ), .A3(\SB4_0/i0_4 ), .ZN(
        \SB4_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3197 ( .A1(\SB4_10/i0_4 ), .A2(\SB4_10/i1_7 ), .A3(\SB4_10/i0[8] ), 
        .ZN(n1323) );
  NAND3_X1 U3198 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0_0 ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3200 ( .A1(\SB3_13/i0[9] ), .A2(\SB3_13/i0_3 ), .A3(
        \SB3_13/i0[10] ), .ZN(\SB3_13/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U3203 ( .A(n1325), .B(n309), .ZN(Ciphertext[176]) );
  NAND4_X1 U3204 ( .A1(\SB4_2/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB4_2/Component_Function_2/NAND4_in[3] ), .A4(
        \SB4_2/Component_Function_2/NAND4_in[0] ), .ZN(n1325) );
  NAND3_X1 U3205 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0_0 ), .A3(
        \SB1_1_9/i0_4 ), .ZN(\SB1_1_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3206 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i0[9] ), .A3(
        \SB1_1_28/i0[8] ), .ZN(\SB1_1_28/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3207 ( .A(n1326), .B(n322), .ZN(Ciphertext[174]) );
  NAND4_X1 U3208 ( .A1(\SB4_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_2/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_2/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_2/Component_Function_0/NAND4_in[0] ), .ZN(n1326) );
  NAND3_X1 U3209 ( .A1(n841), .A2(\SB4_11/i0_0 ), .A3(n551), .ZN(
        \SB4_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3210 ( .A1(\SB4_26/i0_3 ), .A2(\SB4_26/i0_4 ), .A3(\SB4_26/i0[10] ), .ZN(\SB4_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3211 ( .A1(n1949), .A2(n780), .A3(\SB4_27/i0_0 ), .ZN(
        \SB4_27/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U3212 ( .A1(\SB1_3_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_9/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_9/Component_Function_5/NAND4_in[0] ), .A4(n1327), .ZN(
        \RI3[3][137] ) );
  NAND3_X1 U3213 ( .A1(\SB1_3_9/i0_3 ), .A2(\SB1_3_9/i1[9] ), .A3(
        \SB1_3_9/i0_4 ), .ZN(n1327) );
  NAND4_X1 U3215 ( .A1(\SB4_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_16/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_16/Component_Function_0/NAND4_in[0] ), .A4(n1328), .ZN(n1414) );
  NAND3_X1 U3216 ( .A1(\SB4_16/i0[6] ), .A2(\SB4_16/i0[8] ), .A3(
        \SB4_16/i0[7] ), .ZN(n1328) );
  NAND3_X1 U3217 ( .A1(\SB4_1/i0_4 ), .A2(\SB4_1/i1_7 ), .A3(\SB4_1/i0[8] ), 
        .ZN(n1329) );
  NAND3_X1 U3219 ( .A1(n1671), .A2(\SB4_26/i0_4 ), .A3(\SB4_26/i1[9] ), .ZN(
        \SB4_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3220 ( .A1(\SB2_0_14/i0_3 ), .A2(\SB2_0_14/i0[9] ), .A3(
        \SB2_0_14/i0[10] ), .ZN(\SB2_0_14/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3221 ( .A1(\SB3_22/i0_3 ), .A2(\SB3_22/i0[9] ), .A3(
        \SB3_22/i0[10] ), .ZN(\SB3_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3222 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i0[9] ), .A3(
        \SB1_3_19/i0[8] ), .ZN(\SB1_3_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3225 ( .A1(\SB4_21/i0_4 ), .A2(\SB4_21/i1_7 ), .A3(\SB4_21/i0[8] ), 
        .ZN(n1332) );
  XNOR2_X1 U3226 ( .A(n1333), .B(n269), .ZN(Ciphertext[182]) );
  NAND3_X1 U3229 ( .A1(\SB4_18/i0_4 ), .A2(\SB4_18/i1_5 ), .A3(\SB4_18/i0_0 ), 
        .ZN(n1335) );
  NAND3_X1 U3230 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i0[9] ), .A3(
        \SB1_3_6/i0[8] ), .ZN(\SB1_3_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3231 ( .A1(\SB1_1_4/i1_7 ), .A2(\SB1_1_4/i0_4 ), .A3(
        \SB1_1_4/i0[8] ), .ZN(\SB1_1_4/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U3232 ( .A1(\SB2_2_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_8/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_8/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_8/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[143] ) );
  NAND3_X1 U3235 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i1[9] ), .A3(
        \SB1_0_28/i0_4 ), .ZN(\SB1_0_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3236 ( .A1(\SB1_2_7/i0_3 ), .A2(\SB1_2_7/i0[9] ), .A3(
        \SB1_2_7/i0[8] ), .ZN(\SB1_2_7/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U3237 ( .A(\RI1[1][173] ), .ZN(\SB1_1_3/i0_3 ) );
  NAND3_X1 U3239 ( .A1(\SB4_23/i0_4 ), .A2(n848), .A3(\SB4_23/i1[9] ), .ZN(
        \SB4_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3240 ( .A1(\SB4_2/i0_4 ), .A2(\SB4_2/i0_3 ), .A3(\SB4_2/i1[9] ), 
        .ZN(\SB4_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3241 ( .A1(\SB4_28/i0_4 ), .A2(n866), .A3(\SB4_28/i0[10] ), .ZN(
        \SB4_28/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U3244 ( .A1(\SB1_0_26/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_26/Component_Function_5/NAND4_in[3] ), .A4(n1336), .ZN(
        \RI3[0][35] ) );
  NAND3_X1 U3245 ( .A1(\SB1_2_20/i0_3 ), .A2(\SB1_2_20/i0[9] ), .A3(
        \SB1_2_20/i0[8] ), .ZN(\SB1_2_20/Component_Function_2/NAND4_in[2] ) );
  OR3_X1 U3246 ( .A1(\RI1[3][90] ), .A2(\RI1[3][91] ), .A3(\RI1[3][94] ), .ZN(
        \SB1_3_16/Component_Function_5/NAND4_in[3] ) );
  XNOR2_X1 U3247 ( .A(\MC_ARK_ARC_1_3/temp5[29] ), .B(
        \MC_ARK_ARC_1_3/temp6[29] ), .ZN(\RI1[4][29] ) );
  INV_X2 U3248 ( .A(\RI1[3][47] ), .ZN(\SB1_3_24/i0_3 ) );
  XNOR2_X1 U3249 ( .A(\MC_ARK_ARC_1_2/temp5[47] ), .B(
        \MC_ARK_ARC_1_2/temp6[47] ), .ZN(\RI1[3][47] ) );
  XNOR2_X1 U3252 ( .A(n1338), .B(n362), .ZN(Ciphertext[168]) );
  XNOR2_X1 U3253 ( .A(n1339), .B(n310), .ZN(Ciphertext[25]) );
  NAND3_X1 U3254 ( .A1(\SB3_7/i0_0 ), .A2(\SB3_7/i0[7] ), .A3(\SB3_7/i0_3 ), 
        .ZN(n1340) );
  NAND3_X1 U3255 ( .A1(\SB4_21/i0_3 ), .A2(\SB4_21/i0[10] ), .A3(\SB4_21/i0_4 ), .ZN(\SB4_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3256 ( .A1(\SB4_10/i0_3 ), .A2(\SB4_10/i0[10] ), .A3(\SB4_10/i0_4 ), .ZN(\SB4_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3257 ( .A1(\SB1_0_12/i1[9] ), .A2(\SB1_0_12/i0[10] ), .A3(n381), 
        .ZN(\SB1_0_12/Component_Function_2/NAND4_in[0] ) );
  XNOR2_X1 U3258 ( .A(n1342), .B(n1341), .ZN(\RI1[4][131] ) );
  XNOR2_X1 U3259 ( .A(\MC_ARK_ARC_1_3/temp2[131] ), .B(
        \MC_ARK_ARC_1_3/temp4[131] ), .ZN(n1341) );
  XNOR2_X1 U3260 ( .A(\MC_ARK_ARC_1_3/temp3[131] ), .B(
        \MC_ARK_ARC_1_3/temp1[131] ), .ZN(n1342) );
  NAND4_X1 U3261 ( .A1(\SB1_1_28/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_1_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_5/NAND4_in[0] ), .A4(n1343), .ZN(
        \RI3[1][23] ) );
  NAND3_X1 U3262 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i1[9] ), .A3(
        \SB1_1_28/i0_4 ), .ZN(n1343) );
  NAND4_X1 U3263 ( .A1(\SB1_3_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_19/Component_Function_5/NAND4_in[0] ), .A4(n1344), .ZN(
        \RI3[3][77] ) );
  NAND3_X1 U3264 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i1[9] ), .A3(
        \SB1_3_19/i0_4 ), .ZN(n1344) );
  NAND3_X1 U3265 ( .A1(\SB1_2_22/i0_3 ), .A2(\SB1_2_22/i0_0 ), .A3(
        \SB1_2_22/i0_4 ), .ZN(\SB1_2_22/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U3266 ( .A(\MC_ARK_ARC_1_0/temp5[131] ), .B(
        \MC_ARK_ARC_1_0/temp6[131] ), .ZN(\RI1[1][131] ) );
  NAND3_X1 U3267 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0_4 ), .A3(
        \SB1_0_11/i1[9] ), .ZN(n1371) );
  NAND3_X1 U3268 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i1[9] ), .A3(n805), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3269 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0[9] ), .A3(
        \SB1_0_16/i0[8] ), .ZN(\SB1_0_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3271 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i0_4 ), .A3(
        \SB2_3_2/i1[9] ), .ZN(n1345) );
  NAND3_X1 U3272 ( .A1(\SB1_2_30/i0_3 ), .A2(\SB1_2_30/i0_0 ), .A3(
        \SB1_2_30/i0_4 ), .ZN(\SB1_2_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3273 ( .A1(\SB1_2_11/i0_3 ), .A2(\SB1_2_11/i0[9] ), .A3(
        \SB1_2_11/i0[8] ), .ZN(\SB1_2_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3274 ( .A1(\SB1_3_27/i0_3 ), .A2(\SB1_3_27/i0[9] ), .A3(
        \SB1_3_27/i0[8] ), .ZN(\SB1_3_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3275 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i0[9] ), .A3(
        \SB1_1_19/i0[8] ), .ZN(\SB1_1_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3276 ( .A1(\SB1_3_4/i0_3 ), .A2(\SB1_3_4/i0[9] ), .A3(
        \SB1_3_4/i0[8] ), .ZN(\SB1_3_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3277 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i0[9] ), .A3(
        \SB1_1_7/i0[8] ), .ZN(\SB1_1_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3281 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i0[9] ), .A3(
        \SB3_27/i0[10] ), .ZN(\SB3_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3283 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i0[9] ), .A3(
        \SB1_0_17/i0[8] ), .ZN(\SB1_0_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3284 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0[9] ), .A3(
        \SB1_0_9/i0[8] ), .ZN(\SB1_0_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3286 ( .A1(\SB4_15/i0_4 ), .A2(n871), .A3(\SB4_15/i0[10] ), .ZN(
        \SB4_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3287 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i0[10] ), .A3(\SB4_17/i0_4 ), .ZN(\SB4_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3288 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i0_4 ), .ZN(\SB1_3_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3290 ( .A1(n863), .A2(\SB4_8/i1[9] ), .A3(n1638), .ZN(
        \SB4_8/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3292 ( .A(\MC_ARK_ARC_1_3/temp2[77] ), .B(
        \MC_ARK_ARC_1_3/temp4[77] ), .ZN(n1349) );
  XNOR2_X1 U3293 ( .A(\MC_ARK_ARC_1_3/temp1[77] ), .B(
        \MC_ARK_ARC_1_3/temp3[77] ), .ZN(n1350) );
  NAND3_X1 U3294 ( .A1(\SB1_0_16/i0_4 ), .A2(\SB1_0_16/i1_5 ), .A3(
        \SB1_0_16/i0_0 ), .ZN(\SB1_0_16/Component_Function_2/NAND4_in[3] ) );
  XNOR2_X1 U3295 ( .A(n1351), .B(n243), .ZN(Ciphertext[186]) );
  NAND4_X1 U3296 ( .A1(\SB4_0/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_0/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_0/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_0/Component_Function_0/NAND4_in[1] ), .ZN(n1351) );
  NAND4_X1 U3297 ( .A1(\SB3_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_26/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_26/Component_Function_0/NAND4_in[1] ), .A4(n1352), .ZN(
        \RI3[4][60] ) );
  NAND3_X1 U3300 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0[9] ), .A3(
        \SB1_2_13/i0[8] ), .ZN(\SB1_2_13/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3301 ( .A1(\SB1_1_11/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_11/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_11/Component_Function_5/NAND4_in[0] ), .A4(n1353), .ZN(
        \RI3[1][125] ) );
  NAND3_X1 U3302 ( .A1(\SB1_1_11/i0_3 ), .A2(\SB1_1_11/i1[9] ), .A3(
        \SB1_1_11/i0_4 ), .ZN(n1353) );
  NAND3_X1 U3304 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0_0 ), .A3(
        \SB1_2_13/i0_4 ), .ZN(\SB1_2_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3305 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0_0 ), .A3(
        \SB1_0_29/i0_4 ), .ZN(\SB1_0_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3306 ( .A1(\SB1_0_30/i0_0 ), .A2(\SB1_0_30/i1_5 ), .A3(
        \SB1_0_30/i0_4 ), .ZN(\SB1_0_30/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U3307 ( .A1(\SB1_0_13/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_13/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_0_13/Component_Function_2/NAND4_in[1] ), .A4(n1354), .ZN(
        \RI3[0][128] ) );
  NAND3_X1 U3308 ( .A1(\SB1_0_13/i0_0 ), .A2(\SB1_0_13/i1_5 ), .A3(
        \SB1_0_13/i0_4 ), .ZN(n1354) );
  NAND3_X1 U3309 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0[9] ), .A3(
        \SB1_0_10/i0[8] ), .ZN(\SB1_0_10/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3310 ( .A(\MC_ARK_ARC_1_0/temp2[95] ), .B(
        \MC_ARK_ARC_1_0/temp4[95] ), .ZN(n1355) );
  XNOR2_X1 U3311 ( .A(\MC_ARK_ARC_1_0/temp3[95] ), .B(
        \MC_ARK_ARC_1_0/temp1[95] ), .ZN(n1356) );
  NAND3_X1 U3312 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0[9] ), .A3(
        \SB1_0_0/i0[8] ), .ZN(\SB1_0_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3313 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0[9] ), .A3(
        \SB1_0_29/i0[8] ), .ZN(\SB1_0_29/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3314 ( .A1(\SB1_0_2/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_5/NAND4_in[3] ), .A4(n1357), .ZN(
        \RI3[0][179] ) );
  NAND3_X1 U3315 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0_4 ), .A3(
        \SB1_0_2/i1[9] ), .ZN(n1357) );
  NAND3_X1 U3317 ( .A1(\SB2_0_28/i0_4 ), .A2(\SB2_0_28/i0_3 ), .A3(
        \SB2_0_28/i1[9] ), .ZN(n1358) );
  NAND4_X1 U3318 ( .A1(\SB1_3_0/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_3_0/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_5/NAND4_in[0] ), .A4(n1359), .ZN(
        \RI3[3][191] ) );
  NAND3_X1 U3319 ( .A1(n809), .A2(\SB1_3_0/i1[9] ), .A3(\SB1_3_0/i0_4 ), .ZN(
        n1359) );
  NAND4_X1 U3322 ( .A1(\SB1_2_21/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_21/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_21/Component_Function_5/NAND4_in[0] ), .A4(n1361), .ZN(
        \RI3[2][65] ) );
  NAND3_X1 U3323 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i1[9] ), .A3(
        \SB1_2_21/i0_4 ), .ZN(n1361) );
  NAND3_X1 U3327 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i1_5 ), .A3(\SB4_22/i0_4 ), 
        .ZN(n1363) );
  XNOR2_X1 U3328 ( .A(n1365), .B(n1364), .ZN(\RI1[3][161] ) );
  XNOR2_X1 U3329 ( .A(\MC_ARK_ARC_1_2/temp1[161] ), .B(
        \MC_ARK_ARC_1_2/temp4[161] ), .ZN(n1364) );
  XNOR2_X1 U3330 ( .A(\MC_ARK_ARC_1_2/temp3[161] ), .B(
        \MC_ARK_ARC_1_2/temp2[161] ), .ZN(n1365) );
  NAND4_X1 U3331 ( .A1(\SB1_1_22/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_22/Component_Function_5/NAND4_in[0] ), .A4(n1366), .ZN(
        \RI3[1][59] ) );
  NAND3_X1 U3332 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0[9] ), .A3(
        \SB1_3_8/i0[8] ), .ZN(\SB1_3_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3333 ( .A1(\SB1_2_1/i0_3 ), .A2(\SB1_2_1/i0[9] ), .A3(
        \SB1_2_1/i0[8] ), .ZN(\SB1_2_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3335 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0_4 ), .A3(
        \SB1_1_30/i1[9] ), .ZN(\SB1_1_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3337 ( .A1(\SB1_0_1/i0_3 ), .A2(\SB1_0_1/i0_0 ), .A3(
        \SB1_0_1/i0_4 ), .ZN(\SB1_0_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3340 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i0_0 ), .A3(\SB4_16/i0[7] ), 
        .ZN(\SB4_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3341 ( .A1(\SB2_0_30/i0_3 ), .A2(\RI3[0][6] ), .A3(
        \SB2_0_30/i0[8] ), .ZN(\SB2_0_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3342 ( .A1(\SB1_0_30/i0_3 ), .A2(\SB1_0_30/i1[9] ), .A3(
        \SB1_0_30/i0_4 ), .ZN(\SB1_0_30/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U3343 ( .A(\RI1[2][83] ), .ZN(\SB1_2_18/i0_3 ) );
  NAND3_X1 U3344 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0[9] ), .A3(
        \SB1_0_7/i0[8] ), .ZN(\SB1_0_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3345 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0[9] ), .A3(
        \SB1_0_2/i0[8] ), .ZN(\SB1_0_2/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U3346 ( .A(\RI1[1][191] ), .ZN(\SB1_1_0/i0_3 ) );
  NAND3_X1 U3348 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i0_4 ), .A3(\SB4_16/i1[9] ), 
        .ZN(\SB4_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3349 ( .A1(n1949), .A2(\SB4_27/i1[9] ), .A3(n780), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3350 ( .A(n1370), .B(\MC_ARK_ARC_1_1/temp6[125] ), .ZN(
        \RI1[2][125] ) );
  XNOR2_X1 U3351 ( .A(\MC_ARK_ARC_1_1/temp1[125] ), .B(
        \MC_ARK_ARC_1_1/temp2[125] ), .ZN(n1370) );
  NAND3_X1 U3352 ( .A1(\SB1_0_4/i0_3 ), .A2(\SB1_0_4/i0_0 ), .A3(
        \SB1_0_4/i0_4 ), .ZN(\SB1_0_4/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U3353 ( .A1(\SB1_0_11/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_11/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_0_11/Component_Function_5/NAND4_in[0] ), .A4(n1371), .ZN(
        \RI3[0][125] ) );
  NAND3_X1 U3356 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i0[9] ), .A3(
        \SB1_3_1/i0[8] ), .ZN(\SB1_3_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3359 ( .A1(\SB2_2_22/i0_4 ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i1[9] ), .ZN(\SB2_2_22/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3362 ( .A1(\SB4_4/i0_3 ), .A2(\SB4_4/i0_4 ), .A3(\SB4_4/i0[10] ), 
        .ZN(\SB4_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3363 ( .A1(n1664), .A2(\SB1_0_8/i0[9] ), .A3(\SB1_0_8/i0[8] ), 
        .ZN(\SB1_0_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3364 ( .A1(n1657), .A2(\SB1_2_9/i0[9] ), .A3(\SB1_2_9/i0[8] ), 
        .ZN(\SB1_2_9/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3365 ( .A(n1375), .B(n1376), .ZN(\RI1[3][17] ) );
  XNOR2_X1 U3366 ( .A(\MC_ARK_ARC_1_2/temp1[17] ), .B(
        \MC_ARK_ARC_1_2/temp4[17] ), .ZN(n1375) );
  XNOR2_X1 U3367 ( .A(\MC_ARK_ARC_1_2/temp3[17] ), .B(
        \MC_ARK_ARC_1_2/temp2[17] ), .ZN(n1376) );
  NAND3_X1 U3368 ( .A1(\SB2_0_4/i0_4 ), .A2(\SB2_0_4/i1_7 ), .A3(
        \SB2_0_4/i0[8] ), .ZN(\SB2_0_4/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 U3369 ( .A1(\SB1_1_4/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_4/Component_Function_5/NAND4_in[0] ), .A4(n1377), .ZN(
        \RI3[1][167] ) );
  NAND3_X1 U3370 ( .A1(\SB1_1_4/i0_3 ), .A2(\SB1_1_4/i1[9] ), .A3(
        \SB1_1_4/i0_4 ), .ZN(n1377) );
  NAND4_X1 U3371 ( .A1(\SB1_2_29/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_2_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_5/NAND4_in[0] ), .A4(n1378), .ZN(
        \RI3[2][17] ) );
  NAND3_X1 U3372 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0_0 ), .A3(
        \SB1_0_6/i0_4 ), .ZN(\SB1_0_6/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U3375 ( .A1(\SB3_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_0/NAND4_in[0] ), .A4(n1380), .ZN(
        \RI3[4][126] ) );
  NAND3_X1 U3376 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i0[7] ), .A3(\SB3_15/i0_3 ), 
        .ZN(n1380) );
  NAND3_X1 U3378 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0[9] ), .A3(
        \SB2_2_30/i0[10] ), .ZN(\SB2_2_30/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3379 ( .A1(n1949), .A2(n780), .A3(\SB4_27/i0[10] ), .ZN(
        \SB4_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3380 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i1[9] ), .A3(
        \SB1_0_13/i0_4 ), .ZN(\SB1_0_13/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3382 ( .A(n1382), .B(n224), .ZN(Ciphertext[134]) );
  NAND4_X1 U3383 ( .A1(\SB4_9/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_9/Component_Function_2/NAND4_in[1] ), .A3(
        \SB4_9/Component_Function_2/NAND4_in[3] ), .A4(
        \SB4_9/Component_Function_2/NAND4_in[0] ), .ZN(n1382) );
  NAND3_X1 U3384 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0[9] ), .A3(
        \SB1_0_28/i0[8] ), .ZN(\SB1_0_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3385 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0[9] ), .A3(
        \SB1_0_15/i0[8] ), .ZN(\SB1_0_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3386 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[9] ), .A3(
        \SB1_1_22/i0[8] ), .ZN(\SB1_1_22/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3388 ( .A1(\SB1_1_0/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_0/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_0/Component_Function_5/NAND4_in[0] ), .A4(n1383), .ZN(
        \RI3[1][191] ) );
  NAND3_X1 U3389 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i1[9] ), .A3(
        \SB1_1_0/i0_4 ), .ZN(n1383) );
  NAND3_X1 U3390 ( .A1(\SB1_3_2/i0_3 ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i0_4 ), .ZN(\SB1_3_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3391 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i1[9] ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3392 ( .A1(\SB4_25/i0_3 ), .A2(n821), .A3(\SB4_25/i0_0 ), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3393 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i0_0 ), .A3(\SB4_25/i0_4 ), 
        .ZN(\SB4_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3395 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0_0 ), .A3(n844), .ZN(
        \SB4_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3398 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i0_4 ), .A3(\SB3_13/i1[9] ), 
        .ZN(\SB3_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3399 ( .A1(\SB1_3_9/i0_3 ), .A2(\SB1_3_9/i0[9] ), .A3(
        \SB1_3_9/i0[8] ), .ZN(\SB1_3_9/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3400 ( .A1(\SB1_0_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_0_1/Component_Function_2/NAND4_in[1] ), .A4(n1385), .ZN(
        \RI3[0][8] ) );
  NAND3_X1 U3401 ( .A1(\SB1_0_1/i0_0 ), .A2(\SB1_0_1/i1_5 ), .A3(
        \SB1_0_1/i0_4 ), .ZN(n1385) );
  NAND3_X1 U3403 ( .A1(\SB2_0_8/i0_4 ), .A2(\SB2_0_8/i0_3 ), .A3(
        \SB2_0_8/i1[9] ), .ZN(n1386) );
  NAND4_X1 U3407 ( .A1(\SB1_3_27/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_3_27/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_27/Component_Function_5/NAND4_in[0] ), .A4(n1389), .ZN(
        \RI3[3][29] ) );
  NAND3_X1 U3408 ( .A1(\SB1_3_27/i0_3 ), .A2(\SB1_3_27/i1[9] ), .A3(
        \SB1_3_27/i0_4 ), .ZN(n1389) );
  NAND4_X1 U3409 ( .A1(\SB1_1_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_8/Component_Function_5/NAND4_in[0] ), .A4(n1390), .ZN(
        \RI3[1][143] ) );
  NAND3_X1 U3410 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i1[9] ), .A3(
        \SB1_1_8/i0_4 ), .ZN(n1390) );
  NAND3_X1 U3411 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i0_0 ), .A3(
        \SB1_2_5/i0_4 ), .ZN(\SB1_2_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3412 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0_0 ), .A3(
        \SB1_0_5/i0_4 ), .ZN(\SB1_0_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3413 ( .A1(\SB2_2_3/i0[8] ), .A2(\SB2_2_3/i1_5 ), .A3(
        \SB2_2_3/i3[0] ), .ZN(\SB2_2_3/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U3414 ( .A1(\SB3_18/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_18/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_18/Component_Function_0/NAND4_in[1] ), .A4(n1391), .ZN(
        \RI3[4][108] ) );
  NAND3_X1 U3415 ( .A1(\SB3_18/i0_0 ), .A2(\SB3_18/i0[7] ), .A3(\SB3_18/i0_3 ), 
        .ZN(n1391) );
  XNOR2_X1 U3416 ( .A(n1392), .B(n320), .ZN(Ciphertext[92]) );
  NAND3_X1 U3418 ( .A1(\SB4_20/i0_3 ), .A2(n844), .A3(\SB4_20/i1[9] ), .ZN(
        \SB4_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3419 ( .A1(\SB4_12/i0_3 ), .A2(\SB4_12/i0_4 ), .A3(\SB4_12/i0[10] ), .ZN(\SB4_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3420 ( .A1(\SB4_22/i0_3 ), .A2(n779), .A3(\SB4_22/i0[10] ), .ZN(
        \SB4_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3421 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i1[9] ), .A3(
        \SB1_0_17/i0_4 ), .ZN(\SB1_0_17/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3422 ( .A(n1393), .B(n200), .ZN(Ciphertext[110]) );
  NAND3_X1 U3424 ( .A1(\SB1_0_3/i0_3 ), .A2(\SB1_0_3/i0[9] ), .A3(
        \SB1_0_3/i0[8] ), .ZN(\SB1_0_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3425 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[9] ), .A3(
        \SB1_3_21/i0[8] ), .ZN(\SB1_3_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3426 ( .A1(\SB2_0_31/i0_3 ), .A2(\SB2_0_31/i0[9] ), .A3(
        \SB2_0_31/i0[8] ), .ZN(\SB2_0_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3428 ( .A1(\SB4_29/i0_3 ), .A2(n2131), .A3(\SB4_29/i0[10] ), .ZN(
        \SB4_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3429 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i0[10] ), .A3(n799), .ZN(
        \SB4_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3430 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0[9] ), .A3(
        \SB1_0_20/i0[8] ), .ZN(\SB1_0_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3431 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[9] ), .A3(
        \SB1_0_25/i0[8] ), .ZN(\SB1_0_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3433 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i0[9] ), .A3(
        \SB1_2_3/i0[8] ), .ZN(\SB1_2_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3435 ( .A1(\SB1_0_23/i0_0 ), .A2(\SB1_0_23/i1_5 ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3440 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i0[9] ), .A3(
        \SB1_2_18/i0[8] ), .ZN(\SB1_2_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3441 ( .A1(\SB2_0_13/i0_4 ), .A2(\SB2_0_13/i0_3 ), .A3(
        \SB2_0_13/i1[9] ), .ZN(n1397) );
  XNOR2_X1 U3442 ( .A(n1398), .B(n203), .ZN(Ciphertext[41]) );
  NAND4_X1 U3443 ( .A1(\SB4_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_25/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_25/Component_Function_5/NAND4_in[0] ), .ZN(n1398) );
  INV_X2 U3444 ( .A(\RI1[2][125] ), .ZN(\SB1_2_11/i0_3 ) );
  XNOR2_X1 U3448 ( .A(n1401), .B(n311), .ZN(Ciphertext[66]) );
  NAND3_X1 U3449 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i0[10] ), .A3(\SB4_22/i0_4 ), .ZN(\SB4_22/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U3453 ( .A1(\SB1_1_27/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_27/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_27/Component_Function_5/NAND4_in[0] ), .A4(n1404), .ZN(
        \RI3[1][29] ) );
  NAND3_X1 U3454 ( .A1(\SB1_1_27/i0_3 ), .A2(\SB1_1_27/i1[9] ), .A3(
        \SB1_1_27/i0_4 ), .ZN(n1404) );
  NAND4_X1 U3457 ( .A1(\SB3_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_0/NAND4_in[0] ), .A4(n1406), .ZN(
        \RI3[4][156] ) );
  NAND3_X1 U3458 ( .A1(\SB3_10/i0_0 ), .A2(\SB3_10/i0[7] ), .A3(\SB3_10/i0_3 ), 
        .ZN(n1406) );
  XNOR2_X1 U3459 ( .A(n1407), .B(n315), .ZN(Ciphertext[38]) );
  NAND4_X1 U3460 ( .A1(\SB4_25/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB4_25/Component_Function_2/NAND4_in[3] ), .A4(
        \SB4_25/Component_Function_2/NAND4_in[0] ), .ZN(n1407) );
  NAND3_X1 U3461 ( .A1(\SB3_30/i0[7] ), .A2(\SB3_30/i0_0 ), .A3(\SB3_30/i0_3 ), 
        .ZN(\SB3_30/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U3462 ( .A1(\SB3_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_0/NAND4_in[0] ), .A4(n1408), .ZN(
        \RI3[4][72] ) );
  NAND3_X1 U3463 ( .A1(\SB3_24/i0[7] ), .A2(\SB3_24/i0_0 ), .A3(\SB3_24/i0_3 ), 
        .ZN(n1408) );
  NAND3_X1 U3464 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i0[9] ), .A3(
        \SB1_0_19/i0[8] ), .ZN(\SB1_0_19/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3468 ( .A1(\SB1_2_0/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_0/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_0/Component_Function_5/NAND4_in[0] ), .A4(n1411), .ZN(
        \RI3[2][191] ) );
  NAND3_X1 U3469 ( .A1(\SB1_2_0/i0_3 ), .A2(\SB1_2_0/i1[9] ), .A3(
        \SB1_2_0/i0_4 ), .ZN(n1411) );
  NAND3_X1 U3472 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i1[9] ), .A3(
        \SB1_3_6/i0_4 ), .ZN(\SB1_3_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3473 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i1[9] ), .A3(
        \SB1_3_18/i0_4 ), .ZN(\SB1_3_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3476 ( .A1(\SB1_1_27/i0_3 ), .A2(\SB1_1_27/i0[9] ), .A3(
        \SB1_1_27/i0[8] ), .ZN(\SB1_1_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3477 ( .A1(\SB2_0_16/i0_4 ), .A2(\SB2_0_16/i0_3 ), .A3(
        \SB2_0_16/i1[9] ), .ZN(\SB2_0_16/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3478 ( .A(n1414), .B(n334), .ZN(Ciphertext[90]) );
  NAND3_X1 U3481 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0[9] ), .A3(
        \SB1_0_20/i0[10] ), .ZN(\SB1_0_20/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3482 ( .A1(\SB1_0_16/i0[10] ), .A2(\SB1_0_16/i1[9] ), .A3(
        \SB1_0_16/i1_7 ), .ZN(\SB1_0_16/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U3483 ( .A1(\SB3_29/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_0/NAND4_in[0] ), .A4(n1416), .ZN(
        \RI3[4][42] ) );
  NAND3_X1 U3484 ( .A1(\SB3_29/i0[7] ), .A2(\SB3_29/i0_0 ), .A3(\SB3_29/i0_3 ), 
        .ZN(n1416) );
  XNOR2_X1 U3485 ( .A(n1417), .B(n275), .ZN(Ciphertext[44]) );
  NAND3_X1 U3487 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0[9] ), .A3(
        \SB1_1_15/i0[8] ), .ZN(\SB1_1_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3489 ( .A1(\SB2_0_9/i0_4 ), .A2(\SB2_0_9/i0_3 ), .A3(
        \SB2_0_9/i1[9] ), .ZN(n1418) );
  NAND4_X1 U3491 ( .A1(\SB1_3_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_12/Component_Function_5/NAND4_in[0] ), .A4(n1419), .ZN(
        \RI3[3][119] ) );
  NAND3_X1 U3492 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i1[9] ), .A3(
        \SB1_3_12/i0_4 ), .ZN(n1419) );
  NAND3_X1 U3493 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0[9] ), .A3(
        \SB1_0_18/i0[8] ), .ZN(\SB1_0_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3495 ( .A1(\SB2_1_21/i0_3 ), .A2(\SB2_1_21/i0_4 ), .A3(
        \SB2_1_21/i1[9] ), .ZN(\SB2_1_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3496 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i1[9] ), .A3(
        \SB1_1_21/i0_4 ), .ZN(\SB1_1_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3501 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i0[9] ), .A3(
        \SB1_3_12/i0[8] ), .ZN(\SB1_3_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3502 ( .A1(\SB1_3_7/i0_3 ), .A2(\SB1_3_7/i0[9] ), .A3(
        \SB1_3_7/i0[8] ), .ZN(\SB1_3_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3503 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i0[9] ), .A3(
        \SB1_3_13/i0[8] ), .ZN(\SB1_3_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3504 ( .A1(\SB2_0_4/i0_4 ), .A2(\SB2_0_4/i0_3 ), .A3(
        \SB2_0_4/i1[9] ), .ZN(\SB2_0_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3506 ( .A1(\SB2_0_13/i0_3 ), .A2(\SB2_0_13/i0[9] ), .A3(
        \SB2_0_13/i0[8] ), .ZN(\SB2_0_13/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3507 ( .A(\MC_ARK_ARC_1_0/temp5[177] ), .B(n1423), .ZN(
        \RI1[1][177] ) );
  XNOR2_X1 U3508 ( .A(\MC_ARK_ARC_1_0/temp3[177] ), .B(
        \MC_ARK_ARC_1_0/temp4[177] ), .ZN(n1423) );
  NAND3_X1 U3509 ( .A1(n851), .A2(\SB4_22/i0_4 ), .A3(\SB4_22/i0_0 ), .ZN(
        \SB4_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3510 ( .A1(\SB1_0_0/i1_7 ), .A2(\SB1_0_0/i0[10] ), .A3(
        \SB1_0_0/i1[9] ), .ZN(\SB1_0_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3511 ( .A1(\SB1_0_3/i0_3 ), .A2(\SB1_0_3/i0_0 ), .A3(
        \SB1_0_3/i0_4 ), .ZN(\SB1_0_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3512 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i0_0 ), .A3(
        \SB1_3_13/i0_4 ), .ZN(\SB1_3_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3513 ( .A1(\SB2_0_30/i0[8] ), .A2(\SB2_0_30/i1_5 ), .A3(
        \SB2_0_30/i3[0] ), .ZN(\SB2_0_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3514 ( .A1(\SB3_22/i1_7 ), .A2(\SB3_22/i0[8] ), .A3(\SB3_22/i0_3 ), 
        .ZN(\SB3_22/Component_Function_1/NAND4_in[1] ) );
  NAND4_X1 U3515 ( .A1(\SB3_17/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_17/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_17/Component_Function_0/NAND4_in[1] ), .A4(n1424), .ZN(
        \RI3[4][114] ) );
  NAND3_X1 U3516 ( .A1(\SB3_17/i0_0 ), .A2(\SB3_17/i0[7] ), .A3(n867), .ZN(
        n1424) );
  XNOR2_X1 U3518 ( .A(n1426), .B(n226), .ZN(Ciphertext[24]) );
  NAND4_X1 U3519 ( .A1(\SB4_27/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_27/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_27/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_27/Component_Function_0/NAND4_in[0] ), .ZN(n1426) );
  NAND3_X1 U3522 ( .A1(\SB1_0_15/i0[10] ), .A2(\SB1_0_15/i1[9] ), .A3(
        \SB1_0_15/i1_7 ), .ZN(\SB1_0_15/Component_Function_3/NAND4_in[2] ) );
  XNOR2_X1 U3523 ( .A(n1428), .B(n267), .ZN(Ciphertext[100]) );
  NAND4_X1 U3524 ( .A1(\SB4_15/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_15/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_15/Component_Function_4/NAND4_in[1] ), .ZN(n1428) );
  XNOR2_X1 U3525 ( .A(n1429), .B(n319), .ZN(Ciphertext[10]) );
  NAND4_X1 U3526 ( .A1(\SB4_30/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_30/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_30/Component_Function_4/NAND4_in[1] ), .ZN(n1429) );
  NAND4_X1 U3529 ( .A1(\SB1_1_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_12/Component_Function_5/NAND4_in[0] ), .A4(n1431), .ZN(
        \RI3[1][119] ) );
  NAND3_X1 U3530 ( .A1(\SB1_1_12/i0_3 ), .A2(\SB1_1_12/i1[9] ), .A3(
        \SB1_1_12/i0_4 ), .ZN(n1431) );
  NAND4_X1 U3531 ( .A1(\SB1_3_29/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_29/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_29/Component_Function_5/NAND4_in[0] ), .A4(n1432), .ZN(
        \RI3[3][17] ) );
  NAND3_X1 U3532 ( .A1(\SB1_3_29/i0_3 ), .A2(\SB1_3_29/i1[9] ), .A3(
        \SB1_3_29/i0_4 ), .ZN(n1432) );
  XNOR2_X1 U3535 ( .A(n1434), .B(n356), .ZN(Ciphertext[114]) );
  NAND4_X1 U3536 ( .A1(\SB4_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_12/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_12/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_12/Component_Function_0/NAND4_in[0] ), .ZN(n1434) );
  NAND3_X1 U3537 ( .A1(\SB2_3_13/i0_3 ), .A2(n2107), .A3(\SB2_3_13/i0[10] ), 
        .ZN(\SB2_3_13/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U3538 ( .A(n1435), .B(n261), .ZN(Ciphertext[46]) );
  NAND4_X1 U3539 ( .A1(\SB4_24/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_24/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_24/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_24/Component_Function_4/NAND4_in[1] ), .ZN(n1435) );
  XNOR2_X1 U3540 ( .A(n1436), .B(n233), .ZN(Ciphertext[119]) );
  NAND4_X1 U3541 ( .A1(\SB4_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_12/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_12/Component_Function_5/NAND4_in[0] ), .ZN(n1436) );
  XNOR2_X1 U3542 ( .A(n1437), .B(n336), .ZN(Ciphertext[172]) );
  NAND4_X1 U3543 ( .A1(\SB4_3/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_3/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_3/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_3/Component_Function_4/NAND4_in[1] ), .ZN(n1437) );
  NAND3_X1 U3544 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i0_4 ), .A3(
        \SB2_0_20/i1[9] ), .ZN(n1438) );
  NAND4_X1 U3547 ( .A1(\SB1_0_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_20/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_0_20/Component_Function_5/NAND4_in[0] ), .A4(n1440), .ZN(
        \RI3[0][71] ) );
  NAND3_X1 U3548 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i1[9] ), .A3(
        \SB1_0_20/i0_4 ), .ZN(n1440) );
  NAND3_X1 U3549 ( .A1(\SB2_0_31/i0[8] ), .A2(\SB2_0_31/i1_5 ), .A3(
        \SB2_0_31/i3[0] ), .ZN(\SB2_0_31/Component_Function_3/NAND4_in[3] ) );
  XNOR2_X1 U3550 ( .A(n1441), .B(n214), .ZN(Ciphertext[108]) );
  NAND3_X1 U3551 ( .A1(\SB4_5/i0_3 ), .A2(\SB4_5/i1[9] ), .A3(n834), .ZN(
        \SB4_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3552 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i1[9] ), .A3(
        \SB1_2_5/i0_4 ), .ZN(\SB1_2_5/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3555 ( .A(n1443), .B(n369), .ZN(Ciphertext[112]) );
  NAND4_X1 U3556 ( .A1(\SB4_13/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_13/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_13/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_13/Component_Function_4/NAND4_in[1] ), .ZN(n1443) );
  NAND3_X1 U3557 ( .A1(\SB1_3_28/i0_3 ), .A2(\SB1_3_28/i0[9] ), .A3(
        \SB1_3_28/i0[8] ), .ZN(\SB1_3_28/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U3559 ( .A(\RI1[1][119] ), .ZN(\SB1_1_12/i0_3 ) );
  NAND3_X1 U3560 ( .A1(\SB2_0_26/i0_4 ), .A2(\RI3[0][30] ), .A3(
        \SB2_0_26/i0[6] ), .ZN(n1445) );
  XNOR2_X1 U3561 ( .A(n1446), .B(n220), .ZN(Ciphertext[162]) );
  NAND3_X1 U3562 ( .A1(\SB1_3_14/i0_3 ), .A2(\SB1_3_14/i0[9] ), .A3(
        \SB1_3_14/i0[8] ), .ZN(\SB1_3_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3563 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0[9] ), .A3(
        \SB1_3_26/i0[8] ), .ZN(\SB1_3_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3564 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0[9] ), .A3(
        \SB1_1_6/i0[8] ), .ZN(\SB1_1_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3565 ( .A1(\SB1_3_22/i0_3 ), .A2(\SB1_3_22/i0[9] ), .A3(
        \SB1_3_22/i0[8] ), .ZN(\SB1_3_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3566 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i0[9] ), .A3(
        \SB1_3_17/i0[8] ), .ZN(\SB1_3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3567 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i0[9] ), .A3(
        \SB1_2_14/i0[8] ), .ZN(\SB1_2_14/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3568 ( .A1(\SB1_2_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_20/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_20/Component_Function_5/NAND4_in[0] ), .A4(n1447), .ZN(
        \RI3[2][71] ) );
  NAND3_X1 U3569 ( .A1(\SB1_2_20/i0_3 ), .A2(\SB1_2_20/i1[9] ), .A3(
        \SB1_2_20/i0_4 ), .ZN(n1447) );
  NAND3_X1 U3570 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i1[9] ), .A3(
        \SB1_2_8/i0_4 ), .ZN(\SB1_2_8/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3571 ( .A(n1448), .B(n284), .ZN(Ciphertext[70]) );
  NAND4_X1 U3572 ( .A1(\SB4_20/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_20/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_20/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_20/Component_Function_4/NAND4_in[1] ), .ZN(n1448) );
  XNOR2_X1 U3573 ( .A(n1449), .B(n301), .ZN(Ciphertext[40]) );
  NAND3_X1 U3576 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0[9] ), .A3(
        \SB1_1_0/i0[8] ), .ZN(\SB1_1_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3577 ( .A1(\SB1_3_29/i0_3 ), .A2(\SB1_3_29/i0[9] ), .A3(
        \SB1_3_29/i0[8] ), .ZN(\SB1_3_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3578 ( .A1(\SB1_3_2/i0_3 ), .A2(\SB1_3_2/i0[9] ), .A3(
        \SB1_3_2/i0[8] ), .ZN(\SB1_3_2/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3583 ( .A1(\SB1_2_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_3/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_3/Component_Function_5/NAND4_in[0] ), .A4(n1453), .ZN(
        \RI3[2][173] ) );
  XNOR2_X1 U3584 ( .A(n1454), .B(n248), .ZN(Ciphertext[48]) );
  NAND4_X1 U3585 ( .A1(\SB4_23/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_23/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_23/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_23/Component_Function_0/NAND4_in[0] ), .ZN(n1454) );
  NAND3_X1 U3586 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i0_4 ), .ZN(\SB1_3_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3587 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i0[9] ), .A3(
        \SB2_0_6/i0[10] ), .ZN(\SB2_0_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3588 ( .A1(\SB1_0_28/i0[10] ), .A2(\SB1_0_28/i1[9] ), .A3(
        \SB1_0_28/i1_7 ), .ZN(\SB1_0_28/Component_Function_3/NAND4_in[2] ) );
  XNOR2_X1 U3589 ( .A(n1455), .B(n216), .ZN(Ciphertext[190]) );
  NAND4_X1 U3590 ( .A1(\SB4_0/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_0/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_0/Component_Function_4/NAND4_in[1] ), .ZN(n1455) );
  NAND3_X1 U3593 ( .A1(n809), .A2(\SB1_3_0/i0[9] ), .A3(\SB1_3_0/i0[8] ), .ZN(
        \SB1_3_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3594 ( .A1(n814), .A2(\SB1_2_29/i0[9] ), .A3(\SB1_2_29/i0[8] ), 
        .ZN(\SB1_2_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3595 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0[9] ), .A3(
        \SB1_1_9/i0[8] ), .ZN(\SB1_1_9/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3596 ( .A(n1457), .B(n352), .ZN(Ciphertext[142]) );
  NAND4_X1 U3597 ( .A1(\SB4_8/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_8/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_8/Component_Function_4/NAND4_in[1] ), .ZN(n1457) );
  XNOR2_X1 U3598 ( .A(n1459), .B(n1458), .ZN(\RI1[1][38] ) );
  XNOR2_X1 U3599 ( .A(\MC_ARK_ARC_1_0/temp3[38] ), .B(
        \MC_ARK_ARC_1_0/temp1[38] ), .ZN(n1458) );
  XNOR2_X1 U3600 ( .A(\MC_ARK_ARC_1_0/temp4[38] ), .B(
        \MC_ARK_ARC_1_0/temp2[38] ), .ZN(n1459) );
  NAND3_X1 U3601 ( .A1(\SB1_0_24/i0_3 ), .A2(\SB1_0_24/i0_0 ), .A3(
        \SB1_0_24/i0_4 ), .ZN(\SB1_0_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3602 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0_0 ), .A3(
        \SB1_0_7/i0_4 ), .ZN(\SB1_0_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3603 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i0_0 ), .A3(
        \SB1_3_25/i0_4 ), .ZN(\SB1_3_25/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U3604 ( .A(n1460), .B(n208), .ZN(Ciphertext[54]) );
  NAND4_X1 U3605 ( .A1(\SB4_22/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_22/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_22/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_22/Component_Function_0/NAND4_in[0] ), .ZN(n1460) );
  NAND3_X1 U3607 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i1[9] ), .A3(
        \SB1_3_5/i0_4 ), .ZN(\SB1_3_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3608 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i1[9] ), .A3(
        \SB1_3_16/i0_4 ), .ZN(\SB1_3_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3609 ( .A1(n2106), .A2(\SB4_31/i1[9] ), .A3(\SB4_31/i0_4 ), .ZN(
        \SB4_31/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U3610 ( .A(n1462), .B(n250), .ZN(Ciphertext[130]) );
  NAND4_X1 U3611 ( .A1(\SB4_10/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_10/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_10/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_10/Component_Function_4/NAND4_in[1] ), .ZN(n1462) );
  XNOR2_X1 U3612 ( .A(n1463), .B(n199), .ZN(Ciphertext[28]) );
  NAND4_X1 U3613 ( .A1(\SB4_27/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_27/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_27/Component_Function_4/NAND4_in[1] ), .ZN(n1463) );
  XNOR2_X1 U3615 ( .A(n1465), .B(n240), .ZN(Ciphertext[22]) );
  NAND4_X1 U3616 ( .A1(\SB4_28/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_28/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_28/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_28/Component_Function_4/NAND4_in[1] ), .ZN(n1465) );
  XNOR2_X1 U3617 ( .A(n1466), .B(n358), .ZN(Ciphertext[4]) );
  NAND3_X1 U3618 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i0[9] ), .A3(
        \SB1_3_16/i0[8] ), .ZN(\SB1_3_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3619 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i0[9] ), .A3(
        \SB1_3_11/i0[8] ), .ZN(\SB1_3_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3620 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0[9] ), .A3(
        \SB1_2_12/i0[8] ), .ZN(\SB1_2_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3621 ( .A1(\SB1_2_28/i0_3 ), .A2(\SB1_2_28/i0[9] ), .A3(
        \SB1_2_28/i0[8] ), .ZN(\SB1_2_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3622 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i0[9] ), .A3(
        \SB1_2_8/i0[8] ), .ZN(\SB1_2_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3623 ( .A1(\SB1_3_20/i0_3 ), .A2(\SB1_3_20/i0[9] ), .A3(
        \SB1_3_20/i0[8] ), .ZN(\SB1_3_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3624 ( .A1(\SB1_2_23/i0_3 ), .A2(\SB1_2_23/i0[9] ), .A3(
        \SB1_2_23/i0[8] ), .ZN(\SB1_2_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3625 ( .A1(\SB1_2_17/i0_3 ), .A2(\SB1_2_17/i0[9] ), .A3(
        \SB1_2_17/i0[8] ), .ZN(\SB1_2_17/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U3626 ( .A(\RI1[3][35] ), .ZN(\SB1_3_26/i0_3 ) );
  XNOR2_X1 U3627 ( .A(\MC_ARK_ARC_1_2/temp5[35] ), .B(
        \MC_ARK_ARC_1_2/temp6[35] ), .ZN(\RI1[3][35] ) );
  NAND3_X1 U3628 ( .A1(\SB2_0_30/i0_4 ), .A2(\SB2_0_30/i0[9] ), .A3(
        \SB2_0_30/i0[6] ), .ZN(n1467) );
  NAND3_X1 U3629 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i0_4 ), 
        .ZN(\SB3_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3630 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i1[9] ), .A3(\SB3_19/i0_4 ), 
        .ZN(\SB3_19/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U3631 ( .A1(\SB2_0_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_3/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_0_3/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_0_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][1] ) );
  NAND4_X2 U3632 ( .A1(\SB1_3_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_12/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][124] ) );
  NAND4_X2 U3634 ( .A1(\SB2_3_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_23/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][73] ) );
  NAND4_X2 U3635 ( .A1(\SB2_3_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_23/Component_Function_0/NAND4_in[2] ), .ZN(\RI5[3][78] ) );
  NAND4_X2 U3636 ( .A1(\SB2_3_24/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_24/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][67] ) );
  NAND4_X2 U3637 ( .A1(\SB2_3_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_24/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][57] ) );
  NAND4_X2 U3638 ( .A1(\SB2_3_25/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_25/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_3_25/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][46] ) );
  NAND4_X2 U3639 ( .A1(\SB2_3_25/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_25/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_3_25/Component_Function_0/NAND4_in[2] ), .ZN(\RI5[3][66] ) );
  NAND4_X2 U3640 ( .A1(\SB2_3_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_25/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][61] ) );
  NAND4_X2 U3642 ( .A1(\SB2_3_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][79] ) );
  NAND4_X2 U3644 ( .A1(\SB2_3_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_26/Component_Function_0/NAND4_in[2] ), .ZN(\RI5[3][60] ) );
  NAND4_X2 U3645 ( .A1(\SB2_3_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_26/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][55] ) );
  NAND4_X2 U3647 ( .A1(\SB2_3_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_19/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][97] ) );
  NAND4_X2 U3648 ( .A1(\SB2_3_19/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_19/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_19/Component_Function_2/NAND4_in[0] ), .ZN(\RI5[3][92] ) );
  NAND4_X2 U3649 ( .A1(\SB2_3_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_19/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][87] ) );
  NAND4_X2 U3650 ( .A1(\SB2_3_19/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_19/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_19/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_3_19/Component_Function_4/NAND4_in[1] ), .ZN(\RI5[3][82] ) );
  NAND4_X2 U3653 ( .A1(\SB2_3_16/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_16/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][120] ) );
  NAND4_X2 U3654 ( .A1(\SB2_3_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_16/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_16/Component_Function_1/NAND4_in[1] ), .ZN(\RI5[3][115] ) );
  NAND4_X2 U3655 ( .A1(\SB2_3_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_17/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][94] ) );
  NAND4_X2 U3656 ( .A1(\SB2_3_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_17/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][109] ) );
  NAND4_X2 U3657 ( .A1(\SB2_3_21/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_21/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][90] ) );
  NAND4_X2 U3658 ( .A1(\SB2_3_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_21/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][85] ) );
  NAND4_X2 U3660 ( .A1(\SB2_3_15/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_15/Component_Function_1/NAND4_in[0] ), .ZN(\RI5[3][121] ) );
  NAND4_X2 U3661 ( .A1(\SB2_3_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_11/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][145] ) );
  NAND4_X2 U3662 ( .A1(\SB2_3_11/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_3_11/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_11/Component_Function_2/NAND4_in[0] ), .ZN(\RI5[3][140] ) );
  NAND4_X2 U3664 ( .A1(\SB2_3_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_11/Component_Function_0/NAND4_in[2] ), .ZN(\RI5[3][150] ) );
  NAND4_X2 U3665 ( .A1(\SB2_3_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_12/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][139] ) );
  NAND4_X2 U3666 ( .A1(\SB2_3_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][133] ) );
  NAND4_X2 U3667 ( .A1(\SB2_3_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_14/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][127] ) );
  NAND4_X2 U3669 ( .A1(\SB2_3_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_7/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][159] ) );
  NAND4_X2 U3670 ( .A1(\SB2_3_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_8/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][163] ) );
  NAND4_X2 U3671 ( .A1(\SB2_3_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_8/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_8/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][153] ) );
  NAND4_X2 U3674 ( .A1(\SB2_3_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_9/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][157] ) );
  NAND4_X2 U3675 ( .A1(\SB2_3_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_10/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][156] ) );
  NAND4_X2 U3676 ( .A1(\SB2_3_10/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_10/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][151] ) );
  NAND4_X2 U3677 ( .A1(\SB2_3_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_3/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][1] ) );
  NAND4_X2 U3678 ( .A1(\SB2_3_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_3/Component_Function_0/NAND4_in[1] ), .ZN(\RI5[3][6] ) );
  NAND4_X2 U3679 ( .A1(\SB2_3_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][187] ) );
  NAND4_X2 U3680 ( .A1(\SB2_3_4/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_4/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][0] ) );
  NAND4_X2 U3681 ( .A1(\SB2_3_5/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_5/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][171] ) );
  NAND4_X2 U3682 ( .A1(\SB2_3_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_5/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_5/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][186] ) );
  NAND4_X2 U3683 ( .A1(\SB2_3_5/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_5/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_5/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][181] ) );
  NAND4_X2 U3685 ( .A1(\SB2_3_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_1/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_1/Component_Function_0/NAND4_in[1] ), .ZN(\RI5[3][18] ) );
  NAND4_X2 U3686 ( .A1(\SB2_3_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_1/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][13] ) );
  NAND4_X2 U3687 ( .A1(\SB2_3_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_2/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][7] ) );
  NAND4_X2 U3688 ( .A1(\SB2_3_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_6/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_6/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_6/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][160] ) );
  NAND4_X2 U3689 ( .A1(\SB2_3_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_6/Component_Function_0/NAND4_in[2] ), .ZN(\RI5[3][180] ) );
  NAND4_X2 U3690 ( .A1(\SB2_3_6/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_6/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][175] ) );
  NAND4_X2 U3691 ( .A1(\SB2_3_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_29/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][37] ) );
  NAND4_X2 U3692 ( .A1(\SB2_3_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_29/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_29/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][27] ) );
  NAND4_X2 U3693 ( .A1(\SB2_3_30/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_30/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_30/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][31] ) );
  NAND4_X2 U3694 ( .A1(\SB2_3_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_30/Component_Function_0/NAND4_in[1] ), .ZN(\RI5[3][36] ) );
  NAND4_X2 U3695 ( .A1(\SB2_3_31/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_31/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_3_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_31/Component_Function_0/NAND4_in[1] ), .ZN(\RI5[3][30] ) );
  NAND4_X2 U3696 ( .A1(\SB2_3_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_31/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_31/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_3_31/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][25] ) );
  NAND4_X2 U3697 ( .A1(\SB2_3_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_27/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][54] ) );
  NAND4_X2 U3698 ( .A1(\SB2_3_28/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_3_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_28/Component_Function_2/NAND4_in[0] ), .ZN(\RI5[3][38] ) );
  NAND4_X2 U3699 ( .A1(\SB2_3_28/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_28/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][48] ) );
  NAND4_X2 U3700 ( .A1(\SB2_3_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_28/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][43] ) );
  NAND4_X2 U3701 ( .A1(\SB2_3_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_0/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][9] ) );
  NAND4_X2 U3702 ( .A1(\SB2_3_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_0/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][24] ) );
  NAND4_X2 U3703 ( .A1(\SB2_3_0/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_0/Component_Function_1/NAND4_in[0] ), .ZN(\RI5[3][19] ) );
  CLKBUF_X1 U3704 ( .A(Key[161]), .Z(n392) );
  BUF_X2 U852 ( .A(\RI5[3][131] ), .Z(n801) );
  BUF_X2 \SB1_1_3/BUF_3  ( .A(\RI1[1][171] ), .Z(\SB1_1_3/i0[8] ) );
  BUF_X1 U608 ( .A(\RI1[4][119] ), .Z(\SB3_12/i1_5 ) );
  BUF_X2 \SB2_1_11/BUF_1  ( .A(\RI3[1][121] ), .Z(\SB2_1_11/i0[6] ) );
  BUF_X2 \SB2_1_19/BUF_0  ( .A(\RI3[1][72] ), .Z(\SB2_1_19/i0[9] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_158  ( .A(\RI5[2][158] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[158] ) );
  BUF_X2 \SB1_2_22/BUF_3  ( .A(\RI1[2][57] ), .Z(\SB1_2_22/i0[8] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_3/BUF_14  ( .A(\RI5[3][14] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[14] ) );
  BUF_X2 U633 ( .A(\RI1[2][176] ), .Z(\SB1_2_2/i1[9] ) );
  BUF_X2 \SB4_18/BUF_1  ( .A(\RI3[4][79] ), .Z(\SB4_18/i0[6] ) );
  INV_X1 \SB1_0_31/INV_5  ( .A(n187), .ZN(\SB1_0_31/i0_3 ) );
  INV_X1 U631 ( .A(n67), .ZN(\SB1_0_11/i0_3 ) );
  BUF_X2 U628 ( .A(\RI1[1][75] ), .Z(\SB1_1_19/i0[8] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_3/BUF_154  ( .A(\RI5[3][154] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[154] ) );
  BUF_X2 \SB2_0_6/BUF_0  ( .A(\RI3[0][150] ), .Z(\SB2_0_6/i0[9] ) );
  BUF_X1 \SB1_1_29/BUF_1  ( .A(\RI1[1][13] ), .Z(\SB1_1_29/i1_7 ) );
  BUF_X2 U650 ( .A(\RI3[0][137] ), .Z(\SB2_0_9/i0_3 ) );
  BUF_X2 \SB2_3_30/BUF_0  ( .A(\RI3[3][6] ), .Z(\SB2_3_30/i0[9] ) );
  BUF_X2 \SB2_2_13/BUF_0  ( .A(\RI3[2][108] ), .Z(\SB2_2_13/i0[9] ) );
  BUF_X2 \SB2_0_8/BUF_2  ( .A(\RI3[0][140] ), .Z(\SB2_0_8/i0_0 ) );
  INV_X1 U623 ( .A(n91), .ZN(\SB1_0_15/i0_3 ) );
  BUF_X2 \SB4_13/BUF_0  ( .A(\RI3[4][108] ), .Z(\SB4_13/i0[9] ) );
  INV_X1 U187 ( .A(n444), .ZN(n320) );
  INV_X1 U502 ( .A(n458), .ZN(n302) );
  BUF_X1 \SB1_2_20/BUF_0  ( .A(\RI1[2][66] ), .Z(\SB1_2_20/i3[0] ) );
  BUF_X2 \SB2_0_19/BUF_1  ( .A(\RI3[0][73] ), .Z(\SB2_0_19/i0[6] ) );
  INV_X1 \SB1_1_30/INV_4  ( .A(\RI1[1][10] ), .ZN(\SB1_1_30/i0_4 ) );
  BUF_X2 \SB2_0_17/BUF_3  ( .A(\RI3[0][87] ), .Z(\SB2_0_17/i0[10] ) );
  BUF_X1 \SB1_2_17/BUF_1  ( .A(\RI1[2][85] ), .Z(\SB1_2_17/i1_7 ) );
  BUF_X2 \SB1_1_16/BUF_2  ( .A(\RI1[1][92] ), .Z(\SB1_1_16/i1[9] ) );
  BUF_X2 \SB4_9/BUF_1  ( .A(\RI3[4][133] ), .Z(\SB4_9/i0[6] ) );
  NAND4_X2 U1693 ( .A1(\SB2_0_30/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_30/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_30/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_30/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[21] ) );
  BUF_X2 \SB2_0_25/BUF_5  ( .A(\RI3[0][41] ), .Z(\SB2_0_25/i0_3 ) );
  BUF_X2 \SB2_0_8/BUF_3  ( .A(\RI3[0][141] ), .Z(\SB2_0_8/i0[10] ) );
  BUF_X2 \SB2_0_30/BUF_5  ( .A(\RI3[0][11] ), .Z(\SB2_0_30/i0_3 ) );
  BUF_X2 \SB2_2_3/BUF_0  ( .A(\RI3[2][168] ), .Z(\SB2_2_3/i0[9] ) );
  BUF_X1 \SB3_26/BUF_0  ( .A(\RI1[4][30] ), .Z(\SB3_26/i3[0] ) );
  NAND4_X2 U3299 ( .A1(\SB2_0_31/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_0_31/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_0_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[5] ) );
  INV_X1 \SB1_0_8/INV_5  ( .A(n49), .ZN(\SB1_0_8/i0_3 ) );
  BUF_X1 \SB1_3_7/BUF_1  ( .A(\RI1[3][145] ), .Z(\SB1_3_7/i1_7 ) );
  BUF_X2 \SB2_0_17/BUF_0  ( .A(\RI3[0][84] ), .Z(\SB2_0_17/i0[9] ) );
  INV_X1 \SB1_0_22/INV_5  ( .A(n133), .ZN(\SB1_0_22/i0_3 ) );
  BUF_X1 \SB1_2_15/BUF_1  ( .A(\RI1[2][97] ), .Z(\SB1_2_15/i1_7 ) );
  BUF_X2 \SB1_0_13/BUF_2  ( .A(n82), .Z(\SB1_0_13/i1[9] ) );
  BUF_X2 U568 ( .A(\RI3[0][134] ), .Z(\SB2_0_9/i0_0 ) );
  INV_X1 U190 ( .A(n450), .ZN(n292) );
  BUF_X2 U558 ( .A(\RI3[2][174] ), .Z(\SB2_2_2/i0[9] ) );
  BUF_X2 \SB2_1_26/BUF_0  ( .A(\RI3[1][30] ), .Z(\SB2_1_26/i0[9] ) );
  BUF_X2 \SB2_0_1/BUF_1  ( .A(\RI3[0][181] ), .Z(\SB2_0_1/i0[6] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_64  ( .A(\RI5[0][64] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[64] ) );
  BUF_X1 U1558 ( .A(\RI5[3][113] ), .Z(n796) );
  INV_X1 \SB1_0_9/INV_5  ( .A(n55), .ZN(\SB1_0_9/i0_3 ) );
  BUF_X1 \SB3_12/BUF_0  ( .A(\RI1[4][114] ), .Z(\SB3_12/i3[0] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_61  ( .A(\RI5[2][61] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[61] ) );
  BUF_X1 \SB3_17/BUF_0  ( .A(\RI1[4][84] ), .Z(\SB3_17/i3[0] ) );
  BUF_X1 \SB1_3_24/BUF_1  ( .A(\RI1[3][43] ), .Z(\SB1_3_24/i1_7 ) );
  BUF_X1 \SB1_2_10/BUF_1  ( .A(\RI1[2][127] ), .Z(\SB1_2_10/i1_7 ) );
  INV_X1 U153 ( .A(\MC_ARK_ARC_1_0/buf_keyinput[40] ), .ZN(n286) );
  BUF_X2 \SB2_0_3/BUF_1  ( .A(\RI3[0][169] ), .Z(\SB2_0_3/i0[6] ) );
  BUF_X1 \SB3_9/BUF_0  ( .A(\RI1[4][132] ), .Z(\SB3_9/i3[0] ) );
  NAND4_X2 U2763 ( .A1(\SB2_0_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_21/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_21/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[65] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_80  ( .A(\RI5[0][80] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[80] ) );
  BUF_X2 U648 ( .A(\RI3[1][155] ), .Z(\SB2_1_6/i0_3 ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_94  ( .A(\RI5[2][94] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[94] ) );
  INV_X1 \SB1_0_3/INV_5  ( .A(n19), .ZN(\SB1_0_3/i0_3 ) );
  INV_X1 \SB1_3_21/INV_2  ( .A(\RI1[3][62] ), .ZN(\SB1_3_21/i0_0 ) );
  INV_X1 \SB1_2_5/INV_0  ( .A(\RI1[2][156] ), .ZN(\SB1_2_5/i0[9] ) );
  BUF_X1 \SB1_2_28/BUF_1  ( .A(\RI1[2][19] ), .Z(\SB1_2_28/i1_7 ) );
  INV_X1 U632 ( .A(n127), .ZN(\SB1_0_21/i0_3 ) );
  BUF_X1 \SB3_27/BUF_0  ( .A(\RI1[4][24] ), .Z(\SB3_27/i3[0] ) );
  BUF_X2 \SB2_0_13/BUF_0  ( .A(\RI3[0][108] ), .Z(\SB2_0_13/i0[9] ) );
  BUF_X1 U766 ( .A(n11), .Z(\SB1_0_1/i1_7 ) );
  BUF_X2 \SB2_0_28/BUF_3  ( .A(\RI3[0][21] ), .Z(\SB2_0_28/i0[10] ) );
  BUF_X2 \SB2_0_28/BUF_2  ( .A(\RI3[0][20] ), .Z(\SB2_0_28/i0_0 ) );
  INV_X1 \SB1_2_31/INV_3  ( .A(\RI1[2][3] ), .ZN(\SB1_2_31/i0[10] ) );
  INV_X1 \SB1_0_8/INV_4  ( .A(n50), .ZN(\SB1_0_8/i0_4 ) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_106  ( .A(\RI5[0][106] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[106] ) );
  INV_X1 U201 ( .A(n451), .ZN(n247) );
  INV_X1 U102 ( .A(Key[139]), .ZN(n243) );
  INV_X1 U229 ( .A(\MC_ARK_ARC_1_3/buf_keyinput[179] ), .ZN(n220) );
  BUF_X2 U639 ( .A(\RI3[0][143] ), .Z(\SB2_0_8/i0_3 ) );
  NAND4_X2 U745 ( .A1(\SB2_2_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_21/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[65] ) );
  INV_X1 U188 ( .A(n484), .ZN(n206) );
  BUF_X2 \SB2_0_28/BUF_0  ( .A(\RI3[0][18] ), .Z(\SB2_0_28/i0[9] ) );
  INV_X1 U626 ( .A(n97), .ZN(\SB1_0_16/i0_3 ) );
  BUF_X1 \SB1_2_3/BUF_1  ( .A(\RI1[2][169] ), .Z(\SB1_2_3/i1_7 ) );
  BUF_X1 \SB1_1_16/BUF_1  ( .A(\RI1[1][91] ), .Z(\SB1_1_16/i1_7 ) );
  BUF_X1 \SB1_1_7/BUF_1  ( .A(\RI1[1][145] ), .Z(\SB1_1_7/i1_7 ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_86  ( .A(\RI5[1][86] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[86] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_181  ( .A(\RI5[2][181] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[181] ) );
  BUF_X2 \SB4_31/BUF_0  ( .A(\RI3[4][0] ), .Z(\SB4_31/i0[9] ) );
  BUF_X2 \SB2_0_21/BUF_0  ( .A(\RI3[0][60] ), .Z(\SB2_0_21/i0[9] ) );
  INV_X2 U689 ( .A(n7), .ZN(\SB1_0_1/i0_3 ) );
  BUF_X2 \SB2_3_3/BUF_1  ( .A(\RI3[3][169] ), .Z(\SB2_3_3/i0[6] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_8  ( .A(\RI5[0][8] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[8] ) );
  INV_X1 U686 ( .A(n157), .ZN(\SB1_0_26/i0_3 ) );
  BUF_X1 \SB1_2_6/BUF_1  ( .A(\RI1[2][151] ), .Z(\SB1_2_6/i1_7 ) );
  BUF_X1 \SB3_29/BUF_0  ( .A(\RI1[4][12] ), .Z(\SB3_29/i3[0] ) );
  BUF_X1 \SB1_3_22/BUF_1  ( .A(\RI1[3][55] ), .Z(\SB1_3_22/i1_7 ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_190  ( .A(\RI5[0][190] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[190] ) );
  NAND4_X2 U1747 ( .A1(n996), .A2(\SB2_2_16/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_2_16/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[95] ) );
  INV_X1 \SB1_0_19/INV_4  ( .A(n116), .ZN(\SB1_0_19/i0_4 ) );
  INV_X1 \SB1_1_8/INV_4  ( .A(\RI1[1][142] ), .ZN(\SB1_1_8/i0_4 ) );
  BUF_X1 \SB1_3_21/BUF_1  ( .A(\RI1[3][61] ), .Z(\SB1_3_21/i1_7 ) );
  BUF_X1 \SB1_3_18/BUF_1  ( .A(\RI1[3][79] ), .Z(\SB1_3_18/i1_7 ) );
  BUF_X2 \SB2_0_14/BUF_3  ( .A(\RI3[0][105] ), .Z(\SB2_0_14/i0[10] ) );
  BUF_X2 U670 ( .A(\RI3[3][115] ), .Z(\SB2_3_12/i0[6] ) );
  NAND4_X2 U2070 ( .A1(\SB2_1_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_19/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[77] ) );
  BUF_X1 \SB1_3_20/BUF_1  ( .A(\RI1[3][67] ), .Z(\SB1_3_20/i1_7 ) );
  BUF_X1 \SB3_4/BUF_0  ( .A(\RI1[4][162] ), .Z(\SB3_4/i3[0] ) );
  BUF_X2 \SB2_0_24/BUF_5  ( .A(\RI3[0][47] ), .Z(\SB2_0_24/i0_3 ) );
  NAND4_X2 U3242 ( .A1(\SB2_1_9/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_9/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_9/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[137] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_130  ( .A(\RI5[0][130] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[130] ) );
  BUF_X2 \SB2_3_3/BUF_2  ( .A(\RI3[3][170] ), .Z(\SB2_3_3/i0_0 ) );
  NAND4_X4 U1069 ( .A1(\SB2_3_24/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_24/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_24/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_24/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[52] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_164  ( .A(\RI5[2][164] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[164] ) );
  INV_X1 U297 ( .A(n508), .ZN(n200) );
  BUF_X2 \SB2_0_24/BUF_0  ( .A(\RI3[0][42] ), .Z(\SB2_0_24/i0[9] ) );
  BUF_X2 \SB4_26/BUF_1  ( .A(\RI3[4][31] ), .Z(\SB4_26/i0[6] ) );
  INV_X1 \SB1_1_20/INV_3  ( .A(\RI1[1][69] ), .ZN(\SB1_1_20/i0[10] ) );
  BUF_X1 \SB1_3_26/BUF_1  ( .A(\RI1[3][31] ), .Z(\SB1_3_26/i1_7 ) );
  BUF_X1 U798 ( .A(\RI1[2][115] ), .Z(\SB1_2_12/i1_7 ) );
  NAND4_X2 U759 ( .A1(\SB2_0_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_5/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_5/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[161] ) );
  BUF_X2 \SB2_1_27/BUF_0  ( .A(\RI3[1][24] ), .Z(\SB2_1_27/i0[9] ) );
  BUF_X1 U1616 ( .A(\RI3[4][125] ), .Z(\SB4_11/i0_3 ) );
  CLKBUF_X1 U24 ( .A(Key[188]), .Z(n498) );
  CLKBUF_X1 U39 ( .A(Key[104]), .Z(n477) );
  INV_X1 U236 ( .A(\MC_ARK_ARC_1_1/buf_keyinput[8] ), .ZN(n329) );
  CLKBUF_X1 U45 ( .A(Key[152]), .Z(n485) );
  CLKBUF_X1 U34 ( .A(Key[100]), .Z(n463) );
  CLKBUF_X1 U80 ( .A(Key[44]), .Z(n475) );
  CLKBUF_X1 U719 ( .A(Key[156]), .Z(n377) );
  CLKBUF_X1 U6 ( .A(Key[184]), .Z(n474) );
  CLKBUF_X1 U123 ( .A(Key[107]), .Z(n388) );
  CLKBUF_X1 U32 ( .A(Key[135]), .Z(n510) );
  CLKBUF_X1 U63 ( .A(Key[68]), .Z(n486) );
  CLKBUF_X1 U72 ( .A(Key[39]), .Z(n472) );
  BUF_X1 U69 ( .A(Key[81]), .Z(n488) );
  CLKBUF_X1 U76 ( .A(Key[172]), .Z(n470) );
  CLKBUF_X1 U1 ( .A(Key[52]), .Z(n375) );
  CLKBUF_X1 U22 ( .A(Key[45]), .Z(n453) );
  CLKBUF_X1 U23 ( .A(Key[38]), .Z(n480) );
  CLKBUF_X1 U99 ( .A(Key[56]), .Z(n437) );
  CLKBUF_X1 U54 ( .A(Key[26]), .Z(n466) );
  CLKBUF_X1 U90 ( .A(Key[28]), .Z(n448) );
  INV_X1 \SB1_0_25/INV_4  ( .A(n152), .ZN(\SB1_0_25/i0_4 ) );
  BUF_X1 \SB1_0_5/BUF_3  ( .A(n33), .Z(\SB1_0_5/i0[8] ) );
  INV_X1 \SB1_0_29/INV_4  ( .A(n176), .ZN(\SB1_0_29/i0_4 ) );
  INV_X1 \SB1_0_0/INV_0  ( .A(n6), .ZN(\SB1_0_0/i0[9] ) );
  BUF_X1 U763 ( .A(n63), .Z(\SB1_0_10/i0[8] ) );
  INV_X1 \SB1_0_10/INV_4  ( .A(n62), .ZN(\SB1_0_10/i0_4 ) );
  INV_X1 \SB1_0_23/INV_3  ( .A(n141), .ZN(\SB1_0_23/i0[10] ) );
  INV_X1 \SB1_0_21/INV_4  ( .A(n128), .ZN(\SB1_0_21/i0_4 ) );
  BUF_X1 \SB1_0_9/BUF_2  ( .A(n58), .Z(\SB1_0_9/i1[9] ) );
  INV_X1 \SB1_0_16/INV_4  ( .A(n98), .ZN(\SB1_0_16/i0_4 ) );
  INV_X1 \SB1_0_12/INV_2  ( .A(n76), .ZN(\SB1_0_12/i0_0 ) );
  BUF_X1 \SB1_0_18/BUF_3  ( .A(n111), .Z(\SB1_0_18/i0[8] ) );
  INV_X1 \SB1_0_23/INV_4  ( .A(n140), .ZN(\SB1_0_23/i0_4 ) );
  INV_X1 U769 ( .A(n83), .ZN(\SB1_0_13/i0[6] ) );
  INV_X1 U672 ( .A(n43), .ZN(\SB1_0_7/i0_3 ) );
  INV_X1 U143 ( .A(n388), .ZN(n273) );
  BUF_X1 \SB1_0_23/BUF_3  ( .A(n141), .Z(\SB1_0_23/i0[8] ) );
  BUF_X1 \SB2_0_3/BUF_0  ( .A(\RI3[0][168] ), .Z(\SB2_0_3/i0[9] ) );
  BUF_X1 \SB2_0_7/BUF_0  ( .A(\RI3[0][144] ), .Z(\SB2_0_7/i0[9] ) );
  BUF_X1 U776 ( .A(\RI3[0][102] ), .Z(\SB2_0_14/i0[9] ) );
  NAND4_X1 U1555 ( .A1(n1230), .A2(\SB2_0_1/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_1/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_1/Component_Function_5/NAND4_in[0] ), .ZN(n794) );
  NAND4_X2 U1098 ( .A1(n965), .A2(\SB2_0_27/Component_Function_4/NAND4_in[3] ), 
        .A3(\SB2_0_27/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_27/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[34] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_32  ( .A(\RI5[0][32] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[32] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_168  ( .A(\RI5[0][168] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[168] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_36  ( .A(\RI5[0][36] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[36] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_187  ( .A(\RI5[0][187] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[187] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_12  ( .A(\RI5[0][12] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[12] ) );
  INV_X1 \SB1_1_3/INV_4  ( .A(\RI1[1][172] ), .ZN(\SB1_1_3/i0_4 ) );
  BUF_X1 \SB1_1_15/BUF_3  ( .A(\RI1[1][99] ), .Z(\SB1_1_15/i0[8] ) );
  INV_X1 \SB1_1_4/INV_1  ( .A(\RI1[1][163] ), .ZN(\SB1_1_4/i0[6] ) );
  BUF_X1 \SB2_1_13/BUF_0  ( .A(\RI3[1][108] ), .Z(\SB2_1_13/i0[9] ) );
  BUF_X1 \SB2_1_18/BUF_1  ( .A(\RI3[1][79] ), .Z(\SB2_1_18/i0[6] ) );
  BUF_X1 \SB2_1_3/BUF_0  ( .A(\RI3[1][168] ), .Z(\SB2_1_3/i0[9] ) );
  BUF_X1 \SB2_1_28/BUF_1  ( .A(\RI3[1][19] ), .Z(\SB2_1_28/i0[6] ) );
  BUF_X1 \SB2_1_29/BUF_0  ( .A(\RI3[1][12] ), .Z(\SB2_1_29/i0[9] ) );
  BUF_X1 U785 ( .A(\RI3[1][126] ), .Z(\SB2_1_10/i0[9] ) );
  BUF_X1 U531 ( .A(\RI3[1][1] ), .Z(\SB2_1_31/i0[6] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_44  ( .A(\RI5[1][44] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[44] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_127  ( .A(\RI5[1][127] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[127] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_156  ( .A(\RI5[1][156] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[156] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_31  ( .A(\RI5[1][31] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[31] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_150  ( .A(\RI5[1][150] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[150] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_187  ( .A(\RI5[1][187] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[187] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_181  ( .A(\RI5[1][181] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[181] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_139  ( .A(\RI5[1][139] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[139] ) );
  INV_X1 \SB1_2_16/INV_0  ( .A(\RI1[2][90] ), .ZN(\SB1_2_16/i0[9] ) );
  BUF_X2 \SB1_2_6/BUF_3  ( .A(\RI1[2][153] ), .Z(\SB1_2_6/i0[8] ) );
  BUF_X1 U801 ( .A(\RI3[2][1] ), .Z(\SB2_2_31/i0[6] ) );
  BUF_X1 \SB2_2_29/BUF_0  ( .A(\RI3[2][12] ), .Z(\SB2_2_29/i0[9] ) );
  BUF_X1 \SB2_2_14/BUF_1  ( .A(\RI3[2][103] ), .Z(\SB2_2_14/i0[6] ) );
  BUF_X1 \SB2_2_27/BUF_0  ( .A(\RI3[2][24] ), .Z(\SB2_2_27/i0[9] ) );
  BUF_X1 U746 ( .A(\RI3[2][84] ), .Z(\SB2_2_17/i0[9] ) );
  INV_X1 \SB2_2_7/INV_2  ( .A(\RI3[2][146] ), .ZN(\SB2_2_7/i1[9] ) );
  NAND4_X2 U544 ( .A1(\SB2_2_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_30/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_30/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][21] ) );
  NAND4_X2 U1756 ( .A1(\SB2_2_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_24/Component_Function_3/NAND4_in[2] ), .A4(n1065), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[57] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_146  ( .A(\RI5[2][146] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[146] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_140  ( .A(\RI5[2][140] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[140] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_115  ( .A(\RI5[2][115] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[115] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_124  ( .A(\RI5[2][124] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[124] ) );
  BUF_X2 U742 ( .A(\RI5[2][19] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[19] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_25  ( .A(\RI5[2][25] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[25] ) );
  BUF_X1 U619 ( .A(\RI1[3][122] ), .Z(\SB1_3_11/i1[9] ) );
  INV_X1 \SB1_3_15/INV_3  ( .A(\RI1[3][99] ), .ZN(\SB1_3_15/i0[10] ) );
  BUF_X1 \SB2_3_15/BUF_0  ( .A(\RI3[3][96] ), .Z(\SB2_3_15/i0[9] ) );
  BUF_X1 \SB2_3_13/BUF_1  ( .A(\RI3[3][109] ), .Z(\SB2_3_13/i0[6] ) );
  BUF_X1 \SB2_3_11/BUF_1  ( .A(\RI3[3][121] ), .Z(\SB2_3_11/i0[6] ) );
  BUF_X1 U642 ( .A(\RI3[3][145] ), .Z(\SB2_3_7/i0[6] ) );
  BUF_X1 \SB2_3_4/BUF_1  ( .A(\RI3[3][163] ), .Z(\SB2_3_4/i0[6] ) );
  BUF_X1 \SB2_3_27/BUF_0  ( .A(\RI3[3][24] ), .Z(\SB2_3_27/i0[9] ) );
  BUF_X2 U645 ( .A(\MC_ARK_ARC_1_3/buf_datainput[125] ), .Z(n521) );
  CLKBUF_X1 \SB3_26/BUF_4  ( .A(\RI1[4][34] ), .Z(\SB3_26/i0[7] ) );
  BUF_X2 \SB2_3_28/BUF_2  ( .A(\RI3[3][20] ), .Z(\SB2_3_28/i0_0 ) );
  CLKBUF_X3 U546 ( .A(\RI5[3][141] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[141] )
         );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_152  ( .A(\RI5[2][152] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[152] ) );
  BUF_X1 \SB1_0_2/BUF_3  ( .A(n15), .Z(\SB1_0_2/i0[8] ) );
  BUF_X1 U773 ( .A(n105), .Z(\SB1_0_17/i0[8] ) );
  BUF_X1 \SB1_0_29/BUF_5  ( .A(n175), .Z(\SB1_0_29/i1_5 ) );
  BUF_X1 \SB1_0_7/BUF_3  ( .A(n45), .Z(\SB1_0_7/i0[8] ) );
  NAND4_X2 \SB2_0_26/Component_Function_0/N5  ( .A1(
        \SB2_0_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_26/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][60] ) );
  NAND4_X2 \SB2_0_9/Component_Function_1/N5  ( .A1(
        \SB2_0_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_9/Component_Function_1/NAND4_in[2] ), .ZN(\RI5[0][157] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_128  ( .A(\RI5[0][128] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[128] ) );
  BUF_X1 \SB1_1_24/BUF_3  ( .A(\RI1[1][45] ), .Z(\SB1_1_24/i0[8] ) );
  BUF_X1 \SB1_1_8/BUF_3  ( .A(\RI1[1][141] ), .Z(\SB1_1_8/i0[8] ) );
  NAND4_X2 \SB2_1_4/Component_Function_3/N5  ( .A1(
        \SB2_1_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][177] ) );
  NAND4_X2 \SB2_1_12/Component_Function_3/N5  ( .A1(
        \SB2_1_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_12/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][129] ) );
  BUF_X1 \SB1_2_29/BUF_5  ( .A(\RI1[2][17] ), .Z(\SB1_2_29/i1_5 ) );
  BUF_X1 \SB1_2_21/BUF_3  ( .A(\RI1[2][63] ), .Z(\SB1_2_21/i0[8] ) );
  BUF_X1 \SB1_2_1/BUF_3  ( .A(\RI1[2][183] ), .Z(\SB1_2_1/i0[8] ) );
  NAND4_X2 \SB2_2_13/Component_Function_3/N5  ( .A1(
        \SB2_2_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][123] ) );
  NAND4_X2 \SB2_3_1/Component_Function_3/N5  ( .A1(
        \SB2_3_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_1/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_1/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][3] ) );
  NAND4_X2 \SB2_3_23/Component_Function_3/N5  ( .A1(
        \SB2_3_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][63] ) );
  BUF_X1 \SB3_4/BUF_3  ( .A(\RI1[4][165] ), .Z(\SB3_4/i0[8] ) );
  BUF_X1 \SB3_30/BUF_2  ( .A(\RI1[4][8] ), .Z(\SB3_30/i1[9] ) );
  BUF_X1 \SB3_3/BUF_2  ( .A(\RI1[4][170] ), .Z(\SB3_3/i1[9] ) );
  BUF_X1 \SB3_16/BUF_2  ( .A(\RI1[4][92] ), .Z(\SB3_16/i1[9] ) );
  BUF_X1 U557 ( .A(\RI1[4][63] ), .Z(\SB3_21/i0[8] ) );
  BUF_X1 \SB3_13/BUF_3  ( .A(\RI1[4][111] ), .Z(\SB3_13/i0[8] ) );
  BUF_X1 U4 ( .A(\RI1[4][44] ), .Z(\SB3_24/i1[9] ) );
  CLKBUF_X2 U8 ( .A(\RI3[3][8] ), .Z(\SB2_3_30/i0_0 ) );
  BUF_X1 U9 ( .A(\RI3[3][133] ), .Z(\SB2_3_9/i0[6] ) );
  BUF_X2 U112 ( .A(\RI1[3][74] ), .Z(\SB1_3_19/i1[9] ) );
  BUF_X2 U117 ( .A(\RI1[3][75] ), .Z(\SB1_3_19/i0[8] ) );
  BUF_X1 U171 ( .A(\RI3[2][181] ), .Z(\SB2_2_1/i0[6] ) );
  CLKBUF_X2 U178 ( .A(\RI1[2][33] ), .Z(\SB1_2_26/i0[8] ) );
  BUF_X1 U241 ( .A(\RI1[2][27] ), .Z(\SB1_2_27/i0[8] ) );
  BUF_X2 U253 ( .A(\RI1[1][104] ), .Z(\SB1_1_14/i1[9] ) );
  BUF_X1 U300 ( .A(n99), .Z(\SB1_0_16/i0[8] ) );
  NAND4_X2 U523 ( .A1(\SB2_3_16/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_16/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_16/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[100] ) );
  BUF_X1 U537 ( .A(\RI1[1][12] ), .Z(\SB1_1_29/i3[0] ) );
  NAND4_X2 U549 ( .A1(\SB2_1_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_13/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_13/Component_Function_5/NAND4_in[0] ), .ZN(n807) );
  BUF_X2 U567 ( .A(\RI5[3][149] ), .Z(n850) );
  NAND4_X2 U576 ( .A1(\SB2_3_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_9/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][147] ) );
  NAND4_X1 U610 ( .A1(\SB2_0_27/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_27/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_27/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[29] ) );
  NAND4_X1 U616 ( .A1(\SB2_2_13/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_13/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_13/Component_Function_4/NAND4_in[0] ), .A4(n1706), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[118] ) );
  CLKBUF_X1 U621 ( .A(\MC_ARK_ARC_1_0/buf_datainput[44] ), .Z(n1473) );
  BUF_X1 U629 ( .A(\MC_ARK_ARC_1_0/buf_datainput[44] ), .Z(n1474) );
  BUF_X1 U635 ( .A(\MC_ARK_ARC_1_0/buf_datainput[44] ), .Z(n1475) );
  NAND4_X1 U636 ( .A1(\SB2_0_27/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_27/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_27/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_27/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[44] ) );
  NAND4_X1 U655 ( .A1(\SB2_1_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][171] ) );
  CLKBUF_X1 U656 ( .A(n133), .Z(\SB1_0_22/i1_5 ) );
  BUF_X1 U661 ( .A(\MC_ARK_ARC_1_0/buf_datainput[107] ), .Z(n1480) );
  NAND4_X1 U681 ( .A1(\SB2_0_14/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_14/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_0_14/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_14/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[107] ) );
  BUF_X1 U701 ( .A(\MC_ARK_ARC_1_0/buf_datainput[41] ), .Z(n1483) );
  NAND4_X1 U704 ( .A1(n1399), .A2(\SB2_0_25/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_25/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_25/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[41] ) );
  INV_X1 U709 ( .A(Key[27]), .ZN(n348) );
  BUF_X1 U712 ( .A(\RI5[1][183] ), .Z(n1486) );
  NAND4_X1 U714 ( .A1(\SB2_1_3/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_3/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_3/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][183] ) );
  NAND4_X1 U720 ( .A1(n1052), .A2(\SB2_1_3/Component_Function_4/NAND4_in[0] ), 
        .A3(\SB2_1_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_3/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[178] ) );
  NAND4_X1 U731 ( .A1(\SB2_2_10/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_10/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_10/Component_Function_3/NAND4_in[2] ), .A4(n1214), .ZN(
        \RI5[2][141] ) );
  NAND4_X1 U741 ( .A1(\SB2_0_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_2/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_2/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_2/Component_Function_3/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[189] ) );
  NAND4_X1 U814 ( .A1(n1422), .A2(\SB2_1_25/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_1_25/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_25/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[41] ) );
  BUF_X1 U853 ( .A(\MC_ARK_ARC_1_2/buf_datainput[89] ), .Z(n1501) );
  NAND4_X1 U855 ( .A1(\SB2_2_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_17/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_17/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_17/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[89] ) );
  NAND4_X1 U863 ( .A1(\SB2_2_20/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_20/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_20/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[71] ) );
  BUF_X1 U866 ( .A(\MC_ARK_ARC_1_1/buf_datainput[71] ), .Z(n1505) );
  NAND4_X1 U868 ( .A1(\SB2_1_20/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_20/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_20/Component_Function_5/NAND4_in[3] ), .A4(n1718), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[71] ) );
  CLKBUF_X1 U874 ( .A(\RI1[4][101] ), .Z(\SB3_15/i1_5 ) );
  BUF_X1 U894 ( .A(\MC_ARK_ARC_1_0/buf_datainput[35] ), .Z(n1508) );
  CLKBUF_X1 U895 ( .A(\MC_ARK_ARC_1_0/buf_datainput[35] ), .Z(n1509) );
  NAND4_X1 U896 ( .A1(\SB2_0_26/Component_Function_5/NAND4_in[2] ), .A2(n1445), 
        .A3(n1141), .A4(\SB2_0_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[35] ) );
  CLKBUF_X3 U907 ( .A(\RI5[2][183] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[183] )
         );
  INV_X2 U946 ( .A(\RI1[3][59] ), .ZN(\SB1_3_22/i0_3 ) );
  BUF_X1 U963 ( .A(\RI1[1][1] ), .Z(\SB1_1_31/i1_7 ) );
  BUF_X2 U975 ( .A(\RI1[3][183] ), .Z(\SB1_3_1/i0[8] ) );
  INV_X1 U994 ( .A(n181), .ZN(\SB1_0_30/i0_3 ) );
  BUF_X1 U995 ( .A(n181), .Z(\SB1_0_30/i1_5 ) );
  BUF_X2 U997 ( .A(\RI3[4][175] ), .Z(\SB4_2/i0[6] ) );
  INV_X2 U1015 ( .A(\RI1[2][143] ), .ZN(\SB1_2_8/i0_3 ) );
  CLKBUF_X1 U1029 ( .A(n139), .Z(\SB1_0_23/i1_5 ) );
  BUF_X1 U1035 ( .A(\RI5[3][11] ), .Z(n1650) );
  NAND4_X2 U1048 ( .A1(\SB2_3_22/Component_Function_5/NAND4_in[1] ), .A2(n585), 
        .A3(\SB2_3_22/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_22/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[59] ) );
  NAND4_X1 U1051 ( .A1(\SB2_3_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_8/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_8/Component_Function_5/NAND4_in[0] ), .ZN(n1661) );
  BUF_X1 U1056 ( .A(\RI3[3][19] ), .Z(\SB2_3_28/i0[6] ) );
  BUF_X2 U1058 ( .A(\RI1[3][116] ), .Z(\SB1_3_12/i1[9] ) );
  BUF_X2 U1075 ( .A(\RI1[3][171] ), .Z(\SB1_3_3/i0[8] ) );
  CLKBUF_X3 U1081 ( .A(\RI5[2][32] ), .Z(n1511) );
  BUF_X2 U1087 ( .A(\RI3[2][159] ), .Z(\SB2_2_5/i0[10] ) );
  NAND4_X1 U1088 ( .A1(\SB1_2_7/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_7/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_7/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_7/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[2][174] ) );
  BUF_X2 U1104 ( .A(\RI1[2][50] ), .Z(\SB1_2_23/i1[9] ) );
  INV_X1 U1105 ( .A(\RI1[2][120] ), .ZN(\SB1_2_11/i0[9] ) );
  BUF_X2 U1107 ( .A(\RI5[1][103] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[103] ) );
  BUF_X2 U1108 ( .A(\RI5[1][144] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[144] ) );
  BUF_X2 U1109 ( .A(\RI5[1][157] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[157] ) );
  AND2_X1 U1123 ( .A1(\RI3[1][172] ), .A2(\RI3[1][168] ), .ZN(n1556) );
  INV_X1 U1126 ( .A(\RI1[1][66] ), .ZN(\SB1_1_20/i0[9] ) );
  BUF_X2 U1133 ( .A(\RI5[0][42] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[42] ) );
  NAND4_X1 U1152 ( .A1(\SB2_0_16/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_0_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_16/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_0_16/Component_Function_5/NAND4_in[0] ), .ZN(n875) );
  BUF_X2 U1162 ( .A(\RI3[0][158] ), .Z(\SB2_0_5/i0_0 ) );
  BUF_X1 U1163 ( .A(n117), .Z(\SB1_0_19/i0[8] ) );
  INV_X1 U1188 ( .A(n42), .ZN(\SB1_0_6/i0[9] ) );
  BUF_X1 U1197 ( .A(n171), .Z(\SB1_0_28/i0[8] ) );
  BUF_X1 U1213 ( .A(n81), .Z(\SB1_0_13/i0[8] ) );
  BUF_X1 U1221 ( .A(n136), .Z(\SB1_0_22/i1[9] ) );
  INV_X1 U1224 ( .A(n12), .ZN(\SB1_0_1/i0[9] ) );
  INV_X1 U1244 ( .A(n44), .ZN(\SB1_0_7/i0_4 ) );
  CLKBUF_X1 U1245 ( .A(n47), .Z(\SB1_0_7/i1_7 ) );
  INV_X1 U1246 ( .A(n158), .ZN(\SB1_0_26/i0_4 ) );
  CLKBUF_X1 U1247 ( .A(n163), .Z(\SB1_0_27/i1_5 ) );
  BUF_X1 U1249 ( .A(\RI3[0][180] ), .Z(\SB2_0_1/i0[9] ) );
  NAND4_X1 U1251 ( .A1(n1230), .A2(\SB2_0_1/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_1/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_1/Component_Function_5/NAND4_in[0] ), .ZN(n795) );
  BUF_X1 U1262 ( .A(\RI3[1][66] ), .Z(\SB2_1_20/i0[9] ) );
  BUF_X1 U1282 ( .A(\RI3[1][60] ), .Z(\SB2_1_21/i0[9] ) );
  BUF_X1 U1287 ( .A(\RI3[1][90] ), .Z(\SB2_1_16/i0[9] ) );
  BUF_X1 U1289 ( .A(\RI3[1][102] ), .Z(\SB2_1_14/i0[9] ) );
  BUF_X1 U1291 ( .A(\RI3[1][0] ), .Z(\SB2_1_31/i0[9] ) );
  NAND4_X1 U1294 ( .A1(\SB2_1_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_13/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_13/Component_Function_5/NAND4_in[0] ), .ZN(n808) );
  XNOR2_X1 U1295 ( .A(n807), .B(n493), .ZN(\MC_ARK_ARC_1_1/temp4[77] ) );
  CLKBUF_X1 U1297 ( .A(\RI1[2][91] ), .Z(\SB1_2_16/i1_7 ) );
  BUF_X1 U1313 ( .A(\RI3[2][138] ), .Z(\SB2_2_8/i0[9] ) );
  INV_X1 U1314 ( .A(\RI3[2][27] ), .ZN(\SB2_2_27/i0[8] ) );
  NAND4_X1 U1337 ( .A1(\SB1_2_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_4/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_4/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_4/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[2][0] ) );
  BUF_X1 U1352 ( .A(\RI3[2][60] ), .Z(\SB2_2_21/i0[9] ) );
  XNOR2_X1 U1353 ( .A(n846), .B(n512), .ZN(\MC_ARK_ARC_1_2/temp4[5] ) );
  CLKBUF_X1 U1358 ( .A(\RI1[3][25] ), .Z(\SB1_3_27/i1_7 ) );
  CLKBUF_X1 U1361 ( .A(\RI1[3][52] ), .Z(\SB1_3_23/i0[7] ) );
  AND4_X1 U1362 ( .A1(\SB1_3_27/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_27/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_27/Component_Function_5/NAND4_in[0] ), .A4(n1389), .ZN(n1630)
         );
  XNOR2_X1 U1364 ( .A(\MC_ARK_ARC_1_3/buf_datainput[137] ), .B(
        \MC_ARK_ARC_1_1/buf_keyinput[189] ), .ZN(\MC_ARK_ARC_1_3/temp4[101] )
         );
  BUF_X1 U1365 ( .A(\RI1[4][9] ), .Z(\SB3_30/i0[8] ) );
  CLKBUF_X1 U1366 ( .A(\RI1[4][78] ), .Z(\SB3_18/i3[0] ) );
  CLKBUF_X1 U1374 ( .A(\RI1[4][112] ), .Z(\SB3_13/i0[7] ) );
  CLKBUF_X1 U1375 ( .A(\RI1[4][160] ), .Z(\SB3_5/i0[7] ) );
  INV_X1 U1399 ( .A(n453), .ZN(n332) );
  INV_X1 U1400 ( .A(n495), .ZN(n275) );
  INV_X1 U1417 ( .A(n475), .ZN(n333) );
  INV_X1 U1430 ( .A(n492), .ZN(n257) );
  INV_X1 U1444 ( .A(n375), .ZN(n325) );
  INV_X1 U1448 ( .A(\MC_ARK_ARC_1_2/buf_keyinput[107] ), .ZN(n258) );
  INV_X1 U1449 ( .A(n390), .ZN(n290) );
  INV_X1 U1454 ( .A(n379), .ZN(n361) );
  INV_X1 U1455 ( .A(Key[145]), .ZN(n238) );
  INV_X1 U1458 ( .A(n487), .ZN(n242) );
  INV_X1 U1460 ( .A(n404), .ZN(n313) );
  INV_X1 U1461 ( .A(Key[18]), .ZN(n357) );
  INV_X1 U1475 ( .A(n490), .ZN(n291) );
  AND4_X1 U1476 ( .A1(\SB3_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_4/NAND4_in[3] ), .ZN(n1512) );
  AND4_X1 U1477 ( .A1(\SB1_3_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_4/NAND4_in[3] ), .ZN(n1513) );
  INV_X1 U1478 ( .A(\MC_ARK_ARC_1_1/buf_keyinput[125] ), .ZN(n354) );
  INV_X1 U1481 ( .A(Key[31]), .ZN(n344) );
  NAND4_X1 U1491 ( .A1(\SB1_1_4/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_4/Component_Function_4/NAND4_in[3] ), .A4(n1514), .ZN(
        \RI3[1][172] ) );
  NAND3_X1 U1494 ( .A1(n2149), .A2(\SB1_1_4/i0[10] ), .A3(\SB1_1_4/i0[9] ), 
        .ZN(n1514) );
  NAND4_X1 U1495 ( .A1(n663), .A2(\SB3_24/Component_Function_3/NAND4_in[1] ), 
        .A3(\SB3_24/Component_Function_3/NAND4_in[2] ), .A4(n1515), .ZN(
        \RI3[4][57] ) );
  NAND3_X1 U1499 ( .A1(\SB3_24/i1[9] ), .A2(\SB3_24/i0[6] ), .A3(n872), .ZN(
        n1515) );
  NAND4_X1 U1500 ( .A1(\SB3_10/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_5/NAND4_in[0] ), .A4(n1516), .ZN(
        \RI3[4][131] ) );
  NAND3_X1 U1501 ( .A1(\SB3_10/i0_3 ), .A2(\SB3_10/i1[9] ), .A3(\SB3_10/i0_4 ), 
        .ZN(n1516) );
  NAND4_X1 U1502 ( .A1(\SB2_2_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_16/Component_Function_3/NAND4_in[1] ), .A4(n1517), .ZN(
        \RI5[2][105] ) );
  NAND3_X1 U1503 ( .A1(\SB2_2_16/i3[0] ), .A2(\SB2_2_16/i1_5 ), .A3(
        \SB2_2_16/i0[8] ), .ZN(n1517) );
  XNOR2_X1 U1504 ( .A(\MC_ARK_ARC_1_3/temp6[43] ), .B(n1518), .ZN(\RI1[4][43] ) );
  XNOR2_X1 U1506 ( .A(\MC_ARK_ARC_1_3/temp2[43] ), .B(
        \MC_ARK_ARC_1_3/temp1[43] ), .ZN(n1518) );
  XNOR2_X1 U1507 ( .A(\MC_ARK_ARC_1_3/temp5[92] ), .B(n1519), .ZN(\RI1[4][92] ) );
  XNOR2_X1 U1511 ( .A(\MC_ARK_ARC_1_3/temp3[92] ), .B(
        \MC_ARK_ARC_1_3/temp4[92] ), .ZN(n1519) );
  NAND4_X2 U1513 ( .A1(\SB2_3_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_3_13/Component_Function_2/NAND4_in[2] ), .A3(n1520), .A4(
        \SB2_3_13/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[128] ) );
  NAND3_X1 U1530 ( .A1(\SB2_3_13/i0_0 ), .A2(\SB2_3_13/i1_5 ), .A3(
        \SB2_3_13/i0_4 ), .ZN(n1520) );
  XNOR2_X1 U1562 ( .A(n1522), .B(n347), .ZN(Ciphertext[129]) );
  NAND4_X1 U1565 ( .A1(n1909), .A2(\SB4_10/Component_Function_3/NAND4_in[0] ), 
        .A3(n1880), .A4(\SB4_10/Component_Function_3/NAND4_in[3] ), .ZN(n1522)
         );
  INV_X1 U1567 ( .A(\RI1[4][124] ), .ZN(\SB3_11/i0_4 ) );
  XNOR2_X1 U1571 ( .A(\MC_ARK_ARC_1_3/temp5[124] ), .B(
        \MC_ARK_ARC_1_3/temp6[124] ), .ZN(\RI1[4][124] ) );
  NAND4_X1 U1572 ( .A1(\SB1_0_27/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_27/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_0_27/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_0_27/Component_Function_4/NAND4_in[1] ), .ZN(\RI3[0][34] ) );
  NAND3_X1 U1610 ( .A1(n2141), .A2(\SB1_1_11/i0[10] ), .A3(\SB1_1_11/i0_4 ), 
        .ZN(\SB1_1_11/Component_Function_0/NAND4_in[2] ) );
  NAND4_X4 U1611 ( .A1(\SB2_1_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_3/NAND4_in[2] ), .A3(n1032), .A4(n1232), 
        .ZN(\MC_ARK_ARC_1_1/buf_datainput[69] ) );
  NAND4_X2 U1628 ( .A1(\SB2_2_31/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_31/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[15] ) );
  NAND3_X1 U1629 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i1[9] ), .A3(
        \SB2_2_7/i0[6] ), .ZN(\SB2_2_7/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U1630 ( .A1(\SB4_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_24/Component_Function_3/NAND4_in[3] ), .A4(n1523), .ZN(
        \RI4[4][45] ) );
  NAND3_X1 U1637 ( .A1(\SB4_24/i0[10] ), .A2(\SB4_24/i1[9] ), .A3(
        \SB4_24/i1_7 ), .ZN(n1523) );
  XNOR2_X1 U1671 ( .A(n1524), .B(n345), .ZN(Ciphertext[47]) );
  NAND4_X1 U1686 ( .A1(\SB4_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_24/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_24/Component_Function_5/NAND4_in[0] ), .ZN(n1524) );
  NAND4_X1 U1687 ( .A1(\SB1_3_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_31/Component_Function_5/NAND4_in[0] ), .A4(n1525), .ZN(
        \RI3[3][5] ) );
  NAND3_X1 U1688 ( .A1(\SB1_3_31/i1[9] ), .A2(\SB1_3_31/i0_3 ), .A3(
        \SB1_3_31/i0_4 ), .ZN(n1525) );
  NAND4_X1 U1703 ( .A1(\SB1_2_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_2/NAND4_in[2] ), .A4(n1526), .ZN(
        \RI3[2][98] ) );
  NAND3_X1 U1704 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i0_4 ), .A3(
        \SB1_2_18/i1_5 ), .ZN(n1526) );
  NAND4_X2 U1705 ( .A1(\SB2_0_31/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_31/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[15] ) );
  NAND3_X1 U1726 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i1_7 ), .A3(\SB4_7/i0[8] ), 
        .ZN(n1527) );
  NAND4_X1 U1732 ( .A1(\SB1_1_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_7/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_1_7/Component_Function_3/NAND4_in[0] ), .A4(n1529), .ZN(
        \RI3[1][159] ) );
  NAND3_X1 U1759 ( .A1(\SB1_1_7/i1[9] ), .A2(\SB1_1_7/i0[10] ), .A3(
        \SB1_1_7/i1_7 ), .ZN(n1529) );
  NAND3_X1 U1771 ( .A1(\SB2_1_5/i0_4 ), .A2(\SB2_1_5/i1_7 ), .A3(
        \SB2_1_5/i0[8] ), .ZN(\SB2_1_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1772 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i0[10] ), .A3(n805), .ZN(
        \SB4_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1774 ( .A1(\SB1_3_7/i1[9] ), .A2(\SB1_3_7/i0[10] ), .A3(
        \SB1_3_7/i1_7 ), .ZN(\SB1_3_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1775 ( .A1(\SB2_0_10/i0_3 ), .A2(\SB2_0_10/i0[9] ), .A3(
        \SB2_0_10/i0[10] ), .ZN(\SB2_0_10/Component_Function_4/NAND4_in[2] )
         );
  NAND4_X1 U1776 ( .A1(\SB1_1_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_3/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_1_3/Component_Function_5/NAND4_in[0] ), .A4(n1530), .ZN(
        \RI3[1][173] ) );
  NAND3_X1 U1777 ( .A1(\SB1_1_3/i0_4 ), .A2(\SB1_1_3/i0[9] ), .A3(
        \SB1_1_3/i0[6] ), .ZN(n1530) );
  NAND3_X1 U1791 ( .A1(\SB2_1_6/i0_4 ), .A2(\RI3[1][150] ), .A3(
        \SB2_1_6/i0[6] ), .ZN(\SB2_1_6/Component_Function_5/NAND4_in[3] ) );
  NAND4_X1 U1792 ( .A1(\SB2_2_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_24/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_24/Component_Function_2/NAND4_in[1] ), .A4(n1531), .ZN(
        \RI5[2][62] ) );
  NAND3_X1 U1799 ( .A1(\SB2_2_24/i0_0 ), .A2(\SB2_2_24/i0_4 ), .A3(
        \SB2_2_24/i1_5 ), .ZN(n1531) );
  NAND4_X2 U1805 ( .A1(\SB2_0_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_7/Component_Function_3/NAND4_in[0] ), .A3(n1174), .A4(
        \SB2_0_7/Component_Function_3/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[159] ) );
  NAND3_X1 U1816 ( .A1(\SB2_0_6/i0_4 ), .A2(\SB2_0_6/i0_0 ), .A3(
        \SB2_0_6/i1_5 ), .ZN(\SB2_0_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1817 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i0_4 ), .A3(
        \SB1_2_27/i1_5 ), .ZN(n1157) );
  NAND3_X1 U1818 ( .A1(\SB2_2_21/i0[10] ), .A2(\SB2_2_21/i0_0 ), .A3(
        \SB2_2_21/i0[6] ), .ZN(\SB2_2_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1824 ( .A1(\SB1_2_15/i1[9] ), .A2(\SB1_2_15/i0_3 ), .A3(
        \SB1_2_15/i0_4 ), .ZN(n603) );
  NAND3_X1 U1826 ( .A1(\SB2_0_7/i0_4 ), .A2(\SB2_0_7/i0_3 ), .A3(
        \SB2_0_7/i0_0 ), .ZN(\SB2_0_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1829 ( .A1(\SB2_1_18/i0[10] ), .A2(\SB2_1_18/i0_0 ), .A3(
        \SB2_1_18/i0[6] ), .ZN(\SB2_1_18/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U1830 ( .A1(\SB2_0_0/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_0/Component_Function_3/NAND4_in[0] ), .A3(n1692), .A4(n1532), 
        .ZN(\RI5[0][9] ) );
  NAND3_X1 U1831 ( .A1(\SB2_0_0/i3[0] ), .A2(\SB2_0_0/i1_5 ), .A3(
        \SB2_0_0/i0[8] ), .ZN(n1532) );
  NAND3_X1 U1845 ( .A1(\SB2_1_5/i0[8] ), .A2(\SB2_1_5/i1_5 ), .A3(
        \SB2_1_5/i3[0] ), .ZN(\SB2_1_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1846 ( .A1(\SB2_3_3/i0_3 ), .A2(\SB2_3_3/i0[9] ), .A3(
        \SB2_3_3/i0[10] ), .ZN(\SB2_3_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1850 ( .A1(\SB2_0_13/i0[9] ), .A2(\SB2_0_13/i0_3 ), .A3(
        \SB2_0_13/i0[10] ), .ZN(\SB2_0_13/Component_Function_4/NAND4_in[2] )
         );
  XNOR2_X1 U1851 ( .A(n1533), .B(n414), .ZN(Ciphertext[76]) );
  NAND4_X1 U1852 ( .A1(\SB4_19/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_19/Component_Function_4/NAND4_in[3] ), .A3(
        \SB4_19/Component_Function_4/NAND4_in[0] ), .A4(n1860), .ZN(n1533) );
  NAND4_X1 U1853 ( .A1(\SB1_3_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_3/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_3/Component_Function_5/NAND4_in[0] ), .A4(n1534), .ZN(
        \RI3[3][173] ) );
  NAND3_X1 U1866 ( .A1(\SB1_3_3/i1[9] ), .A2(\SB1_3_3/i0_3 ), .A3(
        \SB1_3_3/i0_4 ), .ZN(n1534) );
  OR3_X1 U1868 ( .A1(\RI1[2][151] ), .A2(\RI1[2][152] ), .A3(\RI1[2][153] ), 
        .ZN(\SB1_2_6/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1869 ( .A1(\SB1_2_12/i1[9] ), .A2(\SB1_2_12/i0_3 ), .A3(
        \SB1_2_12/i0_4 ), .ZN(\SB1_2_12/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U1871 ( .A1(\SB2_1_28/i0_0 ), .A2(\SB2_1_28/i3[0] ), .ZN(n1535) );
  OR3_X1 U1874 ( .A1(\RI1[2][116] ), .A2(\RI1[2][115] ), .A3(\RI1[2][117] ), 
        .ZN(\SB1_2_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1875 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i0_4 ), .A3(\SB4_19/i0_3 ), 
        .ZN(\SB4_19/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U1881 ( .A1(\SB2_1_24/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_24/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_24/Component_Function_2/NAND4_in[1] ), .A4(n1536), .ZN(
        \RI5[1][62] ) );
  NAND3_X1 U1890 ( .A1(\SB2_1_24/i0_4 ), .A2(\SB2_1_24/i0_0 ), .A3(
        \SB2_1_24/i1_5 ), .ZN(n1536) );
  NAND4_X4 U1896 ( .A1(\SB2_0_11/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_11/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_11/Component_Function_1/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[145] ) );
  NAND3_X1 U1938 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0_4 ), .A3(
        \SB1_0_29/i0[10] ), .ZN(\SB1_0_29/Component_Function_0/NAND4_in[2] )
         );
  NAND3_X1 U1946 ( .A1(\SB3_11/i0[8] ), .A2(\SB3_11/i1_7 ), .A3(\SB3_11/i0_4 ), 
        .ZN(\SB3_11/Component_Function_1/NAND4_in[3] ) );
  XNOR2_X1 U1966 ( .A(n1538), .B(\MC_ARK_ARC_1_3/temp6[37] ), .ZN(\RI1[4][37] ) );
  XNOR2_X1 U1980 ( .A(\MC_ARK_ARC_1_3/temp1[37] ), .B(
        \MC_ARK_ARC_1_3/temp2[37] ), .ZN(n1538) );
  XNOR2_X1 U1993 ( .A(n1539), .B(n217), .ZN(Ciphertext[39]) );
  NAND4_X1 U1994 ( .A1(\SB4_25/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_25/Component_Function_3/NAND4_in[0] ), .A3(n1757), .A4(
        \SB4_25/Component_Function_3/NAND4_in[3] ), .ZN(n1539) );
  NAND3_X1 U1995 ( .A1(\SB2_2_5/i0_4 ), .A2(\SB2_2_5/i0_0 ), .A3(
        \SB2_2_5/i0_3 ), .ZN(\SB2_2_5/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2000 ( .A(\MC_ARK_ARC_1_1/temp6[158] ), .B(n1540), .ZN(
        \RI1[2][158] ) );
  XNOR2_X1 U2001 ( .A(\MC_ARK_ARC_1_1/temp2[158] ), .B(
        \MC_ARK_ARC_1_1/temp1[158] ), .ZN(n1540) );
  XNOR2_X1 U2003 ( .A(n1541), .B(n223), .ZN(Ciphertext[93]) );
  NAND4_X1 U2004 ( .A1(\SB4_16/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_16/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_16/Component_Function_3/NAND4_in[3] ), .ZN(n1541) );
  NAND3_X1 U2023 ( .A1(\SB2_1_21/i0[9] ), .A2(\SB2_1_21/i0_3 ), .A3(
        \SB2_1_21/i0[10] ), .ZN(\SB2_1_21/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2038 ( .A1(\SB3_25/i0_3 ), .A2(\SB3_25/i1[9] ), .A3(\SB3_25/i0_4 ), 
        .ZN(\SB3_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2039 ( .A1(\SB2_1_4/i0[10] ), .A2(\SB2_1_4/i0_0 ), .A3(
        \SB2_1_4/i0[6] ), .ZN(\SB2_1_4/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2040 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i0[7] ), .A3(
        \SB1_1_26/i0_0 ), .ZN(\SB1_1_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2042 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i1_5 ), .A3(
        \SB2_2_7/i0_4 ), .ZN(\SB2_2_7/Component_Function_2/NAND4_in[3] ) );
  NAND4_X4 U2043 ( .A1(\SB2_3_5/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_5/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_5/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_3_5/Component_Function_2/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[176] ) );
  NAND3_X1 U2053 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i1_5 ), .A3(\SB4_10/i0_4 ), 
        .ZN(n1542) );
  NAND4_X1 U2075 ( .A1(\SB4_26/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_26/Component_Function_4/NAND4_in[3] ), .A3(n744), .A4(n1543), 
        .ZN(n1160) );
  NAND3_X1 U2083 ( .A1(\SB4_26/i0_0 ), .A2(\SB4_26/i0[8] ), .A3(\SB4_26/i0[9] ), .ZN(n1543) );
  NAND4_X1 U2095 ( .A1(\SB4_4/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_4/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_4/Component_Function_2/NAND4_in[0] ), .A4(n1544), .ZN(n1798) );
  NAND3_X1 U2097 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i0_4 ), .A3(\SB4_4/i1_5 ), 
        .ZN(n1544) );
  NAND3_X1 U2106 ( .A1(\SB4_26/i0[6] ), .A2(\SB4_26/i0[8] ), .A3(
        \SB4_26/i0[7] ), .ZN(n1545) );
  XNOR2_X1 U2113 ( .A(n1546), .B(n222), .ZN(Ciphertext[52]) );
  NAND4_X1 U2119 ( .A1(\SB4_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB4_23/Component_Function_4/NAND4_in[2] ), .A3(
        \SB4_23/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_23/Component_Function_4/NAND4_in[1] ), .ZN(n1546) );
  XNOR2_X1 U2127 ( .A(n1547), .B(n207), .ZN(Ciphertext[13]) );
  NAND4_X1 U2128 ( .A1(\SB4_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_29/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_29/Component_Function_1/NAND4_in[0] ), .A4(n1296), .ZN(n1547) );
  NAND3_X1 U2136 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i1_5 ), .A3(
        \SB4_26/i1[9] ), .ZN(n1548) );
  NAND4_X1 U2137 ( .A1(\SB2_3_0/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_0/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_0/Component_Function_2/NAND4_in[1] ), .A4(n1549), .ZN(
        \RI5[3][14] ) );
  NAND3_X1 U2138 ( .A1(\SB2_3_0/i0_4 ), .A2(\SB2_3_0/i0_0 ), .A3(
        \SB2_3_0/i1_5 ), .ZN(n1549) );
  NAND4_X1 U2145 ( .A1(\SB4_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_4/Component_Function_3/NAND4_in[3] ), .A4(n1550), .ZN(n732) );
  NAND3_X1 U2146 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i1[9] ), .A3(\SB4_4/i1_7 ), 
        .ZN(n1550) );
  XNOR2_X1 U2147 ( .A(n1551), .B(n228), .ZN(Ciphertext[106]) );
  NAND4_X2 U2160 ( .A1(\SB2_3_18/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_18/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_18/Component_Function_2/NAND4_in[1] ), .A4(n1552), .ZN(
        \RI5[3][98] ) );
  NAND3_X1 U2164 ( .A1(\SB2_3_18/i0_0 ), .A2(\SB2_3_18/i1_5 ), .A3(
        \SB2_3_18/i0_4 ), .ZN(n1552) );
  NAND4_X1 U2183 ( .A1(\SB1_3_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_17/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_17/Component_Function_5/NAND4_in[0] ), .A4(n1554), .ZN(
        \RI3[3][89] ) );
  NAND3_X1 U2184 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i0[9] ), .A3(
        \SB1_3_17/i0[6] ), .ZN(n1554) );
  NAND4_X4 U2185 ( .A1(n1166), .A2(\SB2_3_0/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_3_0/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[191] ) );
  NAND2_X1 U2197 ( .A1(\SB2_1_3/i0[6] ), .A2(n1556), .ZN(n1555) );
  NAND3_X1 U2198 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i0[10] ), .A3(\SB4_4/i0[6] ), 
        .ZN(\SB4_4/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U2202 ( .A(n1557), .B(n276), .ZN(Ciphertext[85]) );
  NAND4_X1 U2203 ( .A1(\SB4_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_17/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_17/Component_Function_1/NAND4_in[0] ), .ZN(n1557) );
  NAND3_X1 U2209 ( .A1(\SB2_2_10/i0_4 ), .A2(\SB2_2_10/i1_5 ), .A3(
        \SB2_2_10/i1[9] ), .ZN(n1558) );
  XNOR2_X1 U2221 ( .A(n1559), .B(n236), .ZN(Ciphertext[50]) );
  NAND4_X1 U2222 ( .A1(n591), .A2(\SB4_23/Component_Function_2/NAND4_in[2] ), 
        .A3(\SB4_23/Component_Function_2/NAND4_in[0] ), .A4(
        \SB4_23/Component_Function_2/NAND4_in[1] ), .ZN(n1559) );
  XNOR2_X1 U2235 ( .A(n1560), .B(n303), .ZN(Ciphertext[122]) );
  NAND4_X1 U2244 ( .A1(\SB4_11/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_11/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_11/Component_Function_2/NAND4_in[0] ), .A4(n1039), .ZN(n1560) );
  XNOR2_X1 U2247 ( .A(n1562), .B(n1561), .ZN(\RI1[1][53] ) );
  XNOR2_X1 U2255 ( .A(\MC_ARK_ARC_1_0/temp4[53] ), .B(
        \MC_ARK_ARC_1_0/temp1[53] ), .ZN(n1561) );
  XNOR2_X1 U2259 ( .A(\MC_ARK_ARC_1_0/temp2[53] ), .B(
        \MC_ARK_ARC_1_0/temp3[53] ), .ZN(n1562) );
  NAND3_X1 U2268 ( .A1(\SB4_9/i0_3 ), .A2(\SB4_9/i0[9] ), .A3(\SB4_9/i0[10] ), 
        .ZN(n1563) );
  NAND3_X1 U2294 ( .A1(\SB2_3_21/i0_0 ), .A2(\SB2_3_21/i3[0] ), .A3(
        \SB2_3_21/i1_7 ), .ZN(\SB2_3_21/Component_Function_4/NAND4_in[1] ) );
  XNOR2_X1 U2307 ( .A(n1564), .B(n290), .ZN(Ciphertext[124]) );
  NAND4_X1 U2308 ( .A1(\SB4_11/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_11/Component_Function_4/NAND4_in[0] ), .A3(n1287), .A4(
        \SB4_11/Component_Function_4/NAND4_in[1] ), .ZN(n1564) );
  NAND3_X1 U2309 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0[8] ), .A3(\SB4_16/i0[9] ), .ZN(n932) );
  XNOR2_X1 U2310 ( .A(n1565), .B(n342), .ZN(Ciphertext[116]) );
  NAND4_X1 U2332 ( .A1(\SB4_12/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_12/Component_Function_2/NAND4_in[2] ), .A3(n1893), .A4(
        \SB4_12/Component_Function_2/NAND4_in[0] ), .ZN(n1565) );
  NAND4_X1 U2357 ( .A1(\SB3_27/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_27/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_27/Component_Function_5/NAND4_in[0] ), .A4(n1566), .ZN(
        \RI3[4][29] ) );
  NAND3_X1 U2371 ( .A1(\SB3_27/i1[9] ), .A2(\SB3_27/i0_3 ), .A3(\SB3_27/i0_4 ), 
        .ZN(n1566) );
  XNOR2_X1 U2380 ( .A(\MC_ARK_ARC_1_3/temp6[26] ), .B(n1567), .ZN(\RI1[4][26] ) );
  XNOR2_X1 U2382 ( .A(\MC_ARK_ARC_1_3/temp1[26] ), .B(
        \MC_ARK_ARC_1_3/temp2[26] ), .ZN(n1567) );
  NAND4_X1 U2398 ( .A1(\SB3_15/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_15/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_2/NAND4_in[0] ), .A4(n1569), .ZN(
        \RI3[4][116] ) );
  NAND3_X1 U2408 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i1_5 ), .A3(\SB3_15/i0_4 ), 
        .ZN(n1569) );
  NAND4_X1 U2421 ( .A1(\SB1_3_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_20/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_3_20/Component_Function_1/NAND4_in[2] ), .A4(n1570), .ZN(
        \RI3[3][91] ) );
  NAND3_X1 U2429 ( .A1(\SB1_3_20/i0[8] ), .A2(\SB1_3_20/i1_7 ), .A3(
        \SB1_3_20/i0_4 ), .ZN(n1570) );
  NAND3_X1 U2431 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0_4 ), .A3(\SB4_24/i1[9] ), 
        .ZN(\SB4_24/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U2439 ( .A(\MC_ARK_ARC_1_2/temp5[39] ), .B(n1571), .ZN(\RI1[3][39] ) );
  XNOR2_X1 U2440 ( .A(\MC_ARK_ARC_1_2/temp3[39] ), .B(
        \MC_ARK_ARC_1_2/temp4[39] ), .ZN(n1571) );
  NAND3_X1 U2445 ( .A1(\SB4_9/i0_0 ), .A2(\SB4_9/i1_7 ), .A3(\SB4_9/i3[0] ), 
        .ZN(n1572) );
  XNOR2_X1 U2454 ( .A(n1573), .B(n307), .ZN(Ciphertext[94]) );
  NAND4_X1 U2455 ( .A1(\SB4_16/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_16/Component_Function_4/NAND4_in[3] ), .A3(
        \SB4_16/Component_Function_4/NAND4_in[1] ), .A4(n932), .ZN(n1573) );
  NAND3_X1 U2494 ( .A1(\SB2_3_23/i0[8] ), .A2(\SB2_3_23/i3[0] ), .A3(
        \SB2_3_23/i1_5 ), .ZN(\SB2_3_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2495 ( .A1(\SB1_0_24/i0_3 ), .A2(\SB1_0_24/i1[9] ), .A3(
        \SB1_0_24/i0_4 ), .ZN(\SB1_0_24/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U2497 ( .A(\MC_ARK_ARC_1_2/temp5[71] ), .B(n1575), .ZN(\RI1[3][71] ) );
  XNOR2_X1 U2499 ( .A(\MC_ARK_ARC_1_2/temp3[71] ), .B(
        \MC_ARK_ARC_1_2/temp4[71] ), .ZN(n1575) );
  NAND3_X1 U2504 ( .A1(\SB1_0_18/i1_5 ), .A2(\SB1_0_18/i1[9] ), .A3(
        \SB1_0_18/i0_4 ), .ZN(n1576) );
  NAND4_X1 U2507 ( .A1(\SB1_3_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_30/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_30/Component_Function_5/NAND4_in[0] ), .A4(n1577), .ZN(
        \RI3[3][11] ) );
  NAND3_X1 U2525 ( .A1(\SB1_3_30/i1[9] ), .A2(\SB1_3_30/i0_3 ), .A3(
        \SB1_3_30/i0_4 ), .ZN(n1577) );
  XNOR2_X1 U2541 ( .A(\MC_ARK_ARC_1_3/temp5[113] ), .B(
        \MC_ARK_ARC_1_3/temp6[113] ), .ZN(\RI1[4][113] ) );
  NAND3_X1 U2543 ( .A1(\SB2_1_3/i0[10] ), .A2(\SB2_1_3/i1[9] ), .A3(
        \SB2_1_3/i1_7 ), .ZN(\SB2_1_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2544 ( .A1(\SB1_0_21/i0[7] ), .A2(\SB1_0_21/i0_3 ), .A3(
        \SB1_0_21/i0_0 ), .ZN(\SB1_0_21/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U2545 ( .A1(\SB1_3_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_15/Component_Function_5/NAND4_in[0] ), .A4(n1578), .ZN(
        \RI3[3][101] ) );
  NAND3_X1 U2575 ( .A1(\SB1_3_15/i1[9] ), .A2(\SB1_3_15/i0_3 ), .A3(
        \SB1_3_15/i0_4 ), .ZN(n1578) );
  NAND3_X1 U2576 ( .A1(\SB1_2_14/i1[9] ), .A2(\SB1_2_14/i0[10] ), .A3(
        \SB1_2_14/i1_7 ), .ZN(\SB1_2_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2585 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i1_5 ), .A3(
        \SB2_0_3/i1[9] ), .ZN(\SB2_0_3/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U2586 ( .A1(\SB2_3_27/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_27/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_27/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_27/Component_Function_4/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[34] ) );
  NAND3_X1 U2601 ( .A1(\SB2_2_6/i0_0 ), .A2(\RI3[2][154] ), .A3(\SB2_2_6/i1_5 ), .ZN(n1838) );
  NAND3_X1 U2603 ( .A1(\SB4_2/i0[10] ), .A2(n785), .A3(\SB4_2/i0_3 ), .ZN(
        \SB4_2/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U2619 ( .A1(\SB2_0_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_19/Component_Function_2/NAND4_in[1] ), .A4(n1579), .ZN(
        \RI5[0][92] ) );
  NAND3_X1 U2631 ( .A1(\SB2_0_19/i0_0 ), .A2(\SB2_0_19/i0_4 ), .A3(
        \SB2_0_19/i1_5 ), .ZN(n1579) );
  NAND4_X2 U2634 ( .A1(\SB2_0_4/Component_Function_3/NAND4_in[1] ), .A2(n1056), 
        .A3(n1064), .A4(n1581), .ZN(\MC_ARK_ARC_1_0/buf_datainput[177] ) );
  NAND3_X1 U2635 ( .A1(\SB2_0_4/i0[8] ), .A2(\SB2_0_4/i3[0] ), .A3(
        \SB2_0_4/i1_5 ), .ZN(n1581) );
  BUF_X2 U2647 ( .A(\RI1[3][68] ), .Z(\SB1_3_20/i1[9] ) );
  OR3_X1 U2649 ( .A1(\RI1[3][69] ), .A2(\RI1[3][67] ), .A3(\RI1[3][68] ), .ZN(
        \SB1_3_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2653 ( .A1(\SB1_1_5/i0_0 ), .A2(\SB1_1_5/i0_4 ), .A3(
        \SB1_1_5/i1_5 ), .ZN(\SB1_1_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2654 ( .A1(\SB4_22/i0_4 ), .A2(\SB4_22/i1_7 ), .A3(\SB4_22/i0[8] ), 
        .ZN(\SB4_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2676 ( .A1(\SB3_23/i0[10] ), .A2(\SB3_23/i0_3 ), .A3(
        \SB3_23/i0[9] ), .ZN(n1200) );
  NAND3_X1 U2677 ( .A1(\SB2_2_19/i0[8] ), .A2(\SB2_2_19/i1_5 ), .A3(
        \SB2_2_19/i3[0] ), .ZN(\SB2_2_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2679 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i1_5 ), .A3(\SB4_19/i0_4 ), 
        .ZN(n1614) );
  NAND3_X1 U2683 ( .A1(\SB2_1_1/i0[9] ), .A2(\SB2_1_1/i0_3 ), .A3(
        \SB2_1_1/i0[10] ), .ZN(\SB2_1_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2688 ( .A1(n1671), .A2(\SB4_26/i0_0 ), .A3(\SB4_26/i0[7] ), .ZN(
        \SB4_26/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U2689 ( .A(n1583), .B(n1582), .ZN(\RI1[2][177] ) );
  XNOR2_X1 U2692 ( .A(\MC_ARK_ARC_1_1/temp1[177] ), .B(
        \MC_ARK_ARC_1_1/temp4[177] ), .ZN(n1582) );
  XNOR2_X1 U2697 ( .A(\MC_ARK_ARC_1_1/temp3[177] ), .B(
        \MC_ARK_ARC_1_1/temp2[177] ), .ZN(n1583) );
  NAND3_X1 U2727 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i1[9] ), .A3(
        \SB2_2_23/i0[6] ), .ZN(n1584) );
  NAND3_X1 U2728 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i0[9] ), .A3(
        \SB2_2_13/i0[8] ), .ZN(\SB2_2_13/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U2743 ( .A(\MC_ARK_ARC_1_2/temp5[175] ), .B(n1585), .ZN(
        \RI1[3][175] ) );
  XNOR2_X1 U2750 ( .A(\MC_ARK_ARC_1_2/temp4[175] ), .B(
        \MC_ARK_ARC_1_2/temp3[175] ), .ZN(n1585) );
  NAND3_X1 U2751 ( .A1(\SB1_3_21/i1[9] ), .A2(\SB1_3_21/i0[10] ), .A3(
        \SB1_3_21/i1_7 ), .ZN(\SB1_3_21/Component_Function_3/NAND4_in[2] ) );
  XNOR2_X1 U2752 ( .A(n1586), .B(n262), .ZN(Ciphertext[87]) );
  NAND4_X1 U2757 ( .A1(\SB4_17/Component_Function_3/NAND4_in[0] ), .A2(n1839), 
        .A3(n1914), .A4(\SB4_17/Component_Function_3/NAND4_in[3] ), .ZN(n1586)
         );
  NAND3_X1 U2772 ( .A1(\SB2_3_12/i0[10] ), .A2(\SB2_3_12/i1[9] ), .A3(
        \SB2_3_12/i1_7 ), .ZN(\SB2_3_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2776 ( .A1(\SB2_1_11/i0_0 ), .A2(\SB2_1_11/i0[10] ), .A3(
        \SB2_1_11/i0[6] ), .ZN(\SB2_1_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2781 ( .A1(\SB4_7/i0[6] ), .A2(\SB4_7/i1[9] ), .A3(n877), .ZN(
        \SB4_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2790 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i0[10] ), .A3(
        \SB3_14/i0[6] ), .ZN(\SB3_14/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U2799 ( .A(n1588), .B(n237), .ZN(Ciphertext[91]) );
  NAND4_X1 U2801 ( .A1(\SB4_16/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_16/Component_Function_1/NAND4_in[0] ), .A3(n1299), .A4(
        \SB4_16/Component_Function_1/NAND4_in[2] ), .ZN(n1588) );
  NAND3_X1 U2822 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i0[10] ), .A3(
        \SB1_3_11/i0[9] ), .ZN(\SB1_3_11/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U2834 ( .A(n1590), .B(n211), .ZN(Ciphertext[177]) );
  NAND3_X1 U2837 ( .A1(\SB2_3_2/i0[10] ), .A2(\SB2_3_2/i1[9] ), .A3(
        \SB2_3_2/i1_7 ), .ZN(\SB2_3_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2843 ( .A1(\SB2_3_16/i0_0 ), .A2(\SB2_3_16/i1_5 ), .A3(
        \RI3[3][94] ), .ZN(\SB2_3_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2844 ( .A1(\SB4_31/i0_0 ), .A2(n1670), .A3(\SB4_31/i0_4 ), .ZN(
        \SB4_31/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2845 ( .A(n1591), .B(n297), .ZN(Ciphertext[27]) );
  NAND4_X1 U2847 ( .A1(\SB4_27/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_27/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_27/Component_Function_3/NAND4_in[3] ), .ZN(n1591) );
  NAND3_X1 U2848 ( .A1(\SB2_0_13/i0_3 ), .A2(\SB2_0_13/i0_0 ), .A3(
        \SB2_0_13/i0_4 ), .ZN(\SB2_0_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2849 ( .A1(\SB1_3_18/i1[9] ), .A2(\SB1_3_18/i0[10] ), .A3(
        \SB1_3_18/i1_7 ), .ZN(\SB1_3_18/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U2850 ( .A1(\SB3_2/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_2/Component_Function_2/NAND4_in[0] ), .A4(n1592), .ZN(\RI3[4][2] ) );
  NAND3_X1 U2852 ( .A1(\SB3_2/i0_0 ), .A2(\SB3_2/i1_5 ), .A3(\SB3_2/i0_4 ), 
        .ZN(n1592) );
  NAND4_X1 U2872 ( .A1(\SB2_3_10/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_10/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_10/Component_Function_4/NAND4_in[0] ), .A4(n1593), .ZN(
        \RI5[3][136] ) );
  NAND3_X1 U2876 ( .A1(\SB2_3_10/i0_4 ), .A2(\SB2_3_10/i1[9] ), .A3(
        \SB2_3_10/i1_5 ), .ZN(n1593) );
  NAND3_X1 U2877 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i1_5 ), .A3(\SB4_5/i1[9] ), 
        .ZN(\SB4_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2878 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0_4 ), .A3(
        \SB2_3_10/i0_0 ), .ZN(\SB2_3_10/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U2886 ( .A(n1594), .B(n1595), .ZN(\RI1[3][94] ) );
  XNOR2_X1 U2896 ( .A(\MC_ARK_ARC_1_2/temp4[94] ), .B(
        \MC_ARK_ARC_1_2/temp1[94] ), .ZN(n1594) );
  XNOR2_X1 U2900 ( .A(\MC_ARK_ARC_1_2/temp2[94] ), .B(
        \MC_ARK_ARC_1_2/temp3[94] ), .ZN(n1595) );
  NAND3_X1 U2901 ( .A1(\SB4_27/i1_5 ), .A2(\SB4_27/i3[0] ), .A3(\SB4_27/i0[8] ), .ZN(\SB4_27/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U2911 ( .A1(\SB2_2_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_26/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_26/Component_Function_4/NAND4_in[1] ), .A4(n1596), .ZN(
        \RI5[2][40] ) );
  NAND3_X1 U2912 ( .A1(\SB2_2_26/i0_4 ), .A2(\SB2_2_26/i1_5 ), .A3(
        \SB2_2_26/i1[9] ), .ZN(n1596) );
  XNOR2_X1 U2925 ( .A(n1597), .B(n212), .ZN(Ciphertext[26]) );
  NAND4_X1 U2926 ( .A1(\SB4_27/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_2/NAND4_in[1] ), .A3(n1840), .A4(n1725), 
        .ZN(n1597) );
  NAND4_X1 U2934 ( .A1(\SB2_0_9/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_0_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_4/NAND4_in[0] ), .A4(n1598), .ZN(
        \RI5[0][142] ) );
  NAND3_X1 U2935 ( .A1(\SB2_0_9/i0_4 ), .A2(\SB2_0_9/i1[9] ), .A3(
        \SB2_0_9/i1_5 ), .ZN(n1598) );
  XNOR2_X1 U2943 ( .A(\MC_ARK_ARC_1_1/temp5[188] ), .B(n1599), .ZN(
        \RI1[2][188] ) );
  XNOR2_X1 U2958 ( .A(\MC_ARK_ARC_1_1/temp3[188] ), .B(
        \MC_ARK_ARC_1_1/temp4[188] ), .ZN(n1599) );
  NAND4_X1 U2961 ( .A1(\SB2_2_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_0/Component_Function_4/NAND4_in[1] ), .A4(n1600), .ZN(
        \RI5[2][4] ) );
  NAND3_X1 U2966 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0[10] ), .A3(
        \SB2_2_0/i0[9] ), .ZN(n1600) );
  NAND4_X2 U2985 ( .A1(n1211), .A2(\SB2_3_12/Component_Function_5/NAND4_in[1] ), .A3(\SB2_3_12/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[119] ) );
  NAND3_X1 U2988 ( .A1(\SB2_2_16/i0_4 ), .A2(\SB2_2_16/i1_7 ), .A3(
        \SB2_2_16/i0[8] ), .ZN(\SB2_2_16/Component_Function_1/NAND4_in[3] ) );
  XNOR2_X1 U3049 ( .A(n1604), .B(\MC_ARK_ARC_1_3/temp6[72] ), .ZN(\RI1[4][72] ) );
  XNOR2_X1 U3055 ( .A(\MC_ARK_ARC_1_3/temp1[72] ), .B(
        \MC_ARK_ARC_1_3/temp2[72] ), .ZN(n1604) );
  NAND3_X1 U3056 ( .A1(\SB1_1_16/i0_0 ), .A2(\SB1_1_16/i0_4 ), .A3(
        \SB1_1_16/i1_5 ), .ZN(\SB1_1_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3060 ( .A1(\SB1_1_18/i0_3 ), .A2(\SB1_1_18/i0[10] ), .A3(
        \SB1_1_18/i0[9] ), .ZN(\SB1_1_18/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U3077 ( .A1(\SB2_3_7/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_3_7/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_5/NAND4_in[0] ), .A4(n1605), .ZN(
        \RI5[3][149] ) );
  NAND3_X1 U3078 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0_4 ), .A3(
        \SB2_3_7/i1[9] ), .ZN(n1605) );
  NAND3_X1 U3100 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i0[10] ), .A3(\SB3_21/i0_4 ), .ZN(\SB3_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3109 ( .A1(\SB2_3_29/i0[10] ), .A2(n2115), .A3(\SB2_3_29/i0_0 ), 
        .ZN(\SB2_3_29/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U3111 ( .A1(\SB4_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_25/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_25/Component_Function_1/NAND4_in[0] ), .A4(n1607), .ZN(n1849) );
  NAND3_X1 U3114 ( .A1(\SB4_25/i0[9] ), .A2(\SB4_25/i1_5 ), .A3(\SB4_25/i0[6] ), .ZN(n1607) );
  NAND3_X1 U3116 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i0[9] ), .A3(\SB4_6/i0[8] ), 
        .ZN(\SB4_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U3130 ( .A1(\SB2_1_17/i0_4 ), .A2(\SB2_1_17/i0_3 ), .A3(
        \SB2_1_17/i1[9] ), .ZN(\SB2_1_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3139 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0[7] ), .A3(
        \SB1_0_23/i0_0 ), .ZN(\SB1_0_23/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U3140 ( .A1(\SB1_3_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_23/i0_4 ) );
  NAND4_X1 U3148 ( .A1(\SB4_21/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_21/Component_Function_3/NAND4_in[3] ), .A3(
        \SB4_21/Component_Function_3/NAND4_in[0] ), .A4(n1608), .ZN(n1045) );
  NAND3_X1 U3163 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i1[9] ), .A3(
        \SB4_21/i1_7 ), .ZN(n1608) );
  NAND4_X1 U3179 ( .A1(\SB3_23/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_23/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_23/Component_Function_3/NAND4_in[1] ), .A4(n1609), .ZN(
        \RI3[4][63] ) );
  NAND3_X1 U3180 ( .A1(\SB3_23/i3[0] ), .A2(\SB3_23/i1_5 ), .A3(\SB3_23/i0[8] ), .ZN(n1609) );
  NAND3_X1 U3186 ( .A1(\SB2_0_30/i0_4 ), .A2(\SB2_0_30/i1[9] ), .A3(
        \SB2_0_30/i0_3 ), .ZN(\SB2_0_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3195 ( .A1(\SB2_0_31/i0[10] ), .A2(\SB2_0_31/i1_5 ), .A3(
        \SB2_0_31/i1[9] ), .ZN(\SB2_0_31/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U3196 ( .A1(\SB3_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_11/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_5/NAND4_in[0] ), .A4(n1610), .ZN(
        \RI3[4][125] ) );
  NAND3_X1 U3199 ( .A1(\SB3_11/i0[9] ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i0[6] ), .ZN(n1610) );
  NAND3_X1 U3201 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i1_5 ), .A3(\SB3_14/i0_4 ), 
        .ZN(\SB3_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3202 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i1[9] ), .A3(
        \SB4_30/i1_7 ), .ZN(\SB4_30/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U3214 ( .A1(\SB4_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_30/Component_Function_5/NAND4_in[0] ), .A4(n1611), .ZN(n1620) );
  NAND3_X1 U3218 ( .A1(\SB4_30/i0[9] ), .A2(\SB4_30/i0_4 ), .A3(\SB4_30/i0[6] ), .ZN(n1611) );
  NAND4_X1 U3223 ( .A1(\SB3_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_31/Component_Function_2/NAND4_in[1] ), .A4(n1612), .ZN(
        \RI3[4][20] ) );
  NAND3_X1 U3224 ( .A1(\SB3_31/i1_5 ), .A2(\SB3_31/i0_0 ), .A3(\SB3_31/i0_4 ), 
        .ZN(n1612) );
  NAND4_X1 U3278 ( .A1(\SB2_0_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_18/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_18/Component_Function_2/NAND4_in[1] ), .A4(n1615), .ZN(
        \RI5[0][98] ) );
  NAND3_X1 U3282 ( .A1(\SB2_0_18/i0_4 ), .A2(\SB2_0_18/i0_0 ), .A3(
        \SB2_0_18/i1_5 ), .ZN(n1615) );
  NAND3_X1 U3285 ( .A1(\SB2_2_20/i0[8] ), .A2(\SB2_2_20/i3[0] ), .A3(
        \SB2_2_20/i1_5 ), .ZN(n923) );
  NAND3_X1 U3291 ( .A1(\SB2_1_3/i0_3 ), .A2(\SB2_1_3/i1[9] ), .A3(
        \SB2_1_3/i0[6] ), .ZN(\SB2_1_3/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U3298 ( .A1(\SB3_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_15/Component_Function_5/NAND4_in[0] ), .A4(n1616), .ZN(
        \RI3[4][101] ) );
  NAND3_X1 U3303 ( .A1(\SB3_15/i1[9] ), .A2(\SB3_15/i0_3 ), .A3(\SB3_15/i0_4 ), 
        .ZN(n1616) );
  NAND3_X1 U3316 ( .A1(\SB1_3_18/i0[10] ), .A2(\SB1_3_18/i0[9] ), .A3(
        \SB1_3_18/i0_3 ), .ZN(\SB1_3_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3324 ( .A1(\SB4_31/i0_4 ), .A2(n1964), .A3(\SB4_31/i1[9] ), .ZN(
        n620) );
  NAND3_X1 U3325 ( .A1(\SB1_2_3/i1[9] ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i1_7 ), .ZN(\SB1_2_3/Component_Function_3/NAND4_in[2] ) );
  XNOR2_X1 U3334 ( .A(n1617), .B(n260), .ZN(Ciphertext[5]) );
  NAND4_X1 U3338 ( .A1(\SB4_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_31/Component_Function_5/NAND4_in[0] ), .ZN(n1617) );
  NAND4_X1 U3354 ( .A1(\SB2_2_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_1/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_1/Component_Function_1/NAND4_in[0] ), .A4(n1619), .ZN(
        \RI5[2][13] ) );
  NAND3_X1 U3355 ( .A1(\SB2_2_1/i0_4 ), .A2(\SB2_2_1/i1_7 ), .A3(
        \SB2_2_1/i0[8] ), .ZN(n1619) );
  XNOR2_X1 U3357 ( .A(n1620), .B(n221), .ZN(Ciphertext[11]) );
  NAND4_X2 U3358 ( .A1(\SB2_0_31/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_31/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_0_31/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_31/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[20] ) );
  NAND4_X2 U3360 ( .A1(\SB2_0_3/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_3/Component_Function_0/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[6] ) );
  NAND3_X1 U3361 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i3[0] ), .A3(\SB4_11/i1_7 ), 
        .ZN(\SB4_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3377 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0[10] ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3381 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i0_0 ), .A3(\SB3_7/i0[6] ), 
        .ZN(\SB3_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3405 ( .A1(\SB3_30/i0[8] ), .A2(\SB3_30/i1_7 ), .A3(\SB3_30/i0_3 ), 
        .ZN(\SB3_30/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U3406 ( .A1(\SB2_0_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_26/Component_Function_3/NAND4_in[0] ), .A3(n1777), .A4(
        \SB2_0_26/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[0][45] ) );
  NAND4_X1 U3417 ( .A1(\SB1_3_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_0/NAND4_in[3] ), .ZN(n1623) );
  NAND4_X1 U3423 ( .A1(\SB2_1_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_7/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_7/Component_Function_2/NAND4_in[1] ), .A4(n1712), .ZN(n1624) );
  CLKBUF_X1 U3439 ( .A(n121), .Z(\SB1_0_20/i1_5 ) );
  NAND4_X1 U3445 ( .A1(\SB2_3_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_7/Component_Function_2/NAND4_in[2] ), .ZN(n1626) );
  NAND4_X1 U3450 ( .A1(\SB2_3_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_7/Component_Function_2/NAND4_in[2] ), .ZN(n1627) );
  NAND4_X1 U3451 ( .A1(\SB2_3_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_7/Component_Function_2/NAND4_in[2] ), .ZN(\RI5[3][164] ) );
  BUF_X1 U3452 ( .A(\RI1[1][21] ), .Z(\SB1_1_28/i0[8] ) );
  CLKBUF_X1 U3455 ( .A(\RI1[4][82] ), .Z(\SB3_18/i0[7] ) );
  NAND4_X1 U3456 ( .A1(n1367), .A2(\SB2_2_4/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_2_4/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_4/Component_Function_5/NAND4_in[0] ), .ZN(n1628) );
  NAND4_X1 U3465 ( .A1(n1367), .A2(\SB2_2_4/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_2_4/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_4/Component_Function_5/NAND4_in[0] ), .ZN(n1629) );
  NAND4_X1 U3474 ( .A1(n1367), .A2(\SB2_2_4/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_2_4/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[167] ) );
  NAND4_X1 U3475 ( .A1(n767), .A2(\SB2_0_23/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_0_23/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_23/Component_Function_5/NAND4_in[3] ), .ZN(n1631) );
  NAND4_X1 U3480 ( .A1(n767), .A2(\SB2_0_23/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_0_23/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_23/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[53] ) );
  BUF_X1 U3486 ( .A(\RI1[4][188] ), .Z(\SB3_0/i1[9] ) );
  NAND4_X1 U3488 ( .A1(\SB2_2_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_31/Component_Function_5/NAND4_in[0] ), .ZN(n1633) );
  NAND4_X1 U3490 ( .A1(\SB2_2_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_31/Component_Function_5/NAND4_in[0] ), .ZN(n1634) );
  NAND4_X1 U3494 ( .A1(\SB2_2_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[5] ) );
  NAND4_X1 U3498 ( .A1(\SB2_2_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_5/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_5/Component_Function_5/NAND4_in[3] ), .ZN(n1635) );
  NAND4_X1 U3499 ( .A1(\SB2_2_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_5/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_5/Component_Function_5/NAND4_in[3] ), .ZN(n1636) );
  NAND4_X1 U3500 ( .A1(\SB2_2_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_5/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_5/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[161] ) );
  INV_X1 U3505 ( .A(\RI1[2][91] ), .ZN(\SB1_2_16/i0[6] ) );
  NAND4_X2 U3517 ( .A1(\SB2_0_16/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_16/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_16/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[105] ) );
  NAND4_X1 U3520 ( .A1(\SB1_3_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_1/NAND4_in[3] ), .ZN(n1637) );
  NAND4_X2 U3521 ( .A1(\SB2_3_1/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_1/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_1/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_3_1/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[3][8] ) );
  CLKBUF_X1 U3527 ( .A(\RI1[4][40] ), .Z(\SB3_25/i0[7] ) );
  CLKBUF_X1 U3545 ( .A(Key[191]), .Z(n406) );
  CLKBUF_X1 U3546 ( .A(Key[185]), .Z(n454) );
  NAND4_X2 U3553 ( .A1(\SB3_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_4/NAND4_in[3] ), .ZN(n1638) );
  CLKBUF_X1 U3554 ( .A(\RI1[4][142] ), .Z(\SB3_8/i0[7] ) );
  CLKBUF_X1 U3558 ( .A(\RI1[4][46] ), .Z(\SB3_24/i0[7] ) );
  CLKBUF_X1 U3581 ( .A(\RI1[4][70] ), .Z(\SB3_20/i0[7] ) );
  NAND4_X1 U3582 ( .A1(\SB1_3_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_0/NAND4_in[3] ), .ZN(n1639) );
  NAND4_X1 U3592 ( .A1(\SB2_1_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_31/Component_Function_5/NAND4_in[0] ), .ZN(n1640) );
  NAND4_X1 U3614 ( .A1(\SB2_1_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_31/Component_Function_5/NAND4_in[0] ), .ZN(n1641) );
  NAND4_X1 U3646 ( .A1(\SB2_1_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[5] ) );
  NAND4_X1 U3651 ( .A1(\SB2_1_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_5/NAND4_in[3] ), .A4(n563), .ZN(n1642) );
  NAND4_X1 U3652 ( .A1(\SB2_1_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_5/NAND4_in[3] ), .A4(n563), .ZN(n1643) );
  INV_X1 U3659 ( .A(\RI1[2][71] ), .ZN(n1644) );
  NAND4_X1 U3668 ( .A1(\SB2_1_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_5/NAND4_in[3] ), .A4(n563), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[17] ) );
  INV_X1 U3672 ( .A(\RI1[2][71] ), .ZN(\SB1_2_20/i0_3 ) );
  CLKBUF_X1 U3684 ( .A(\RI1[4][59] ), .Z(\SB3_22/i1_5 ) );
  NAND4_X1 U3706 ( .A1(\SB2_1_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_2/NAND4_in[1] ), .A3(n611), .A4(
        \SB2_1_21/Component_Function_2/NAND4_in[3] ), .ZN(n1645) );
  NAND4_X1 U3707 ( .A1(\SB2_1_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_2/NAND4_in[1] ), .A3(n611), .A4(
        \SB2_1_21/Component_Function_2/NAND4_in[3] ), .ZN(n1646) );
  NAND4_X1 U3708 ( .A1(\SB2_1_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_2/NAND4_in[1] ), .A3(n611), .A4(
        \SB2_1_21/Component_Function_2/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[80] ) );
  INV_X1 U3709 ( .A(\RI1[3][101] ), .ZN(n1647) );
  INV_X1 U3710 ( .A(\RI1[3][101] ), .ZN(\SB1_3_15/i0_3 ) );
  INV_X1 U3712 ( .A(\RI1[2][179] ), .ZN(n1648) );
  INV_X1 U3713 ( .A(\RI1[2][179] ), .ZN(\SB1_2_2/i0_3 ) );
  INV_X1 U3714 ( .A(\RI1[2][77] ), .ZN(n1649) );
  INV_X1 U3715 ( .A(\RI1[2][77] ), .ZN(\SB1_2_19/i0_3 ) );
  NAND4_X1 U3716 ( .A1(\SB1_3_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_4/NAND4_in[3] ), .ZN(n1651) );
  NAND4_X1 U3717 ( .A1(\SB1_3_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_4/NAND4_in[3] ), .ZN(n1652) );
  BUF_X2 U3719 ( .A(\RI5[3][23] ), .Z(n1653) );
  CLKBUF_X1 U3720 ( .A(\RI5[3][23] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[23] )
         );
  BUF_X1 U3722 ( .A(\RI1[4][155] ), .Z(\SB3_6/i1_5 ) );
  CLKBUF_X1 U3723 ( .A(\RI1[4][120] ), .Z(\SB3_11/i3[0] ) );
  NAND4_X1 U3725 ( .A1(\SB2_3_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_15/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_15/Component_Function_0/NAND4_in[2] ), .ZN(n1654) );
  NAND4_X1 U3726 ( .A1(\SB2_3_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_15/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_15/Component_Function_0/NAND4_in[2] ), .ZN(\RI5[3][126] ) );
  NAND4_X1 U3727 ( .A1(n988), .A2(\SB2_1_10/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_1_10/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_10/Component_Function_5/NAND4_in[0] ), .ZN(n1655) );
  NAND4_X1 U3728 ( .A1(n988), .A2(\SB2_1_10/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_1_10/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_10/Component_Function_5/NAND4_in[0] ), .ZN(n1656) );
  NAND4_X1 U3730 ( .A1(n988), .A2(\SB2_1_10/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_1_10/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[131] ) );
  NAND4_X1 U3732 ( .A1(\SB2_3_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_20/Component_Function_3/NAND4_in[3] ), .ZN(n1658) );
  NAND4_X1 U3733 ( .A1(\SB2_3_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_20/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][81] ) );
  NAND4_X1 U3734 ( .A1(\SB2_0_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_5/NAND4_in[3] ), .A4(n751), .ZN(n1659) );
  NAND4_X1 U3735 ( .A1(\SB2_0_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_5/NAND4_in[3] ), .A4(n751), .ZN(n1660) );
  NAND4_X1 U3736 ( .A1(\SB2_0_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_5/NAND4_in[3] ), .A4(n751), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[179] ) );
  NAND4_X1 U3738 ( .A1(\SB2_3_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_8/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_8/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[143] ) );
  CLKBUF_X1 U3739 ( .A(\SB2_3_31/i1[9] ), .Z(n1662) );
  BUF_X1 U3740 ( .A(\RI3[4][137] ), .Z(n1663) );
  BUF_X1 U3741 ( .A(\RI3[4][137] ), .Z(\SB4_9/i0_3 ) );
  INV_X1 U3742 ( .A(n49), .ZN(n1664) );
  NAND4_X1 U3743 ( .A1(\SB2_2_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_5/NAND4_in[0] ), .A4(n1866), .ZN(n1665)
         );
  NAND4_X1 U3744 ( .A1(\SB2_2_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_5/NAND4_in[0] ), .A4(n1866), .ZN(n1666)
         );
  NAND4_X1 U3745 ( .A1(\SB2_2_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_5/NAND4_in[0] ), .A4(n1866), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[107] ) );
  BUF_X1 U3746 ( .A(\RI3[4][167] ), .Z(n1667) );
  BUF_X1 U3747 ( .A(\RI3[4][167] ), .Z(\SB4_4/i0_3 ) );
  BUF_X1 U3748 ( .A(\RI3[4][11] ), .Z(n1668) );
  BUF_X1 U3749 ( .A(\RI3[4][11] ), .Z(\SB4_30/i0_3 ) );
  INV_X1 U3750 ( .A(\RI1[4][5] ), .ZN(n1669) );
  NAND4_X1 U3751 ( .A1(\SB3_31/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_5/NAND4_in[3] ), .ZN(n1670) );
  BUF_X1 U3752 ( .A(\RI3[4][35] ), .Z(n1671) );
  BUF_X1 U3753 ( .A(\RI3[4][35] ), .Z(\SB4_26/i0_3 ) );
  BUF_X1 U3754 ( .A(\RI3[4][191] ), .Z(n1672) );
  BUF_X1 U3755 ( .A(\RI3[4][191] ), .Z(\SB4_0/i0_3 ) );
  NAND3_X1 U3757 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0_4 ), .A3(
        \SB1_0_23/i1[9] ), .ZN(n1673) );
  NAND3_X1 U3759 ( .A1(\SB2_0_24/i0_4 ), .A2(\SB2_0_24/i0_3 ), .A3(
        \SB2_0_24/i1[9] ), .ZN(\SB2_0_24/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3760 ( .A1(\SB2_0_22/i0_4 ), .A2(\SB2_0_22/i0_0 ), .A3(
        \SB2_0_22/i1_5 ), .ZN(n1674) );
  NAND4_X2 U3762 ( .A1(\SB2_1_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_24/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_24/Component_Function_5/NAND4_in[1] ), .A4(n1755), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[47] ) );
  NAND3_X1 U3763 ( .A1(\SB1_2_27/i0_3 ), .A2(\SB1_2_27/i0[10] ), .A3(
        \SB1_2_27/i0[9] ), .ZN(\SB1_2_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3764 ( .A1(n1639), .A2(\SB2_3_8/i0[8] ), .A3(\SB2_3_8/i0_3 ), .ZN(
        \SB2_3_8/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U3765 ( .A1(\SB2_0_24/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_24/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_24/Component_Function_4/NAND4_in[0] ), .A4(n1675), .ZN(
        \RI5[0][52] ) );
  NAND3_X1 U3766 ( .A1(\SB2_0_24/i0_4 ), .A2(\SB2_0_24/i1_5 ), .A3(
        \SB2_0_24/i1[9] ), .ZN(n1675) );
  INV_X2 U3767 ( .A(\RI1[3][65] ), .ZN(\SB1_3_21/i0_3 ) );
  XNOR2_X1 U3768 ( .A(\MC_ARK_ARC_1_2/temp6[65] ), .B(
        \MC_ARK_ARC_1_2/temp5[65] ), .ZN(\RI1[3][65] ) );
  NAND3_X1 U3769 ( .A1(\SB2_0_18/i0[6] ), .A2(\SB2_0_18/i0[9] ), .A3(
        \SB2_0_18/i0_4 ), .ZN(\SB2_0_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3770 ( .A1(\SB2_0_12/i0_3 ), .A2(\SB2_0_12/i1[9] ), .A3(
        \SB2_0_12/i0[6] ), .ZN(\SB2_0_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3772 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i0_0 ), .A3(
        \SB1_1_9/i0[6] ), .ZN(\SB1_1_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3773 ( .A1(\SB2_0_26/i0_0 ), .A2(\SB2_0_26/i0[7] ), .A3(
        \SB2_0_26/i0_3 ), .ZN(\SB2_0_26/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U3775 ( .A1(n1742), .A2(\SB2_2_21/Component_Function_2/NAND4_in[1] ), .A3(\SB2_2_21/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_2_21/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[80] ) );
  NAND4_X1 U3776 ( .A1(\SB2_2_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_4/Component_Function_4/NAND4_in[1] ), .A4(n1676), .ZN(
        \RI5[2][172] ) );
  NAND3_X1 U3777 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0[9] ), .A3(
        \SB2_2_4/i0[10] ), .ZN(n1676) );
  NAND4_X1 U3778 ( .A1(\SB2_2_1/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_1/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_1/Component_Function_4/NAND4_in[1] ), .A4(n1677), .ZN(
        \RI5[2][190] ) );
  NAND3_X1 U3779 ( .A1(\SB2_2_1/i0_4 ), .A2(\SB2_2_1/i1_5 ), .A3(
        \SB2_2_1/i1[9] ), .ZN(n1677) );
  NAND3_X1 U3780 ( .A1(\SB2_2_1/i0_0 ), .A2(\RI3[2][184] ), .A3(\SB2_2_1/i1_5 ), .ZN(n587) );
  NAND3_X1 U3781 ( .A1(\SB2_0_1/i0_4 ), .A2(\SB2_0_1/i0_0 ), .A3(
        \SB2_0_1/i1_5 ), .ZN(n568) );
  NAND3_X1 U3782 ( .A1(\SB2_0_14/i0[10] ), .A2(\SB2_0_14/i1_5 ), .A3(
        \SB2_0_14/i1[9] ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U3783 ( .A(\RI1[2][167] ), .ZN(\SB1_2_4/i0_3 ) );
  XNOR2_X1 U3784 ( .A(\MC_ARK_ARC_1_1/temp5[167] ), .B(
        \MC_ARK_ARC_1_1/temp6[167] ), .ZN(\RI1[2][167] ) );
  XNOR2_X1 U3785 ( .A(n922), .B(n1678), .ZN(\RI1[1][27] ) );
  XNOR2_X1 U3786 ( .A(\MC_ARK_ARC_1_0/temp3[27] ), .B(
        \MC_ARK_ARC_1_0/temp4[27] ), .ZN(n1678) );
  NAND4_X2 U3787 ( .A1(\SB2_0_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_7/Component_Function_5/NAND4_in[1] ), .A4(n1679), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[149] ) );
  NAND2_X1 U3788 ( .A1(\SB2_0_7/i0_0 ), .A2(\SB2_0_7/i3[0] ), .ZN(n1679) );
  XNOR2_X1 U3789 ( .A(n1680), .B(n1815), .ZN(\RI1[3][80] ) );
  XNOR2_X1 U3790 ( .A(\MC_ARK_ARC_1_2/temp3[80] ), .B(
        \MC_ARK_ARC_1_2/temp2[80] ), .ZN(n1680) );
  NAND4_X1 U3791 ( .A1(\SB1_1_25/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_25/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_25/Component_Function_5/NAND4_in[0] ), .A4(n1681), .ZN(
        \RI3[1][41] ) );
  NAND3_X1 U3792 ( .A1(\SB1_1_25/i1[9] ), .A2(\SB1_1_25/i0_3 ), .A3(
        \SB1_1_25/i0_4 ), .ZN(n1681) );
  NAND3_X1 U3793 ( .A1(\SB1_1_28/i0_0 ), .A2(\SB1_1_28/i0_4 ), .A3(
        \SB1_1_28/i1_5 ), .ZN(n1845) );
  XNOR2_X1 U3794 ( .A(n1682), .B(\MC_ARK_ARC_1_2/temp6[44] ), .ZN(\RI1[3][44] ) );
  XNOR2_X1 U3795 ( .A(\MC_ARK_ARC_1_2/temp2[44] ), .B(
        \MC_ARK_ARC_1_2/temp1[44] ), .ZN(n1682) );
  NAND2_X1 U3796 ( .A1(\SB2_0_23/i0[9] ), .A2(\SB2_0_23/i0[10] ), .ZN(
        \SB2_0_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3797 ( .A1(\SB2_2_16/i0_0 ), .A2(\SB2_2_16/i0[10] ), .A3(
        \RI3[2][91] ), .ZN(\SB2_2_16/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U3798 ( .A1(\SB2_1_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_14/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_1_14/Component_Function_4/NAND4_in[1] ), .A4(n1683), .ZN(
        \RI5[1][112] ) );
  NAND3_X1 U3799 ( .A1(\SB2_1_14/i0_4 ), .A2(\SB2_1_14/i1_5 ), .A3(
        \SB2_1_14/i1[9] ), .ZN(n1683) );
  NAND3_X1 U3800 ( .A1(\SB1_1_17/i0[9] ), .A2(\SB1_1_17/i0[8] ), .A3(
        \SB1_1_17/i0_3 ), .ZN(\SB1_1_17/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U3801 ( .A(\MC_ARK_ARC_1_0/buf_datainput[84] ), .B(
        \MC_ARK_ARC_1_0/buf_datainput[78] ), .ZN(\MC_ARK_ARC_1_0/temp1[84] )
         );
  NAND4_X2 U3802 ( .A1(\SB2_0_23/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_23/Component_Function_0/NAND4_in[3] ), .A3(n1709), .A4(
        \SB2_0_23/Component_Function_0/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[78] ) );
  NAND3_X1 U3803 ( .A1(\SB3_26/i0_3 ), .A2(\SB3_26/i1[9] ), .A3(\SB3_26/i0_4 ), 
        .ZN(n1688) );
  XNOR2_X1 U3805 ( .A(n1685), .B(n1684), .ZN(\RI1[1][71] ) );
  XNOR2_X1 U3806 ( .A(\MC_ARK_ARC_1_0/temp2[71] ), .B(
        \MC_ARK_ARC_1_0/temp4[71] ), .ZN(n1684) );
  XNOR2_X1 U3807 ( .A(\MC_ARK_ARC_1_0/temp1[71] ), .B(
        \MC_ARK_ARC_1_0/temp3[71] ), .ZN(n1685) );
  NAND2_X1 U3808 ( .A1(\SB2_2_11/i0[6] ), .A2(n1686), .ZN(
        \SB2_2_11/Component_Function_5/NAND4_in[3] ) );
  AND2_X1 U3809 ( .A1(\RI3[2][120] ), .A2(\RI3[2][124] ), .ZN(n1686) );
  NAND3_X1 U3812 ( .A1(\SB2_0_30/i0_4 ), .A2(\SB2_0_30/i1[9] ), .A3(
        \SB2_0_30/i1_5 ), .ZN(n1687) );
  NAND4_X1 U3813 ( .A1(\SB3_26/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_26/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_26/Component_Function_5/NAND4_in[0] ), .A4(n1688), .ZN(
        \RI3[4][35] ) );
  NAND3_X1 U3814 ( .A1(\SB1_3_7/i0[8] ), .A2(\SB1_3_7/i1_7 ), .A3(
        \SB1_3_7/i0_4 ), .ZN(\SB1_3_7/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 U3815 ( .A1(\SB2_0_0/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_0/Component_Function_4/NAND4_in[2] ), .A4(n1689), .ZN(
        \RI5[0][4] ) );
  NAND4_X2 U3819 ( .A1(n1222), .A2(\SB2_0_26/Component_Function_4/NAND4_in[0] ), .A3(\SB2_0_26/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_0_26/Component_Function_4/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[40] ) );
  NAND4_X1 U3820 ( .A1(\SB1_1_4/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_4/Component_Function_2/NAND4_in[2] ), .A4(n1691), .ZN(
        \RI3[1][182] ) );
  NAND3_X1 U3821 ( .A1(\SB1_1_4/i0_4 ), .A2(\SB1_1_4/i0_0 ), .A3(
        \SB1_1_4/i1_5 ), .ZN(n1691) );
  NAND3_X1 U3822 ( .A1(\SB2_3_7/i0_4 ), .A2(\SB2_3_7/i0[9] ), .A3(
        \SB2_3_7/i0[6] ), .ZN(\SB2_3_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3823 ( .A1(\SB1_2_18/i1[9] ), .A2(\SB1_2_18/i1_7 ), .A3(
        \SB1_2_18/i0[10] ), .ZN(\SB1_2_18/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U3824 ( .A1(\SB2_0_0/i0_4 ), .A2(\SB2_0_0/i0_0 ), .A3(
        \SB2_0_0/i0_3 ), .ZN(n1692) );
  NAND3_X1 U3825 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0[9] ), .A3(
        \SB1_3_8/i0[10] ), .ZN(\SB1_3_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3826 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0[10] ), .A3(
        \SB1_0_21/i0[9] ), .ZN(\SB1_0_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3827 ( .A1(\SB2_0_25/i0_4 ), .A2(\SB2_0_25/i0_3 ), .A3(
        \SB2_0_25/i1[9] ), .ZN(n1399) );
  NAND3_X1 U3828 ( .A1(\SB1_1_24/i0_4 ), .A2(\SB1_1_24/i0_0 ), .A3(
        \SB1_1_24/i1_5 ), .ZN(n1729) );
  NAND3_X1 U3829 ( .A1(\SB2_1_1/i0_0 ), .A2(\SB2_1_1/i0[10] ), .A3(
        \SB2_1_1/i0[6] ), .ZN(\SB2_1_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3830 ( .A1(\SB2_0_29/i0[10] ), .A2(\SB2_0_29/i1_5 ), .A3(
        \SB2_0_29/i1[9] ), .ZN(\SB2_0_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3831 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3832 ( .A1(\SB2_2_15/i0_0 ), .A2(\SB2_2_15/i0[10] ), .A3(
        \SB2_2_15/i0[6] ), .ZN(\SB2_2_15/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U3833 ( .A1(\SB2_0_23/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_23/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_0_23/Component_Function_2/NAND4_in[1] ), .A4(n1693), .ZN(
        \RI5[0][68] ) );
  NAND3_X1 U3834 ( .A1(\SB2_0_23/i0_0 ), .A2(\SB2_0_23/i1_5 ), .A3(
        \SB2_0_23/i0_4 ), .ZN(n1693) );
  NAND4_X1 U3835 ( .A1(\SB2_1_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_17/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_1_17/Component_Function_5/NAND4_in[1] ), .A4(n1694), .ZN(
        \RI5[1][89] ) );
  NAND3_X1 U3836 ( .A1(\SB2_1_17/i0[9] ), .A2(\SB2_1_17/i0_4 ), .A3(
        \SB2_1_17/i0[6] ), .ZN(n1694) );
  NAND3_X1 U3837 ( .A1(\SB1_0_26/i0[7] ), .A2(\SB1_0_26/i0_3 ), .A3(
        \SB1_0_26/i0_0 ), .ZN(\SB1_0_26/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U3841 ( .A(\MC_ARK_ARC_1_0/temp1[47] ), .B(
        \MC_ARK_ARC_1_0/temp4[47] ), .ZN(n1696) );
  XNOR2_X1 U3842 ( .A(\MC_ARK_ARC_1_0/temp3[47] ), .B(
        \MC_ARK_ARC_1_0/temp2[47] ), .ZN(n1697) );
  NAND3_X1 U3843 ( .A1(\SB1_2_10/i1[9] ), .A2(\SB1_2_10/i0[10] ), .A3(
        \SB1_2_10/i1_7 ), .ZN(\SB1_2_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3844 ( .A1(\SB1_3_20/i0_0 ), .A2(\SB1_3_20/i0_4 ), .A3(
        \SB1_3_20/i1_5 ), .ZN(n762) );
  NAND4_X1 U3845 ( .A1(\SB1_2_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_22/Component_Function_4/NAND4_in[3] ), .A4(n1698), .ZN(
        \RI3[2][64] ) );
  NAND3_X1 U3846 ( .A1(\SB1_2_22/i0_3 ), .A2(\SB1_2_22/i0[10] ), .A3(
        \SB1_2_22/i0[9] ), .ZN(n1698) );
  NAND4_X1 U3848 ( .A1(\SB2_3_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_24/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_5/NAND4_in[0] ), .A4(n1700), .ZN(
        \RI5[3][47] ) );
  NAND3_X1 U3849 ( .A1(\SB2_3_24/i0_4 ), .A2(\RI3[3][42] ), .A3(
        \SB2_3_24/i0[6] ), .ZN(n1700) );
  NAND3_X1 U3850 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i1[9] ), .A3(
        \SB1_3_24/i1_7 ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3853 ( .A1(\SB1_1_16/i1[9] ), .A2(\SB1_1_16/i0[10] ), .A3(
        \SB1_1_16/i1_7 ), .ZN(\SB1_1_16/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U3854 ( .A1(n676), .A2(\SB2_2_2/Component_Function_4/NAND4_in[2] ), 
        .A3(\SB2_2_2/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_2/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[184] ) );
  INV_X2 U3855 ( .A(\RI1[1][143] ), .ZN(\SB1_1_8/i0_3 ) );
  XNOR2_X1 U3856 ( .A(\MC_ARK_ARC_1_0/temp5[143] ), .B(
        \MC_ARK_ARC_1_0/temp6[143] ), .ZN(\RI1[1][143] ) );
  NAND3_X1 U3857 ( .A1(\SB2_0_12/i0_4 ), .A2(\SB2_0_12/i0_0 ), .A3(
        \SB2_0_12/i1_5 ), .ZN(\SB2_0_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3859 ( .A1(\SB2_3_3/i0_3 ), .A2(\SB2_3_3/i0_4 ), .A3(
        \SB2_3_3/i1[9] ), .ZN(n1702) );
  NAND4_X2 U3860 ( .A1(\SB2_0_20/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_20/Component_Function_2/NAND4_in[1] ), .A3(n885), .A4(n1703), 
        .ZN(\MC_ARK_ARC_1_0/buf_datainput[86] ) );
  NAND3_X1 U3861 ( .A1(\SB2_0_20/i0[10] ), .A2(\SB2_0_20/i1[9] ), .A3(
        \SB2_0_20/i1_5 ), .ZN(n1703) );
  OR3_X1 U3862 ( .A1(\RI1[1][92] ), .A2(\RI1[1][93] ), .A3(\RI1[1][91] ), .ZN(
        \SB1_1_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3863 ( .A1(\SB2_0_1/i0[9] ), .A2(\SB2_0_1/i0_3 ), .A3(
        \SB2_0_1/i0[8] ), .ZN(\SB2_0_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3864 ( .A1(\SB1_1_20/i0[9] ), .A2(\SB1_1_20/i1_5 ), .A3(
        \SB1_1_20/i0[6] ), .ZN(\SB1_1_20/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U3865 ( .A1(\SB2_1_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_7/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_7/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[149] ) );
  NAND3_X1 U3867 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i1[9] ), .A3(
        \SB2_0_6/i0_4 ), .ZN(n1444) );
  NAND3_X1 U3868 ( .A1(\SB1_1_10/i1_5 ), .A2(\SB1_1_10/i0_0 ), .A3(
        \SB1_1_10/i0_4 ), .ZN(n1734) );
  XNOR2_X1 U3869 ( .A(\MC_ARK_ARC_1_1/temp6[120] ), .B(
        \MC_ARK_ARC_1_1/temp5[120] ), .ZN(\RI1[2][120] ) );
  NAND3_X1 U3870 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0[10] ), .A3(
        \SB2_0_16/i0[9] ), .ZN(n1704) );
  NAND4_X1 U3871 ( .A1(\SB1_0_16/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_16/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_0_16/Component_Function_5/NAND4_in[3] ), .A4(n1705), .ZN(
        \RI3[0][95] ) );
  NAND3_X1 U3872 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0_4 ), .A3(
        \SB1_0_16/i1[9] ), .ZN(n1705) );
  NAND4_X2 U3873 ( .A1(\SB2_2_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_11/Component_Function_5/NAND4_in[1] ), .A3(n668), .A4(
        \SB2_2_11/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[125] ) );
  NAND3_X1 U3874 ( .A1(\SB2_0_20/i0[9] ), .A2(\SB2_0_20/i0_4 ), .A3(
        \SB2_0_20/i0[6] ), .ZN(n1263) );
  NAND4_X4 U3875 ( .A1(\SB2_1_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_7/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_7/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[159] ) );
  NAND3_X1 U3876 ( .A1(\SB2_2_13/i0_0 ), .A2(\SB2_2_13/i3[0] ), .A3(
        \SB2_2_13/i1_7 ), .ZN(n1706) );
  NAND3_X1 U3877 ( .A1(\SB2_0_3/i0[6] ), .A2(\SB2_0_3/i0_0 ), .A3(
        \SB2_0_3/i0[10] ), .ZN(\SB2_0_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3880 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0[10] ), .A3(
        \SB1_2_21/i0_4 ), .ZN(\SB1_2_21/Component_Function_0/NAND4_in[2] ) );
  XNOR2_X1 U3882 ( .A(\MC_ARK_ARC_1_0/temp5[66] ), .B(
        \MC_ARK_ARC_1_0/temp6[66] ), .ZN(\RI1[1][66] ) );
  NAND3_X1 U3885 ( .A1(\SB2_0_8/i0_3 ), .A2(\SB2_0_8/i0_0 ), .A3(
        \SB2_0_8/i0[7] ), .ZN(\SB2_0_8/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U3886 ( .A(\MC_ARK_ARC_1_0/buf_datainput[131] ), .B(n875), .ZN(
        \MC_ARK_ARC_1_0/temp3[29] ) );
  NAND3_X1 U3887 ( .A1(\SB1_3_29/i0[10] ), .A2(\SB1_3_29/i1[9] ), .A3(
        \SB1_3_29/i1_7 ), .ZN(\SB1_3_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3888 ( .A1(\SB1_2_22/i1[9] ), .A2(\SB1_2_22/i0[10] ), .A3(
        \SB1_2_22/i1_7 ), .ZN(\SB1_2_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3889 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i0[10] ), .A3(
        \SB2_0_23/i0_4 ), .ZN(n1709) );
  NAND3_X1 U3890 ( .A1(\SB2_3_27/i0[10] ), .A2(\SB2_3_27/i0_0 ), .A3(
        \SB2_3_27/i0[6] ), .ZN(\SB2_3_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3891 ( .A1(\SB2_0_3/i0[7] ), .A2(\SB2_0_3/i0_0 ), .A3(
        \SB2_0_3/i0_3 ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3892 ( .A1(\SB1_1_9/i0[9] ), .A2(\SB1_1_9/i1_5 ), .A3(
        \SB1_1_9/i0[6] ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3893 ( .A1(\SB1_1_29/i0[9] ), .A2(\SB1_1_29/i1_5 ), .A3(
        \SB1_1_29/i0[6] ), .ZN(\SB1_1_29/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U3894 ( .A1(\SB1_0_4/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_4/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_4/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_0_4/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_0_3/i0_4 ) );
  NAND3_X1 U3897 ( .A1(n826), .A2(\SB1_1_10/i0[10] ), .A3(\SB1_1_10/i0_4 ), 
        .ZN(\SB1_1_10/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U3898 ( .A1(\SB2_1_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_5/Component_Function_5/NAND4_in[1] ), .A3(n1711), .A4(n586), 
        .ZN(\MC_ARK_ARC_1_1/buf_datainput[161] ) );
  NAND3_X1 U3899 ( .A1(\SB2_1_5/i0_4 ), .A2(\SB2_1_5/i0[9] ), .A3(
        \SB2_1_5/i0[6] ), .ZN(n1711) );
  NAND3_X1 U3900 ( .A1(\SB2_1_7/i0_0 ), .A2(\SB2_1_7/i0_4 ), .A3(
        \SB2_1_7/i1_5 ), .ZN(n1712) );
  NAND3_X1 U3903 ( .A1(\SB1_2_20/i1_7 ), .A2(\SB1_2_20/i0_4 ), .A3(
        \SB1_2_20/i0[8] ), .ZN(\SB1_2_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3904 ( .A1(\SB1_3_9/i0_3 ), .A2(\SB1_3_9/i1[9] ), .A3(
        \SB1_3_9/i0[6] ), .ZN(\SB1_3_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3905 ( .A1(\SB1_1_18/i0_4 ), .A2(\SB1_1_18/i1[9] ), .A3(
        \SB1_1_18/i1_5 ), .ZN(\SB1_1_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3906 ( .A1(\SB1_2_17/i0_3 ), .A2(\SB1_2_17/i0_0 ), .A3(
        \SB1_2_17/i0_4 ), .ZN(\SB1_2_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3907 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0[7] ), .A3(
        \SB1_1_14/i0_0 ), .ZN(\SB1_1_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3909 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i0_0 ), .A3(
        \SB2_0_23/i0_4 ), .ZN(n1714) );
  NAND3_X1 U3911 ( .A1(\SB2_0_28/i0_4 ), .A2(\SB2_0_28/i0[9] ), .A3(
        \SB2_0_28/i0[6] ), .ZN(\SB2_0_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3913 ( .A1(\SB2_2_15/i0[9] ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i0[8] ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3914 ( .A1(\SB2_1_7/i0[9] ), .A2(\SB2_1_7/i0[10] ), .A3(
        \SB2_1_7/i0_3 ), .ZN(\SB2_1_7/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U3915 ( .A(n1715), .B(\MC_ARK_ARC_1_0/temp5[158] ), .ZN(
        \RI1[1][158] ) );
  XNOR2_X1 U3916 ( .A(\MC_ARK_ARC_1_0/temp4[158] ), .B(
        \MC_ARK_ARC_1_0/temp3[158] ), .ZN(n1715) );
  NAND4_X1 U3919 ( .A1(\SB1_1_1/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_1/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_1/Component_Function_2/NAND4_in[2] ), .A4(n1717), .ZN(
        \RI3[1][8] ) );
  NAND3_X1 U3920 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i0_4 ), .A3(
        \SB1_1_1/i1_5 ), .ZN(n1717) );
  NAND2_X1 U3921 ( .A1(\SB2_1_20/i0_0 ), .A2(\SB2_1_20/i3[0] ), .ZN(n1718) );
  NAND4_X1 U3922 ( .A1(\SB4_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_13/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_13/Component_Function_2/NAND4_in[3] ), .A4(n1719), .ZN(n1393) );
  NAND3_X1 U3923 ( .A1(\SB4_13/i0[10] ), .A2(\SB4_13/i1_5 ), .A3(
        \SB4_13/i1[9] ), .ZN(n1719) );
  NAND4_X1 U3924 ( .A1(\SB4_13/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_13/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_13/Component_Function_3/NAND4_in[3] ), .A4(n1720), .ZN(n557) );
  NAND3_X1 U3925 ( .A1(\SB4_13/i0[10] ), .A2(\SB4_13/i1[9] ), .A3(
        \SB4_13/i1_7 ), .ZN(n1720) );
  NAND4_X1 U3926 ( .A1(\SB2_1_6/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_6/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_6/Component_Function_3/NAND4_in[3] ), .A4(n1721), .ZN(
        \RI5[1][165] ) );
  NAND3_X1 U3927 ( .A1(\SB2_1_6/i0[10] ), .A2(\SB2_1_6/i1_7 ), .A3(
        \SB2_1_6/i1[9] ), .ZN(n1721) );
  NAND4_X1 U3928 ( .A1(\SB1_2_31/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_31/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_31/Component_Function_1/NAND4_in[0] ), .A4(n1722), .ZN(
        \RI3[2][25] ) );
  NAND3_X1 U3929 ( .A1(\SB1_2_31/i0[8] ), .A2(\SB1_2_31/i1_7 ), .A3(
        \SB1_2_31/i0_4 ), .ZN(n1722) );
  NAND3_X1 U3930 ( .A1(\SB4_30/i0[9] ), .A2(\SB4_30/i1_5 ), .A3(\SB4_30/i0[6] ), .ZN(\SB4_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3931 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i0[7] ), .A3(\SB3_12/i0_0 ), 
        .ZN(\SB3_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3932 ( .A1(\SB2_2_28/i0_0 ), .A2(\SB2_2_28/i3[0] ), .A3(
        \SB2_2_28/i1_7 ), .ZN(\SB2_2_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3933 ( .A1(\SB2_0_18/i1_7 ), .A2(\SB2_0_18/i3[0] ), .A3(
        \SB2_0_18/i0_0 ), .ZN(\SB2_0_18/Component_Function_4/NAND4_in[1] ) );
  NAND4_X1 U3934 ( .A1(\SB1_3_12/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_12/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_12/Component_Function_1/NAND4_in[0] ), .A4(n1723), .ZN(
        \RI3[3][139] ) );
  NAND3_X1 U3935 ( .A1(\SB1_3_12/i1_7 ), .A2(\SB1_3_12/i0_4 ), .A3(
        \SB1_3_12/i0[8] ), .ZN(n1723) );
  NAND3_X1 U3936 ( .A1(\SB2_2_16/i0[6] ), .A2(\SB2_2_16/i0_4 ), .A3(
        \SB2_2_16/i0[9] ), .ZN(\SB2_2_16/Component_Function_5/NAND4_in[3] ) );
  NAND4_X1 U3937 ( .A1(\SB1_1_27/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_27/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_27/Component_Function_2/NAND4_in[2] ), .A4(n1724), .ZN(
        \RI3[1][44] ) );
  NAND3_X1 U3938 ( .A1(\SB1_1_27/i0_0 ), .A2(\SB1_1_27/i0_4 ), .A3(
        \SB1_1_27/i1_5 ), .ZN(n1724) );
  NAND3_X1 U3939 ( .A1(\SB4_27/i0_0 ), .A2(\SB4_27/i1_5 ), .A3(n780), .ZN(
        n1725) );
  NAND3_X1 U3940 ( .A1(\SB4_27/i0_0 ), .A2(\SB4_27/i3[0] ), .A3(\SB4_27/i1_7 ), 
        .ZN(\SB4_27/Component_Function_4/NAND4_in[1] ) );
  NAND4_X1 U3941 ( .A1(\SB3_30/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_30/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_30/Component_Function_2/NAND4_in[2] ), .A4(n1726), .ZN(
        \RI3[4][26] ) );
  NAND3_X1 U3942 ( .A1(\SB3_30/i0_0 ), .A2(\SB3_30/i1_5 ), .A3(\SB3_30/i0_4 ), 
        .ZN(n1726) );
  NAND4_X2 U3943 ( .A1(n680), .A2(\SB2_3_16/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB2_3_16/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_3_16/Component_Function_2/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[110] ) );
  XNOR2_X1 U3944 ( .A(n1727), .B(n323), .ZN(Ciphertext[23]) );
  NAND4_X1 U3945 ( .A1(\SB4_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_28/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_28/Component_Function_5/NAND4_in[0] ), .ZN(n1727) );
  NAND4_X1 U3946 ( .A1(\SB4_28/Component_Function_3/NAND4_in[3] ), .A2(
        \SB4_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_28/Component_Function_3/NAND4_in[0] ), .A4(n1728), .ZN(n1289) );
  NAND3_X1 U3947 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i1[9] ), .A3(
        \SB4_28/i1_7 ), .ZN(n1728) );
  NAND3_X1 U3948 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i1[9] ), .A3(
        \SB2_0_20/i0[6] ), .ZN(\SB2_0_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3949 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[8] ), .A3(
        \SB2_2_16/i0[9] ), .ZN(\SB2_2_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3951 ( .A1(\SB2_0_3/i0_4 ), .A2(\SB2_0_3/i1[9] ), .A3(
        \SB2_0_3/i1_5 ), .ZN(\SB2_0_3/Component_Function_4/NAND4_in[3] ) );
  NAND4_X1 U3952 ( .A1(\SB1_1_24/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_24/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_24/Component_Function_2/NAND4_in[2] ), .A4(n1729), .ZN(
        \RI3[1][62] ) );
  NAND4_X2 U3953 ( .A1(\SB2_1_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_12/Component_Function_5/NAND4_in[1] ), .A4(n566), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[119] ) );
  XNOR2_X1 U3954 ( .A(\MC_ARK_ARC_1_0/temp5[179] ), .B(n1730), .ZN(
        \RI1[1][179] ) );
  XNOR2_X1 U3955 ( .A(\MC_ARK_ARC_1_0/temp3[179] ), .B(
        \MC_ARK_ARC_1_0/temp4[179] ), .ZN(n1730) );
  XNOR2_X1 U3958 ( .A(\MC_ARK_ARC_1_0/temp3[41] ), .B(
        \MC_ARK_ARC_1_0/temp2[41] ), .ZN(n1732) );
  NAND4_X1 U3960 ( .A1(\SB2_0_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_14/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_14/Component_Function_2/NAND4_in[1] ), .A4(n1733), .ZN(
        \RI5[0][122] ) );
  NAND3_X1 U3961 ( .A1(\SB2_0_14/i0_0 ), .A2(\SB2_0_14/i0_4 ), .A3(
        \SB2_0_14/i1_5 ), .ZN(n1733) );
  NAND4_X1 U3962 ( .A1(\SB1_1_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_2/NAND4_in[2] ), .A4(n1734), .ZN(
        \RI3[1][146] ) );
  NAND3_X1 U3963 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0_4 ), .A3(
        \SB1_0_7/i1[9] ), .ZN(\SB1_0_7/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U3964 ( .A1(\SB2_1_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_14/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_14/Component_Function_1/NAND4_in[0] ), .A4(n1735), .ZN(
        \RI5[1][127] ) );
  NAND3_X1 U3965 ( .A1(\SB2_1_14/i0_4 ), .A2(\SB2_1_14/i1_7 ), .A3(
        \SB2_1_14/i0[8] ), .ZN(n1735) );
  NAND3_X1 U3966 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i0[10] ), .A3(
        \SB1_1_21/i0[9] ), .ZN(\SB1_1_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3967 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i0_0 ), .A3(
        \SB1_1_28/i0_4 ), .ZN(\SB1_1_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3968 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i1_5 ), .A3(
        \SB2_1_9/i1[9] ), .ZN(\SB2_1_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3969 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i0_3 ), .A3(
        \SB1_3_3/i0[9] ), .ZN(\SB1_3_3/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U3970 ( .A1(\SB2_1_0/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_0/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_0/Component_Function_2/NAND4_in[1] ), .A4(n1736), .ZN(
        \RI5[1][14] ) );
  NAND3_X1 U3971 ( .A1(\SB2_1_0/i0_4 ), .A2(\SB2_1_0/i1_5 ), .A3(
        \SB2_1_0/i0_0 ), .ZN(n1736) );
  NAND3_X1 U3972 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0[10] ), .A3(
        \SB1_0_29/i0[9] ), .ZN(\SB1_0_29/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U3973 ( .A(n1738), .B(n1737), .ZN(\RI1[2][71] ) );
  XNOR2_X1 U3974 ( .A(\MC_ARK_ARC_1_1/temp2[71] ), .B(
        \MC_ARK_ARC_1_1/temp4[71] ), .ZN(n1737) );
  XNOR2_X1 U3975 ( .A(\MC_ARK_ARC_1_1/temp3[71] ), .B(
        \MC_ARK_ARC_1_1/temp1[71] ), .ZN(n1738) );
  NAND4_X1 U3976 ( .A1(\SB1_3_25/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_25/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_25/Component_Function_5/NAND4_in[0] ), .A4(n1739), .ZN(
        \RI3[3][41] ) );
  NAND3_X1 U3977 ( .A1(\SB1_3_25/i1[9] ), .A2(\SB1_3_25/i0_4 ), .A3(
        \SB1_3_25/i0_3 ), .ZN(n1739) );
  NAND4_X1 U3978 ( .A1(\SB2_2_19/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_19/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_19/Component_Function_4/NAND4_in[1] ), .A4(n1740), .ZN(
        \RI5[2][82] ) );
  NAND3_X1 U3979 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0[10] ), .A3(
        \SB2_2_19/i0[9] ), .ZN(n1740) );
  NAND4_X1 U3980 ( .A1(\SB2_0_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_28/Component_Function_2/NAND4_in[1] ), .A4(n1741), .ZN(
        \RI5[0][38] ) );
  NAND3_X1 U3981 ( .A1(\SB2_0_28/i0_4 ), .A2(\SB2_0_28/i1_5 ), .A3(
        \SB2_0_28/i0_0 ), .ZN(n1741) );
  NAND3_X1 U3983 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0[6] ), .A3(
        \SB2_0_21/i1[9] ), .ZN(\SB2_0_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3984 ( .A1(\SB2_2_21/i0[9] ), .A2(\SB2_2_21/i0_3 ), .A3(
        \SB2_2_21/i0[8] ), .ZN(n1742) );
  NAND3_X1 U3985 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0_4 ), .A3(
        \SB2_2_4/i1[9] ), .ZN(n1367) );
  NAND3_X1 U3986 ( .A1(\SB1_2_28/i1[9] ), .A2(\SB1_2_28/i0[10] ), .A3(
        \SB1_2_28/i1_7 ), .ZN(\SB1_2_28/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U3987 ( .A1(\SB1_1_8/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_8/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_1_7/i0_4 ) );
  XNOR2_X1 U3988 ( .A(n1744), .B(n1743), .ZN(\RI1[2][191] ) );
  XNOR2_X1 U3989 ( .A(\MC_ARK_ARC_1_1/temp1[191] ), .B(
        \MC_ARK_ARC_1_1/temp4[191] ), .ZN(n1743) );
  XNOR2_X1 U3990 ( .A(\MC_ARK_ARC_1_1/temp2[191] ), .B(
        \MC_ARK_ARC_1_1/temp3[191] ), .ZN(n1744) );
  NAND3_X1 U3991 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i1[9] ), .A3(
        \SB2_2_2/i1_5 ), .ZN(n676) );
  NAND3_X1 U3992 ( .A1(\SB1_1_0/i0_0 ), .A2(\SB1_1_0/i1_5 ), .A3(
        \SB1_1_0/i0_4 ), .ZN(\SB1_1_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3997 ( .A1(\SB2_0_7/i0[10] ), .A2(\SB2_0_7/i1_5 ), .A3(
        \SB2_0_7/i1[9] ), .ZN(\SB2_0_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3998 ( .A1(\SB1_0_9/i0[10] ), .A2(\SB1_0_9/i0_3 ), .A3(
        \SB1_0_9/i0[9] ), .ZN(\SB1_0_9/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U3999 ( .A1(n1386), .A2(\SB2_0_8/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_8/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_8/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[143] ) );
  NAND4_X1 U4000 ( .A1(\SB2_3_30/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_3_30/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_30/Component_Function_2/NAND4_in[1] ), .A4(n1747), .ZN(
        \RI5[3][26] ) );
  NAND3_X1 U4001 ( .A1(\SB2_3_30/i0[9] ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB2_3_30/i0[8] ), .ZN(n1747) );
  XNOR2_X1 U4003 ( .A(n1749), .B(n232), .ZN(Ciphertext[78]) );
  NAND4_X1 U4004 ( .A1(\SB4_18/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_18/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_18/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_18/Component_Function_0/NAND4_in[0] ), .ZN(n1749) );
  NAND4_X1 U4005 ( .A1(\SB3_3/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_3/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_3/Component_Function_2/NAND4_in[0] ), .A4(n1750), .ZN(
        \RI3[4][188] ) );
  NAND3_X1 U4006 ( .A1(\SB3_3/i0_0 ), .A2(\SB3_3/i0_4 ), .A3(\SB3_3/i1_5 ), 
        .ZN(n1750) );
  NAND3_X1 U4007 ( .A1(n809), .A2(\SB1_3_0/i0[10] ), .A3(\SB1_3_0/i0_4 ), .ZN(
        \SB1_3_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4008 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0[6] ), .A3(
        \SB2_2_1/i0[10] ), .ZN(\SB2_2_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U4009 ( .A1(\SB2_0_5/i0[9] ), .A2(\SB2_0_5/i0_3 ), .A3(
        \SB2_0_5/i0[8] ), .ZN(\SB2_0_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4010 ( .A1(\SB2_0_6/i0[9] ), .A2(\SB2_0_6/i0_4 ), .A3(
        \SB2_0_6/i0[6] ), .ZN(\SB2_0_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4011 ( .A1(\SB2_0_0/i0[10] ), .A2(\SB2_0_0/i1_5 ), .A3(
        \SB2_0_0/i1[9] ), .ZN(\SB2_0_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4012 ( .A1(\SB2_3_8/i0[10] ), .A2(\SB2_3_8/i0_0 ), .A3(
        \SB2_3_8/i0[6] ), .ZN(\SB2_3_8/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U4014 ( .A1(\SB1_1_22/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_22/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_22/Component_Function_2/NAND4_in[2] ), .A4(n1751), .ZN(
        \RI3[1][74] ) );
  NAND3_X1 U4015 ( .A1(\SB1_1_22/i0_0 ), .A2(\SB1_1_22/i0_4 ), .A3(
        \SB1_1_22/i1_5 ), .ZN(n1751) );
  NAND4_X1 U4016 ( .A1(\SB1_1_31/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_31/Component_Function_4/NAND4_in[2] ), .A4(n1752), .ZN(
        \RI3[1][10] ) );
  NAND3_X1 U4017 ( .A1(\SB1_1_31/i1[9] ), .A2(\SB1_1_31/i0_4 ), .A3(
        \SB1_1_31/i1_5 ), .ZN(n1752) );
  NAND3_X1 U4018 ( .A1(\SB2_0_0/i0_4 ), .A2(\SB2_0_0/i0_3 ), .A3(
        \SB2_0_0/i1[9] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4019 ( .A1(\SB4_5/i0_3 ), .A2(\SB4_5/i0_0 ), .A3(n549), .ZN(
        \SB4_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4020 ( .A1(n1657), .A2(\SB1_2_9/i0[10] ), .A3(\SB1_2_9/i0[9] ), 
        .ZN(\SB1_2_9/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4021 ( .A1(\SB1_2_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_9/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_9/Component_Function_5/NAND4_in[0] ), .A4(n1753), .ZN(
        \RI3[2][137] ) );
  NAND3_X1 U4022 ( .A1(n1657), .A2(\SB1_2_9/i1[9] ), .A3(\SB1_2_9/i0_4 ), .ZN(
        n1753) );
  NAND3_X1 U4023 ( .A1(\SB1_2_0/i0_3 ), .A2(\SB1_2_0/i0[10] ), .A3(
        \SB1_2_0/i0[9] ), .ZN(\SB1_2_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4024 ( .A1(\SB1_2_11/i0_3 ), .A2(\SB1_2_11/i0[10] ), .A3(
        \SB1_2_11/i0[9] ), .ZN(\SB1_2_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4025 ( .A1(\SB2_2_5/i0_4 ), .A2(\SB2_2_5/i1[9] ), .A3(
        \SB2_2_5/i0_3 ), .ZN(\SB2_2_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4026 ( .A1(\SB1_2_17/i0_3 ), .A2(\SB1_2_17/i1[9] ), .A3(
        \SB1_2_17/i0_4 ), .ZN(n1797) );
  NAND3_X1 U4027 ( .A1(\SB2_0_23/i0[6] ), .A2(\SB2_0_23/i0_0 ), .A3(
        \SB2_0_23/i0[10] ), .ZN(\SB2_0_23/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U4029 ( .A1(\SB2_0_10/i0_3 ), .A2(\SB2_0_10/i0[9] ), .A3(
        \SB2_0_10/i0[8] ), .ZN(n1754) );
  NAND3_X1 U4030 ( .A1(\SB2_1_9/i0_0 ), .A2(\SB2_1_9/i0_4 ), .A3(
        \SB2_1_9/i1_5 ), .ZN(n894) );
  NAND3_X1 U4031 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0[9] ), .A3(
        \SB1_0_16/i0[10] ), .ZN(\SB1_0_16/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U4032 ( .A1(\SB1_1_18/i0_0 ), .A2(\SB1_1_18/i0_4 ), .A3(
        \SB1_1_18/i1_5 ), .ZN(\SB1_1_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4034 ( .A1(\SB2_3_2/i0[9] ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0[8] ), .ZN(\SB2_3_2/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U4035 ( .A1(\SB2_1_24/i0_0 ), .A2(\SB2_1_24/i3[0] ), .ZN(n1755) );
  NAND3_X1 U4036 ( .A1(\SB1_2_1/i0_3 ), .A2(\SB1_2_1/i1[9] ), .A3(
        \SB1_2_1/i0[6] ), .ZN(\SB1_2_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4037 ( .A1(\SB2_1_5/i0_4 ), .A2(\SB2_1_5/i0_0 ), .A3(
        \SB2_1_5/i1_5 ), .ZN(\SB2_1_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4038 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i1_5 ), .ZN(\SB1_3_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4039 ( .A1(\SB2_0_19/i0[6] ), .A2(\SB2_0_19/i0_0 ), .A3(
        \SB2_0_19/i0[10] ), .ZN(\SB2_0_19/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U4040 ( .A1(\SB2_0_14/i0[6] ), .A2(\SB2_0_14/i1[9] ), .A3(
        \SB2_0_14/i0_3 ), .ZN(\SB2_0_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4041 ( .A1(n2131), .A2(\SB4_29/i1_5 ), .A3(\SB4_29/i1[9] ), .ZN(
        n1921) );
  NAND3_X1 U4042 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i1[9] ), .A3(
        \SB2_0_3/i1_7 ), .ZN(\SB2_0_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4044 ( .A1(\SB2_0_7/i0_4 ), .A2(\SB2_0_7/i1_5 ), .A3(
        \SB2_0_7/i1[9] ), .ZN(n1756) );
  NAND3_X1 U4045 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i1[9] ), .A3(
        \SB4_25/i1_7 ), .ZN(n1757) );
  NAND3_X1 U4046 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i1_7 ), .ZN(\SB1_3_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4047 ( .A1(\SB1_2_17/i0[6] ), .A2(\SB1_2_17/i0_0 ), .A3(
        \SB1_2_17/i0[10] ), .ZN(\SB1_2_17/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U4048 ( .A1(\SB2_1_4/i0[8] ), .A2(\SB2_1_4/i1_5 ), .A3(
        \SB2_1_4/i3[0] ), .ZN(\SB2_1_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4049 ( .A1(\SB2_0_12/i0_3 ), .A2(\SB2_0_12/i0[9] ), .A3(
        \SB2_0_12/i0[8] ), .ZN(\SB2_0_12/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U4050 ( .A1(\SB2_0_12/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_12/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_12/Component_Function_3/NAND4_in[2] ), .A4(n1758), .ZN(
        \RI5[0][129] ) );
  NAND3_X1 U4051 ( .A1(\SB2_0_12/i1_5 ), .A2(\SB2_0_12/i3[0] ), .A3(
        \SB2_0_12/i0[8] ), .ZN(n1758) );
  NAND4_X1 U4052 ( .A1(\SB2_1_27/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_27/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_27/Component_Function_4/NAND4_in[1] ), .A4(n1759), .ZN(
        \RI5[1][34] ) );
  NAND3_X1 U4053 ( .A1(\SB2_1_27/i0_3 ), .A2(\SB2_1_27/i0[9] ), .A3(
        \SB2_1_27/i0[10] ), .ZN(n1759) );
  NAND3_X1 U4056 ( .A1(\SB4_22/i0_4 ), .A2(n779), .A3(\SB4_22/i0[6] ), .ZN(
        \SB4_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4057 ( .A1(\SB4_13/i0_4 ), .A2(\SB4_13/i0[9] ), .A3(\SB4_13/i0[6] ), .ZN(\SB4_13/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U4058 ( .A1(\SB2_3_9/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_9/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_9/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_3_9/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[142] ) );
  NAND4_X2 U4059 ( .A1(\SB2_2_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_24/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_24/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[47] ) );
  NAND4_X1 U4060 ( .A1(\SB2_1_26/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_26/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_26/Component_Function_1/NAND4_in[0] ), .A4(n1761), .ZN(
        \RI5[1][55] ) );
  NAND3_X1 U4061 ( .A1(\SB2_1_26/i0_4 ), .A2(\SB2_1_26/i1_7 ), .A3(
        \SB2_1_26/i0[8] ), .ZN(n1761) );
  INV_X2 U4062 ( .A(\RI1[2][35] ), .ZN(\SB1_2_26/i0_3 ) );
  NAND3_X1 U4068 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0[10] ), .A3(
        \SB1_0_7/i0[9] ), .ZN(\SB1_0_7/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4069 ( .A1(\SB1_2_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_2_1/Component_Function_3/NAND4_in[0] ), .A4(n1763), .ZN(
        \RI3[2][3] ) );
  NAND3_X1 U4070 ( .A1(\SB1_2_1/i3[0] ), .A2(\SB1_2_1/i1_5 ), .A3(
        \SB1_2_1/i0[8] ), .ZN(n1763) );
  NAND3_X1 U4072 ( .A1(\SB2_1_15/i0_4 ), .A2(\RI3[1][96] ), .A3(
        \SB2_1_15/i0[6] ), .ZN(\SB2_1_15/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U4073 ( .A1(\SB2_3_31/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_31/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_3_31/Component_Function_2/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[20] ) );
  NAND3_X1 U4074 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0[10] ), .A3(
        \SB1_1_6/i0[9] ), .ZN(\SB1_1_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4075 ( .A1(\SB2_2_29/i0[9] ), .A2(\SB2_2_29/i0[10] ), .A3(
        \SB2_2_29/i0_3 ), .ZN(\SB2_2_29/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4076 ( .A1(\SB1_3_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_31/Component_Function_2/NAND4_in[2] ), .A4(n1765), .ZN(
        \RI3[3][20] ) );
  NAND3_X1 U4077 ( .A1(\SB1_3_31/i0_0 ), .A2(\SB1_3_31/i1_5 ), .A3(
        \SB1_3_31/i0_4 ), .ZN(n1765) );
  NAND3_X1 U4078 ( .A1(\SB2_1_8/i0_0 ), .A2(\SB2_1_8/i0[6] ), .A3(
        \SB2_1_8/i0[10] ), .ZN(\SB2_1_8/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U4079 ( .A(n1766), .B(n658), .ZN(\RI1[3][155] ) );
  XNOR2_X1 U4080 ( .A(\MC_ARK_ARC_1_2/temp3[155] ), .B(
        \MC_ARK_ARC_1_2/temp2[155] ), .ZN(n1766) );
  XNOR2_X1 U4081 ( .A(n1767), .B(n364), .ZN(Ciphertext[58]) );
  NAND4_X1 U4082 ( .A1(n706), .A2(\SB4_22/Component_Function_4/NAND4_in[2] ), 
        .A3(\SB4_22/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_22/Component_Function_4/NAND4_in[1] ), .ZN(n1767) );
  NAND2_X1 U4083 ( .A1(\SB2_2_15/i0[6] ), .A2(n1768), .ZN(
        \SB2_2_15/Component_Function_5/NAND4_in[3] ) );
  AND2_X1 U4084 ( .A1(\RI3[2][100] ), .A2(\RI3[2][96] ), .ZN(n1768) );
  XNOR2_X1 U4085 ( .A(n1769), .B(n1794), .ZN(\RI1[1][146] ) );
  XNOR2_X1 U4086 ( .A(\MC_ARK_ARC_1_0/temp1[146] ), .B(
        \MC_ARK_ARC_1_0/temp2[146] ), .ZN(n1769) );
  NAND3_X1 U4088 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i1_5 ), .A3(
        \SB4_29/i1[9] ), .ZN(n1770) );
  NAND3_X1 U4089 ( .A1(\SB1_1_15/i1[9] ), .A2(\SB1_1_15/i0[10] ), .A3(
        \SB1_1_15/i1_7 ), .ZN(\SB1_1_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4091 ( .A1(\SB2_1_2/i3[0] ), .A2(\SB2_1_2/i0[8] ), .A3(
        \SB2_1_2/i1_5 ), .ZN(n1771) );
  NAND4_X1 U4092 ( .A1(\SB1_3_18/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_18/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_18/Component_Function_2/NAND4_in[2] ), .A4(n1772), .ZN(
        \RI3[3][98] ) );
  NAND3_X1 U4093 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i0_4 ), .A3(
        \SB1_3_18/i1_5 ), .ZN(n1772) );
  NAND4_X2 U4094 ( .A1(\SB2_1_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_13/Component_Function_3/NAND4_in[2] ), .A4(n1773), .ZN(
        \RI5[1][123] ) );
  NAND3_X1 U4095 ( .A1(\SB2_1_13/i3[0] ), .A2(\SB2_1_13/i0[8] ), .A3(
        \SB2_1_13/i1_5 ), .ZN(n1773) );
  NAND4_X1 U4096 ( .A1(\SB2_3_15/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_15/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_15/Component_Function_2/NAND4_in[1] ), .A4(n1774), .ZN(
        \RI5[3][116] ) );
  NAND3_X1 U4097 ( .A1(\SB2_3_15/i0_0 ), .A2(\SB2_3_15/i1_5 ), .A3(
        \SB2_3_15/i0_4 ), .ZN(n1774) );
  NAND3_X1 U4098 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0_0 ), .A3(
        \SB1_0_16/i0_4 ), .ZN(\SB1_0_16/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U4099 ( .A1(\SB2_0_3/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_3/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_2/NAND4_in[0] ), .A4(n938), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[188] ) );
  NAND3_X1 U4100 ( .A1(\SB2_2_26/i0[9] ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i0[8] ), .ZN(n1284) );
  NAND3_X1 U4101 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i0_4 ), .A3(
        \SB1_3_7/i1_5 ), .ZN(n667) );
  NAND4_X1 U4103 ( .A1(\SB2_1_22/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_22/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_22/Component_Function_4/NAND4_in[1] ), .A4(n1775), .ZN(
        \RI5[1][64] ) );
  NAND3_X1 U4104 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0[10] ), .A3(
        \SB2_1_22/i0[9] ), .ZN(n1775) );
  NAND4_X1 U4106 ( .A1(\SB1_3_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_8/Component_Function_5/NAND4_in[0] ), .A4(n1776), .ZN(
        \RI3[3][143] ) );
  NAND3_X1 U4107 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i1[9] ), .A3(
        \SB1_3_8/i0_4 ), .ZN(n1776) );
  NAND3_X1 U4108 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0[6] ), .A3(
        \SB2_1_26/i0[10] ), .ZN(\SB2_1_26/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X1 U4109 ( .A1(\SB2_0_26/i0[10] ), .A2(\SB2_0_26/i1[9] ), .A3(
        \SB2_0_26/i1_7 ), .ZN(n1777) );
  NAND4_X1 U4110 ( .A1(\SB1_3_28/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_3_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_5/NAND4_in[0] ), .A4(n1778), .ZN(
        \RI3[3][23] ) );
  NAND3_X1 U4111 ( .A1(\SB1_3_28/i1[9] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i0_4 ), .ZN(n1778) );
  NAND3_X1 U4112 ( .A1(\SB4_7/i0[10] ), .A2(\SB4_7/i1_5 ), .A3(\SB4_7/i1[9] ), 
        .ZN(n1779) );
  XNOR2_X1 U4113 ( .A(n1781), .B(n1780), .ZN(\RI1[1][23] ) );
  XNOR2_X1 U4114 ( .A(\MC_ARK_ARC_1_0/temp2[23] ), .B(
        \MC_ARK_ARC_1_0/temp4[23] ), .ZN(n1780) );
  XNOR2_X1 U4115 ( .A(\MC_ARK_ARC_1_0/temp3[23] ), .B(
        \MC_ARK_ARC_1_0/temp1[23] ), .ZN(n1781) );
  NAND3_X1 U4116 ( .A1(\SB1_2_8/i0[7] ), .A2(\SB1_2_8/i0_0 ), .A3(
        \SB1_2_8/i0_3 ), .ZN(\SB1_2_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4117 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i1_5 ), .A3(n834), .ZN(
        \SB4_5/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U4118 ( .A1(\SB1_3_24/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_24/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_24/Component_Function_2/NAND4_in[2] ), .A4(n1782), .ZN(
        \RI3[3][62] ) );
  NAND3_X1 U4119 ( .A1(\SB1_3_24/i0_0 ), .A2(\SB1_3_24/i0_4 ), .A3(
        \SB1_3_24/i1_5 ), .ZN(n1782) );
  NAND3_X1 U4120 ( .A1(\SB2_0_31/i0_4 ), .A2(\SB2_0_31/i0_0 ), .A3(
        \SB2_0_31/i0_3 ), .ZN(\SB2_0_31/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U4121 ( .A(n1783), .B(n273), .ZN(Ciphertext[154]) );
  NAND4_X1 U4122 ( .A1(\SB4_6/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_6/Component_Function_4/NAND4_in[3] ), .A3(
        \SB4_6/Component_Function_4/NAND4_in[0] ), .A4(n747), .ZN(n1783) );
  NAND3_X1 U4123 ( .A1(\SB2_3_27/i0[9] ), .A2(n1630), .A3(\SB2_3_27/i0[6] ), 
        .ZN(\SB2_3_27/Component_Function_1/NAND4_in[2] ) );
  NAND4_X1 U4128 ( .A1(\SB2_0_4/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_0_4/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_4/Component_Function_4/NAND4_in[1] ), .A4(n1786), .ZN(
        \RI5[0][172] ) );
  NAND3_X1 U4129 ( .A1(\SB2_0_4/i0_4 ), .A2(\SB2_0_4/i1[9] ), .A3(
        \SB2_0_4/i1_5 ), .ZN(n1786) );
  XNOR2_X1 U4131 ( .A(n1787), .B(n351), .ZN(Ciphertext[101]) );
  NAND4_X1 U4132 ( .A1(\SB4_15/Component_Function_5/NAND4_in[2] ), .A2(n929), 
        .A3(n1059), .A4(\SB4_15/Component_Function_5/NAND4_in[0] ), .ZN(n1787)
         );
  XNOR2_X1 U4134 ( .A(n1788), .B(n198), .ZN(Ciphertext[179]) );
  NAND4_X1 U4135 ( .A1(\SB4_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_2/Component_Function_5/NAND4_in[3] ), .A3(n1822), .A4(
        \SB4_2/Component_Function_5/NAND4_in[0] ), .ZN(n1788) );
  NAND4_X2 U4136 ( .A1(\SB2_0_22/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_22/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_22/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[69] ) );
  NAND4_X1 U4137 ( .A1(\SB2_1_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_29/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_29/Component_Function_1/NAND4_in[2] ), .A4(n1789), .ZN(
        \RI5[1][37] ) );
  NAND3_X1 U4138 ( .A1(\SB2_1_29/i0_4 ), .A2(\SB2_1_29/i1_7 ), .A3(
        \SB2_1_29/i0[8] ), .ZN(n1789) );
  NAND3_X1 U4139 ( .A1(\SB1_3_15/i0[10] ), .A2(\SB1_3_15/i1_5 ), .A3(
        \SB1_3_15/i1[9] ), .ZN(\SB1_3_15/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4140 ( .A1(\SB3_22/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_2/NAND4_in[0] ), .A4(n1790), .ZN(
        \RI3[4][74] ) );
  NAND3_X1 U4141 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i1_5 ), .A3(\SB3_22/i0_4 ), 
        .ZN(n1790) );
  NAND3_X1 U4144 ( .A1(\SB3_9/i0_0 ), .A2(\SB3_9/i1_5 ), .A3(\SB3_9/i0_4 ), 
        .ZN(\SB3_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4145 ( .A1(\SB1_3_15/i0[10] ), .A2(\SB1_3_15/i1_7 ), .A3(
        \SB1_3_15/i1[9] ), .ZN(\SB1_3_15/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U4146 ( .A1(\SB1_1_10/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_1_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_5/NAND4_in[0] ), .A4(n1792), .ZN(
        \RI3[1][131] ) );
  NAND3_X1 U4147 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i1[9] ), .A3(
        \SB1_1_10/i0_4 ), .ZN(n1792) );
  NAND3_X1 U4148 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0[8] ), .A3(
        \SB2_2_28/i0[9] ), .ZN(n1793) );
  NAND3_X1 U4149 ( .A1(\SB1_2_15/i0_3 ), .A2(\SB1_2_15/i0[9] ), .A3(
        \SB1_2_15/i0[8] ), .ZN(\SB1_2_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4150 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i1[9] ), .A3(
        \SB4_15/i1_7 ), .ZN(\SB4_15/Component_Function_3/NAND4_in[2] ) );
  XNOR2_X1 U4151 ( .A(\MC_ARK_ARC_1_0/temp3[146] ), .B(
        \MC_ARK_ARC_1_0/temp4[146] ), .ZN(n1794) );
  NAND3_X1 U4153 ( .A1(\SB2_0_9/i0_3 ), .A2(\SB2_0_9/i0[10] ), .A3(
        \SB2_0_9/i0[9] ), .ZN(\SB2_0_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4154 ( .A1(\SB2_2_25/i0_4 ), .A2(\SB2_2_25/i1_7 ), .A3(
        \SB2_2_25/i0[8] ), .ZN(\SB2_2_25/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U4155 ( .A1(\SB2_0_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_9/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[147] ) );
  NAND4_X1 U4156 ( .A1(\SB2_1_31/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_31/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_31/Component_Function_4/NAND4_in[1] ), .A4(n1795), .ZN(
        \RI5[1][10] ) );
  NAND3_X1 U4157 ( .A1(\SB2_1_31/i0_3 ), .A2(\RI3[1][0] ), .A3(
        \SB2_1_31/i0[10] ), .ZN(n1795) );
  NAND3_X1 U4158 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i1[9] ), .A3(\SB4_12/i1_5 ), 
        .ZN(\SB4_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4161 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0[10] ), .ZN(\SB2_2_7/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4162 ( .A1(\SB2_2_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_27/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_27/Component_Function_2/NAND4_in[2] ), .A4(n1796), .ZN(
        \RI5[2][44] ) );
  NAND3_X1 U4163 ( .A1(\SB2_2_27/i0_4 ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB2_2_27/i0_0 ), .ZN(n1796) );
  NAND4_X1 U4164 ( .A1(\SB1_2_17/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_17/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_2_17/Component_Function_5/NAND4_in[3] ), .A4(n1797), .ZN(
        \RI3[2][89] ) );
  NAND3_X1 U4165 ( .A1(\SB2_1_14/i0[9] ), .A2(\SB2_1_14/i0_3 ), .A3(
        \SB2_1_14/i0[8] ), .ZN(\SB2_1_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4166 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0_0 ), .A3(
        \SB1_1_16/i0_4 ), .ZN(\SB1_1_16/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U4167 ( .A(n1798), .B(n206), .ZN(Ciphertext[164]) );
  NAND3_X1 U4168 ( .A1(\SB2_0_0/i0[6] ), .A2(\SB2_0_0/i0_0 ), .A3(
        \SB2_0_0/i0[10] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4169 ( .A1(\SB2_0_5/i0[6] ), .A2(\SB2_0_5/i0_4 ), .A3(
        \RI3[0][156] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4170 ( .A1(\SB2_0_23/i3[0] ), .A2(\SB2_0_23/i1_5 ), .A3(
        \SB2_0_23/i0[8] ), .ZN(n1799) );
  NAND3_X1 U4172 ( .A1(\SB2_0_5/i3[0] ), .A2(\SB2_0_5/i1_5 ), .A3(
        \SB2_0_5/i0[8] ), .ZN(n1800) );
  NAND4_X1 U4173 ( .A1(\SB2_2_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_25/Component_Function_4/NAND4_in[1] ), .A4(n1801), .ZN(
        \RI5[2][46] ) );
  NAND3_X1 U4174 ( .A1(\SB2_2_25/i0_4 ), .A2(\SB2_2_25/i1_5 ), .A3(
        \SB2_2_25/i1[9] ), .ZN(n1801) );
  XNOR2_X1 U4175 ( .A(n1802), .B(\MC_ARK_ARC_1_1/temp5[134] ), .ZN(
        \RI1[2][134] ) );
  XNOR2_X1 U4176 ( .A(\MC_ARK_ARC_1_1/temp3[134] ), .B(
        \MC_ARK_ARC_1_1/temp4[134] ), .ZN(n1802) );
  NAND3_X1 U4177 ( .A1(\SB2_0_8/i0_3 ), .A2(\SB2_0_8/i0[9] ), .A3(
        \SB2_0_8/i0[8] ), .ZN(\SB2_0_8/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U4178 ( .A1(\SB4_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_11/Component_Function_3/NAND4_in[3] ), .A3(n1847), .A4(n1803), 
        .ZN(n1841) );
  NAND3_X1 U4179 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i1_7 ), .A3(
        \SB4_11/i1[9] ), .ZN(n1803) );
  NAND3_X1 U4180 ( .A1(\SB2_1_6/i0_4 ), .A2(\SB2_1_6/i0_3 ), .A3(
        \SB2_1_6/i1[9] ), .ZN(\SB2_1_6/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U4181 ( .A1(\SB3_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_3/NAND4_in[3] ), .A3(
        \SB3_28/Component_Function_3/NAND4_in[1] ), .A4(n1804), .ZN(
        \RI3[4][33] ) );
  NAND3_X1 U4182 ( .A1(\SB3_28/i1_7 ), .A2(\SB3_28/i0[10] ), .A3(
        \SB3_28/i1[9] ), .ZN(n1804) );
  NAND4_X1 U4183 ( .A1(\SB4_4/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_4/Component_Function_1/NAND4_in[0] ), .A3(
        \SB4_4/Component_Function_1/NAND4_in[3] ), .A4(n1805), .ZN(n1030) );
  NAND3_X1 U4184 ( .A1(\SB4_4/i0[9] ), .A2(\SB4_4/i1_5 ), .A3(\SB4_4/i0[6] ), 
        .ZN(n1805) );
  NAND3_X1 U4185 ( .A1(\SB4_4/i0[9] ), .A2(\SB4_4/i0_4 ), .A3(\SB4_4/i0[6] ), 
        .ZN(n1806) );
  NAND4_X1 U4186 ( .A1(\SB3_14/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_3/NAND4_in[0] ), .A4(n1807), .ZN(
        \RI3[4][117] ) );
  NAND3_X1 U4187 ( .A1(\SB3_14/i3[0] ), .A2(\SB3_14/i1_5 ), .A3(\SB3_14/i0[8] ), .ZN(n1807) );
  NAND4_X1 U4188 ( .A1(\SB2_2_25/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_25/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_25/Component_Function_2/NAND4_in[1] ), .A4(n1808), .ZN(
        \RI5[2][56] ) );
  NAND3_X1 U4189 ( .A1(\SB2_2_25/i0_4 ), .A2(\SB2_2_25/i1_5 ), .A3(
        \SB2_2_25/i0_0 ), .ZN(n1808) );
  XNOR2_X1 U4190 ( .A(\MC_ARK_ARC_1_3/buf_datainput[12] ), .B(\RI5[3][168] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[102] ) );
  NAND4_X2 U4191 ( .A1(\SB2_3_8/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_8/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_8/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][168] ) );
  NAND3_X1 U4192 ( .A1(\RI3[0][168] ), .A2(\SB2_0_3/i0_4 ), .A3(\RI3[0][169] ), 
        .ZN(\SB2_0_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4193 ( .A1(\SB2_0_9/i0_4 ), .A2(\SB2_0_9/i0[9] ), .A3(
        \SB2_0_9/i0[6] ), .ZN(\SB2_0_9/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U4195 ( .A1(n1418), .A2(\SB2_0_9/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_0_9/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_9/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[137] ) );
  NAND3_X1 U4196 ( .A1(\SB4_22/i1_5 ), .A2(\SB4_22/i1[9] ), .A3(
        \SB4_22/i0[10] ), .ZN(n567) );
  NAND3_X1 U4197 ( .A1(\SB2_2_11/i0[9] ), .A2(\SB2_2_11/i0_3 ), .A3(
        \SB2_2_11/i0[8] ), .ZN(n1210) );
  NAND3_X1 U4198 ( .A1(\SB1_2_17/i3[0] ), .A2(\SB1_2_17/i1_5 ), .A3(
        \SB1_2_17/i0[8] ), .ZN(\SB1_2_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4199 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i1_5 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4200 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0_4 ), .A3(
        \SB2_1_15/i1[9] ), .ZN(\SB2_1_15/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4201 ( .A1(\SB1_2_27/i0_3 ), .A2(\SB1_2_27/i1[9] ), .A3(
        \SB1_2_27/i0_4 ), .ZN(n1809) );
  NAND3_X1 U4202 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0[10] ), .A3(
        \SB1_0_6/i0[9] ), .ZN(\SB1_0_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4203 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0[10] ), .A3(
        \SB1_1_14/i0_4 ), .ZN(\SB1_1_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4204 ( .A1(\SB1_0_2/i0[9] ), .A2(\SB1_0_2/i0[10] ), .A3(
        \SB1_0_2/i0_3 ), .ZN(\SB1_0_2/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4205 ( .A1(\SB1_2_27/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_27/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_2_27/Component_Function_5/NAND4_in[3] ), .A4(n1809), .ZN(
        \RI3[2][29] ) );
  NAND3_X1 U4206 ( .A1(\SB2_1_19/i0[8] ), .A2(\SB2_1_19/i3[0] ), .A3(
        \SB2_1_19/i1_5 ), .ZN(n709) );
  XNOR2_X1 U4207 ( .A(n1811), .B(n1810), .ZN(\RI1[2][77] ) );
  XNOR2_X1 U4208 ( .A(\MC_ARK_ARC_1_1/temp3[77] ), .B(
        \MC_ARK_ARC_1_1/temp4[77] ), .ZN(n1810) );
  XNOR2_X1 U4209 ( .A(\MC_ARK_ARC_1_1/temp1[77] ), .B(
        \MC_ARK_ARC_1_1/temp2[77] ), .ZN(n1811) );
  NAND3_X1 U4210 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i0_4 ), .ZN(\SB1_1_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4211 ( .A1(\SB1_0_5/i0_4 ), .A2(\SB1_0_5/i0_0 ), .A3(
        \SB1_0_5/i1_5 ), .ZN(\SB1_0_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4212 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i0_0 ), .A3(
        \SB1_1_26/i0[6] ), .ZN(\SB1_1_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4213 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i1[9] ), .A3(
        \SB1_0_29/i0_4 ), .ZN(\SB1_0_29/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U4214 ( .A1(\SB1_1_1/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_1/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_1/Component_Function_5/NAND4_in[0] ), .A4(n1812), .ZN(
        \RI3[1][185] ) );
  NAND3_X1 U4215 ( .A1(\SB1_1_1/i1[9] ), .A2(\SB1_1_1/i0_3 ), .A3(
        \SB1_1_1/i0_4 ), .ZN(n1812) );
  XNOR2_X1 U4217 ( .A(\MC_ARK_ARC_1_1/temp1[185] ), .B(
        \MC_ARK_ARC_1_1/temp4[185] ), .ZN(n1813) );
  XNOR2_X1 U4218 ( .A(\MC_ARK_ARC_1_1/temp3[185] ), .B(
        \MC_ARK_ARC_1_1/temp2[185] ), .ZN(n1814) );
  NAND3_X1 U4219 ( .A1(\SB2_0_3/i0_0 ), .A2(\SB2_0_3/i3[0] ), .A3(
        \SB2_0_3/i1_7 ), .ZN(\SB2_0_3/Component_Function_4/NAND4_in[1] ) );
  XNOR2_X1 U4220 ( .A(\MC_ARK_ARC_1_2/temp1[80] ), .B(
        \MC_ARK_ARC_1_2/temp4[80] ), .ZN(n1815) );
  NAND3_X1 U4221 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0_0 ), .A3(
        \SB2_0_21/i0_4 ), .ZN(\SB2_0_21/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U4222 ( .A(n1816), .B(n294), .ZN(Ciphertext[96]) );
  NAND4_X1 U4223 ( .A1(\SB4_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_15/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_15/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_15/Component_Function_0/NAND4_in[1] ), .ZN(n1816) );
  NAND4_X1 U4224 ( .A1(\SB1_2_22/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_22/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_2_22/Component_Function_5/NAND4_in[3] ), .A4(n1817), .ZN(
        \RI3[2][59] ) );
  NAND3_X1 U4225 ( .A1(\SB1_2_22/i0_3 ), .A2(\SB1_2_22/i1[9] ), .A3(
        \SB1_2_22/i0_4 ), .ZN(n1817) );
  NAND3_X1 U4226 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i1[9] ), .A3(
        \SB1_1_20/i0_4 ), .ZN(\SB1_1_20/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U4227 ( .A(n1819), .B(n1818), .ZN(\RI1[2][149] ) );
  XNOR2_X1 U4228 ( .A(\MC_ARK_ARC_1_1/temp1[149] ), .B(
        \MC_ARK_ARC_1_1/temp4[149] ), .ZN(n1818) );
  XNOR2_X1 U4229 ( .A(\MC_ARK_ARC_1_1/temp2[149] ), .B(
        \MC_ARK_ARC_1_1/temp3[149] ), .ZN(n1819) );
  NAND3_X1 U4230 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i0[9] ), .A3(
        \SB2_1_31/i0[8] ), .ZN(\SB2_1_31/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U4231 ( .A(n1820), .B(\MC_ARK_ARC_1_3/temp6[64] ), .ZN(\RI1[4][64] ) );
  XNOR2_X1 U4232 ( .A(\MC_ARK_ARC_1_3/temp2[64] ), .B(
        \MC_ARK_ARC_1_3/temp1[64] ), .ZN(n1820) );
  NAND4_X1 U4233 ( .A1(\SB2_1_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_17/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_17/Component_Function_2/NAND4_in[1] ), .A4(n1821), .ZN(
        \RI5[1][104] ) );
  NAND3_X1 U4234 ( .A1(\SB2_1_17/i0_0 ), .A2(\SB2_1_17/i0_4 ), .A3(
        \SB2_1_17/i1_5 ), .ZN(n1821) );
  NAND3_X1 U4235 ( .A1(\SB2_0_24/i0[10] ), .A2(\SB2_0_24/i1_5 ), .A3(
        \SB2_0_24/i1[9] ), .ZN(\SB2_0_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4236 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i0[6] ), 
        .ZN(n1822) );
  XNOR2_X1 U4237 ( .A(n1823), .B(n272), .ZN(Ciphertext[113]) );
  NAND4_X1 U4238 ( .A1(\SB4_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_13/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_13/Component_Function_5/NAND4_in[3] ), .ZN(n1823) );
  NAND3_X1 U4239 ( .A1(\SB4_11/i1_5 ), .A2(n805), .A3(\SB4_11/i1[9] ), .ZN(
        n1287) );
  NAND4_X2 U4244 ( .A1(\SB2_0_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_8/Component_Function_3/NAND4_in[0] ), .A3(n1121), .A4(
        \SB2_0_8/Component_Function_3/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[153] ) );
  NAND3_X1 U4245 ( .A1(\SB1_0_12/i0_0 ), .A2(n381), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4249 ( .A1(\SB2_0_5/i0_4 ), .A2(\SB2_0_5/i0_3 ), .A3(
        \SB2_0_5/i1[9] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4250 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0[8] ), .A3(
        \SB1_0_18/i1_7 ), .ZN(\SB1_0_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4251 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[10] ), .A3(
        \SB1_1_20/i0[9] ), .ZN(\SB1_1_20/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4252 ( .A1(\SB3_29/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_3/NAND4_in[0] ), .A4(n1827), .ZN(
        \RI3[4][27] ) );
  NAND3_X1 U4253 ( .A1(\SB3_29/i3[0] ), .A2(\SB3_29/i0[8] ), .A3(\SB3_29/i1_5 ), .ZN(n1827) );
  NAND3_X1 U4254 ( .A1(\SB1_3_29/i0[10] ), .A2(\SB1_3_29/i0_3 ), .A3(
        \SB1_3_29/i0[6] ), .ZN(\SB1_3_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U4255 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i0[6] ), .A3(
        \RI3[1][180] ), .ZN(\SB2_1_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4256 ( .A1(n2132), .A2(\SB2_0_26/i0[10] ), .A3(\SB2_0_26/i0_3 ), 
        .ZN(n1222) );
  NAND3_X1 U4257 ( .A1(\SB2_0_24/i3[0] ), .A2(\SB2_0_24/i1_5 ), .A3(
        \SB2_0_24/i0[8] ), .ZN(\SB2_0_24/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U4258 ( .A1(\SB1_3_2/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_2/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_3_2/Component_Function_5/NAND4_in[0] ), .A4(n1828), .ZN(
        \RI3[3][179] ) );
  NAND3_X1 U4259 ( .A1(\SB1_3_2/i0_4 ), .A2(\SB1_3_2/i0[9] ), .A3(
        \SB1_3_2/i0[6] ), .ZN(n1828) );
  NAND3_X1 U4260 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i1_7 ), .A3(
        \SB2_1_2/i1[9] ), .ZN(\SB2_1_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4261 ( .A1(\SB2_1_13/i0_4 ), .A2(\SB2_1_13/i1_7 ), .A3(
        \SB2_1_13/i0[8] ), .ZN(\SB2_1_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4262 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0[9] ), .A3(
        \SB2_1_4/i0[8] ), .ZN(\SB2_1_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4263 ( .A1(\SB2_0_11/i0[9] ), .A2(\SB2_0_11/i0[10] ), .A3(
        \SB2_0_11/i0_3 ), .ZN(\SB2_0_11/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4264 ( .A1(\SB1_0_8/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_8/Component_Function_4/NAND4_in[3] ), .A4(n1829), .ZN(
        \RI3[0][148] ) );
  NAND3_X1 U4265 ( .A1(\SB1_0_8/i1_7 ), .A2(\SB1_0_8/i3[0] ), .A3(
        \SB1_0_8/i0_0 ), .ZN(n1829) );
  NAND3_X1 U4266 ( .A1(\SB2_0_30/i0[10] ), .A2(\SB2_0_30/i1[9] ), .A3(
        \SB2_0_30/i1_7 ), .ZN(\SB2_0_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4267 ( .A1(\SB1_0_5/i0_4 ), .A2(\SB1_0_5/i0_3 ), .A3(
        \SB1_0_5/i1[9] ), .ZN(n582) );
  NAND3_X1 U4268 ( .A1(\SB1_2_29/i1[9] ), .A2(\SB1_2_29/i0_4 ), .A3(
        \SB1_2_29/i0_3 ), .ZN(n1378) );
  NAND3_X1 U4269 ( .A1(\SB4_27/i0[10] ), .A2(\SB4_27/i1[9] ), .A3(
        \SB4_27/i1_7 ), .ZN(\SB4_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4270 ( .A1(\SB1_1_22/i1[9] ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i1_7 ), .ZN(\SB1_1_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4271 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i0_0 ), .A3(
        \SB2_2_27/i0[6] ), .ZN(\SB2_2_27/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U4272 ( .A1(\SB1_0_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_8/Component_Function_3/NAND4_in[3] ), .A4(n1830), .ZN(
        \RI3[0][153] ) );
  NAND3_X1 U4273 ( .A1(\SB1_0_8/i1_7 ), .A2(\SB1_0_8/i1[9] ), .A3(
        \SB1_0_8/i0[10] ), .ZN(n1830) );
  NAND3_X1 U4274 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[9] ), .A3(
        \SB2_0_22/i0[10] ), .ZN(\SB2_0_22/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U4275 ( .A1(\SB1_2_7/i0_3 ), .A2(\SB1_2_7/i0[10] ), .A3(
        \SB1_2_7/i0[9] ), .ZN(\SB1_2_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4276 ( .A1(\SB2_2_4/i0_4 ), .A2(\SB2_2_4/i0[9] ), .A3(
        \SB2_2_4/i0[6] ), .ZN(\SB2_2_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4277 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i0[8] ), .A3(
        \SB1_2_5/i0[9] ), .ZN(\SB1_2_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4278 ( .A1(\SB2_2_14/i0_4 ), .A2(\SB2_2_14/i0_0 ), .A3(
        \SB2_2_14/i0_3 ), .ZN(\SB2_2_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4279 ( .A1(\SB2_0_17/i3[0] ), .A2(\SB2_0_17/i1_5 ), .A3(
        \SB2_0_17/i0[8] ), .ZN(\SB2_0_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4280 ( .A1(\SB2_2_14/i0_4 ), .A2(\SB2_2_14/i1_5 ), .A3(
        \SB2_2_14/i1[9] ), .ZN(n1199) );
  NAND3_X1 U4281 ( .A1(\SB2_1_12/i0_3 ), .A2(\SB2_1_12/i0_4 ), .A3(
        \SB2_1_12/i1[9] ), .ZN(\SB2_1_12/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U4282 ( .A1(\SB2_0_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_0_17/Component_Function_2/NAND4_in[1] ), .A4(n1831), .ZN(
        \RI5[0][104] ) );
  NAND3_X1 U4283 ( .A1(\SB2_0_17/i0[9] ), .A2(\SB2_0_17/i0_3 ), .A3(
        \SB2_0_17/i0[8] ), .ZN(n1831) );
  NAND4_X1 U4284 ( .A1(\SB1_0_21/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_0_21/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_5/NAND4_in[0] ), .A4(n1832), .ZN(
        \RI3[0][65] ) );
  NAND3_X1 U4285 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0_4 ), .A3(
        \SB1_0_21/i1[9] ), .ZN(n1832) );
  NAND4_X1 U4286 ( .A1(\SB1_1_31/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_1_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_5/NAND4_in[0] ), .A4(n1833), .ZN(
        \RI3[1][5] ) );
  NAND3_X1 U4287 ( .A1(\SB1_1_31/i1[9] ), .A2(\SB1_1_31/i0_3 ), .A3(
        \SB1_1_31/i0_4 ), .ZN(n1833) );
  NAND4_X1 U4288 ( .A1(\SB1_0_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_0_19/Component_Function_3/NAND4_in[1] ), .A4(n1834), .ZN(
        \RI3[0][87] ) );
  NAND3_X1 U4289 ( .A1(\SB1_0_19/i1_7 ), .A2(\SB1_0_19/i0[10] ), .A3(
        \SB1_0_19/i1[9] ), .ZN(n1834) );
  NAND3_X1 U4290 ( .A1(\SB1_0_1/i1_5 ), .A2(\SB1_0_1/i0[9] ), .A3(
        \SB1_0_1/i0[6] ), .ZN(n1270) );
  INV_X2 U4293 ( .A(\RI1[2][59] ), .ZN(\SB1_2_22/i0_3 ) );
  XNOR2_X1 U4294 ( .A(n721), .B(\MC_ARK_ARC_1_1/temp6[59] ), .ZN(\RI1[2][59] )
         );
  NAND3_X1 U4295 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i0_4 ), .A3(
        \SB1_1_30/i1_5 ), .ZN(n1920) );
  XNOR2_X1 U4296 ( .A(n1836), .B(n350), .ZN(Ciphertext[60]) );
  NAND4_X1 U4297 ( .A1(\SB4_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_21/Component_Function_0/NAND4_in[3] ), .A3(n1105), .A4(
        \SB4_21/Component_Function_0/NAND4_in[0] ), .ZN(n1836) );
  XNOR2_X1 U4298 ( .A(n1837), .B(n324), .ZN(Ciphertext[64]) );
  NAND4_X1 U4299 ( .A1(\SB4_21/Component_Function_4/NAND4_in[2] ), .A2(n679), 
        .A3(\SB4_21/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_21/Component_Function_4/NAND4_in[1] ), .ZN(n1837) );
  NAND3_X1 U4300 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i0[10] ), .A3(
        \SB1_0_13/i0[9] ), .ZN(\SB1_0_13/Component_Function_4/NAND4_in[2] ) );
  INV_X2 U4301 ( .A(\RI1[3][71] ), .ZN(\SB1_3_20/i0_3 ) );
  NAND4_X1 U4302 ( .A1(n1161), .A2(\SB2_2_6/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB2_2_6/Component_Function_2/NAND4_in[1] ), .A4(n1838), .ZN(
        \RI5[2][170] ) );
  NAND3_X1 U4303 ( .A1(\SB2_3_20/i1[9] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i0[6] ), .ZN(\SB2_3_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4304 ( .A1(\SB4_17/i0_0 ), .A2(\SB4_17/i0_3 ), .A3(\SB4_17/i0_4 ), 
        .ZN(n1839) );
  NAND3_X1 U4305 ( .A1(\SB4_27/i0[10] ), .A2(\SB4_27/i1_5 ), .A3(
        \SB4_27/i1[9] ), .ZN(n1840) );
  XNOR2_X1 U4306 ( .A(n1841), .B(n205), .ZN(Ciphertext[123]) );
  NAND3_X1 U4307 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i1_5 ), .ZN(\SB1_3_3/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4310 ( .A1(\SB1_3_2/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_2/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_2/Component_Function_2/NAND4_in[2] ), .A4(n1843), .ZN(
        \RI3[3][2] ) );
  NAND3_X1 U4311 ( .A1(\SB1_3_2/i0_0 ), .A2(\SB1_3_2/i0_4 ), .A3(
        \SB1_3_2/i1_5 ), .ZN(n1843) );
  NAND4_X1 U4312 ( .A1(\SB1_1_23/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_23/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_1_23/Component_Function_5/NAND4_in[3] ), .A4(n1844), .ZN(
        \RI3[1][53] ) );
  NAND3_X1 U4313 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i1[9] ), .A3(
        \SB1_1_23/i0_4 ), .ZN(n1844) );
  NAND3_X1 U4314 ( .A1(\SB2_2_17/i0_0 ), .A2(\SB2_2_17/i0[10] ), .A3(
        \SB2_2_17/i0[6] ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4315 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB2_2_27/i0[6] ), .ZN(\SB2_2_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U4316 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i1[9] ), .ZN(n1295) );
  NAND3_X1 U4317 ( .A1(\SB2_0_30/i0[6] ), .A2(\SB2_0_30/i0_0 ), .A3(
        \SB2_0_30/i0[10] ), .ZN(\SB2_0_30/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U4318 ( .A1(\SB4_6/i0_4 ), .A2(n858), .A3(\SB4_6/i1[9] ), .ZN(
        \SB4_6/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U4319 ( .A1(\SB1_1_28/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_2/NAND4_in[0] ), .A4(n1845), .ZN(
        \RI3[1][38] ) );
  NAND3_X1 U4320 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i0_3 ), .A3(
        \SB1_3_2/i0[9] ), .ZN(n1123) );
  NAND4_X1 U4321 ( .A1(\SB3_24/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_24/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_5/NAND4_in[0] ), .A4(n1846), .ZN(
        \RI3[4][47] ) );
  NAND3_X1 U4322 ( .A1(\SB3_24/i1[9] ), .A2(\SB3_24/i0_4 ), .A3(\SB3_24/i0_3 ), 
        .ZN(n1846) );
  NAND3_X1 U4324 ( .A1(\SB2_1_8/i0[9] ), .A2(\SB2_1_8/i0[8] ), .A3(
        \SB2_1_8/i0_0 ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U4325 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[10] ), .A3(
        \SB1_0_25/i0[9] ), .ZN(\SB1_0_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4326 ( .A1(\SB4_11/i0_0 ), .A2(n841), .A3(n805), .ZN(n1847) );
  XNOR2_X1 U4329 ( .A(n1849), .B(n231), .ZN(Ciphertext[37]) );
  NAND4_X1 U4330 ( .A1(\SB1_3_30/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_30/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_30/Component_Function_3/NAND4_in[2] ), .A4(n1850), .ZN(
        \RI3[3][21] ) );
  NAND3_X1 U4331 ( .A1(\SB1_3_30/i3[0] ), .A2(\SB1_3_30/i1_5 ), .A3(
        \SB1_3_30/i0[8] ), .ZN(n1850) );
  XNOR2_X1 U4332 ( .A(n1851), .B(n288), .ZN(Ciphertext[42]) );
  NAND4_X1 U4333 ( .A1(\SB4_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_24/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_24/Component_Function_0/NAND4_in[0] ), .A4(n951), .ZN(n1851) );
  NAND3_X1 U4334 ( .A1(n2141), .A2(\SB1_1_11/i0[10] ), .A3(\SB1_1_11/i0[9] ), 
        .ZN(\SB1_1_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4335 ( .A1(\SB1_3_30/i0_3 ), .A2(\SB1_3_30/i0[9] ), .A3(
        \SB1_3_30/i0[10] ), .ZN(\SB1_3_30/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U4336 ( .A1(\SB2_1_6/i0[9] ), .A2(\SB2_1_6/i0_3 ), .A3(
        \SB2_1_6/i0[8] ), .ZN(\SB2_1_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4337 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0[10] ), .A3(
        \SB1_0_0/i0[9] ), .ZN(\SB1_0_0/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U4338 ( .A1(\SB1_1_11/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_11/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_11/Component_Function_2/NAND4_in[2] ), .A4(n1852), .ZN(
        \RI3[1][140] ) );
  NAND3_X1 U4339 ( .A1(\SB1_1_11/i0_0 ), .A2(\SB1_1_11/i0_4 ), .A3(
        \SB1_1_11/i1_5 ), .ZN(n1852) );
  NAND4_X1 U4340 ( .A1(\SB4_24/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_24/Component_Function_2/NAND4_in[3] ), .A4(n1853), .ZN(n1417) );
  NAND3_X1 U4341 ( .A1(\SB4_24/i0[10] ), .A2(\SB4_24/i1_5 ), .A3(
        \SB4_24/i1[9] ), .ZN(n1853) );
  XNOR2_X1 U4342 ( .A(\MC_ARK_ARC_1_3/buf_datainput[132] ), .B(\RI5[3][96] ), 
        .ZN(\MC_ARK_ARC_1_3/temp3[30] ) );
  NAND4_X2 U4343 ( .A1(\SB2_3_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_20/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_20/Component_Function_0/NAND4_in[0] ), .ZN(\RI5[3][96] ) );
  NAND3_X1 U4344 ( .A1(\SB1_3_30/i0_3 ), .A2(\SB1_3_30/i0[9] ), .A3(
        \SB1_3_30/i0[8] ), .ZN(\SB1_3_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4345 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i0_0 ), .A3(\SB3_12/i0_4 ), 
        .ZN(\SB3_12/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U4347 ( .A1(\SB2_0_0/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_0/Component_Function_2/NAND4_in[0] ), .A3(n917), .A4(n1855), 
        .ZN(\RI5[0][14] ) );
  NAND3_X1 U4348 ( .A1(\SB2_0_0/i0[9] ), .A2(\SB2_0_0/i0_3 ), .A3(
        \SB2_0_0/i0[8] ), .ZN(n1855) );
  NAND3_X1 U4349 ( .A1(\SB1_2_17/i0_4 ), .A2(\SB1_2_17/i1[9] ), .A3(
        \SB1_2_17/i1_5 ), .ZN(\SB1_2_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4351 ( .A1(\SB1_1_29/i0[10] ), .A2(\SB1_1_29/i0_0 ), .A3(
        \SB1_1_29/i0[6] ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4352 ( .A1(\SB3_30/i1[9] ), .A2(\SB3_30/i0[10] ), .A3(
        \SB3_30/i1_7 ), .ZN(\SB3_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4353 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i1_5 ), .A3(
        \SB4_28/i1[9] ), .ZN(\SB4_28/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4354 ( .A1(\SB1_3_11/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_3_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_3/NAND4_in[0] ), .A4(n1856), .ZN(
        \RI3[3][135] ) );
  NAND3_X1 U4355 ( .A1(\SB1_3_11/i0[8] ), .A2(\SB1_3_11/i3[0] ), .A3(
        \SB1_3_11/i1_5 ), .ZN(n1856) );
  NAND3_X1 U4356 ( .A1(\SB1_1_29/i0[10] ), .A2(\SB1_1_29/i1[9] ), .A3(
        \SB1_1_29/i1_7 ), .ZN(\SB1_1_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4357 ( .A1(\SB2_1_27/i0[10] ), .A2(\SB2_1_27/i0_0 ), .A3(
        \SB2_1_27/i0[6] ), .ZN(\SB2_1_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4358 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i0_0 ), .A3(
        \SB2_1_10/i0[6] ), .ZN(\SB2_1_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4359 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0_4 ), .A3(
        \SB2_1_24/i1[9] ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4360 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i0_3 ), .A3(
        \SB2_1_2/i1[9] ), .ZN(\SB2_1_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4361 ( .A1(n2106), .A2(\SB4_31/i0[7] ), .A3(\SB4_31/i0_0 ), .ZN(
        \SB4_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4362 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0[9] ), .A3(
        \SB2_2_20/i0[8] ), .ZN(\SB2_2_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4363 ( .A1(\SB1_0_29/i1_7 ), .A2(\SB1_0_29/i0_4 ), .A3(
        \SB1_0_29/i0[8] ), .ZN(\SB1_0_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4365 ( .A1(\SB2_0_24/i0_4 ), .A2(\SB2_0_24/i0_0 ), .A3(
        \SB2_0_24/i1_5 ), .ZN(n1857) );
  NAND4_X1 U4366 ( .A1(\SB1_2_16/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_16/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_16/Component_Function_2/NAND4_in[1] ), .A4(n1858), .ZN(
        \RI3[2][110] ) );
  NAND3_X1 U4369 ( .A1(\SB1_1_30/i1[9] ), .A2(\SB1_1_30/i0[10] ), .A3(
        \SB1_1_30/i1_7 ), .ZN(\SB1_1_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4370 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i0[9] ), .A3(
        \SB1_1_8/i0[8] ), .ZN(\SB1_1_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4371 ( .A1(\SB1_2_9/i0_0 ), .A2(\SB1_2_9/i0_4 ), .A3(
        \SB1_2_9/i1_5 ), .ZN(n903) );
  NAND3_X1 U4372 ( .A1(\SB1_1_18/i0_3 ), .A2(\SB1_1_18/i0[10] ), .A3(
        \SB1_1_18/i0_4 ), .ZN(\SB1_1_18/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U4373 ( .A1(\SB2_1_15/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_15/Component_Function_4/NAND4_in[1] ), .A4(n1859), .ZN(
        \RI5[1][106] ) );
  NAND3_X1 U4374 ( .A1(\SB2_1_15/i0_4 ), .A2(\SB2_1_15/i1_5 ), .A3(
        \SB2_1_15/i1[9] ), .ZN(n1859) );
  NAND3_X1 U4375 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i3[0] ), .A3(\SB4_19/i1_7 ), 
        .ZN(n1860) );
  XNOR2_X1 U4376 ( .A(n1862), .B(n1861), .ZN(\RI1[3][101] ) );
  XNOR2_X1 U4377 ( .A(\MC_ARK_ARC_1_2/temp1[101] ), .B(
        \MC_ARK_ARC_1_2/temp4[101] ), .ZN(n1861) );
  XNOR2_X1 U4378 ( .A(\MC_ARK_ARC_1_2/temp2[101] ), .B(
        \MC_ARK_ARC_1_2/temp3[101] ), .ZN(n1862) );
  XNOR2_X1 U4379 ( .A(n984), .B(n1863), .ZN(\RI1[2][89] ) );
  XNOR2_X1 U4380 ( .A(\MC_ARK_ARC_1_1/temp2[89] ), .B(
        \MC_ARK_ARC_1_1/temp4[89] ), .ZN(n1863) );
  NAND3_X1 U4381 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i0_4 ), .A3(
        \SB1_2_2/i1_5 ), .ZN(\SB1_2_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4382 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB2_3_25/i0_4 ), .A3(
        \SB2_3_25/i1[9] ), .ZN(\SB2_3_25/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U4384 ( .A(n1865), .B(n1864), .ZN(\RI1[2][155] ) );
  XNOR2_X1 U4385 ( .A(\MC_ARK_ARC_1_1/temp3[155] ), .B(
        \MC_ARK_ARC_1_1/temp4[155] ), .ZN(n1864) );
  XNOR2_X1 U4386 ( .A(\MC_ARK_ARC_1_1/temp1[155] ), .B(
        \MC_ARK_ARC_1_1/temp2[155] ), .ZN(n1865) );
  NAND3_X1 U4387 ( .A1(\SB4_22/i1_5 ), .A2(n779), .A3(\SB4_22/i0[6] ), .ZN(
        n1036) );
  NAND3_X1 U4389 ( .A1(\SB2_1_12/i0[8] ), .A2(\SB2_1_12/i1_5 ), .A3(
        \SB2_1_12/i3[0] ), .ZN(\SB2_1_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4390 ( .A1(\SB1_0_4/i0[6] ), .A2(\SB1_0_4/i0[9] ), .A3(
        \SB1_0_4/i0_4 ), .ZN(\SB1_0_4/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U4391 ( .A1(\SB2_2_14/i0[6] ), .A2(n1867), .ZN(n1866) );
  AND2_X1 U4392 ( .A1(\RI3[2][106] ), .A2(\RI3[2][102] ), .ZN(n1867) );
  XNOR2_X1 U4393 ( .A(n1868), .B(n416), .ZN(Ciphertext[109]) );
  NAND4_X1 U4394 ( .A1(\SB4_13/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_13/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_13/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_13/Component_Function_1/NAND4_in[2] ), .ZN(n1868) );
  NAND4_X1 U4395 ( .A1(\SB1_0_25/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_25/Component_Function_5/NAND4_in[3] ), .A4(n1869), .ZN(
        \RI3[0][41] ) );
  NAND3_X1 U4396 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0_4 ), .A3(
        \SB1_0_25/i1[9] ), .ZN(n1869) );
  NAND4_X1 U4399 ( .A1(\SB1_3_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_23/Component_Function_1/NAND4_in[0] ), .A4(n1871), .ZN(
        \RI3[3][73] ) );
  NAND3_X1 U4400 ( .A1(\SB1_3_23/i1_7 ), .A2(\SB1_3_23/i0_4 ), .A3(
        \SB1_3_23/i0[8] ), .ZN(n1871) );
  NAND3_X1 U4401 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i1[9] ), .A3(
        \SB1_3_19/i0[6] ), .ZN(\SB1_3_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4402 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i1[9] ), .A3(
        \SB1_1_8/i0[6] ), .ZN(\SB1_1_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4403 ( .A1(\SB2_1_21/i0_3 ), .A2(\SB2_1_21/i0_4 ), .A3(
        \SB2_1_21/i0_0 ), .ZN(\SB2_1_21/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U4404 ( .A1(\SB2_2_17/i0[6] ), .A2(n1872), .ZN(
        \SB2_2_17/Component_Function_5/NAND4_in[3] ) );
  AND2_X1 U4405 ( .A1(\RI3[2][88] ), .A2(\RI3[2][84] ), .ZN(n1872) );
  XNOR2_X1 U4406 ( .A(n1873), .B(n417), .ZN(Ciphertext[171]) );
  NAND4_X1 U4407 ( .A1(\SB4_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_3/Component_Function_3/NAND4_in[3] ), .ZN(n1873) );
  NAND4_X1 U4408 ( .A1(\SB4_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_1/Component_Function_3/NAND4_in[3] ), .A3(
        \SB4_1/Component_Function_3/NAND4_in[0] ), .A4(n1874), .ZN(
        \RI4[4][183] ) );
  NAND3_X1 U4409 ( .A1(\SB4_1/i0[10] ), .A2(\SB4_1/i1[9] ), .A3(\SB4_1/i1_7 ), 
        .ZN(n1874) );
  NAND4_X1 U4410 ( .A1(\SB3_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_14/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_14/Component_Function_0/NAND4_in[1] ), .A4(n1875), .ZN(
        \RI3[4][132] ) );
  NAND3_X1 U4411 ( .A1(\SB3_14/i0[7] ), .A2(\SB3_14/i0_0 ), .A3(n860), .ZN(
        n1875) );
  NAND4_X1 U4412 ( .A1(\SB1_1_2/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_2/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_1_2/Component_Function_4/NAND4_in[0] ), .A4(n1876), .ZN(
        \RI3[1][184] ) );
  NAND3_X1 U4413 ( .A1(\SB1_1_2/i0_3 ), .A2(\SB1_1_2/i0[10] ), .A3(
        \SB1_1_2/i0[9] ), .ZN(n1876) );
  NAND4_X2 U4414 ( .A1(\SB2_3_10/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_10/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_3_10/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_3_10/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[146] ) );
  NAND4_X1 U4415 ( .A1(\SB2_2_18/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_18/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_18/Component_Function_2/NAND4_in[0] ), .A4(n1877), .ZN(
        \RI5[2][98] ) );
  NAND3_X1 U4416 ( .A1(\SB2_2_18/i0_4 ), .A2(\SB2_2_18/i1_5 ), .A3(
        \SB2_2_18/i0_0 ), .ZN(n1877) );
  NAND3_X1 U4417 ( .A1(\SB2_1_30/i0_4 ), .A2(\SB2_1_30/i1_7 ), .A3(
        \SB2_1_30/i0[8] ), .ZN(\SB2_1_30/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 U4418 ( .A1(\SB2_3_1/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_3_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_1/Component_Function_5/NAND4_in[0] ), .A4(n1878), .ZN(
        \RI5[3][185] ) );
  NAND3_X1 U4419 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i1[9] ), .A3(
        \SB2_3_1/i0_4 ), .ZN(n1878) );
  XNOR2_X1 U4420 ( .A(n1879), .B(n235), .ZN(Ciphertext[9]) );
  NAND4_X1 U4421 ( .A1(\SB4_30/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_30/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_30/Component_Function_3/NAND4_in[3] ), .A4(
        \SB4_30/Component_Function_3/NAND4_in[2] ), .ZN(n1879) );
  NAND3_X1 U4422 ( .A1(n2131), .A2(\SB4_29/i0_3 ), .A3(\SB4_29/i0_0 ), .ZN(
        \SB4_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4423 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i1[9] ), .A3(
        \SB4_10/i1_7 ), .ZN(n1880) );
  NAND3_X1 U4424 ( .A1(\SB4_18/i0_3 ), .A2(\SB4_18/i0_0 ), .A3(\SB4_18/i0[7] ), 
        .ZN(\SB4_18/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U4425 ( .A(\MC_ARK_ARC_1_3/temp6[82] ), .B(n1881), .ZN(\RI1[4][82] ) );
  XNOR2_X1 U4426 ( .A(\MC_ARK_ARC_1_3/temp2[82] ), .B(
        \MC_ARK_ARC_1_3/temp1[82] ), .ZN(n1881) );
  XNOR2_X1 U4427 ( .A(\MC_ARK_ARC_1_1/temp6[51] ), .B(n1882), .ZN(\RI1[2][51] ) );
  XNOR2_X1 U4428 ( .A(\MC_ARK_ARC_1_1/temp1[51] ), .B(
        \MC_ARK_ARC_1_1/temp2[51] ), .ZN(n1882) );
  NAND3_X1 U4430 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i1_7 ), .A3(\SB4_16/i3[0] ), 
        .ZN(\SB4_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4432 ( .A1(\SB2_1_7/i0_3 ), .A2(\SB2_1_7/i0_4 ), .A3(
        \SB2_1_7/i1[9] ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4433 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i1[9] ), .A3(
        \SB1_1_7/i0_4 ), .ZN(n1912) );
  NAND3_X1 U4434 ( .A1(\SB2_1_30/i0[10] ), .A2(\SB2_1_30/i0_0 ), .A3(
        \SB2_1_30/i0[6] ), .ZN(\SB2_1_30/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4435 ( .A1(\SB4_6/i0_4 ), .A2(\SB4_6/i0_3 ), .A3(\SB4_6/i0_0 ), 
        .ZN(\SB4_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4436 ( .A1(\SB4_18/i0_4 ), .A2(\SB4_18/i0_0 ), .A3(\SB4_18/i0_3 ), 
        .ZN(\SB4_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4437 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i1_5 ), .A3(
        \SB2_0_27/i1[9] ), .ZN(\SB2_0_27/Component_Function_2/NAND4_in[0] ) );
  OR3_X1 U4438 ( .A1(\RI1[2][84] ), .A2(\RI1[2][85] ), .A3(\RI1[2][88] ), .ZN(
        \SB1_2_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4439 ( .A1(\SB2_0_15/i0_3 ), .A2(\SB2_0_15/i0[10] ), .A3(
        \SB2_0_15/i0[9] ), .ZN(\SB2_0_15/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4440 ( .A1(n2148), .A2(\SB4_13/i1[9] ), .A3(\SB4_13/i0_4 ), .ZN(
        \SB4_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4441 ( .A1(\SB1_2_21/i0_4 ), .A2(\SB1_2_21/i1_7 ), .A3(
        \SB1_2_21/i0[8] ), .ZN(\SB1_2_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4442 ( .A1(\SB1_0_1/i0_3 ), .A2(\SB1_0_1/i0[10] ), .A3(
        \SB1_0_1/i0[9] ), .ZN(\SB1_0_1/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U4443 ( .A(n1884), .B(n258), .ZN(Ciphertext[115]) );
  NAND4_X1 U4444 ( .A1(\SB4_12/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_12/Component_Function_1/NAND4_in[0] ), .A3(n1923), .A4(
        \SB4_12/Component_Function_1/NAND4_in[2] ), .ZN(n1884) );
  NAND3_X1 U4445 ( .A1(\SB1_2_0/i0_3 ), .A2(\SB1_2_0/i0[9] ), .A3(
        \SB1_2_0/i0[8] ), .ZN(\SB1_2_0/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U4446 ( .A(n1885), .B(n251), .ZN(Ciphertext[20]) );
  XNOR2_X1 U4447 ( .A(n1886), .B(n308), .ZN(Ciphertext[135]) );
  NAND4_X1 U4448 ( .A1(\SB4_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_9/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_9/Component_Function_3/NAND4_in[3] ), .A4(
        \SB4_9/Component_Function_3/NAND4_in[2] ), .ZN(n1886) );
  NAND3_X1 U4450 ( .A1(\SB1_0_4/i0[6] ), .A2(\SB1_0_4/i1_5 ), .A3(
        \SB1_0_4/i0[9] ), .ZN(\SB1_0_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4451 ( .A1(\SB4_11/i0_0 ), .A2(n805), .A3(\SB4_11/i1_5 ), .ZN(
        n1039) );
  XNOR2_X1 U4452 ( .A(n1887), .B(n277), .ZN(Ciphertext[126]) );
  NAND4_X1 U4453 ( .A1(\SB4_10/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_10/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_10/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_10/Component_Function_0/NAND4_in[0] ), .ZN(n1887) );
  NAND3_X1 U4454 ( .A1(\SB3_28/i0[10] ), .A2(\SB3_28/i0_0 ), .A3(
        \SB3_28/i0[6] ), .ZN(\SB3_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4455 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0[10] ), .A3(
        \SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U4456 ( .A(n1889), .B(n1888), .ZN(\RI1[1][161] ) );
  XNOR2_X1 U4457 ( .A(\MC_ARK_ARC_1_0/temp1[161] ), .B(
        \MC_ARK_ARC_1_0/temp4[161] ), .ZN(n1888) );
  XNOR2_X1 U4458 ( .A(\MC_ARK_ARC_1_0/temp3[161] ), .B(
        \MC_ARK_ARC_1_0/temp2[161] ), .ZN(n1889) );
  XNOR2_X1 U4460 ( .A(n1891), .B(n209), .ZN(Ciphertext[95]) );
  NAND4_X1 U4461 ( .A1(\SB4_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_16/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_16/Component_Function_5/NAND4_in[0] ), .ZN(n1891) );
  INV_X1 U4462 ( .A(\RI1[4][88] ), .ZN(\SB3_17/i0_4 ) );
  XNOR2_X1 U4463 ( .A(\MC_ARK_ARC_1_3/temp6[88] ), .B(
        \MC_ARK_ARC_1_3/temp5[88] ), .ZN(\RI1[4][88] ) );
  NAND3_X1 U4466 ( .A1(\SB1_0_11/i0[7] ), .A2(\SB1_0_11/i0_0 ), .A3(
        \SB1_0_11/i0_3 ), .ZN(\SB1_0_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4467 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i1_5 ), .A3(\SB4_12/i0_0 ), 
        .ZN(n1893) );
  NAND3_X1 U4468 ( .A1(n1964), .A2(\SB4_31/i0[10] ), .A3(\SB4_31/i1[9] ), .ZN(
        n1894) );
  NAND3_X1 U4469 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0_0 ), .A3(
        \SB2_1_30/i0_4 ), .ZN(\SB2_1_30/Component_Function_3/NAND4_in[1] ) );
  XNOR2_X1 U4470 ( .A(n1895), .B(n201), .ZN(Ciphertext[151]) );
  NAND4_X1 U4471 ( .A1(\SB4_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_6/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_6/Component_Function_1/NAND4_in[2] ), .ZN(n1895) );
  NAND3_X1 U4472 ( .A1(\SB1_2_19/i0_3 ), .A2(\SB1_2_19/i0[9] ), .A3(
        \SB1_2_19/i0[8] ), .ZN(\SB1_2_19/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U4473 ( .A1(\SB1_1_6/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_6/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_6/Component_Function_5/NAND4_in[0] ), .A4(n1896), .ZN(
        \RI3[1][155] ) );
  NAND3_X1 U4474 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0_4 ), .A3(
        \SB1_1_6/i1[9] ), .ZN(n1896) );
  NAND3_X1 U4475 ( .A1(\SB4_9/i0_3 ), .A2(\RI3[4][136] ), .A3(\SB4_9/i0[10] ), 
        .ZN(\SB4_9/Component_Function_0/NAND4_in[2] ) );
  XNOR2_X1 U4477 ( .A(n1897), .B(n280), .ZN(Ciphertext[57]) );
  NAND4_X1 U4478 ( .A1(\SB4_22/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_22/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_22/Component_Function_3/NAND4_in[3] ), .A4(
        \SB4_22/Component_Function_3/NAND4_in[2] ), .ZN(n1897) );
  NAND3_X1 U4479 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0[10] ), .A3(
        \SB1_0_22/i0[9] ), .ZN(\SB1_0_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4480 ( .A1(\SB2_2_28/i3[0] ), .A2(\SB2_2_28/i1_5 ), .A3(
        \SB2_2_28/i0[8] ), .ZN(\SB2_2_28/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U4482 ( .A(\RI1[1][92] ), .ZN(\SB1_1_16/i0_0 ) );
  XNOR2_X1 U4483 ( .A(\MC_ARK_ARC_1_0/temp5[92] ), .B(
        \MC_ARK_ARC_1_0/temp6[92] ), .ZN(\RI1[1][92] ) );
  INV_X2 U4484 ( .A(\RI1[3][11] ), .ZN(\SB1_3_30/i0_3 ) );
  XNOR2_X1 U4485 ( .A(\MC_ARK_ARC_1_2/temp6[11] ), .B(
        \MC_ARK_ARC_1_2/temp5[11] ), .ZN(\RI1[3][11] ) );
  NAND4_X1 U4486 ( .A1(\SB1_2_10/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_10/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_10/Component_Function_0/NAND4_in[1] ), .A4(n1898), .ZN(
        \RI3[2][156] ) );
  NAND3_X1 U4487 ( .A1(\SB1_2_10/i0_3 ), .A2(\SB1_2_10/i0[10] ), .A3(
        \SB1_2_10/i0_4 ), .ZN(n1898) );
  NAND4_X1 U4488 ( .A1(\SB1_1_16/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_16/Component_Function_4/NAND4_in[2] ), .A4(n1899), .ZN(
        \RI3[1][100] ) );
  NAND3_X1 U4489 ( .A1(\SB1_1_16/i1[9] ), .A2(\SB1_1_16/i1_5 ), .A3(
        \SB1_1_16/i0_4 ), .ZN(n1899) );
  NAND3_X1 U4490 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0[10] ), .A3(
        \SB1_0_15/i0_4 ), .ZN(\SB1_0_15/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U4491 ( .A1(\SB1_3_19/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_3_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_3/NAND4_in[0] ), .A4(n1900), .ZN(
        \RI3[3][87] ) );
  NAND3_X1 U4492 ( .A1(\SB1_3_19/i3[0] ), .A2(\SB1_3_19/i1_5 ), .A3(
        \SB1_3_19/i0[8] ), .ZN(n1900) );
  XNOR2_X1 U4493 ( .A(n1901), .B(n415), .ZN(Ciphertext[104]) );
  NAND4_X1 U4494 ( .A1(\SB4_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_14/Component_Function_2/NAND4_in[1] ), .A3(n769), .A4(
        \SB4_14/Component_Function_2/NAND4_in[0] ), .ZN(n1901) );
  XNOR2_X1 U4495 ( .A(n1350), .B(n1349), .ZN(\RI1[4][77] ) );
  NAND3_X1 U4496 ( .A1(\SB1_0_30/i0_3 ), .A2(\SB1_0_30/i0[9] ), .A3(
        \SB1_0_30/i0[8] ), .ZN(\SB1_0_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4497 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i0[10] ), .A3(
        \SB1_1_8/i0[9] ), .ZN(\SB1_1_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4498 ( .A1(\SB1_0_11/i1_7 ), .A2(\SB1_0_11/i0_4 ), .A3(
        \SB1_0_11/i0[8] ), .ZN(\SB1_0_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4499 ( .A1(\SB2_1_13/i0_3 ), .A2(\RI3[1][108] ), .A3(
        \SB2_1_13/i0[8] ), .ZN(\SB2_1_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4500 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i1_5 ), .A3(
        \SB2_1_5/i1[9] ), .ZN(\SB2_1_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4502 ( .A1(\SB2_0_10/i3[0] ), .A2(\SB2_0_10/i1_5 ), .A3(
        \SB2_0_10/i0[8] ), .ZN(n1902) );
  XNOR2_X1 U4503 ( .A(\MC_ARK_ARC_1_2/temp5[63] ), .B(n1903), .ZN(\RI1[3][63] ) );
  XNOR2_X1 U4504 ( .A(\MC_ARK_ARC_1_2/temp3[63] ), .B(
        \MC_ARK_ARC_1_2/temp4[63] ), .ZN(n1903) );
  NAND4_X1 U4505 ( .A1(\SB2_2_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_20/Component_Function_3/NAND4_in[2] ), .A3(n923), .A4(n1904), 
        .ZN(\RI5[2][81] ) );
  NAND3_X1 U4506 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0_0 ), .A3(
        \SB2_2_20/i0_4 ), .ZN(n1904) );
  XNOR2_X1 U4507 ( .A(n1905), .B(n292), .ZN(Ciphertext[14]) );
  NAND3_X1 U4508 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0_0 ), .A3(
        \SB1_0_11/i0_4 ), .ZN(\SB1_0_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4509 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0_3 ), .A3(
        \SB3_31/i0[10] ), .ZN(\SB3_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4510 ( .A1(\SB1_0_26/i1_5 ), .A2(\SB1_0_26/i1[9] ), .A3(
        \SB1_0_26/i0_4 ), .ZN(\SB1_0_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4511 ( .A1(\SB1_0_31/i0_3 ), .A2(\SB1_0_31/i1[9] ), .A3(
        \SB1_0_31/i0_4 ), .ZN(\SB1_0_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4512 ( .A1(\SB4_6/i0_4 ), .A2(\SB4_6/i1[9] ), .A3(\SB4_6/i1_5 ), 
        .ZN(\SB4_6/Component_Function_4/NAND4_in[3] ) );
  NAND4_X1 U4513 ( .A1(\SB4_16/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_16/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_16/Component_Function_2/NAND4_in[3] ), .A4(n1906), .ZN(n1392) );
  NAND3_X1 U4514 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i1_5 ), .A3(
        \SB4_16/i1[9] ), .ZN(n1906) );
  NAND4_X1 U4515 ( .A1(\SB4_18/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_18/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_18/Component_Function_5/NAND4_in[0] ), .A4(n1907), .ZN(n765) );
  NAND3_X1 U4516 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i0_0 ), .A3(
        \SB4_18/i0[6] ), .ZN(n1907) );
  NAND3_X1 U4517 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0[9] ), .A3(
        \SB2_2_19/i0[8] ), .ZN(\SB2_2_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4518 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0[9] ), .A3(
        \SB2_1_30/i0[8] ), .ZN(\SB2_1_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4519 ( .A1(\SB2_0_15/i0_3 ), .A2(\SB2_0_15/i1[9] ), .A3(
        \SB2_0_15/i0[6] ), .ZN(\SB2_0_15/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U4520 ( .A1(\SB2_0_8/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_8/Component_Function_4/NAND4_in[1] ), .A4(n1908), .ZN(
        \RI5[0][148] ) );
  NAND3_X1 U4521 ( .A1(\SB2_0_8/i0_3 ), .A2(\SB2_0_8/i0[9] ), .A3(
        \SB2_0_8/i0[10] ), .ZN(n1908) );
  NAND3_X1 U4522 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i0_3 ), .A3(\SB4_10/i0_4 ), 
        .ZN(n1909) );
  NAND3_X1 U4525 ( .A1(\SB2_1_15/i0[10] ), .A2(\SB2_1_15/i1_5 ), .A3(
        \SB2_1_15/i1[9] ), .ZN(\SB2_1_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4526 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i0_4 ), .A3(
        \SB2_0_23/i1[9] ), .ZN(n767) );
  NAND3_X1 U4527 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0[9] ), .A3(\SB3_19/i0[8] ), .ZN(\SB3_19/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U4528 ( .A1(\SB1_0_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_22/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_22/Component_Function_1/NAND4_in[0] ), .A4(n1911), .ZN(
        \RI3[0][79] ) );
  NAND3_X1 U4529 ( .A1(\SB1_0_22/i1_7 ), .A2(\SB1_0_22/i0_4 ), .A3(
        \SB1_0_22/i0[8] ), .ZN(n1911) );
  NAND4_X1 U4530 ( .A1(\SB1_1_7/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_1_7/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_5/NAND4_in[0] ), .A4(n1912), .ZN(
        \RI3[1][149] ) );
  NAND3_X1 U4531 ( .A1(\SB2_3_18/i0[10] ), .A2(\SB2_3_18/i0_3 ), .A3(
        \SB2_3_18/i0[9] ), .ZN(\SB2_3_18/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U4532 ( .A(n1913), .B(n316), .ZN(Ciphertext[79]) );
  NAND4_X1 U4533 ( .A1(\SB4_18/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_18/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_18/Component_Function_1/NAND4_in[0] ), .ZN(n1913) );
  NAND3_X1 U4534 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i1[9] ), .A3(
        \SB4_17/i1_7 ), .ZN(n1914) );
  NAND3_X1 U4535 ( .A1(\SB1_1_31/i0_3 ), .A2(\SB1_1_31/i0[10] ), .A3(
        \SB1_1_31/i0[9] ), .ZN(\SB1_1_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4537 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i1_7 ), .A3(\SB4_5/i3[0] ), 
        .ZN(n1915) );
  NAND4_X1 U4538 ( .A1(\SB4_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_8/Component_Function_1/NAND4_in[0] ), .A3(n1320), .A4(n1916), 
        .ZN(n914) );
  NAND3_X1 U4539 ( .A1(\SB4_8/i0[9] ), .A2(\SB4_8/i1_5 ), .A3(\SB4_8/i0[6] ), 
        .ZN(n1916) );
  NAND3_X1 U4540 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i3[0] ), .A3(\SB4_10/i1_7 ), 
        .ZN(\SB4_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4541 ( .A1(\SB1_0_4/i0_3 ), .A2(\SB1_0_4/i0[10] ), .A3(
        \SB1_0_4/i0[9] ), .ZN(\SB1_0_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4542 ( .A1(\SB4_11/i0[6] ), .A2(\SB4_11/i0[9] ), .A3(n805), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U4543 ( .A1(\SB3_12/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_12/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_12/Component_Function_4/NAND4_in[3] ), .A4(
        \SB3_12/Component_Function_4/NAND4_in[1] ), .ZN(n805) );
  NAND4_X2 U4544 ( .A1(\SB2_3_17/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_17/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[104] ) );
  NAND3_X1 U4545 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[9] ), .A3(
        \SB1_3_31/i0[8] ), .ZN(\SB1_3_31/Component_Function_2/NAND4_in[2] ) );
  XNOR2_X1 U4546 ( .A(n1918), .B(n1917), .ZN(\RI1[3][77] ) );
  XNOR2_X1 U4547 ( .A(\MC_ARK_ARC_1_2/temp2[77] ), .B(
        \MC_ARK_ARC_1_2/temp4[77] ), .ZN(n1917) );
  XNOR2_X1 U4548 ( .A(\MC_ARK_ARC_1_2/temp1[77] ), .B(
        \MC_ARK_ARC_1_2/temp3[77] ), .ZN(n1918) );
  NAND3_X1 U4550 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i1[9] ), .A3(
        \SB1_1_0/i1_7 ), .ZN(\SB1_1_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4552 ( .A1(\SB2_1_2/i0[9] ), .A2(\SB2_1_2/i0_3 ), .A3(
        \SB2_1_2/i0[8] ), .ZN(\SB2_1_2/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U4553 ( .A1(\SB1_1_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_30/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_2/NAND4_in[2] ), .A4(n1920), .ZN(
        \RI3[1][26] ) );
  NAND3_X1 U4554 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0_0 ), .A3(
        \SB1_0_25/i0_4 ), .ZN(\SB1_0_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4555 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i1[9] ), .A3(
        \SB1_1_4/i1_5 ), .ZN(\SB1_1_4/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4556 ( .A1(\SB4_29/Component_Function_4/NAND4_in[2] ), .A2(n773), 
        .A3(\SB4_29/Component_Function_4/NAND4_in[1] ), .A4(n1921), .ZN(n1924)
         );
  NAND4_X1 U4557 ( .A1(\SB4_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_3/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_3/Component_Function_5/NAND4_in[0] ), .A4(n1922), .ZN(n1003) );
  NAND3_X1 U4558 ( .A1(\SB4_3/i0[10] ), .A2(\SB4_3/i0_0 ), .A3(\SB4_3/i0[6] ), 
        .ZN(n1922) );
  NAND3_X1 U4559 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i0[8] ), .A3(\SB4_12/i1_7 ), 
        .ZN(n1923) );
  NAND3_X1 U4560 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0_4 ), .A3(
        \SB1_0_9/i1[9] ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4561 ( .A1(\SB3_12/i0[10] ), .A2(\SB3_12/i0_3 ), .A3(\SB3_12/i0_4 ), .ZN(\SB3_12/Component_Function_0/NAND4_in[2] ) );
  XNOR2_X1 U4562 ( .A(n1924), .B(n279), .ZN(Ciphertext[16]) );
  NAND4_X2 U4563 ( .A1(\SB1_0_24/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_24/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_0_24/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_0_24/Component_Function_4/NAND4_in[0] ), .ZN(\SB2_0_23/i0_4 ) );
  NAND3_X1 U4564 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i1[9] ), .A3(\SB4_13/i0[6] ), .ZN(\SB4_13/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U4565 ( .A1(\SB2_2_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_18/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[2][108] ) );
  NAND4_X2 U4566 ( .A1(\SB1_3_17/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_17/Component_Function_4/NAND4_in[0] ), .A3(n734), .A4(
        \SB1_3_17/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[3][94] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_3/BUF_88  ( .A(\RI5[3][88] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[88] ) );
  BUF_X2 U924 ( .A(\RI3[3][173] ), .Z(\SB2_3_3/i0_3 ) );
  BUF_X2 \SB2_3_2/BUF_5  ( .A(\RI3[3][179] ), .Z(\SB2_3_2/i0_3 ) );
  BUF_X2 U933 ( .A(\RI3[1][173] ), .Z(\SB2_1_3/i0_3 ) );
  BUF_X2 \SB2_2_26/BUF_1  ( .A(\RI3[2][31] ), .Z(\SB2_2_26/i0[6] ) );
  NAND4_X4 \SB2_1_11/Component_Function_3/N5  ( .A1(
        \SB2_1_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_11/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][135] ) );
  NAND4_X4 U1064 ( .A1(\SB2_1_8/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_8/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_1_8/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_8/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[148] ) );
  INV_X1 U516 ( .A(n427), .ZN(n363) );
  NAND4_X2 U1549 ( .A1(\SB3_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_1/Component_Function_1/NAND4_in[3] ), .ZN(n791) );
  BUF_X1 \SB1_1_28/BUF_1  ( .A(\RI1[1][19] ), .Z(\SB1_1_28/i1_7 ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_122  ( .A(\RI5[2][122] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[122] ) );
  BUF_X2 \SB1_2_16/BUF_3  ( .A(\RI1[2][93] ), .Z(\SB1_2_16/i0[8] ) );
  BUF_X2 \SB2_0_16/BUF_0  ( .A(\RI3[0][90] ), .Z(\SB2_0_16/i0[9] ) );
  NAND4_X2 U4481 ( .A1(\SB2_1_16/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_16/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_16/Component_Function_3/NAND4_in[2] ), .A4(n771), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[105] ) );
  BUF_X2 U1248 ( .A(\RI3[0][156] ), .Z(\SB2_0_5/i0[9] ) );
  BUF_X2 \SB2_3_3/BUF_0  ( .A(\RI3[3][168] ), .Z(\SB2_3_3/i0[9] ) );
  BUF_X1 \SB1_3_23/BUF_1  ( .A(\RI1[3][49] ), .Z(\SB1_3_23/i1_7 ) );
  BUF_X1 U1357 ( .A(\RI1[3][169] ), .Z(\SB1_3_3/i1_7 ) );
  BUF_X2 \SB2_3_31/BUF_1  ( .A(\RI3[3][1] ), .Z(\SB2_3_31/i0[6] ) );
  BUF_X2 \SB2_0_0/BUF_0  ( .A(\RI3[0][186] ), .Z(\SB2_0_0/i0[9] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_86  ( .A(\RI5[2][86] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[86] ) );
  NAND4_X2 U2269 ( .A1(\SB2_3_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_18/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[83] ) );
  INV_X1 U144 ( .A(\MC_ARK_ARC_1_0/buf_keyinput[95] ), .ZN(n285) );
  BUF_X1 \SB1_3_31/BUF_1  ( .A(\RI1[3][1] ), .Z(\SB1_3_31/i1_7 ) );
  BUF_X2 \SB2_0_18/BUF_1  ( .A(\RI3[0][79] ), .Z(\SB2_0_18/i0[6] ) );
  BUF_X1 U602 ( .A(\MC_ARK_ARC_1_1/buf_datainput[191] ), .Z(n514) );
  BUF_X2 U1349 ( .A(\RI3[2][133] ), .Z(\SB2_2_9/i0[6] ) );
  BUF_X2 \SB1_1_26/BUF_3  ( .A(\RI1[1][33] ), .Z(\SB1_1_26/i0[8] ) );
  BUF_X2 \SB2_2_24/BUF_0  ( .A(\RI3[2][42] ), .Z(\SB2_2_24/i0[9] ) );
  BUF_X2 U972 ( .A(\RI1[3][2] ), .Z(\SB1_3_31/i1[9] ) );
  BUF_X1 \SB1_0_8/BUF_1  ( .A(n53), .Z(\SB1_0_8/i1_7 ) );
  BUF_X2 \SB4_1/BUF_0  ( .A(\RI3[4][180] ), .Z(\SB4_1/i0[9] ) );
  INV_X1 U1215 ( .A(n154), .ZN(\SB1_0_25/i0_0 ) );
  NAND4_X2 U2680 ( .A1(\SB2_1_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_21/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[65] ) );
  INV_X1 \SB1_0_10/INV_5  ( .A(n61), .ZN(\SB1_0_10/i0_3 ) );
  INV_X1 U1421 ( .A(n398), .ZN(n364) );
  INV_X1 U223 ( .A(\MC_ARK_ARC_1_0/buf_keyinput[187] ), .ZN(n221) );
  INV_X1 U231 ( .A(n496), .ZN(n326) );
  INV_X1 U511 ( .A(n462), .ZN(n331) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_136  ( .A(\RI5[0][136] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[136] ) );
  BUF_X1 U3718 ( .A(Key[173]), .Z(n405) );
  BUF_X2 \SB2_2_22/BUF_0  ( .A(\RI3[2][54] ), .Z(\SB2_2_22/i0[9] ) );
  INV_X1 U304 ( .A(n460), .ZN(n343) );
  BUF_X2 \SB2_3_31/BUF_2  ( .A(\RI3[3][2] ), .Z(\SB2_3_31/i0_0 ) );
  BUF_X1 \SB1_2_6/BUF_4  ( .A(\RI1[2][154] ), .Z(\SB1_2_6/i0[7] ) );
  BUF_X1 \SB1_1_20/BUF_1  ( .A(\RI1[1][67] ), .Z(\SB1_1_20/i1_7 ) );
  BUF_X2 \SB2_3_23/BUF_0  ( .A(\RI3[3][48] ), .Z(\SB2_3_23/i0[9] ) );
  BUF_X2 \SB2_0_9/BUF_1  ( .A(\RI3[0][133] ), .Z(\SB2_0_9/i0[6] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_118  ( .A(\RI5[0][118] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[118] ) );
  BUF_X2 U1627 ( .A(\RI5[3][149] ), .Z(n849) );
  BUF_X1 \SB1_1_18/BUF_1  ( .A(\RI1[1][79] ), .Z(\SB1_1_18/i1_7 ) );
  NAND4_X4 U2891 ( .A1(\SB2_3_23/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_23/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_23/Component_Function_5/NAND4_in[1] ), .A4(n1246), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[53] ) );
  BUF_X2 \SB2_0_15/BUF_0  ( .A(\RI3[0][96] ), .Z(\SB2_0_15/i0[9] ) );
  NAND4_X2 U1879 ( .A1(\SB2_0_11/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_11/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_0_11/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_11/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[140] ) );
  BUF_X2 \SB2_0_26/BUF_1  ( .A(\RI3[0][31] ), .Z(\SB2_0_26/i0[6] ) );
  BUF_X2 U1255 ( .A(\RI1[1][189] ), .Z(\SB1_1_0/i0[8] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_100  ( .A(\RI5[2][100] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[100] ) );
  BUF_X1 \SB1_2_19/BUF_1  ( .A(\RI1[2][73] ), .Z(\SB1_2_19/i1_7 ) );
  NAND4_X4 \SB2_2_22/Component_Function_3/N5  ( .A1(
        \SB2_2_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_22/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][69] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_33  ( .A(\RI5[0][33] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[33] ) );
  BUF_X2 U1674 ( .A(\RI3[4][149] ), .Z(n877) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_93  ( .A(\RI5[0][93] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[93] ) );
  NAND4_X4 \SB2_2_7/Component_Function_3/N5  ( .A1(
        \SB2_2_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_7/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_7/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][159] ) );
  NAND4_X2 \SB2_2_27/Component_Function_3/N5  ( .A1(
        \SB2_2_27/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_27/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_27/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][39] ) );
  NAND4_X2 U693 ( .A1(\SB2_1_4/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_4/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_4/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[167] ) );
  BUF_X1 U780 ( .A(\MC_ARK_ARC_1_1/buf_datainput[41] ), .Z(n1497) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_142  ( .A(\RI5[2][142] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[142] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_44  ( .A(\RI5[2][44] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[44] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_171  ( .A(\RI5[0][171] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[171] ) );
  NAND4_X2 U1677 ( .A1(\SB2_1_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_16/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[95] ) );
  BUF_X1 \SB1_1_24/BUF_0  ( .A(\RI1[1][42] ), .Z(\SB1_1_24/i3[0] ) );
  NAND4_X4 U932 ( .A1(n1172), .A2(\SB2_1_22/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_1_22/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_22/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[59] ) );
  NAND4_X2 U1860 ( .A1(n1397), .A2(\SB2_0_13/Component_Function_5/NAND4_in[3] ), .A3(\SB2_0_13/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_13/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[113] ) );
  NAND4_X2 U3771 ( .A1(\SB2_1_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_8/Component_Function_3/NAND4_in[2] ), .A4(n1047), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[153] ) );
  INV_X1 U113 ( .A(Key[121]), .ZN(n259) );
  CLKBUF_X1 U255 ( .A(Key[141]), .Z(n513) );
  CLKBUF_X1 U1186 ( .A(Key[111]), .Z(n509) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_177_0  ( .A(Key[132]), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[177] ) );
  CLKBUF_X1 U78 ( .A(Key[116]), .Z(n467) );
  CLKBUF_X1 U94 ( .A(Key[178]), .Z(n436) );
  CLKBUF_X1 U556 ( .A(Key[189]), .Z(\MC_ARK_ARC_1_0/buf_keyinput[136] ) );
  CLKBUF_X1 U51 ( .A(Key[106]), .Z(n446) );
  CLKBUF_X1 U95 ( .A(Key[105]), .Z(n495) );
  CLKBUF_X1 U267 ( .A(Key[40]), .Z(n469) );
  CLKBUF_X1 U273 ( .A(Key[75]), .Z(n502) );
  INV_X1 U210 ( .A(n456), .ZN(n365) );
  BUF_X1 U928 ( .A(n64), .Z(\SB1_0_10/i1[9] ) );
  INV_X1 \SB1_0_13/INV_4  ( .A(n80), .ZN(\SB1_0_13/i0_4 ) );
  INV_X1 \SB1_0_0/INV_4  ( .A(n2), .ZN(\SB1_0_0/i0_4 ) );
  BUF_X1 \SB1_0_25/BUF_3  ( .A(n153), .Z(\SB1_0_25/i0[8] ) );
  BUF_X1 \SB1_0_0/BUF_3  ( .A(n3), .Z(\SB1_0_0/i0[8] ) );
  BUF_X1 \SB1_0_25/BUF_2  ( .A(n154), .Z(\SB1_0_25/i1[9] ) );
  INV_X1 \SB1_0_12/INV_0  ( .A(n78), .ZN(\SB1_0_12/i0[9] ) );
  BUF_X1 U700 ( .A(n39), .Z(\SB1_0_6/i0[8] ) );
  INV_X1 \SB1_0_23/INV_0  ( .A(n144), .ZN(\SB1_0_23/i0[9] ) );
  INV_X1 \SB1_0_12/INV_4  ( .A(n74), .ZN(\SB1_0_12/i0_4 ) );
  INV_X1 \SB1_0_23/INV_2  ( .A(n142), .ZN(\SB1_0_23/i0_0 ) );
  BUF_X1 \SB1_0_23/BUF_2  ( .A(n142), .Z(\SB1_0_23/i1[9] ) );
  NAND4_X1 \SB1_0_16/Component_Function_0/N5  ( .A1(
        \SB1_0_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_16/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_16/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_16/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][120] ) );
  BUF_X1 \SB2_0_11/BUF_0  ( .A(\RI3[0][120] ), .Z(\SB2_0_11/i0[9] ) );
  BUF_X1 \SB2_0_15/BUF_1  ( .A(\RI3[0][97] ), .Z(\SB2_0_15/i0[6] ) );
  BUF_X1 \SB2_0_30/BUF_1  ( .A(\RI3[0][7] ), .Z(\SB2_0_30/i0[6] ) );
  BUF_X1 U542 ( .A(\RI3[0][139] ), .Z(\SB2_0_8/i0[6] ) );
  BUF_X1 \SB2_0_2/BUF_1  ( .A(\RI3[0][175] ), .Z(\SB2_0_2/i0[6] ) );
  BUF_X2 \SB2_0_14/BUF_4  ( .A(\RI3[0][106] ), .Z(\SB2_0_14/i0_4 ) );
  BUF_X1 \SB2_0_14/BUF_1  ( .A(\RI3[0][103] ), .Z(\SB2_0_14/i0[6] ) );
  BUF_X1 U1161 ( .A(\RI3[0][145] ), .Z(\SB2_0_7/i0[6] ) );
  BUF_X1 \SB2_0_29/BUF_1  ( .A(\RI3[0][13] ), .Z(\SB2_0_29/i0[6] ) );
  BUF_X1 \SB2_0_21/BUF_1  ( .A(\RI3[0][61] ), .Z(\SB2_0_21/i0[6] ) );
  BUF_X1 \SB2_0_6/BUF_1  ( .A(\RI3[0][151] ), .Z(\SB2_0_6/i0[6] ) );
  BUF_X2 \SB2_0_1/BUF_3  ( .A(\RI3[0][183] ), .Z(\SB2_0_1/i0[10] ) );
  BUF_X1 \SB2_0_25/BUF_1  ( .A(\RI3[0][37] ), .Z(\SB2_0_25/i0[6] ) );
  NAND4_X2 U3866 ( .A1(n1358), .A2(\SB2_0_28/Component_Function_5/NAND4_in[3] ), .A3(\SB2_0_28/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[23] ) );
  NAND4_X1 U3479 ( .A1(n767), .A2(\SB2_0_23/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_0_23/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_23/Component_Function_5/NAND4_in[3] ), .ZN(n1632) );
  NAND4_X2 \SB2_0_3/Component_Function_4/N5  ( .A1(
        \SB2_0_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_3/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_3/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_0_3/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][178] ) );
  NAND4_X2 U2595 ( .A1(n1704), .A2(\SB2_0_16/Component_Function_4/NAND4_in[0] ), .A3(\SB2_0_16/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_0_16/Component_Function_4/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[100] ) );
  NAND4_X2 U3758 ( .A1(\SB2_0_22/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_22/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_22/Component_Function_2/NAND4_in[0] ), .A4(n1674), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[74] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_129  ( .A(\RI5[0][129] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[129] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_22  ( .A(\RI5[0][22] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[22] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_172  ( .A(\RI5[0][172] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[172] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_134  ( .A(\RI5[0][134] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[134] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_148  ( .A(\RI5[0][148] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[148] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_92  ( .A(\RI5[0][92] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[92] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_176  ( .A(\RI5[0][176] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[176] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_7  ( .A(\RI5[0][7] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[7] ) );
  BUF_X1 \SB1_1_18/BUF_3  ( .A(\RI1[1][81] ), .Z(\SB1_1_18/i0[8] ) );
  BUF_X1 U657 ( .A(\RI1[1][62] ), .Z(\SB1_1_21/i1[9] ) );
  BUF_X1 U1125 ( .A(\RI1[1][57] ), .Z(\SB1_1_22/i0[8] ) );
  BUF_X1 \SB1_1_1/BUF_2  ( .A(\RI1[1][182] ), .Z(\SB1_1_1/i1[9] ) );
  BUF_X1 \SB1_1_5/BUF_2  ( .A(\RI1[1][158] ), .Z(\SB1_1_5/i1[9] ) );
  BUF_X1 U250 ( .A(\RI1[1][183] ), .Z(\SB1_1_1/i0[8] ) );
  BUF_X1 \SB1_1_10/BUF_3  ( .A(\RI1[1][129] ), .Z(\SB1_1_10/i0[8] ) );
  INV_X1 \SB1_1_20/INV_1  ( .A(\RI1[1][67] ), .ZN(\SB1_1_20/i0[6] ) );
  BUF_X1 \SB2_1_6/BUF_0  ( .A(\RI3[1][150] ), .Z(\SB2_1_6/i0[9] ) );
  BUF_X1 \SB2_1_8/BUF_1  ( .A(\RI3[1][139] ), .Z(\SB2_1_8/i0[6] ) );
  INV_X1 \SB2_1_31/INV_2  ( .A(\RI3[1][2] ), .ZN(\SB2_1_31/i1[9] ) );
  BUF_X1 \SB2_1_15/BUF_1  ( .A(\RI3[1][97] ), .Z(\SB2_1_15/i0[6] ) );
  BUF_X1 U687 ( .A(\RI3[1][78] ), .Z(\SB2_1_18/i0[9] ) );
  BUF_X1 U247 ( .A(\RI3[1][157] ), .Z(\SB2_1_5/i0[6] ) );
  BUF_X1 \SB2_1_7/BUF_1  ( .A(\RI3[1][145] ), .Z(\SB2_1_7/i0[6] ) );
  BUF_X1 \SB2_1_20/BUF_1  ( .A(\RI3[1][67] ), .Z(\SB2_1_20/i0[6] ) );
  BUF_X1 \SB2_1_24/BUF_0  ( .A(\RI3[1][42] ), .Z(\SB2_1_24/i0[9] ) );
  BUF_X1 \SB2_1_0/BUF_0  ( .A(\RI3[1][186] ), .Z(\SB2_1_0/i0[9] ) );
  BUF_X1 \SB2_1_5/BUF_0  ( .A(\RI3[1][156] ), .Z(\SB2_1_5/i0[9] ) );
  BUF_X1 \SB2_1_2/BUF_0  ( .A(\RI3[1][174] ), .Z(\SB2_1_2/i0[9] ) );
  BUF_X1 \SB2_1_4/BUF_0  ( .A(\RI3[1][162] ), .Z(\SB2_1_4/i0[9] ) );
  NAND4_X2 U2061 ( .A1(n1009), .A2(\SB2_1_16/Component_Function_2/NAND4_in[1] ), .A3(\SB2_1_16/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_16/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[110] ) );
  NAND4_X2 U4105 ( .A1(\SB2_1_31/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_31/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_31/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[20] ) );
  NAND4_X1 U1609 ( .A1(\SB2_1_23/Component_Function_5/NAND4_in[3] ), .A2(n1307), .A3(\SB2_1_23/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_23/Component_Function_5/NAND4_in[0] ), .ZN(n837) );
  BUF_X2 U707 ( .A(\RI5[1][2] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[2] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_14  ( .A(\RI5[1][14] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[14] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_104  ( .A(\RI5[1][104] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[104] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_182  ( .A(\RI5[1][182] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[182] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_74  ( .A(\RI5[1][74] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[74] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_62  ( .A(\RI5[1][62] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[62] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_39  ( .A(\RI5[1][39] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[39] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_152  ( .A(\RI5[1][152] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[152] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_118  ( .A(\RI5[1][118] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[118] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_3  ( .A(\RI5[1][3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[3] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_26  ( .A(\RI5[1][26] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[26] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_63  ( .A(\RI5[1][63] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[63] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_61  ( .A(\RI5[1][61] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[61] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_43  ( .A(\RI5[1][43] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[43] ) );
  BUF_X2 U753 ( .A(\RI5[1][87] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[87] ) );
  BUF_X2 U871 ( .A(\RI5[1][179] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[179] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_58  ( .A(\RI5[1][58] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[58] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_142  ( .A(\RI5[1][142] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[142] ) );
  BUF_X2 U787 ( .A(\MC_ARK_ARC_1_1/buf_datainput[41] ), .Z(n1498) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_52  ( .A(\RI5[1][52] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[52] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_130  ( .A(\RI5[1][130] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[130] ) );
  BUF_X2 U604 ( .A(\MC_ARK_ARC_1_1/buf_datainput[191] ), .Z(n515) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_124  ( .A(\RI5[1][124] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[124] ) );
  BUF_X1 U294 ( .A(\RI1[2][159] ), .Z(\SB1_2_5/i0[8] ) );
  BUF_X1 U1099 ( .A(\RI1[2][189] ), .Z(\SB1_2_0/i0[8] ) );
  BUF_X1 U797 ( .A(\RI1[2][15] ), .Z(\SB1_2_29/i0[8] ) );
  BUF_X1 U3081 ( .A(\RI1[2][81] ), .Z(\SB1_2_18/i0[8] ) );
  BUF_X1 \SB1_2_10/BUF_2  ( .A(\RI1[2][128] ), .Z(\SB1_2_10/i1[9] ) );
  BUF_X1 U710 ( .A(\RI1[2][129] ), .Z(\SB1_2_10/i0[8] ) );
  BUF_X1 \SB1_2_13/BUF_3  ( .A(\RI1[2][111] ), .Z(\SB1_2_13/i0[8] ) );
  BUF_X1 U1019 ( .A(\RI1[2][141] ), .Z(\SB1_2_8/i0[8] ) );
  INV_X1 \SB1_2_26/INV_0  ( .A(\RI1[2][30] ), .ZN(\SB1_2_26/i0[9] ) );
  INV_X1 \SB1_2_5/INV_5  ( .A(\RI1[2][161] ), .ZN(\SB1_2_5/i0_3 ) );
  NAND4_X1 U1308 ( .A1(\SB1_2_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_8/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_8/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_8/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[2][168] ) );
  BUF_X1 \SB2_2_10/BUF_0  ( .A(\RI3[2][126] ), .Z(\SB2_2_10/i0[9] ) );
  BUF_X1 \SB2_2_20/BUF_0  ( .A(\RI3[2][66] ), .Z(\SB2_2_20/i0[9] ) );
  BUF_X1 \SB2_2_31/BUF_0  ( .A(\RI3[2][0] ), .Z(\SB2_2_31/i0[9] ) );
  BUF_X1 \SB2_2_19/BUF_0  ( .A(\RI3[2][72] ), .Z(\SB2_2_19/i0[9] ) );
  BUF_X1 U159 ( .A(\RI3[2][49] ), .Z(\SB2_2_23/i0[6] ) );
  BUF_X1 \SB2_2_23/BUF_0  ( .A(\RI3[2][48] ), .Z(\SB2_2_23/i0[9] ) );
  BUF_X1 \SB2_2_10/BUF_1  ( .A(\RI3[2][127] ), .Z(\SB2_2_10/i0[6] ) );
  BUF_X1 \SB2_2_12/BUF_0  ( .A(\RI3[2][114] ), .Z(\SB2_2_12/i0[9] ) );
  BUF_X2 U910 ( .A(\RI3[2][119] ), .Z(\SB2_2_12/i0_3 ) );
  BUF_X1 \SB2_2_4/BUF_0  ( .A(\RI3[2][162] ), .Z(\SB2_2_4/i0[9] ) );
  CLKBUF_X2 \SB2_2_0/BUF_0  ( .A(\RI3[2][186] ), .Z(\SB2_2_0/i0[9] ) );
  BUF_X1 U624 ( .A(\RI3[2][67] ), .Z(\SB2_2_20/i0[6] ) );
  BUF_X1 U856 ( .A(\RI3[2][55] ), .Z(\SB2_2_22/i0[6] ) );
  NAND4_X2 U269 ( .A1(\SB2_2_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_1/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_1/Component_Function_3/NAND4_in[2] ), .A4(n961), .ZN(
        \RI5[2][3] ) );
  NAND4_X1 U1536 ( .A1(n1225), .A2(\SB2_2_23/Component_Function_5/NAND4_in[3] ), .A3(\SB2_2_23/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_23/Component_Function_5/NAND4_in[0] ), .ZN(n781) );
  NAND4_X2 U951 ( .A1(\SB2_2_1/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_1/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_1/Component_Function_2/NAND4_in[0] ), .A4(n587), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[8] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_9  ( .A(\RI5[2][9] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[9] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_148  ( .A(\RI5[2][148] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[148] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_45  ( .A(\RI5[2][45] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[45] ) );
  BUF_X2 U873 ( .A(\RI5[2][62] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[62] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_106  ( .A(\RI5[2][106] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[106] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_112  ( .A(\RI5[2][112] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[112] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_81  ( .A(\RI5[2][81] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[81] ) );
  BUF_X2 U885 ( .A(\RI5[2][188] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[188] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_52  ( .A(\RI5[2][52] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[52] ) );
  BUF_X2 U904 ( .A(\RI5[2][33] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[33] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_1  ( .A(\RI5[2][1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[1] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_43  ( .A(\RI5[2][43] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[43] ) );
  BUF_X2 U862 ( .A(\MC_ARK_ARC_1_2/buf_datainput[71] ), .Z(n1502) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_14  ( .A(\RI5[2][14] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[14] ) );
  INV_X1 \SB1_3_13/INV_5  ( .A(\RI1[3][113] ), .ZN(\SB1_3_13/i0_3 ) );
  BUF_X1 \SB1_3_9/BUF_2  ( .A(\RI1[3][134] ), .Z(\SB1_3_9/i1[9] ) );
  BUF_X1 \SB1_3_29/BUF_3  ( .A(\RI1[3][15] ), .Z(\SB1_3_29/i0[8] ) );
  BUF_X1 U740 ( .A(\RI1[3][20] ), .Z(\SB1_3_28/i1[9] ) );
  BUF_X2 U973 ( .A(\RI1[3][177] ), .Z(\SB1_3_2/i0[8] ) );
  BUF_X1 U959 ( .A(\RI1[3][117] ), .Z(\SB1_3_12/i0[8] ) );
  INV_X1 U3434 ( .A(\RI1[3][23] ), .ZN(\SB1_3_28/i0_3 ) );
  BUF_X1 \SB1_3_23/BUF_3  ( .A(\RI1[3][51] ), .Z(\SB1_3_23/i0[8] ) );
  BUF_X1 U739 ( .A(\RI1[3][123] ), .Z(\SB1_3_11/i0[8] ) );
  BUF_X1 \SB1_3_14/BUF_2  ( .A(\RI1[3][104] ), .Z(\SB1_3_14/i1[9] ) );
  CLKBUF_X1 \SB1_3_8/BUF_4  ( .A(\RI1[3][142] ), .Z(\SB1_3_8/i0[7] ) );
  BUF_X1 \SB1_3_9/BUF_3  ( .A(\RI1[3][135] ), .Z(\SB1_3_9/i0[8] ) );
  BUF_X1 U682 ( .A(\RI1[3][165] ), .Z(\SB1_3_4/i0[8] ) );
  BUF_X1 \SB1_3_14/BUF_3  ( .A(\RI1[3][105] ), .Z(\SB1_3_14/i0[8] ) );
  BUF_X1 U135 ( .A(\RI1[3][57] ), .Z(\SB1_3_22/i0[8] ) );
  BUF_X1 \SB1_3_13/BUF_3  ( .A(\RI1[3][111] ), .Z(\SB1_3_13/i0[8] ) );
  BUF_X1 U614 ( .A(\RI1[3][110] ), .Z(\SB1_3_13/i1[9] ) );
  BUF_X1 U1067 ( .A(\RI1[3][92] ), .Z(\SB1_3_16/i1[9] ) );
  NAND4_X1 U1542 ( .A1(\SB1_3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_4/NAND4_in[3] ), .ZN(n786) );
  BUF_X1 U126 ( .A(\RI3[3][25] ), .Z(\SB2_3_27/i0[6] ) );
  BUF_X1 \SB2_3_2/BUF_0  ( .A(\RI3[3][174] ), .Z(\SB2_3_2/i0[9] ) );
  BUF_X1 \SB2_3_20/BUF_1  ( .A(\RI3[3][67] ), .Z(\SB2_3_20/i0[6] ) );
  BUF_X1 U748 ( .A(\RI3[3][175] ), .Z(\SB2_3_2/i0[6] ) );
  BUF_X1 U668 ( .A(\RI3[3][61] ), .Z(\SB2_3_21/i0[6] ) );
  BUF_X1 U816 ( .A(\RI3[3][55] ), .Z(\SB2_3_22/i0[6] ) );
  BUF_X1 U107 ( .A(\RI3[3][132] ), .Z(n546) );
  BUF_X1 \SB2_3_10/BUF_0  ( .A(\RI3[3][126] ), .Z(\SB2_3_10/i0[9] ) );
  BUF_X1 \SB2_3_25/BUF_1  ( .A(\RI3[3][37] ), .Z(\SB2_3_25/i0[6] ) );
  BUF_X1 \SB2_3_21/BUF_0  ( .A(\RI3[3][60] ), .Z(\SB2_3_21/i0[9] ) );
  BUF_X1 U680 ( .A(\RI3[3][7] ), .Z(\SB2_3_30/i0[6] ) );
  NAND4_X2 U3673 ( .A1(\SB2_3_9/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_9/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_9/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_9/Component_Function_2/NAND4_in[0] ), .ZN(\RI5[3][152] ) );
  NAND4_X2 \SB2_3_25/Component_Function_2/N5  ( .A1(
        \SB2_3_25/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_3_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_25/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_25/Component_Function_2/NAND4_in[0] ), .ZN(\RI5[3][56] ) );
  NAND4_X2 U586 ( .A1(\SB2_3_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_20/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[3][86] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_21  ( .A(\RI5[3][21] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[21] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_174  ( .A(\RI5[3][174] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[174] ) );
  BUF_X2 U1617 ( .A(\RI5[3][47] ), .Z(n842) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_106  ( .A(\RI5[3][106] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[106] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_111  ( .A(\RI5[3][111] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[111] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_114  ( .A(\RI5[3][114] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[114] ) );
  CLKBUF_X1 U533 ( .A(\RI1[4][124] ), .Z(\SB3_11/i0[7] ) );
  BUF_X1 U3 ( .A(\RI1[4][153] ), .Z(\SB3_6/i0[8] ) );
  BUF_X1 \SB3_29/BUF_2  ( .A(\RI1[4][14] ), .Z(\SB3_29/i1[9] ) );
  NAND4_X1 U1532 ( .A1(\SB3_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_0/NAND4_in[0] ), .A4(n1035), .ZN(n779) );
  NAND4_X1 U838 ( .A1(\SB3_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_2/Component_Function_0/NAND4_in[0] ), .A4(n960), .ZN(n790) );
  BUF_X1 \SB4_20/BUF_0  ( .A(\RI3[4][66] ), .Z(\SB4_20/i0[9] ) );
  BUF_X1 \SB4_11/BUF_0  ( .A(\RI3[4][120] ), .Z(\SB4_11/i0[9] ) );
  BUF_X1 U727 ( .A(\RI3[4][59] ), .Z(\SB4_22/i0_3 ) );
  BUF_X1 \SB4_24/BUF_0  ( .A(\RI3[4][42] ), .Z(\SB4_24/i0[9] ) );
  BUF_X1 U3082 ( .A(\RI3[4][90] ), .Z(\SB4_16/i0[9] ) );
  BUF_X1 \SB4_9/BUF_0  ( .A(\RI3[4][132] ), .Z(\SB4_9/i0[9] ) );
  CLKBUF_X1 U84 ( .A(Key[64]), .Z(n455) );
  BUF_X1 U1184 ( .A(Key[103]), .Z(n378) );
  CLKBUF_X1 U67 ( .A(Key[110]), .Z(n501) );
  CLKBUF_X1 U11 ( .A(Key[130]), .Z(n471) );
  CLKBUF_X1 U127 ( .A(Key[17]), .Z(n393) );
  CLKBUF_X1 U1181 ( .A(Key[70]), .Z(n459) );
  BUF_X1 U25 ( .A(Key[10]), .Z(n456) );
  CLKBUF_X1 U97 ( .A(Key[112]), .Z(n435) );
  CLKBUF_X1 U119 ( .A(Key[167]), .Z(n385) );
  CLKBUF_X1 U2 ( .A(Key[136]), .Z(n376) );
  BUF_X1 U601 ( .A(n75), .Z(\SB1_0_12/i0[8] ) );
  INV_X1 U679 ( .A(n151), .ZN(\SB1_0_25/i0_3 ) );
  BUF_X1 \SB2_0_31/BUF_0  ( .A(\RI3[0][0] ), .Z(\SB2_0_31/i0[9] ) );
  BUF_X2 \SB2_0_1/BUF_2  ( .A(\RI3[0][182] ), .Z(\SB2_0_1/i0_0 ) );
  BUF_X1 U761 ( .A(\RI3[0][1] ), .Z(\SB2_0_31/i0[6] ) );
  CLKBUF_X2 \SB2_0_23/BUF_2  ( .A(\RI3[0][50] ), .Z(\SB2_0_23/i0_0 ) );
  BUF_X1 \SB2_0_8/BUF_0  ( .A(\RI3[0][138] ), .Z(\SB2_0_8/i0[9] ) );
  CLKBUF_X2 \SB2_0_6/BUF_3  ( .A(\RI3[0][153] ), .Z(\SB2_0_6/i0[10] ) );
  BUF_X1 U1250 ( .A(\RI3[0][24] ), .Z(\SB2_0_27/i0[9] ) );
  BUF_X1 \SB2_0_18/BUF_0  ( .A(\RI3[0][78] ), .Z(\SB2_0_18/i0[9] ) );
  BUF_X1 \SB2_0_10/BUF_0  ( .A(\RI3[0][126] ), .Z(\SB2_0_10/i0[9] ) );
  BUF_X1 \SB2_0_2/BUF_0  ( .A(\RI3[0][174] ), .Z(\SB2_0_2/i0[9] ) );
  BUF_X1 \SB2_0_20/BUF_0  ( .A(\RI3[0][66] ), .Z(\SB2_0_20/i0[9] ) );
  BUF_X1 \SB2_0_4/BUF_1  ( .A(\RI3[0][163] ), .Z(\SB2_0_4/i0[6] ) );
  NAND4_X2 U4102 ( .A1(\SB2_0_25/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_25/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_25/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_25/Component_Function_3/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[51] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_142  ( .A(\RI5[0][142] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[142] ) );
  CLKBUF_X1 U889 ( .A(\MC_ARK_ARC_1_0/buf_datainput[35] ), .Z(n1507) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_122  ( .A(\RI5[0][122] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[122] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_91  ( .A(\RI5[0][91] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[91] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_96  ( .A(\RI5[0][96] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[96] ) );
  BUF_X1 U609 ( .A(\MC_ARK_ARC_1_0/buf_datainput[29] ), .Z(n1470) );
  BUF_X1 \SB1_1_5/BUF_3  ( .A(\RI1[1][159] ), .Z(\SB1_1_5/i0[8] ) );
  BUF_X1 \SB1_1_17/BUF_3  ( .A(\RI1[1][87] ), .Z(\SB1_1_17/i0[8] ) );
  BUF_X1 \SB1_1_14/BUF_3  ( .A(\RI1[1][105] ), .Z(\SB1_1_14/i0[8] ) );
  BUF_X1 \SB1_1_22/BUF_2  ( .A(\RI1[1][56] ), .Z(\SB1_1_22/i1[9] ) );
  CLKBUF_X2 \SB2_1_17/BUF_0  ( .A(\RI3[1][84] ), .Z(\SB2_1_17/i0[9] ) );
  CLKBUF_X2 \SB2_1_6/BUF_3  ( .A(\RI3[1][153] ), .Z(\SB2_1_6/i0[10] ) );
  BUF_X1 \SB2_1_26/BUF_1  ( .A(\RI3[1][31] ), .Z(\SB2_1_26/i0[6] ) );
  BUF_X1 \SB2_1_30/BUF_0  ( .A(\RI3[1][6] ), .Z(\SB2_1_30/i0[9] ) );
  CLKBUF_X2 \SB2_1_2/BUF_2  ( .A(\RI3[1][176] ), .Z(\SB2_1_2/i0_0 ) );
  BUF_X1 \SB2_1_25/BUF_0  ( .A(\RI3[1][36] ), .Z(\SB2_1_25/i0[9] ) );
  CLKBUF_X2 \SB2_1_14/BUF_2  ( .A(\RI3[1][104] ), .Z(\SB2_1_14/i0_0 ) );
  BUF_X1 \SB2_1_3/BUF_1  ( .A(\RI3[1][169] ), .Z(\SB2_1_3/i0[6] ) );
  NAND4_X2 U574 ( .A1(\SB2_1_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_9/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][147] ) );
  NAND4_X2 U3497 ( .A1(\SB2_1_5/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_5/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_5/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_5/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[176] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_111  ( .A(\RI5[1][111] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[111] ) );
  BUF_X1 \SB1_2_19/BUF_3  ( .A(\RI1[2][75] ), .Z(\SB1_2_19/i0[8] ) );
  CLKBUF_X1 \SB1_2_14/BUF_0  ( .A(\RI1[2][102] ), .Z(\SB1_2_14/i3[0] ) );
  CLKBUF_X2 \SB2_2_28/BUF_3  ( .A(\RI3[2][21] ), .Z(\SB2_2_28/i0[10] ) );
  BUF_X1 \SB2_2_28/BUF_0  ( .A(\RI3[2][18] ), .Z(\SB2_2_28/i0[9] ) );
  CLKBUF_X2 \SB2_2_17/BUF_2  ( .A(\RI3[2][86] ), .Z(\SB2_2_17/i0_0 ) );
  BUF_X1 U948 ( .A(\RI3[2][115] ), .Z(\SB2_2_12/i0[6] ) );
  CLKBUF_X2 \SB2_2_12/BUF_3  ( .A(\RI3[2][117] ), .Z(\SB2_2_12/i0[10] ) );
  BUF_X1 \SB2_2_8/BUF_4  ( .A(\RI3[2][142] ), .Z(\SB2_2_8/i0_4 ) );
  BUF_X2 U566 ( .A(\MC_ARK_ARC_1_2/buf_datainput[71] ), .Z(n1503) );
  BUF_X1 \SB1_3_25/BUF_2  ( .A(\RI1[3][38] ), .Z(\SB1_3_25/i1[9] ) );
  BUF_X2 U810 ( .A(\RI1[3][189] ), .Z(\SB1_3_0/i0[8] ) );
  BUF_X1 U664 ( .A(\RI1[3][159] ), .Z(\SB1_3_5/i0[8] ) );
  BUF_X1 \SB1_3_18/BUF_3  ( .A(\RI1[3][81] ), .Z(\SB1_3_18/i0[8] ) );
  BUF_X2 U662 ( .A(\RI1[3][80] ), .Z(\SB1_3_18/i1[9] ) );
  BUF_X1 U738 ( .A(\RI1[3][26] ), .Z(\SB1_3_27/i1[9] ) );
  BUF_X1 \SB2_3_25/BUF_0  ( .A(\RI3[3][36] ), .Z(\SB2_3_25/i0[9] ) );
  BUF_X1 \SB4_15/BUF_0  ( .A(\RI3[4][96] ), .Z(\SB4_15/i0[9] ) );
  BUF_X1 \SB4_19/BUF_0  ( .A(\RI3[4][72] ), .Z(\SB4_19/i0[9] ) );
  BUF_X1 \SB4_12/BUF_1  ( .A(\RI3[4][115] ), .Z(\SB4_12/i0[6] ) );
  BUF_X2 U1208 ( .A(n4), .Z(\SB1_0_0/i1[9] ) );
  BUF_X2 \SB1_3_16/BUF_3  ( .A(\RI1[3][93] ), .Z(\SB1_3_16/i0[8] ) );
  BUF_X2 U245 ( .A(\RI1[2][147] ), .Z(\SB1_2_7/i0[8] ) );
  BUF_X2 \SB2_3_24/BUF_1  ( .A(\RI3[3][43] ), .Z(\SB2_3_24/i0[6] ) );
  BUF_X2 \SB1_0_12/BUF_2  ( .A(n76), .Z(\SB1_0_12/i1[9] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_46  ( .A(\RI5[0][46] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[46] ) );
  BUF_X2 U1209 ( .A(n88), .Z(\SB1_0_14/i1[9] ) );
  BUF_X2 \SB2_2_7/BUF_0  ( .A(\RI3[2][144] ), .Z(\SB2_2_7/i0[9] ) );
  BUF_X2 \SB1_0_17/BUF_2  ( .A(n106), .Z(\SB1_0_17/i1[9] ) );
  CLKBUF_X3 U1539 ( .A(\RI5[3][117] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[117] )
         );
  CLKBUF_X3 U747 ( .A(\RI5[1][165] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[165] )
         );
  BUF_X2 \SB2_2_12/BUF_2  ( .A(\RI3[2][116] ), .Z(\SB2_2_12/i0_0 ) );
  CLKBUF_X3 \MC_ARK_ARC_1_1/BUF_134  ( .A(\RI5[1][134] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[134] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_134  ( .A(\RI5[2][134] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[134] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_154  ( .A(\RI5[2][154] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[154] ) );
  CLKBUF_X3 U634 ( .A(\RI5[2][74] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[74] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_3/BUF_101  ( .A(\RI5[3][101] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[101] ) );
  BUF_X2 U1254 ( .A(\RI1[1][32] ), .Z(\SB1_1_26/i1[9] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_190  ( .A(\RI5[2][190] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[190] ) );
  BUF_X2 U1653 ( .A(n37), .Z(\SB1_0_6/i1_5 ) );
  BUF_X2 U697 ( .A(\RI3[0][25] ), .Z(\SB2_0_27/i0[6] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_1/BUF_128  ( .A(\RI5[1][128] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[128] ) );
  BUF_X2 U667 ( .A(n172), .Z(\SB1_0_28/i1[9] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_40  ( .A(\RI5[1][40] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[40] ) );
  BUF_X2 \SB2_0_3/BUF_2  ( .A(\RI3[0][170] ), .Z(\SB2_0_3/i0_0 ) );
  CLKBUF_X3 \MC_ARK_ARC_1_1/BUF_170  ( .A(\RI5[1][170] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[170] ) );
  BUF_X2 U1645 ( .A(\RI3[4][102] ), .Z(\SB4_14/i0[9] ) );
  BUF_X2 \SB2_2_26/BUF_0  ( .A(\RI3[2][30] ), .Z(\SB2_2_26/i0[9] ) );
  INV_X2 \SB1_2_4/INV_4  ( .A(\RI1[2][166] ), .ZN(\SB1_2_4/i0_4 ) );
  BUF_X2 \SB4_12/BUF_0  ( .A(\RI3[4][114] ), .Z(\SB4_12/i0[9] ) );
  BUF_X1 \SB1_1_26/BUF_1  ( .A(\RI1[1][31] ), .Z(\SB1_1_26/i1_7 ) );
  BUF_X2 \SB1_0_6/BUF_2  ( .A(n40), .Z(\SB1_0_6/i1[9] ) );
  BUF_X2 \SB2_0_7/BUF_4  ( .A(\RI3[0][148] ), .Z(\SB2_0_7/i0_4 ) );
  CLKBUF_X3 U917 ( .A(\RI5[3][17] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[17] ) );
  BUF_X2 \SB2_0_5/BUF_1  ( .A(\RI3[0][157] ), .Z(\SB2_0_5/i0[6] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_116  ( .A(\RI5[2][116] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[116] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_88  ( .A(\RI5[2][88] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[88] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_0/BUF_25  ( .A(\RI5[0][25] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[25] ) );
  BUF_X2 \SB1_0_31/BUF_2  ( .A(n190), .Z(\SB1_0_31/i1[9] ) );
  BUF_X2 \SB2_1_22/BUF_1  ( .A(\RI3[1][55] ), .Z(\SB2_1_22/i0[6] ) );
  BUF_X2 U654 ( .A(\RI1[3][27] ), .Z(\SB1_3_27/i0[8] ) );
  BUF_X2 \SB2_3_22/BUF_0  ( .A(\RI3[3][54] ), .Z(\SB2_3_22/i0[9] ) );
  OR3_X2 U3959 ( .A1(\SB1_2_6/i0[7] ), .A2(\RI1[2][150] ), .A3(\RI1[2][151] ), 
        .ZN(n1118) );
  INV_X2 \SB1_1_9/INV_0  ( .A(\RI1[1][132] ), .ZN(\SB1_1_9/i0[9] ) );
  BUF_X2 U3711 ( .A(\RI3[2][91] ), .Z(\SB2_2_16/i0[6] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_92  ( .A(\RI5[2][92] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[92] ) );
  BUF_X2 \SB2_1_22/BUF_0  ( .A(\RI3[1][54] ), .Z(\SB2_1_22/i0[9] ) );
  BUF_X2 \SB1_1_27/BUF_3  ( .A(\RI1[1][27] ), .Z(\SB1_1_27/i0[8] ) );
  CLKBUF_X3 U839 ( .A(\RI5[3][89] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[89] ) );
  BUF_X2 \SB2_0_23/BUF_3  ( .A(\RI3[0][51] ), .Z(\SB2_0_23/i0[10] ) );
  BUF_X2 U174 ( .A(\RI1[3][129] ), .Z(\SB1_3_10/i0[8] ) );
  BUF_X2 \SB1_0_18/BUF_2  ( .A(n112), .Z(\SB1_0_18/i1[9] ) );
  CLKBUF_X3 \MC_ARK_ARC_1_2/BUF_50  ( .A(\RI5[2][50] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[50] ) );
  BUF_X2 U1625 ( .A(\RI3[4][53] ), .Z(n848) );
  BUF_X2 U1106 ( .A(\RI1[2][123] ), .Z(\SB1_2_11/i0[8] ) );
  BUF_X2 U138 ( .A(\RI1[3][170] ), .Z(\SB1_3_3/i1[9] ) );
  BUF_X2 \SB2_0_0/BUF_1  ( .A(\RI3[0][187] ), .Z(\SB2_0_0/i0[6] ) );
  BUF_X2 U665 ( .A(\RI1[1][38] ), .Z(\SB1_1_25/i1[9] ) );
  BUF_X1 \SB1_0_8/BUF_5  ( .A(n49), .Z(\SB1_0_8/i1_5 ) );
  CLKBUF_X2 U764 ( .A(n183), .Z(\SB1_0_30/i0[8] ) );
  NAND4_X2 \SB2_0_20/Component_Function_4/N5  ( .A1(
        \SB2_0_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][76] ) );
  NAND4_X2 \SB2_0_13/Component_Function_3/N5  ( .A1(
        \SB2_0_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_13/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[0][123] ) );
  NAND4_X2 \SB2_0_6/Component_Function_3/N5  ( .A1(
        \SB2_0_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[0][165] ) );
  NAND4_X2 \SB2_0_7/Component_Function_1/N5  ( .A1(
        \SB2_0_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_7/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][169] ) );
  NAND4_X2 \SB2_0_11/Component_Function_0/N5  ( .A1(
        \SB2_0_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_11/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][150] ) );
  NAND4_X2 \SB2_0_2/Component_Function_4/N5  ( .A1(
        \SB2_0_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_2/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][184] ) );
  NAND4_X2 \SB2_0_6/Component_Function_2/N5  ( .A1(
        \SB2_0_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[0][170] ) );
  NAND4_X2 U4364 ( .A1(\SB2_0_24/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_24/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_24/Component_Function_2/NAND4_in[0] ), .A4(n1857), .ZN(
        \RI5[0][62] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_90  ( .A(\RI5[0][90] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[90] ) );
  NAND4_X2 \SB2_0_14/Component_Function_4/N5  ( .A1(
        \SB2_0_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_14/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_14/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[0][112] ) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_99  ( .A(\RI5[0][99] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[99] ) );
  BUF_X1 U49 ( .A(Key[9]), .Z(n503) );
  BUF_X2 U1257 ( .A(\RI1[1][128] ), .Z(\SB1_1_10/i1[9] ) );
  BUF_X2 U938 ( .A(\RI1[1][146] ), .Z(\SB1_1_7/i1[9] ) );
  BUF_X2 U1018 ( .A(\RI1[1][44] ), .Z(\SB1_1_24/i1[9] ) );
  BUF_X1 \SB1_1_13/BUF_3  ( .A(\RI1[1][111] ), .Z(\SB1_1_13/i0[8] ) );
  NAND4_X2 \SB2_1_25/Component_Function_2/N5  ( .A1(
        \SB2_1_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_1_25/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[1][56] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_140  ( .A(\RI5[1][140] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[140] ) );
  NAND4_X2 \SB2_1_24/Component_Function_3/N5  ( .A1(
        \SB2_1_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_24/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][57] ) );
  NAND4_X2 U2946 ( .A1(\SB2_1_0/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_0/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_0/Component_Function_3/NAND4_in[2] ), .A4(n1261), .ZN(
        \RI5[1][9] ) );
  BUF_X1 \SB1_2_8/BUF_2  ( .A(\RI1[2][140] ), .Z(\SB1_2_8/i1[9] ) );
  BUF_X1 U286 ( .A(\RI3[2][145] ), .Z(\SB2_2_7/i0[6] ) );
  NAND4_X2 \SB2_2_5/Component_Function_3/N5  ( .A1(
        \SB2_2_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_5/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][171] ) );
  NAND4_X2 \SB2_2_19/Component_Function_3/N5  ( .A1(
        \SB2_2_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_19/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][87] ) );
  NAND4_X2 \SB2_2_4/Component_Function_1/N5  ( .A1(
        \SB2_2_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][187] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_75  ( .A(\RI5[2][75] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[75] ) );
  NAND4_X2 \SB2_2_4/Component_Function_3/N5  ( .A1(
        \SB2_2_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][177] ) );
  NAND4_X2 \SB2_2_14/Component_Function_3/N5  ( .A1(
        \SB2_2_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][117] ) );
  BUF_X2 \MC_ARK_ARC_1_2/BUF_165  ( .A(\RI5[2][165] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[165] ) );
  BUF_X1 U812 ( .A(\RI1[3][62] ), .Z(\SB1_3_21/i1[9] ) );
  BUF_X1 \SB1_3_7/BUF_3  ( .A(\RI1[3][147] ), .Z(\SB1_3_7/i0[8] ) );
  CLKBUF_X2 U979 ( .A(\RI1[3][39] ), .Z(\SB1_3_25/i0[8] ) );
  BUF_X1 \SB1_3_28/BUF_3  ( .A(\RI1[3][21] ), .Z(\SB1_3_28/i0[8] ) );
  BUF_X1 U55 ( .A(\RI3[3][79] ), .Z(\SB2_3_18/i0[6] ) );
  NAND4_X2 \SB2_3_26/Component_Function_3/N5  ( .A1(
        \SB2_3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_26/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[3][45] ) );
  NAND4_X2 \SB2_3_3/Component_Function_2/N5  ( .A1(
        \SB2_3_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_3/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_3/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[3][188] ) );
  NAND4_X2 \SB2_3_2/Component_Function_4/N5  ( .A1(
        \SB2_3_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_2/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][184] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_47  ( .A(\RI5[3][47] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[47] ) );
  BUF_X2 U1613 ( .A(\RI5[3][185] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[185] ) );
  BUF_X2 \MC_ARK_ARC_1_3/BUF_64  ( .A(\RI5[3][64] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[64] ) );
  BUF_X1 \SB3_23/BUF_2  ( .A(\RI1[4][50] ), .Z(\SB3_23/i1[9] ) );
  BUF_X1 \SB3_2/BUF_2  ( .A(\RI1[4][176] ), .Z(\SB3_2/i1[9] ) );
  BUF_X1 \SB3_5/BUF_2  ( .A(\RI1[4][158] ), .Z(\SB3_5/i1[9] ) );
  CLKBUF_X2 U30 ( .A(\RI1[3][8] ), .Z(\SB1_3_30/i1[9] ) );
  CLKBUF_X2 U41 ( .A(\RI1[3][56] ), .Z(\SB1_3_22/i1[9] ) );
  BUF_X1 U52 ( .A(\RI1[3][32] ), .Z(\SB1_3_26/i1[9] ) );
  BUF_X2 U57 ( .A(\RI1[3][86] ), .Z(\SB1_3_17/i1[9] ) );
  BUF_X2 U96 ( .A(\RI1[3][44] ), .Z(\SB1_3_24/i1[9] ) );
  BUF_X2 U100 ( .A(\RI1[3][45] ), .Z(\SB1_3_24/i0[8] ) );
  BUF_X2 U111 ( .A(\RI5[2][98] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[98] ) );
  BUF_X2 U121 ( .A(\RI3[2][43] ), .Z(\SB2_2_24/i0[6] ) );
  BUF_X2 U130 ( .A(\RI3[2][19] ), .Z(\SB2_2_28/i0[6] ) );
  BUF_X2 U131 ( .A(\RI3[2][151] ), .Z(\SB2_2_6/i0[6] ) );
  BUF_X2 U139 ( .A(\RI3[2][187] ), .Z(\SB2_2_0/i0[6] ) );
  BUF_X1 U152 ( .A(\RI1[2][99] ), .Z(\SB1_2_15/i0[8] ) );
  CLKBUF_X2 U162 ( .A(\RI1[2][177] ), .Z(\SB1_2_2/i0[8] ) );
  CLKBUF_X2 U165 ( .A(\RI1[2][165] ), .Z(\SB1_2_4/i0[8] ) );
  CLKBUF_X2 U169 ( .A(\RI1[2][104] ), .Z(\SB1_2_14/i1[9] ) );
  CLKBUF_X2 U170 ( .A(\RI1[2][134] ), .Z(\SB1_2_9/i1[9] ) );
  CLKBUF_X2 U172 ( .A(\RI1[2][86] ), .Z(\SB1_2_17/i1[9] ) );
  CLKBUF_X2 U181 ( .A(\RI1[2][80] ), .Z(\SB1_2_18/i1[9] ) );
  BUF_X2 U185 ( .A(\RI1[2][38] ), .Z(\SB1_2_25/i1[9] ) );
  BUF_X2 U196 ( .A(\RI1[2][182] ), .Z(\SB1_2_1/i1[9] ) );
  BUF_X1 U205 ( .A(\RI1[2][21] ), .Z(\SB1_2_28/i0[8] ) );
  BUF_X2 U206 ( .A(\RI5[1][45] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[45] ) );
  BUF_X1 U208 ( .A(\RI5[1][183] ), .Z(n1958) );
  BUF_X2 U216 ( .A(\RI5[1][68] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[68] ) );
  BUF_X2 U254 ( .A(\RI3[1][37] ), .Z(\SB2_1_25/i0[6] ) );
  BUF_X2 U259 ( .A(\RI3[1][13] ), .Z(\SB2_1_29/i0[6] ) );
  BUF_X2 U270 ( .A(\RI3[1][18] ), .Z(\SB2_1_28/i0[9] ) );
  BUF_X1 U296 ( .A(\RI3[1][151] ), .Z(\SB2_1_6/i0[6] ) );
  BUF_X1 U298 ( .A(\RI3[1][49] ), .Z(\SB2_1_23/i0[6] ) );
  BUF_X2 U305 ( .A(\RI1[1][117] ), .Z(\SB1_1_12/i0[8] ) );
  CLKBUF_X2 U307 ( .A(\RI1[1][165] ), .Z(\SB1_1_4/i0[8] ) );
  CLKBUF_X2 U308 ( .A(\RI1[1][39] ), .Z(\SB1_1_25/i0[8] ) );
  CLKBUF_X2 U309 ( .A(\RI1[1][170] ), .Z(\SB1_1_3/i1[9] ) );
  CLKBUF_X2 U310 ( .A(\RI1[1][74] ), .Z(\SB1_1_19/i1[9] ) );
  CLKBUF_X2 U527 ( .A(\RI1[1][68] ), .Z(\SB1_1_20/i1[9] ) );
  CLKBUF_X2 U528 ( .A(\RI1[1][14] ), .Z(\SB1_1_29/i1[9] ) );
  CLKBUF_X2 U532 ( .A(\RI1[1][140] ), .Z(\SB1_1_8/i1[9] ) );
  BUF_X2 U535 ( .A(\RI1[1][110] ), .Z(\SB1_1_13/i1[9] ) );
  BUF_X2 U536 ( .A(\RI1[1][50] ), .Z(\SB1_1_23/i1[9] ) );
  BUF_X2 U538 ( .A(\MC_ARK_ARC_1_0/buf_datainput[116] ), .Z(n1941) );
  BUF_X2 U539 ( .A(\RI5[0][104] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[104] ) );
  NAND4_X2 U540 ( .A1(n1799), .A2(n1714), .A3(
        \SB2_0_23/Component_Function_3/NAND4_in[2] ), .A4(n2046), .ZN(
        \RI5[0][63] ) );
  NAND4_X2 U543 ( .A1(\SB2_0_9/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_9/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_9/Component_Function_2/NAND4_in[0] ), .A4(n2169), .ZN(
        \RI5[0][152] ) );
  BUF_X2 U550 ( .A(\RI3[0][109] ), .Z(\SB2_0_13/i0[6] ) );
  BUF_X1 U552 ( .A(n21), .Z(\SB1_0_3/i0[8] ) );
  NAND4_X4 U553 ( .A1(\SB2_0_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_0/Component_Function_5/NAND4_in[1] ), .A3(n1155), .A4(
        \SB2_0_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[191] ) );
  BUF_X2 U570 ( .A(\RI5[0][38] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[38] ) );
  BUF_X2 U581 ( .A(\RI1[2][62] ), .Z(\SB1_2_21/i1[9] ) );
  BUF_X2 U600 ( .A(\RI1[2][69] ), .Z(\SB1_2_20/i0[8] ) );
  BUF_X1 U605 ( .A(\RI1[1][149] ), .Z(\SB1_1_7/i1_5 ) );
  BUF_X2 U612 ( .A(n165), .Z(\SB1_0_27/i0[8] ) );
  BUF_X1 U613 ( .A(\RI1[4][173] ), .Z(\SB3_3/i1_5 ) );
  BUF_X2 U615 ( .A(\RI1[2][26] ), .Z(\SB1_2_27/i1[9] ) );
  BUF_X1 U617 ( .A(\RI1[2][191] ), .Z(\SB1_2_0/i1_5 ) );
  BUF_X2 U620 ( .A(n34), .Z(\SB1_0_5/i1[9] ) );
  BUF_X2 U622 ( .A(\RI1[3][3] ), .Z(\SB1_3_31/i0[8] ) );
  BUF_X2 U638 ( .A(\RI1[1][152] ), .Z(\SB1_1_6/i1[9] ) );
  BUF_X2 U640 ( .A(\RI3[1][101] ), .Z(\SB2_1_15/i0_3 ) );
  BUF_X1 U641 ( .A(\RI1[4][64] ), .Z(\SB3_21/i0[7] ) );
  NAND4_X2 U647 ( .A1(\SB2_2_26/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_26/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_26/Component_Function_5/NAND4_in[3] ), .A4(n1189), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[35] ) );
  BUF_X2 U649 ( .A(\RI5[1][171] ), .Z(n1954) );
  BUF_X2 U651 ( .A(\RI1[2][158] ), .Z(\SB1_2_5/i1[9] ) );
  NAND4_X2 U652 ( .A1(\SB2_0_7/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_7/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][174] ) );
  NAND4_X2 U653 ( .A1(\SB2_0_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_10/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[0][156] ) );
  NAND4_X2 U658 ( .A1(\SB2_1_30/Component_Function_5/NAND4_in[2] ), .A2(n561), 
        .A3(\SB2_1_30/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_30/Component_Function_5/NAND4_in[0] ), .ZN(n2105) );
  NAND4_X2 U660 ( .A1(\SB2_2_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_22/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_22/Component_Function_5/NAND4_in[0] ), .ZN(n792) );
  NAND4_X2 U666 ( .A1(n1089), .A2(\SB2_2_28/Component_Function_4/NAND4_in[0] ), 
        .A3(\SB2_2_28/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_2_28/Component_Function_4/NAND4_in[1] ), .ZN(n2142) );
  NAND4_X2 U669 ( .A1(\SB2_2_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_2/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_2/Component_Function_2/NAND4_in[1] ), .A4(n1072), .ZN(
        \RI5[2][2] ) );
  NAND4_X2 U671 ( .A1(\SB2_3_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_27/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[3][49] ) );
  BUF_X2 U677 ( .A(\RI5[3][148] ), .Z(n1510) );
  NAND4_X2 U678 ( .A1(\SB2_3_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_9/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][162] ) );
  CLKBUF_X3 U684 ( .A(\RI5[0][87] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[87] ) );
  CLKBUF_X3 U692 ( .A(\RI5[2][105] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[105] )
         );
  BUF_X2 U694 ( .A(\RI3[1][127] ), .Z(\SB2_1_10/i0[6] ) );
  CLKBUF_X1 U696 ( .A(\MC_ARK_ARC_1_1/buf_datainput[23] ), .Z(n1925) );
  BUF_X1 U703 ( .A(\MC_ARK_ARC_1_1/buf_datainput[23] ), .Z(n1926) );
  CLKBUF_X1 U705 ( .A(\MC_ARK_ARC_1_1/buf_datainput[23] ), .Z(n1927) );
  NAND4_X1 U706 ( .A1(\SB2_1_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_28/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_28/Component_Function_5/NAND4_in[1] ), .A4(n1535), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[23] ) );
  CLKBUF_X1 U708 ( .A(\MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(n1928) );
  BUF_X1 U711 ( .A(\MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(n1929) );
  CLKBUF_X1 U713 ( .A(\MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(n1930) );
  NAND4_X1 U715 ( .A1(\SB2_3_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_14/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_14/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[122] ) );
  CLKBUF_X3 U716 ( .A(\RI1[2][105] ), .Z(\SB1_2_14/i0[8] ) );
  BUF_X1 U717 ( .A(\MC_ARK_ARC_1_2/buf_datainput[136] ), .Z(n1932) );
  BUF_X1 U718 ( .A(\MC_ARK_ARC_1_2/buf_datainput[136] ), .Z(n1933) );
  NAND4_X1 U721 ( .A1(n1558), .A2(\SB2_2_10/Component_Function_4/NAND4_in[0] ), 
        .A3(\SB2_2_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_10/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[136] ) );
  BUF_X2 U722 ( .A(\RI1[3][63] ), .Z(\SB1_3_21/i0[8] ) );
  CLKBUF_X3 U723 ( .A(\RI1[3][140] ), .Z(\SB1_3_8/i1[9] ) );
  CLKBUF_X3 U724 ( .A(\RI1[3][141] ), .Z(\SB1_3_8/i0[8] ) );
  CLKBUF_X1 U725 ( .A(\RI5[1][189] ), .Z(n1934) );
  BUF_X2 U726 ( .A(\RI5[1][189] ), .Z(n1935) );
  NAND4_X1 U729 ( .A1(\SB2_1_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_2/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_2/Component_Function_3/NAND4_in[2] ), .A4(n1771), .ZN(
        \RI5[1][189] ) );
  CLKBUF_X3 U732 ( .A(\RI5[3][68] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[68] ) );
  CLKBUF_X3 U733 ( .A(\RI5[2][26] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[26] ) );
  CLKBUF_X3 U735 ( .A(\RI5[1][38] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[38] ) );
  BUF_X2 U744 ( .A(\RI1[1][15] ), .Z(\SB1_1_29/i0[8] ) );
  BUF_X2 U749 ( .A(n10), .Z(\SB1_0_1/i1[9] ) );
  CLKBUF_X1 U752 ( .A(\MC_ARK_ARC_1_1/buf_datainput[173] ), .Z(n1936) );
  BUF_X2 U755 ( .A(\MC_ARK_ARC_1_1/buf_datainput[173] ), .Z(n1937) );
  NAND4_X1 U756 ( .A1(\SB2_1_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_3/Component_Function_5/NAND4_in[1] ), .A3(n906), .A4(n1555), 
        .ZN(\MC_ARK_ARC_1_1/buf_datainput[173] ) );
  CLKBUF_X3 U757 ( .A(\RI5[2][141] ), .Z(n1951) );
  NAND4_X2 U758 ( .A1(\SB2_2_17/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_17/Component_Function_3/NAND4_in[0] ), .A3(n1311), .A4(
        \SB2_2_17/Component_Function_3/NAND4_in[2] ), .ZN(\RI5[2][99] ) );
  INV_X2 U765 ( .A(\RI1[3][179] ), .ZN(\SB1_3_2/i0_3 ) );
  CLKBUF_X3 U771 ( .A(\RI5[1][89] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[89] ) );
  INV_X2 U786 ( .A(n145), .ZN(\SB1_0_24/i0_3 ) );
  NAND4_X2 U822 ( .A1(\SB2_2_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_25/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][51] ) );
  CLKBUF_X3 U840 ( .A(\RI5[3][76] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[76] ) );
  CLKBUF_X3 U841 ( .A(\RI5[0][27] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[27] ) );
  CLKBUF_X3 U850 ( .A(\RI5[2][110] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[110] )
         );
  CLKBUF_X3 U857 ( .A(\RI5[1][21] ), .Z(\MC_ARK_ARC_1_1/buf_datainput[21] ) );
  BUF_X2 U858 ( .A(\RI1[1][98] ), .Z(\SB1_1_15/i1[9] ) );
  CLKBUF_X2 U859 ( .A(\RI1[2][20] ), .Z(\SB1_2_28/i1[9] ) );
  BUF_X2 U860 ( .A(\RI1[3][188] ), .Z(\SB1_3_0/i1[9] ) );
  CLKBUF_X3 U861 ( .A(\RI1[1][63] ), .Z(\SB1_1_21/i0[8] ) );
  CLKBUF_X3 U865 ( .A(\RI3[1][29] ), .Z(\SB2_1_27/i0_3 ) );
  CLKBUF_X3 U867 ( .A(\RI5[0][3] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[3] ) );
  BUF_X2 U881 ( .A(\RI3[2][40] ), .Z(\SB2_2_25/i0_4 ) );
  CLKBUF_X3 U883 ( .A(\RI5[2][182] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[182] )
         );
  CLKBUF_X2 U888 ( .A(\RI1[2][146] ), .Z(\SB1_2_7/i1[9] ) );
  CLKBUF_X3 U893 ( .A(\RI1[2][135] ), .Z(\SB1_2_9/i0[8] ) );
  CLKBUF_X3 U897 ( .A(\RI1[2][9] ), .Z(\SB1_2_30/i0[8] ) );
  CLKBUF_X3 U905 ( .A(\RI3[2][173] ), .Z(\SB2_2_3/i0_3 ) );
  CLKBUF_X3 U906 ( .A(\RI1[2][110] ), .Z(\SB1_2_13/i1[9] ) );
  INV_X2 U908 ( .A(\RI1[3][119] ), .ZN(\SB1_3_12/i0_3 ) );
  CLKBUF_X3 U909 ( .A(\RI5[2][22] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[22] ) );
  CLKBUF_X2 U925 ( .A(\RI1[3][182] ), .Z(\SB1_3_1/i1[9] ) );
  CLKBUF_X1 U926 ( .A(\MC_ARK_ARC_1_0/buf_datainput[125] ), .Z(n1938) );
  CLKBUF_X3 U929 ( .A(\MC_ARK_ARC_1_0/buf_datainput[125] ), .Z(n1939) );
  NAND4_X1 U941 ( .A1(\SB2_0_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_11/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_11/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_11/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[125] ) );
  BUF_X2 U944 ( .A(\RI3[0][165] ), .Z(\SB2_0_4/i0[10] ) );
  CLKBUF_X3 U952 ( .A(\RI3[1][59] ), .Z(\SB2_1_22/i0_3 ) );
  CLKBUF_X3 U960 ( .A(\RI5[3][40] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[40] ) );
  BUF_X2 U966 ( .A(\RI1[2][171] ), .Z(\SB1_2_3/i0[8] ) );
  CLKBUF_X2 U974 ( .A(\RI1[1][188] ), .Z(\SB1_1_0/i1[9] ) );
  BUF_X2 U980 ( .A(\RI3[2][157] ), .Z(\SB2_2_5/i0[6] ) );
  INV_X2 U991 ( .A(\RI1[3][173] ), .ZN(\SB1_3_3/i0_3 ) );
  NAND4_X2 U993 ( .A1(\SB2_3_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_24/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][72] ) );
  INV_X2 U1002 ( .A(\RI1[3][155] ), .ZN(\SB1_3_6/i0_3 ) );
  BUF_X2 U1003 ( .A(\RI3[2][85] ), .Z(\SB2_2_17/i0[6] ) );
  CLKBUF_X1 U1011 ( .A(\MC_ARK_ARC_1_0/buf_datainput[116] ), .Z(n1940) );
  NAND4_X1 U1016 ( .A1(\SB2_0_15/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_15/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_0_15/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_15/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[116] ) );
  BUF_X2 U1024 ( .A(\RI3[3][139] ), .Z(\SB2_3_8/i0[6] ) );
  CLKBUF_X1 U1025 ( .A(\RI5[3][130] ), .Z(n1942) );
  CLKBUF_X1 U1027 ( .A(\RI5[3][130] ), .Z(n1943) );
  BUF_X1 U1028 ( .A(\RI5[3][130] ), .Z(n1944) );
  NAND4_X1 U1032 ( .A1(\SB2_3_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_11/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_11/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_11/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][130] ) );
  BUF_X2 U1034 ( .A(\RI1[2][87] ), .Z(\SB1_2_17/i0[8] ) );
  BUF_X2 U1036 ( .A(\MC_ARK_ARC_1_1/buf_datainput[35] ), .Z(n519) );
  BUF_X2 U1039 ( .A(\RI3[2][163] ), .Z(\SB2_2_4/i0[6] ) );
  BUF_X2 U1040 ( .A(\RI3[1][187] ), .Z(\SB2_1_0/i0[6] ) );
  CLKBUF_X3 U1043 ( .A(\RI3[1][185] ), .Z(\SB2_1_1/i0_3 ) );
  CLKBUF_X2 U1046 ( .A(\RI1[3][164] ), .Z(\SB1_3_4/i1[9] ) );
  BUF_X2 U1059 ( .A(\RI1[2][164] ), .Z(\SB1_2_4/i1[9] ) );
  CLKBUF_X3 U1073 ( .A(\RI3[1][161] ), .Z(\SB2_1_5/i0_3 ) );
  BUF_X2 U1074 ( .A(\RI3[2][136] ), .Z(\SB2_2_9/i0_4 ) );
  INV_X2 U1082 ( .A(n175), .ZN(\SB1_0_29/i0_3 ) );
  CLKBUF_X3 U1083 ( .A(\RI3[3][107] ), .Z(\SB2_3_14/i0_3 ) );
  BUF_X2 U1097 ( .A(\RI3[1][103] ), .Z(\SB2_1_14/i0[6] ) );
  CLKBUF_X3 U1118 ( .A(\RI1[2][74] ), .Z(\SB1_2_19/i1[9] ) );
  CLKBUF_X3 U1119 ( .A(\RI1[3][87] ), .Z(\SB1_3_17/i0[8] ) );
  CLKBUF_X3 U1153 ( .A(\RI1[3][128] ), .Z(\SB1_3_10/i1[9] ) );
  CLKBUF_X3 U1166 ( .A(n118), .Z(\SB1_0_19/i1[9] ) );
  BUF_X1 U1167 ( .A(n786), .Z(n1945) );
  BUF_X2 U1170 ( .A(\RI3[3][38] ), .Z(\SB2_3_25/i0_0 ) );
  CLKBUF_X3 U1191 ( .A(\RI3[2][131] ), .Z(\SB2_2_10/i0_3 ) );
  BUF_X2 U1204 ( .A(\RI3[3][49] ), .Z(\SB2_3_23/i0[6] ) );
  BUF_X2 U1252 ( .A(\RI3[3][140] ), .Z(\SB2_3_8/i0_0 ) );
  BUF_X2 U1264 ( .A(\RI3[2][90] ), .Z(\SB2_2_16/i0[9] ) );
  BUF_X2 U1273 ( .A(\RI1[1][176] ), .Z(\SB1_1_2/i1[9] ) );
  BUF_X2 U1274 ( .A(\RI3[3][73] ), .Z(\SB2_3_19/i0[6] ) );
  BUF_X2 U1277 ( .A(\RI3[2][121] ), .Z(\SB2_2_11/i0[6] ) );
  CLKBUF_X1 U1290 ( .A(\MC_ARK_ARC_1_3/buf_datainput[167] ), .Z(n1946) );
  BUF_X1 U1298 ( .A(\MC_ARK_ARC_1_3/buf_datainput[167] ), .Z(n1947) );
  CLKBUF_X1 U1321 ( .A(\MC_ARK_ARC_1_3/buf_datainput[167] ), .Z(n1948) );
  NAND4_X1 U1323 ( .A1(n2205), .A2(\SB2_3_4/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_3_4/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[167] ) );
  CLKBUF_X2 U1324 ( .A(\RI3[1][85] ), .Z(\SB2_1_17/i0[6] ) );
  BUF_X2 U1345 ( .A(\RI3[3][135] ), .Z(\SB2_3_9/i0[10] ) );
  BUF_X2 U1363 ( .A(\RI3[3][187] ), .Z(\SB2_3_0/i0[6] ) );
  CLKBUF_X3 U1368 ( .A(\RI1[2][122] ), .Z(\SB1_2_11/i1[9] ) );
  BUF_X2 U1369 ( .A(\RI3[3][182] ), .Z(\SB2_3_1/i0_0 ) );
  BUF_X2 U1377 ( .A(\RI1[2][152] ), .Z(\SB1_2_6/i1[9] ) );
  CLKBUF_X1 U1385 ( .A(\RI1[4][77] ), .Z(\SB3_19/i1_5 ) );
  INV_X1 U1425 ( .A(\RI1[4][77] ), .ZN(\SB3_19/i0_3 ) );
  CLKBUF_X3 U1427 ( .A(\RI1[3][50] ), .Z(\SB1_3_23/i1[9] ) );
  BUF_X2 U1428 ( .A(\RI3[3][146] ), .Z(\SB2_3_7/i0_0 ) );
  CLKBUF_X3 U1429 ( .A(\RI1[3][14] ), .Z(\SB1_3_29/i1[9] ) );
  BUF_X2 U1431 ( .A(\RI3[4][186] ), .Z(\SB4_0/i0[9] ) );
  BUF_X2 U1432 ( .A(\RI3[2][97] ), .Z(\SB2_2_15/i0[6] ) );
  BUF_X2 U1440 ( .A(\RI3[3][31] ), .Z(\SB2_3_26/i0[6] ) );
  BUF_X2 U1441 ( .A(\RI3[1][109] ), .Z(\SB2_1_13/i0[6] ) );
  BUF_X2 U1442 ( .A(\RI1[3][98] ), .Z(\SB1_3_15/i1[9] ) );
  BUF_X2 U1452 ( .A(\RI3[3][104] ), .Z(\SB2_3_14/i0_0 ) );
  BUF_X2 U1453 ( .A(\RI3[4][97] ), .Z(\SB4_15/i0[6] ) );
  CLKBUF_X3 U1463 ( .A(\RI1[4][26] ), .Z(\SB3_27/i1[9] ) );
  INV_X2 U1523 ( .A(n169), .ZN(\SB1_0_28/i0_3 ) );
  INV_X1 U1524 ( .A(\RI1[4][173] ), .ZN(\SB3_3/i0_3 ) );
  BUF_X2 U1533 ( .A(\RI1[2][170] ), .Z(\SB1_2_3/i1[9] ) );
  BUF_X2 U1541 ( .A(\RI1[1][93] ), .Z(\SB1_1_16/i0[8] ) );
  BUF_X2 U1550 ( .A(\RI3[3][85] ), .Z(\SB2_3_17/i0[6] ) );
  BUF_X2 U1552 ( .A(\RI3[3][122] ), .Z(\SB2_3_11/i0_0 ) );
  BUF_X2 U1556 ( .A(\RI1[1][8] ), .Z(\SB1_1_30/i1[9] ) );
  BUF_X2 U1574 ( .A(\RI1[3][69] ), .Z(\SB1_3_20/i0[8] ) );
  CLKBUF_X1 U1575 ( .A(\RI1[4][179] ), .Z(\SB3_2/i1_5 ) );
  INV_X1 U1584 ( .A(\RI1[4][179] ), .ZN(\SB3_2/i0_3 ) );
  BUF_X2 U1585 ( .A(\RI3[4][29] ), .Z(n1949) );
  CLKBUF_X2 U1592 ( .A(\RI5[3][158] ), .Z(n1955) );
  BUF_X2 U1594 ( .A(\RI5[2][111] ), .Z(n1950) );
  BUF_X2 U1604 ( .A(\RI1[2][32] ), .Z(\SB1_2_26/i1[9] ) );
  BUF_X2 U1615 ( .A(\MC_ARK_ARC_1_1/buf_datainput[71] ), .Z(n1952) );
  NAND4_X2 U1626 ( .A1(n1236), .A2(\SB2_1_15/Component_Function_2/NAND4_in[1] ), .A3(\SB2_1_15/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_15/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[116] ) );
  BUF_X2 U1636 ( .A(\MC_ARK_ARC_1_1/buf_datainput[178] ), .Z(n1953) );
  CLKBUF_X2 U1678 ( .A(\RI3[1][14] ), .Z(\SB2_1_29/i0_0 ) );
  BUF_X2 U1711 ( .A(\RI1[1][135] ), .Z(\SB1_1_9/i0[8] ) );
  CLKBUF_X2 U1712 ( .A(\MC_ARK_ARC_1_0/buf_datainput[41] ), .Z(n1961) );
  BUF_X2 U1714 ( .A(\MC_ARK_ARC_1_0/buf_datainput[189] ), .Z(n1495) );
  BUF_X1 U1718 ( .A(\RI3[0][54] ), .Z(\SB2_0_22/i0[9] ) );
  BUF_X1 U1722 ( .A(Key[91]), .Z(n423) );
  BUF_X1 U1728 ( .A(Key[142]), .Z(n461) );
  BUF_X1 U1750 ( .A(\RI3[4][145] ), .Z(\SB4_7/i0[6] ) );
  AND4_X1 U1760 ( .A1(\SB3_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_2/NAND4_in[3] ), .ZN(n2113) );
  BUF_X2 U1780 ( .A(\RI5[3][136] ), .Z(\MC_ARK_ARC_1_3/buf_datainput[136] ) );
  NAND4_X2 U1786 ( .A1(\SB2_3_12/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_12/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_12/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_12/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[124] ) );
  NAND4_X1 U1795 ( .A1(n1242), .A2(\SB2_3_16/Component_Function_5/NAND4_in[3] ), .A3(\SB2_3_16/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_16/Component_Function_5/NAND4_in[0] ), .ZN(n2145) );
  NAND4_X2 U1796 ( .A1(\SB2_3_31/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_31/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_31/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_31/Component_Function_4/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[10] ) );
  BUF_X2 U1800 ( .A(\RI1[3][152] ), .Z(\SB1_3_6/i1[9] ) );
  BUF_X2 U1812 ( .A(\RI1[3][176] ), .Z(\SB1_3_2/i1[9] ) );
  BUF_X2 U1813 ( .A(\RI5[2][128] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[128] ) );
  BUF_X2 U1815 ( .A(\RI5[2][56] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[56] ) );
  BUF_X2 U1821 ( .A(\RI5[2][42] ), .Z(\MC_ARK_ARC_1_2/buf_datainput[42] ) );
  BUF_X2 U1822 ( .A(\MC_ARK_ARC_1_2/buf_datainput[89] ), .Z(n1956) );
  BUF_X2 U1823 ( .A(\MC_ARK_ARC_1_2/buf_datainput[118] ), .Z(n1957) );
  NAND4_X1 U1827 ( .A1(n1584), .A2(\SB2_2_23/Component_Function_3/NAND4_in[1] ), .A3(\SB2_2_23/Component_Function_3/NAND4_in[2] ), .A4(n1014), .ZN(n2101) );
  BUF_X2 U1833 ( .A(\RI3[2][152] ), .Z(\SB2_2_6/i0_0 ) );
  AND4_X1 U1834 ( .A1(\SB1_2_1/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_1/Component_Function_2/NAND4_in[2] ), .A4(n704), .ZN(n2118) );
  BUF_X2 U1841 ( .A(\RI1[2][116] ), .Z(\SB1_2_12/i1[9] ) );
  BUF_X2 U1848 ( .A(\RI1[2][188] ), .Z(\SB1_2_0/i1[9] ) );
  NAND4_X2 U1870 ( .A1(\SB2_1_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_2/NAND4_in[3] ), .A4(n2209), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[50] ) );
  NAND4_X2 U1880 ( .A1(n743), .A2(\SB2_1_10/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB2_1_10/Component_Function_2/NAND4_in[3] ), .A4(n2021), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[146] ) );
  BUF_X1 U1894 ( .A(\RI1[1][26] ), .Z(\SB1_1_27/i1[9] ) );
  BUF_X2 U1897 ( .A(\RI5[0][55] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[55] ) );
  BUF_X2 U1901 ( .A(\RI5[0][30] ), .Z(\MC_ARK_ARC_1_0/buf_datainput[30] ) );
  BUF_X2 U1906 ( .A(\MC_ARK_ARC_1_0/buf_datainput[189] ), .Z(n1959) );
  BUF_X2 U1915 ( .A(\MC_ARK_ARC_1_0/buf_datainput[29] ), .Z(n1960) );
  NAND4_X2 U1916 ( .A1(n2024), .A2(\SB2_0_31/Component_Function_4/NAND4_in[3] ), .A3(\SB2_0_31/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_31/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[10] ) );
  BUF_X2 U1932 ( .A(\MC_ARK_ARC_1_0/buf_datainput[107] ), .Z(n1962) );
  BUF_X2 U1943 ( .A(\RI3[0][127] ), .Z(\SB2_0_10/i0[6] ) );
  INV_X1 U1944 ( .A(n11), .ZN(\SB1_0_1/i0[6] ) );
  BUF_X1 U1967 ( .A(n87), .Z(\SB1_0_14/i0[8] ) );
  CLKBUF_X1 U1981 ( .A(n143), .Z(\SB1_0_23/i1_7 ) );
  BUF_X1 U1982 ( .A(n147), .Z(\SB1_0_24/i0[8] ) );
  BUF_X1 U1996 ( .A(n148), .Z(\SB1_0_24/i1[9] ) );
  BUF_X1 U1997 ( .A(n135), .Z(\SB1_0_22/i0[8] ) );
  CLKBUF_X1 U2024 ( .A(n43), .Z(\SB1_0_7/i1_5 ) );
  BUF_X1 U2049 ( .A(n46), .Z(\SB1_0_7/i1[9] ) );
  BUF_X1 U2050 ( .A(\RI3[0][48] ), .Z(\SB2_0_23/i0[9] ) );
  CLKBUF_X1 U2051 ( .A(\RI1[1][163] ), .Z(\SB1_1_4/i1_7 ) );
  CLKBUF_X3 U2052 ( .A(\RI1[1][3] ), .Z(\SB1_1_31/i0[8] ) );
  BUF_X1 U2065 ( .A(\RI1[1][131] ), .Z(\SB1_1_10/i1_5 ) );
  BUF_X1 U2076 ( .A(\RI1[1][134] ), .Z(\SB1_1_9/i1[9] ) );
  CLKBUF_X3 U2080 ( .A(\RI1[1][177] ), .Z(\SB1_1_2/i0[8] ) );
  BUF_X1 U2098 ( .A(\RI3[1][180] ), .Z(\SB2_1_1/i0[9] ) );
  BUF_X1 U2121 ( .A(\RI3[1][96] ), .Z(\SB2_1_15/i0[9] ) );
  BUF_X1 U2129 ( .A(\RI3[1][144] ), .Z(\SB2_1_7/i0[9] ) );
  BUF_X1 U2148 ( .A(\MC_ARK_ARC_1_1/buf_datainput[35] ), .Z(n517) );
  NAND4_X2 U2152 ( .A1(\SB2_1_20/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_20/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_20/Component_Function_3/NAND4_in[2] ), .A4(n1046), .ZN(
        \RI5[1][81] ) );
  BUF_X1 U2153 ( .A(\RI1[2][179] ), .Z(\SB1_2_2/i1_5 ) );
  BUF_X1 U2154 ( .A(\RI3[2][96] ), .Z(\SB2_2_15/i0[9] ) );
  BUF_X1 U2159 ( .A(\RI3[2][120] ), .Z(\SB2_2_11/i0[9] ) );
  BUF_X1 U2162 ( .A(\RI1[3][99] ), .Z(\SB1_3_15/i0[8] ) );
  BUF_X1 U2165 ( .A(\RI3[3][0] ), .Z(\SB2_3_31/i0[9] ) );
  CLKBUF_X1 U2167 ( .A(\RI1[4][138] ), .Z(\SB3_8/i3[0] ) );
  BUF_X1 U2168 ( .A(\RI3[4][59] ), .Z(n851) );
  BUF_X1 U2175 ( .A(\RI3[4][156] ), .Z(\SB4_5/i0[9] ) );
  INV_X1 U2178 ( .A(\MC_ARK_ARC_1_3/buf_keyinput[44] ), .ZN(n256) );
  INV_X1 U2182 ( .A(\MC_ARK_ARC_1_1/buf_keyinput[183] ), .ZN(n208) );
  INV_X1 U2188 ( .A(\MC_ARK_ARC_1_0/buf_keyinput[136] ), .ZN(n195) );
  INV_X1 U2200 ( .A(n403), .ZN(n346) );
  INV_X1 U2204 ( .A(n397), .ZN(n307) );
  INV_X1 U2210 ( .A(n391), .ZN(n250) );
  INV_X1 U2213 ( .A(n435), .ZN(n268) );
  INV_X1 U2226 ( .A(n467), .ZN(n264) );
  INV_X1 U2260 ( .A(n455), .ZN(n314) );
  INV_X1 U2263 ( .A(Key[153]), .ZN(n230) );
  AND4_X1 U2288 ( .A1(\SB3_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_30/Component_Function_4/NAND4_in[3] ), .ZN(n1963) );
  AND4_X1 U2290 ( .A1(\SB3_31/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_5/NAND4_in[3] ), .ZN(n1964) );
  AND4_X1 U2312 ( .A1(\SB1_3_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_19/Component_Function_1/NAND4_in[3] ), .ZN(n1965) );
  INV_X1 U2313 ( .A(\MC_ARK_ARC_1_1/buf_keyinput[107] ), .ZN(n281) );
  NAND3_X1 U2326 ( .A1(\SB1_1_18/i3[0] ), .A2(\SB1_1_18/i0_0 ), .A3(
        \SB1_1_18/i1_7 ), .ZN(\SB1_1_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2341 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i1_5 ), .A3(
        \SB2_0_10/i1[9] ), .ZN(\SB2_0_10/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U2342 ( .A1(\SB3_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_19/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_5/NAND4_in[0] ), .A4(n1966), .ZN(
        \RI3[4][77] ) );
  NAND3_X1 U2349 ( .A1(\SB3_19/i0[9] ), .A2(\SB3_19/i0_4 ), .A3(\SB3_19/i0[6] ), .ZN(n1966) );
  NAND4_X2 U2356 ( .A1(\SB1_3_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_26/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_3_26/Component_Function_4/NAND4_in[1] ), .A4(n1967), .ZN(
        \SB2_3_25/i0_4 ) );
  NAND3_X1 U2363 ( .A1(\SB1_3_26/i1[9] ), .A2(\SB1_3_26/i1_5 ), .A3(
        \SB1_3_26/i0_4 ), .ZN(n1967) );
  NAND4_X1 U2364 ( .A1(\SB1_1_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_19/Component_Function_5/NAND4_in[0] ), .A4(n1968), .ZN(
        \RI3[1][77] ) );
  NAND3_X1 U2386 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i1[9] ), .A3(
        \SB1_1_19/i0_4 ), .ZN(n1968) );
  NAND4_X1 U2397 ( .A1(\SB3_29/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_29/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_29/Component_Function_2/NAND4_in[3] ), .A4(n1969), .ZN(
        \RI3[4][32] ) );
  NAND3_X1 U2399 ( .A1(\SB3_29/i0[9] ), .A2(\SB3_29/i0[8] ), .A3(\SB3_29/i0_3 ), .ZN(n1969) );
  NAND3_X1 U2412 ( .A1(\SB1_2_16/i1[9] ), .A2(\SB1_2_16/i0_4 ), .A3(
        \SB1_2_16/i1_5 ), .ZN(\SB1_2_16/Component_Function_4/NAND4_in[3] ) );
  NAND4_X1 U2415 ( .A1(\SB2_2_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_21/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_21/Component_Function_4/NAND4_in[1] ), .A4(n1970), .ZN(
        \RI5[2][70] ) );
  NAND3_X1 U2416 ( .A1(\SB2_2_21/i0_4 ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB2_2_21/i1[9] ), .ZN(n1970) );
  NAND4_X1 U2417 ( .A1(\SB1_1_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_20/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_1_20/Component_Function_5/NAND4_in[0] ), .A4(n1971), .ZN(
        \RI3[1][71] ) );
  NAND3_X1 U2422 ( .A1(\SB1_1_20/i0[6] ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i0[9] ), .ZN(n1971) );
  NAND3_X1 U2428 ( .A1(\SB2_3_12/i0_0 ), .A2(\SB2_3_12/i3[0] ), .A3(
        \SB2_3_12/i1_7 ), .ZN(\SB2_3_12/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U2432 ( .A1(\SB2_0_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_21/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[75] ) );
  NAND4_X1 U2435 ( .A1(\SB3_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_5/NAND4_in[0] ), .A4(n1972), .ZN(
        \RI3[4][41] ) );
  NAND3_X1 U2443 ( .A1(\SB3_25/i0[9] ), .A2(\SB3_25/i0[6] ), .A3(\SB3_25/i0_4 ), .ZN(n1972) );
  NAND4_X2 U2450 ( .A1(\SB2_3_21/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_21/Component_Function_4/NAND4_in[1] ), .A4(n1973), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[70] ) );
  NAND3_X1 U2464 ( .A1(\SB2_3_21/i1_5 ), .A2(\SB2_3_21/i1[9] ), .A3(
        \RI3[3][64] ), .ZN(n1973) );
  XNOR2_X1 U2465 ( .A(n1974), .B(n418), .ZN(Ciphertext[180]) );
  NAND4_X1 U2468 ( .A1(\SB4_1/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_1/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_1/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_1/Component_Function_0/NAND4_in[0] ), .ZN(n1974) );
  NAND4_X1 U2469 ( .A1(\SB2_2_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_9/Component_Function_4/NAND4_in[1] ), .A4(n1975), .ZN(
        \RI5[2][142] ) );
  NAND3_X1 U2474 ( .A1(\SB2_2_9/i0_4 ), .A2(\SB2_2_9/i1[9] ), .A3(
        \SB2_2_9/i1_5 ), .ZN(n1975) );
  XNOR2_X1 U2480 ( .A(n1976), .B(n328), .ZN(Ciphertext[36]) );
  NAND4_X1 U2482 ( .A1(\SB4_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_25/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_25/Component_Function_0/NAND4_in[1] ), .ZN(n1976) );
  NAND3_X1 U2491 ( .A1(\SB2_0_0/i0_4 ), .A2(\SB2_0_0/i1[9] ), .A3(
        \SB2_0_0/i1_5 ), .ZN(n1689) );
  NAND3_X1 U2492 ( .A1(\SB4_26/i0_0 ), .A2(\SB4_26/i1_5 ), .A3(\SB4_26/i0_4 ), 
        .ZN(n1996) );
  NAND3_X1 U2500 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0[10] ), .A3(
        \SB2_2_28/i0[6] ), .ZN(n2064) );
  NAND3_X1 U2548 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i1[9] ), .A3(
        \SB2_1_24/i1_7 ), .ZN(\SB2_1_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2549 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i1_5 ), .A3(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2559 ( .A1(\SB1_3_22/i0[10] ), .A2(\SB1_3_22/i0[9] ), .A3(
        \SB1_3_22/i0_3 ), .ZN(\SB1_3_22/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U2560 ( .A1(\SB2_1_6/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_6/Component_Function_4/NAND4_in[1] ), .A4(n1977), .ZN(
        \RI5[1][160] ) );
  NAND3_X1 U2561 ( .A1(\SB2_1_6/i0[9] ), .A2(\SB2_1_6/i0[10] ), .A3(
        \SB2_1_6/i0_3 ), .ZN(n1977) );
  NAND3_X1 U2567 ( .A1(\SB3_29/i0_0 ), .A2(\SB3_29/i1_5 ), .A3(\SB3_29/i0_4 ), 
        .ZN(\SB3_29/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U2568 ( .A1(\SB1_1_1/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_1/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_1_1/Component_Function_0/NAND4_in[1] ), .A4(n1978), .ZN(
        \RI3[1][18] ) );
  NAND3_X1 U2579 ( .A1(\SB1_1_1/i0[7] ), .A2(\SB1_1_1/i0_0 ), .A3(
        \SB1_1_1/i0_3 ), .ZN(n1978) );
  NAND3_X1 U2580 ( .A1(\SB2_0_28/i0[9] ), .A2(\SB2_0_28/i0_3 ), .A3(
        \SB2_0_28/i0[10] ), .ZN(\SB2_0_28/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2590 ( .A1(\SB2_1_2/i0[9] ), .A2(\SB2_1_2/i0_3 ), .A3(
        \SB2_1_2/i0[10] ), .ZN(\SB2_1_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2597 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i0[10] ), .A3(
        \SB1_3_1/i0[9] ), .ZN(\SB1_3_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2610 ( .A1(\SB1_1_10/i1[9] ), .A2(\SB1_1_10/i0[10] ), .A3(
        \SB1_1_10/i1_7 ), .ZN(\SB1_1_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2611 ( .A1(\SB2_3_3/i0_0 ), .A2(\SB2_3_3/i1_7 ), .A3(
        \SB2_3_3/i3[0] ), .ZN(\SB2_3_3/Component_Function_4/NAND4_in[1] ) );
  XNOR2_X1 U2632 ( .A(n1979), .B(n354), .ZN(Ciphertext[32]) );
  NAND4_X1 U2633 ( .A1(\SB4_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_26/Component_Function_2/NAND4_in[1] ), .A3(n1548), .A4(n1996), 
        .ZN(n1979) );
  NAND4_X2 U2645 ( .A1(\SB2_3_3/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_3/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_3/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_3_3/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[178] ) );
  NAND4_X2 U2646 ( .A1(\SB2_3_3/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_3/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_3/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_3_3/Component_Function_3/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[183] ) );
  NAND3_X1 U2655 ( .A1(\SB2_2_26/i0_3 ), .A2(\SB2_2_26/i1[9] ), .A3(
        \SB2_2_26/i0[6] ), .ZN(\SB2_2_26/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U2656 ( .A1(\SB1_3_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_8/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_8/Component_Function_1/NAND4_in[0] ), .A4(n1980), .ZN(
        \RI3[3][163] ) );
  NAND3_X1 U2663 ( .A1(\SB1_3_8/i1_7 ), .A2(\SB1_3_8/i0_4 ), .A3(
        \SB1_3_8/i0[8] ), .ZN(n1980) );
  NAND4_X1 U2664 ( .A1(\SB4_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_2/Component_Function_3/NAND4_in[3] ), .A4(n1981), .ZN(n1590) );
  NAND3_X1 U2698 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i1[9] ), .A3(\SB4_2/i1_7 ), 
        .ZN(n1981) );
  NAND3_X1 U2699 ( .A1(\SB3_4/i0_0 ), .A2(\SB3_4/i0_4 ), .A3(\SB3_4/i0_3 ), 
        .ZN(\SB3_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2712 ( .A1(\SB2_0_8/i0[6] ), .A2(\SB2_0_8/i0_0 ), .A3(
        \SB2_0_8/i0[10] ), .ZN(\SB2_0_8/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U2719 ( .A1(\SB1_3_8/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_8/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_8/Component_Function_2/NAND4_in[2] ), .A4(n1982), .ZN(
        \RI3[3][158] ) );
  NAND3_X1 U2729 ( .A1(\SB1_3_8/i0_0 ), .A2(\SB1_3_8/i0_4 ), .A3(
        \SB1_3_8/i1_5 ), .ZN(n1982) );
  NAND3_X1 U2734 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0[10] ), .A3(
        \SB1_0_28/i0[9] ), .ZN(\SB1_0_28/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U2735 ( .A1(\SB1_3_3/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_3/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_3/Component_Function_2/NAND4_in[2] ), .A4(n1983), .ZN(
        \RI3[3][188] ) );
  NAND3_X1 U2744 ( .A1(\SB1_3_3/i0_0 ), .A2(\SB1_3_3/i0_4 ), .A3(
        \SB1_3_3/i1_5 ), .ZN(n1983) );
  NAND4_X1 U2761 ( .A1(\SB3_8/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_8/Component_Function_4/NAND4_in[1] ), .A4(n1984), .ZN(
        \RI3[4][148] ) );
  NAND3_X1 U2762 ( .A1(\SB3_8/i0[9] ), .A2(\SB3_8/i0[10] ), .A3(\SB3_8/i0_3 ), 
        .ZN(n1984) );
  NAND3_X1 U2786 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i1[9] ), .A3(
        \SB2_2_27/i0[6] ), .ZN(\SB2_2_27/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U2791 ( .A1(\SB4_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_7/Component_Function_2/NAND4_in[2] ), .A3(n1779), .A4(n1985), 
        .ZN(n2242) );
  NAND3_X1 U2794 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i0_0 ), .A3(\SB4_7/i1_5 ), 
        .ZN(n1985) );
  NAND4_X1 U2795 ( .A1(\SB1_2_26/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_26/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_26/Component_Function_5/NAND4_in[0] ), .A4(n1986), .ZN(
        \RI3[2][35] ) );
  NAND3_X1 U2825 ( .A1(\SB1_2_26/i1[9] ), .A2(\SB1_2_26/i0_3 ), .A3(
        \SB1_2_26/i0_4 ), .ZN(n1986) );
  NAND3_X1 U2826 ( .A1(\SB1_1_4/i1[9] ), .A2(\SB1_1_4/i0[10] ), .A3(
        \SB1_1_4/i1_7 ), .ZN(\SB1_1_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2830 ( .A1(\SB2_2_15/i0[9] ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i0[10] ), .ZN(\SB2_2_15/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2831 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i0[9] ), .A3(\SB4_19/i0[8] ), .ZN(\SB4_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2835 ( .A1(\SB2_0_21/i0[10] ), .A2(\SB2_0_21/i1[9] ), .A3(
        \SB2_0_21/i1_7 ), .ZN(\SB2_0_21/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U2853 ( .A1(\SB1_3_20/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_3_20/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_5/NAND4_in[0] ), .A4(n1987), .ZN(
        \RI3[3][71] ) );
  NAND3_X1 U2879 ( .A1(\SB1_3_20/i1[9] ), .A2(\SB1_3_20/i0_3 ), .A3(
        \SB1_3_20/i0_4 ), .ZN(n1987) );
  NAND3_X1 U2910 ( .A1(\SB1_0_3/i1_7 ), .A2(\SB1_0_3/i0[10] ), .A3(
        \SB1_0_3/i1[9] ), .ZN(\SB1_0_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2939 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0_0 ), .A3(
        \SB2_0_4/i0[7] ), .ZN(\SB2_0_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2940 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0[6] ), .A3(
        \SB2_1_30/i0[10] ), .ZN(\SB2_1_30/Component_Function_2/NAND4_in[1] )
         );
  NAND4_X1 U2968 ( .A1(\SB4_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_6/Component_Function_2/NAND4_in[3] ), .A3(
        \SB4_6/Component_Function_2/NAND4_in[2] ), .A4(n1988), .ZN(n2047) );
  NAND3_X1 U2982 ( .A1(\SB4_6/i0[10] ), .A2(\SB4_6/i1_5 ), .A3(\SB4_6/i1[9] ), 
        .ZN(n1988) );
  NAND4_X1 U2983 ( .A1(\SB1_2_28/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_2_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_5/NAND4_in[0] ), .A4(n1989), .ZN(
        \RI3[2][23] ) );
  NAND3_X1 U2984 ( .A1(\SB1_2_28/i1[9] ), .A2(\SB1_2_28/i0_3 ), .A3(
        \SB1_2_28/i0_4 ), .ZN(n1989) );
  NAND3_X1 U2986 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0[9] ), .A3(
        \SB2_1_30/i0[10] ), .ZN(n2070) );
  NAND4_X1 U3010 ( .A1(\SB1_1_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_5/NAND4_in[0] ), .A4(n1990), .ZN(
        \RI3[1][11] ) );
  NAND3_X1 U3017 ( .A1(\SB1_1_30/i0_4 ), .A2(\SB1_1_30/i0[9] ), .A3(
        \SB1_1_30/i0[6] ), .ZN(n1990) );
  NAND4_X2 U3022 ( .A1(\SB2_2_5/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_2_5/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_5/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_2_5/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[176] ) );
  NAND4_X2 U3025 ( .A1(\SB2_0_16/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_16/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_0_16/Component_Function_2/NAND4_in[3] ), .A4(n1991), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[110] ) );
  NAND3_X1 U3040 ( .A1(\SB2_0_16/i0[10] ), .A2(\SB2_0_16/i0_3 ), .A3(
        \SB2_0_16/i0[6] ), .ZN(n1991) );
  OR3_X1 U3043 ( .A1(\RI1[1][9] ), .A2(\RI1[1][7] ), .A3(\RI1[1][8] ), .ZN(
        \SB1_1_30/Component_Function_5/NAND4_in[1] ) );
  NAND4_X1 U3048 ( .A1(\SB3_2/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_2/Component_Function_5/NAND4_in[2] ), .A3(
        \SB3_2/Component_Function_5/NAND4_in[0] ), .A4(n1992), .ZN(
        \RI3[4][179] ) );
  NAND3_X1 U3067 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i0[9] ), .A3(\SB3_2/i0_4 ), 
        .ZN(n1992) );
  NAND4_X1 U3069 ( .A1(\SB1_0_19/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_19/Component_Function_1/NAND4_in[0] ), .A4(n1993), .ZN(
        \RI3[0][97] ) );
  NAND3_X1 U3083 ( .A1(\SB1_0_19/i0[9] ), .A2(\SB1_0_19/i1_5 ), .A3(
        \SB1_0_19/i0[6] ), .ZN(n1993) );
  NAND4_X1 U3084 ( .A1(\SB3_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_8/Component_Function_5/NAND4_in[0] ), .A4(n1994), .ZN(
        \RI3[4][143] ) );
  NAND3_X1 U3087 ( .A1(\SB3_8/i1[9] ), .A2(\SB3_8/i0_4 ), .A3(\SB3_8/i0_3 ), 
        .ZN(n1994) );
  NAND3_X1 U3090 ( .A1(\SB2_0_9/i0[10] ), .A2(\SB2_0_9/i1_5 ), .A3(
        \SB2_0_9/i1[9] ), .ZN(\SB2_0_9/Component_Function_2/NAND4_in[0] ) );
  XNOR2_X1 U3094 ( .A(n1995), .B(n348), .ZN(Ciphertext[170]) );
  NAND4_X1 U3098 ( .A1(\SB4_3/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_3/Component_Function_2/NAND4_in[1] ), .A3(n2244), .A4(n2010), 
        .ZN(n1995) );
  NAND4_X4 U3115 ( .A1(n1243), .A2(\SB2_1_27/Component_Function_5/NAND4_in[3] ), .A3(\SB2_1_27/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[29] ) );
  NAND3_X1 U3117 ( .A1(\SB1_3_3/i0[8] ), .A2(\SB1_3_3/i0_4 ), .A3(
        \SB1_3_3/i1_7 ), .ZN(\SB1_3_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3126 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0[8] ), .A3(
        \SB1_0_23/i0[9] ), .ZN(\SB1_0_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3160 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB2_3_9/i0_0 ), .A3(
        \SB2_3_9/i0[7] ), .ZN(\SB2_3_9/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U3161 ( .A1(\SB1_1_25/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_25/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_25/Component_Function_2/NAND4_in[2] ), .A4(n1997), .ZN(
        \RI3[1][56] ) );
  NAND3_X1 U3227 ( .A1(\SB1_1_25/i0_0 ), .A2(\SB1_1_25/i0_4 ), .A3(
        \SB1_1_25/i1_5 ), .ZN(n1997) );
  NAND3_X1 U3228 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i1[9] ), .A3(
        \SB2_0_27/i1_7 ), .ZN(\SB2_0_27/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U3233 ( .A1(n1209), .A2(\SB2_1_1/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_1_1/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[185] ) );
  NAND3_X1 U3234 ( .A1(\SB2_0_13/i0[6] ), .A2(\SB2_0_13/i0[10] ), .A3(
        \SB2_0_13/i0_0 ), .ZN(\SB2_0_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3238 ( .A1(\SB2_0_28/i0[9] ), .A2(\SB2_0_28/i0_3 ), .A3(
        \SB2_0_28/i0[8] ), .ZN(\SB2_0_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3243 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0_4 ), .A3(
        \SB2_1_18/i0_0 ), .ZN(\SB2_1_18/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U3250 ( .A1(n1345), .A2(\SB2_3_2/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_3_2/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[179] ) );
  NAND3_X1 U3251 ( .A1(\SB1_0_6/i0[10] ), .A2(\SB1_0_6/i0_0 ), .A3(
        \SB1_0_6/i0[6] ), .ZN(\SB1_0_6/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U3270 ( .A(n1999), .B(n1998), .ZN(\RI1[4][146] ) );
  XNOR2_X1 U3279 ( .A(\MC_ARK_ARC_1_3/temp2[146] ), .B(
        \MC_ARK_ARC_1_3/temp4[146] ), .ZN(n1998) );
  XNOR2_X1 U3280 ( .A(\MC_ARK_ARC_1_3/temp1[146] ), .B(
        \MC_ARK_ARC_1_3/temp3[146] ), .ZN(n1999) );
  NAND3_X1 U3289 ( .A1(\SB2_3_31/i0_0 ), .A2(\SB2_3_31/i1_5 ), .A3(n1651), 
        .ZN(\SB2_3_31/Component_Function_2/NAND4_in[3] ) );
  INV_X2 U3320 ( .A(\RI1[1][185] ), .ZN(\SB1_1_1/i0_3 ) );
  XNOR2_X1 U3321 ( .A(n736), .B(\MC_ARK_ARC_1_0/temp5[185] ), .ZN(
        \RI1[1][185] ) );
  XNOR2_X1 U3326 ( .A(n2000), .B(n245), .ZN(Ciphertext[117]) );
  NAND4_X1 U3336 ( .A1(\SB4_12/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_12/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_12/Component_Function_3/NAND4_in[3] ), .ZN(n2000) );
  NAND4_X1 U3339 ( .A1(\SB2_0_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_3/NAND4_in[2] ), .A3(n1800), .A4(n2001), 
        .ZN(\RI5[0][171] ) );
  NAND3_X1 U3347 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0_4 ), .A3(
        \SB2_0_5/i0_0 ), .ZN(n2001) );
  XNOR2_X1 U3373 ( .A(\MC_ARK_ARC_1_0/temp6[118] ), .B(n2002), .ZN(
        \RI1[1][118] ) );
  XNOR2_X1 U3374 ( .A(\MC_ARK_ARC_1_0/temp2[118] ), .B(
        \MC_ARK_ARC_1_0/temp1[118] ), .ZN(n2002) );
  NAND4_X1 U3387 ( .A1(\SB2_0_22/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_0_22/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_22/Component_Function_4/NAND4_in[1] ), .A4(n2003), .ZN(
        \RI5[0][64] ) );
  NAND3_X1 U3394 ( .A1(\SB2_0_22/i0_4 ), .A2(\SB2_0_22/i1_5 ), .A3(
        \SB2_0_22/i1[9] ), .ZN(n2003) );
  XNOR2_X1 U3396 ( .A(n2004), .B(n234), .ZN(Ciphertext[160]) );
  NAND4_X1 U3397 ( .A1(\SB4_5/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_5/Component_Function_4/NAND4_in[0] ), .A3(n1146), .A4(n1915), 
        .ZN(n2004) );
  NAND4_X1 U3402 ( .A1(\SB1_1_12/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_12/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_12/Component_Function_1/NAND4_in[0] ), .A4(n2005), .ZN(
        \RI3[1][139] ) );
  NAND3_X1 U3404 ( .A1(\SB1_1_12/i1_7 ), .A2(\SB1_1_12/i0_4 ), .A3(
        \SB1_1_12/i0[8] ), .ZN(n2005) );
  NAND3_X1 U3427 ( .A1(\SB1_3_23/i1[9] ), .A2(\SB1_3_23/i0_4 ), .A3(
        \SB1_3_23/i1_5 ), .ZN(\SB1_3_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3432 ( .A1(\SB2_0_16/i0_0 ), .A2(\SB2_0_16/i3[0] ), .A3(
        \SB2_0_16/i1_7 ), .ZN(\SB2_0_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3436 ( .A1(\SB1_0_18/i0[10] ), .A2(\SB1_0_18/i0_0 ), .A3(
        \SB1_0_18/i0[6] ), .ZN(\SB1_0_18/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3437 ( .A1(\SB1_3_27/i1[9] ), .A2(\SB1_3_27/i0_4 ), .A3(
        \SB1_3_27/i1_5 ), .ZN(\SB1_3_27/Component_Function_4/NAND4_in[3] ) );
  NAND4_X4 U3438 ( .A1(n1295), .A2(\SB2_3_26/Component_Function_5/NAND4_in[1] ), .A3(\SB2_3_26/Component_Function_5/NAND4_in[3] ), .A4(n2006), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[35] ) );
  NAND2_X1 U3446 ( .A1(\SB2_3_26/i0_0 ), .A2(\SB2_3_26/i3[0] ), .ZN(n2006) );
  NAND4_X4 U3447 ( .A1(\SB2_0_30/Component_Function_4/NAND4_in[2] ), .A2(n1687), .A3(\SB2_0_30/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_30/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[16] ) );
  NAND4_X2 U3466 ( .A1(\SB2_1_18/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_18/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_18/Component_Function_2/NAND4_in[0] ), .A4(n2007), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[98] ) );
  NAND3_X1 U3467 ( .A1(\SB2_1_18/i0_4 ), .A2(\SB2_1_18/i0_0 ), .A3(
        \SB2_1_18/i1_5 ), .ZN(n2007) );
  NAND4_X1 U3470 ( .A1(\SB2_1_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_28/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_28/Component_Function_4/NAND4_in[1] ), .A4(n2008), .ZN(
        \RI5[1][28] ) );
  NAND3_X1 U3471 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0[10] ), .A3(
        \SB2_1_28/i0[9] ), .ZN(n2008) );
  NAND4_X1 U3528 ( .A1(\SB2_3_10/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_3_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_10/Component_Function_5/NAND4_in[0] ), .A4(n2009), .ZN(
        \RI5[3][131] ) );
  NAND3_X1 U3533 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0_4 ), .A3(
        \SB2_3_10/i1[9] ), .ZN(n2009) );
  NAND3_X1 U3534 ( .A1(\SB4_3/i0_4 ), .A2(\SB4_3/i0_0 ), .A3(\SB4_3/i1_5 ), 
        .ZN(n2010) );
  NAND4_X1 U3574 ( .A1(\SB1_1_29/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_29/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_29/Component_Function_5/NAND4_in[0] ), .A4(n2011), .ZN(
        \RI3[1][17] ) );
  NAND3_X1 U3575 ( .A1(\SB1_1_29/i1[9] ), .A2(\SB1_1_29/i0_3 ), .A3(
        \SB1_1_29/i0_4 ), .ZN(n2011) );
  NAND3_X1 U3579 ( .A1(\SB1_0_4/i0[7] ), .A2(\SB1_0_4/i0_3 ), .A3(
        \SB1_0_4/i0_0 ), .ZN(\SB1_0_4/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U3580 ( .A1(\SB2_1_31/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_31/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_31/Component_Function_1/NAND4_in[0] ), .A4(n2012), .ZN(
        \RI5[1][25] ) );
  NAND3_X1 U3591 ( .A1(\SB2_1_31/i0_4 ), .A2(\SB2_1_31/i1_7 ), .A3(
        \SB2_1_31/i0[8] ), .ZN(n2012) );
  NAND4_X1 U3606 ( .A1(\SB2_2_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_3/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_3/Component_Function_2/NAND4_in[3] ), .A4(n2013), .ZN(
        \RI5[2][188] ) );
  NAND3_X1 U3633 ( .A1(\SB2_2_3/i0[9] ), .A2(\SB2_2_3/i0_3 ), .A3(
        \SB2_2_3/i0[8] ), .ZN(n2013) );
  NAND4_X2 U3641 ( .A1(n1203), .A2(\SB2_0_21/Component_Function_4/NAND4_in[0] ), .A3(\SB2_0_21/Component_Function_4/NAND4_in[1] ), .A4(n2014), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[70] ) );
  NAND3_X1 U3643 ( .A1(\SB2_0_21/i0_4 ), .A2(\SB2_0_21/i1[9] ), .A3(
        \SB2_0_21/i1_5 ), .ZN(n2014) );
  NAND3_X1 U3663 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0_4 ), .A3(
        \SB2_3_23/i1[9] ), .ZN(\SB2_3_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3705 ( .A1(\SB1_1_4/i0[7] ), .A2(\SB1_1_4/i0_0 ), .A3(
        \SB1_1_4/i0_3 ), .ZN(\SB1_1_4/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U3721 ( .A1(\SB2_2_12/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_12/Component_Function_4/NAND4_in[1] ), .A4(n2015), .ZN(
        \RI5[2][124] ) );
  NAND3_X1 U3724 ( .A1(\SB2_2_12/i0_4 ), .A2(\SB2_2_12/i1[9] ), .A3(
        \SB2_2_12/i1_5 ), .ZN(n2015) );
  NAND3_X1 U3729 ( .A1(\SB1_3_29/i1[9] ), .A2(\SB1_3_29/i0_4 ), .A3(
        \SB1_3_29/i1_5 ), .ZN(\SB1_3_29/Component_Function_4/NAND4_in[3] ) );
  NAND4_X1 U3731 ( .A1(\SB2_2_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_3/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_3/Component_Function_4/NAND4_in[1] ), .A4(n2016), .ZN(
        \RI5[2][178] ) );
  NAND3_X1 U3737 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0[10] ), .A3(
        \RI3[2][168] ), .ZN(n2016) );
  NAND3_X1 U3756 ( .A1(\SB2_0_11/i0[9] ), .A2(\SB2_0_11/i0[8] ), .A3(
        \SB2_0_11/i0_0 ), .ZN(\SB2_0_11/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U3761 ( .A1(\SB2_1_31/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_31/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_31/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_1_31/Component_Function_3/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[15] ) );
  NAND3_X1 U3774 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0[10] ), .A3(
        \SB1_0_18/i0[9] ), .ZN(\SB1_0_18/Component_Function_4/NAND4_in[2] ) );
  INV_X2 U3804 ( .A(\RI1[1][11] ), .ZN(\SB1_1_30/i0_3 ) );
  XNOR2_X1 U3810 ( .A(n654), .B(n653), .ZN(\RI1[1][11] ) );
  NAND4_X1 U3811 ( .A1(\SB2_1_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_8/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_8/Component_Function_2/NAND4_in[1] ), .A4(n2017), .ZN(
        \RI5[1][158] ) );
  NAND3_X1 U3816 ( .A1(\SB2_1_8/i0_4 ), .A2(\SB2_1_8/i0_0 ), .A3(
        \SB2_1_8/i1_5 ), .ZN(n2017) );
  NAND4_X1 U3817 ( .A1(\SB1_2_4/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_4/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_4/Component_Function_5/NAND4_in[0] ), .A4(n2018), .ZN(
        \RI3[2][167] ) );
  NAND3_X1 U3818 ( .A1(\SB1_2_4/i1[9] ), .A2(\SB1_2_4/i0_3 ), .A3(
        \SB1_2_4/i0_4 ), .ZN(n2018) );
  NAND3_X1 U3838 ( .A1(\SB1_0_9/i0[6] ), .A2(\SB1_0_9/i1_5 ), .A3(
        \SB1_0_9/i0[9] ), .ZN(\SB1_0_9/Component_Function_1/NAND4_in[2] ) );
  XNOR2_X1 U3839 ( .A(\MC_ARK_ARC_1_0/temp5[125] ), .B(n2019), .ZN(
        \RI1[1][125] ) );
  XNOR2_X1 U3840 ( .A(\MC_ARK_ARC_1_0/temp4[125] ), .B(
        \MC_ARK_ARC_1_0/temp3[125] ), .ZN(n2019) );
  NAND4_X1 U3847 ( .A1(\SB1_0_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_3/NAND4_in[1] ), .A3(n2023), .A4(n2020), 
        .ZN(\RI3[0][21] ) );
  NAND3_X1 U3851 ( .A1(\SB1_0_30/i1_7 ), .A2(\SB1_0_30/i0[10] ), .A3(
        \SB1_0_30/i1[9] ), .ZN(n2020) );
  NAND3_X1 U3852 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0_4 ), .A3(
        \SB1_0_12/i1[9] ), .ZN(\SB1_0_12/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3858 ( .A1(\SB2_3_1/i0_0 ), .A2(\SB2_3_1/i0_4 ), .A3(
        \SB2_3_1/i1_5 ), .ZN(\SB2_3_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3878 ( .A1(\SB1_2_14/i0_0 ), .A2(\SB1_2_14/i0_4 ), .A3(
        \SB1_2_14/i0_3 ), .ZN(\SB1_2_14/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U3879 ( .A1(\SB2_0_17/Component_Function_5/NAND4_in[2] ), .A2(n1290), .A3(\SB2_0_17/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[89] ) );
  NAND3_X1 U3881 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i1_5 ), .A3(
        \SB2_1_10/i1[9] ), .ZN(n2021) );
  NAND4_X1 U3883 ( .A1(\SB2_1_15/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_15/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_15/Component_Function_1/NAND4_in[0] ), .A4(n2022), .ZN(
        \RI5[1][121] ) );
  NAND3_X1 U3884 ( .A1(\SB2_1_15/i0_4 ), .A2(\SB2_1_15/i1_7 ), .A3(
        \SB2_1_15/i0[8] ), .ZN(n2022) );
  NAND3_X1 U3895 ( .A1(\SB1_0_30/i3[0] ), .A2(\SB1_0_30/i1_5 ), .A3(
        \SB1_0_30/i0[8] ), .ZN(n2023) );
  NAND3_X1 U3896 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i3[0] ), .A3(
        \SB2_2_10/i1_7 ), .ZN(\SB2_2_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3901 ( .A1(\SB2_0_7/i0_4 ), .A2(\SB2_0_7/i1_5 ), .A3(
        \SB2_0_7/i0_0 ), .ZN(n909) );
  NAND3_X1 U3902 ( .A1(\SB2_1_27/i0_3 ), .A2(\SB2_1_27/i0_4 ), .A3(
        \SB2_1_27/i0_0 ), .ZN(\SB2_1_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3908 ( .A1(\SB2_0_31/i0[10] ), .A2(\SB2_0_31/i0_3 ), .A3(
        \SB2_0_31/i0[9] ), .ZN(n2024) );
  NAND3_X1 U3910 ( .A1(\SB2_1_17/i0[10] ), .A2(\SB2_1_17/i1[9] ), .A3(
        \SB2_1_17/i1_7 ), .ZN(\SB2_1_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3912 ( .A1(\SB2_0_23/i0[9] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0[8] ), .ZN(\SB2_0_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3917 ( .A1(\SB2_3_1/i0_4 ), .A2(\SB2_3_1/i1[9] ), .A3(
        \SB2_3_1/i1_5 ), .ZN(\SB2_3_1/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U3918 ( .A1(n2217), .A2(n1756), .A3(
        \SB2_0_7/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_7/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[154] ) );
  NAND3_X1 U3950 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i0_3 ), .A3(
        \SB2_1_31/i0_4 ), .ZN(\SB2_1_31/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U3956 ( .A1(\SB2_3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_15/Component_Function_4/NAND4_in[3] ), .A4(n2025), .ZN(
        \RI5[3][106] ) );
  NAND3_X1 U3957 ( .A1(\SB2_3_15/i0[10] ), .A2(\SB2_3_15/i0[9] ), .A3(
        \SB2_3_15/i0_3 ), .ZN(n2025) );
  NAND3_X1 U3982 ( .A1(\SB2_0_26/i0[10] ), .A2(\SB2_0_26/i1_5 ), .A3(
        \SB2_0_26/i1[9] ), .ZN(\SB2_0_26/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U3993 ( .A1(\SB2_2_29/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_29/Component_Function_3/NAND4_in[0] ), .A3(n1109), .A4(
        \SB2_2_29/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[27] ) );
  XNOR2_X1 U3994 ( .A(n2026), .B(n992), .ZN(\RI1[3][14] ) );
  XNOR2_X1 U3995 ( .A(\MC_ARK_ARC_1_2/temp1[14] ), .B(
        \MC_ARK_ARC_1_2/temp2[14] ), .ZN(n2026) );
  NAND4_X2 U3996 ( .A1(\SB2_3_29/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_29/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_29/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_29/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[22] ) );
  NAND4_X2 U4002 ( .A1(\SB2_1_17/Component_Function_3/NAND4_in[0] ), .A2(n915), 
        .A3(\SB2_1_17/Component_Function_3/NAND4_in[2] ), .A4(n1194), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[99] ) );
  NAND3_X1 U4013 ( .A1(\SB1_0_26/i0[9] ), .A2(\SB1_0_26/i0_3 ), .A3(
        \SB1_0_26/i0[10] ), .ZN(\SB1_0_26/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U4028 ( .A1(\SB1_1_23/i1[9] ), .A2(\SB1_1_23/i0_4 ), .A3(
        \SB1_1_23/i1_5 ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[3] ) );
  NAND4_X1 U4033 ( .A1(\SB2_1_22/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_22/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_22/Component_Function_2/NAND4_in[1] ), .A4(n2027), .ZN(
        \RI5[1][74] ) );
  NAND3_X1 U4043 ( .A1(\SB2_1_22/i0_4 ), .A2(\SB2_1_22/i0_0 ), .A3(
        \SB2_1_22/i1_5 ), .ZN(n2027) );
  XNOR2_X1 U4054 ( .A(\MC_ARK_ARC_1_1/temp6[128] ), .B(n2028), .ZN(
        \RI1[2][128] ) );
  XNOR2_X1 U4055 ( .A(\MC_ARK_ARC_1_1/temp2[128] ), .B(
        \MC_ARK_ARC_1_1/temp1[128] ), .ZN(n2028) );
  NAND4_X2 U4063 ( .A1(\SB2_0_25/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_25/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_25/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[56] ) );
  BUF_X2 U4064 ( .A(\RI3[1][138] ), .Z(\SB2_1_8/i0[9] ) );
  XNOR2_X1 U4065 ( .A(n2029), .B(n295), .ZN(Ciphertext[137]) );
  NAND4_X1 U4066 ( .A1(\SB4_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_9/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_9/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_9/Component_Function_5/NAND4_in[0] ), .ZN(n2029) );
  NAND4_X1 U4067 ( .A1(\SB1_3_22/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_22/Component_Function_5/NAND4_in[0] ), .A4(n2030), .ZN(
        \RI3[3][59] ) );
  NAND3_X1 U4071 ( .A1(\SB1_3_22/i1[9] ), .A2(\SB1_3_22/i0_3 ), .A3(
        \SB1_3_22/i0_4 ), .ZN(n2030) );
  NAND4_X2 U4087 ( .A1(\SB3_10/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_10/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_10/Component_Function_4/NAND4_in[1] ), .A4(n1114), .ZN(
        \RI3[4][136] ) );
  NAND3_X1 U4090 ( .A1(\SB3_10/i0[9] ), .A2(\SB3_10/i0_3 ), .A3(
        \SB3_10/i0[10] ), .ZN(n1114) );
  NAND3_X1 U4124 ( .A1(\SB2_2_23/i0_4 ), .A2(\SB2_2_23/i1[9] ), .A3(
        \SB2_2_23/i1_5 ), .ZN(\SB2_2_23/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U4125 ( .A1(\SB2_3_22/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_22/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_22/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[74] ) );
  NAND4_X2 U4126 ( .A1(n682), .A2(\SB1_3_5/Component_Function_4/NAND4_in[1] ), 
        .A3(\SB1_3_5/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_3_5/Component_Function_4/NAND4_in[0] ), .ZN(\SB2_3_4/i0_4 ) );
  NAND3_X1 U4127 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i0_3 ), .A3(
        \SB1_3_10/i0[6] ), .ZN(\SB1_3_10/Component_Function_2/NAND4_in[1] ) );
  XNOR2_X1 U4130 ( .A(n2031), .B(n215), .ZN(Ciphertext[149]) );
  NAND4_X1 U4133 ( .A1(n2034), .A2(\SB4_7/Component_Function_5/NAND4_in[3] ), 
        .A3(n1182), .A4(\SB4_7/Component_Function_5/NAND4_in[0] ), .ZN(n2031)
         );
  NAND4_X1 U4142 ( .A1(\SB2_2_5/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_5/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_5/Component_Function_4/NAND4_in[1] ), .A4(n2032), .ZN(
        \RI5[2][166] ) );
  NAND3_X1 U4143 ( .A1(\SB2_2_5/i0_4 ), .A2(\SB2_2_5/i1_5 ), .A3(
        \SB2_2_5/i1[9] ), .ZN(n2032) );
  NAND4_X1 U4152 ( .A1(\SB1_2_11/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_11/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_11/Component_Function_5/NAND4_in[0] ), .A4(n2033), .ZN(
        \RI3[2][125] ) );
  NAND3_X1 U4159 ( .A1(\SB1_2_11/i1[9] ), .A2(\SB1_2_11/i0_3 ), .A3(
        \SB1_2_11/i0_4 ), .ZN(n2033) );
  NAND3_X1 U4160 ( .A1(\SB4_7/i0_4 ), .A2(n877), .A3(\SB4_7/i1[9] ), .ZN(n2034) );
  XNOR2_X1 U4171 ( .A(\MC_ARK_ARC_1_1/buf_datainput[59] ), .B(n838), .ZN(
        \MC_ARK_ARC_1_1/temp1[59] ) );
  NAND4_X2 U4194 ( .A1(n1307), .A2(\SB2_1_23/Component_Function_5/NAND4_in[3] ), .A3(\SB2_1_23/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_23/Component_Function_5/NAND4_in[0] ), .ZN(n838) );
  NAND3_X1 U4216 ( .A1(\SB2_2_12/i0_0 ), .A2(\SB2_2_12/i1_5 ), .A3(
        \RI3[2][118] ), .ZN(\SB2_2_12/Component_Function_2/NAND4_in[3] ) );
  XNOR2_X1 U4240 ( .A(n2035), .B(n229), .ZN(Ciphertext[147]) );
  NAND4_X1 U4241 ( .A1(\SB4_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_7/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_7/Component_Function_3/NAND4_in[3] ), .ZN(n2035) );
  NAND3_X1 U4242 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[9] ), .A3(
        \SB2_1_24/i0[10] ), .ZN(\SB2_1_24/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U4243 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i1[9] ), .A3(
        \SB2_0_25/i0[6] ), .ZN(\SB2_0_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4246 ( .A1(\SB4_1/i0_4 ), .A2(n857), .A3(\SB4_1/i1[9] ), .ZN(
        \SB4_1/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U4247 ( .A1(\SB2_0_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_26/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_26/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[50] ) );
  NAND4_X1 U4248 ( .A1(\SB3_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_12/Component_Function_5/NAND4_in[0] ), .A4(n2036), .ZN(
        \RI3[4][119] ) );
  NAND3_X1 U4291 ( .A1(\SB3_12/i1[9] ), .A2(\SB3_12/i0_4 ), .A3(\SB3_12/i0_3 ), 
        .ZN(n2036) );
  NAND3_X1 U4292 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0_0 ), .A3(
        \SB2_0_11/i0[7] ), .ZN(\SB2_0_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4308 ( .A1(\SB2_2_2/i0_0 ), .A2(\SB2_2_2/i3[0] ), .A3(
        \SB2_2_2/i1_7 ), .ZN(\SB2_2_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4309 ( .A1(\SB2_3_17/i0[10] ), .A2(\SB2_3_17/i1_5 ), .A3(
        \SB2_3_17/i1[9] ), .ZN(\SB2_3_17/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4323 ( .A1(\SB1_2_5/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_5/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_5/Component_Function_2/NAND4_in[2] ), .A4(n2037), .ZN(
        \RI3[2][176] ) );
  NAND3_X1 U4327 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i0_4 ), .A3(
        \SB1_2_5/i1_5 ), .ZN(n2037) );
  NAND3_X1 U4328 ( .A1(\SB2_0_22/i0_3 ), .A2(\RI3[0][55] ), .A3(
        \SB2_0_22/i1[9] ), .ZN(\SB2_0_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4346 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i1[9] ), .A3(\SB4_22/i0[6] ), .ZN(\SB4_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4350 ( .A1(\SB2_2_4/i0[8] ), .A2(\SB2_2_4/i3[0] ), .A3(
        \SB2_2_4/i1_5 ), .ZN(\SB2_2_4/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U4367 ( .A1(\SB4_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_0/Component_Function_3/NAND4_in[1] ), .A3(n761), .A4(n2038), .ZN(
        n2156) );
  NAND3_X1 U4368 ( .A1(\SB4_0/i1_5 ), .A2(\SB4_0/i3[0] ), .A3(\SB4_0/i0[8] ), 
        .ZN(n2038) );
  NAND4_X1 U4383 ( .A1(\SB3_29/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_5/NAND4_in[0] ), .A4(n2039), .ZN(
        \RI3[4][17] ) );
  NAND3_X1 U4388 ( .A1(\SB3_29/i1[9] ), .A2(\SB3_29/i0_4 ), .A3(\SB3_29/i0_3 ), 
        .ZN(n2039) );
  XNOR2_X1 U4397 ( .A(n2040), .B(n367), .ZN(Ciphertext[181]) );
  NAND4_X1 U4398 ( .A1(n1329), .A2(\SB4_1/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB4_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_1/Component_Function_1/NAND4_in[0] ), .ZN(n2040) );
  NAND4_X1 U4429 ( .A1(\SB2_1_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_19/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_19/Component_Function_1/NAND4_in[2] ), .A4(n2041), .ZN(
        \RI5[1][97] ) );
  NAND3_X1 U4431 ( .A1(\SB2_1_19/i0_4 ), .A2(\SB2_1_19/i1_7 ), .A3(
        \SB2_1_19/i0[8] ), .ZN(n2041) );
  NAND4_X1 U4449 ( .A1(\SB3_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_30/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_30/Component_Function_5/NAND4_in[0] ), .A4(n2042), .ZN(
        \RI3[4][11] ) );
  NAND3_X1 U4459 ( .A1(\SB3_30/i1[9] ), .A2(\SB3_30/i0_3 ), .A3(\SB3_30/i0_4 ), 
        .ZN(n2042) );
  NAND3_X1 U4464 ( .A1(\SB1_3_4/i0[10] ), .A2(\SB1_3_4/i0[9] ), .A3(
        \SB1_3_4/i0_3 ), .ZN(\SB1_3_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4465 ( .A1(n1668), .A2(\SB4_30/i0_4 ), .A3(\SB4_30/i1[9] ), .ZN(
        \SB4_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4476 ( .A1(\SB2_3_3/i0_4 ), .A2(\SB2_3_3/i0[9] ), .A3(
        \RI3[3][169] ), .ZN(\SB2_3_3/Component_Function_5/NAND4_in[3] ) );
  XNOR2_X1 U4501 ( .A(n2044), .B(n2043), .ZN(\RI1[4][130] ) );
  XNOR2_X1 U4523 ( .A(\MC_ARK_ARC_1_3/temp4[130] ), .B(
        \MC_ARK_ARC_1_3/temp2[130] ), .ZN(n2043) );
  XNOR2_X1 U4524 ( .A(\MC_ARK_ARC_1_3/temp3[130] ), .B(
        \MC_ARK_ARC_1_3/temp1[130] ), .ZN(n2044) );
  XNOR2_X1 U4536 ( .A(n2045), .B(n263), .ZN(Ciphertext[128]) );
  NAND4_X1 U4549 ( .A1(\SB4_10/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_10/Component_Function_2/NAND4_in[2] ), .A3(n1542), .A4(n691), 
        .ZN(n2045) );
  NAND4_X2 U4551 ( .A1(n1702), .A2(\SB2_3_3/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_3_3/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[173] ) );
  NAND3_X1 U4567 ( .A1(\SB2_0_23/i0[6] ), .A2(\SB2_0_23/i1[9] ), .A3(
        \SB2_0_23/i0_3 ), .ZN(n2046) );
  NAND3_X1 U4568 ( .A1(\SB1_3_16/i0_4 ), .A2(\SB1_3_16/i0_0 ), .A3(
        \SB1_3_16/i1_5 ), .ZN(\SB1_3_16/Component_Function_2/NAND4_in[3] ) );
  XNOR2_X1 U4569 ( .A(n2047), .B(n286), .ZN(Ciphertext[152]) );
  NAND3_X1 U4570 ( .A1(\SB2_1_25/i0_4 ), .A2(\SB2_1_25/i1_7 ), .A3(
        \SB2_1_25/i0[8] ), .ZN(\SB2_1_25/Component_Function_1/NAND4_in[3] ) );
  XNOR2_X1 U4571 ( .A(\MC_ARK_ARC_1_3/temp6[182] ), .B(n2048), .ZN(
        \RI1[4][182] ) );
  XNOR2_X1 U4572 ( .A(\MC_ARK_ARC_1_3/temp2[182] ), .B(
        \MC_ARK_ARC_1_3/temp1[182] ), .ZN(n2048) );
  NAND3_X1 U4573 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0[7] ), .A3(
        \SB1_0_28/i0_0 ), .ZN(\SB1_0_28/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U4574 ( .A1(\SB4_30/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_2/NAND4_in[1] ), .A3(n661), .A4(n2049), 
        .ZN(n2096) );
  NAND3_X1 U4575 ( .A1(\SB4_30/i0_0 ), .A2(\SB4_30/i0_4 ), .A3(\SB4_30/i1_5 ), 
        .ZN(n2049) );
  NAND4_X1 U4576 ( .A1(n1673), .A2(\SB1_0_23/Component_Function_5/NAND4_in[1] ), .A3(\SB1_0_23/Component_Function_5/NAND4_in[3] ), .A4(n2050), .ZN(
        \RI3[0][53] ) );
  NAND2_X1 U4577 ( .A1(\SB1_0_23/i3[0] ), .A2(\SB1_0_23/i0_0 ), .ZN(n2050) );
  NAND3_X1 U4578 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i0[10] ), .ZN(\SB2_2_31/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U4579 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i1[9] ), .A3(
        \SB1_2_31/i0_4 ), .ZN(n2055) );
  NAND3_X1 U4580 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[7] ), .A3(
        \SB1_0_25/i0_0 ), .ZN(n1267) );
  XNOR2_X1 U4581 ( .A(n2051), .B(n346), .ZN(Ciphertext[88]) );
  NAND4_X1 U4582 ( .A1(\SB4_17/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_17/Component_Function_4/NAND4_in[3] ), .A3(n2232), .A4(n2223), 
        .ZN(n2051) );
  NAND4_X1 U4583 ( .A1(\SB3_17/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_17/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_5/NAND4_in[0] ), .A4(n2052), .ZN(
        \RI3[4][89] ) );
  NAND3_X1 U4584 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i1[9] ), .A3(\SB3_17/i0_4 ), 
        .ZN(n2052) );
  NAND4_X2 U4585 ( .A1(\SB2_0_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_7/Component_Function_2/NAND4_in[2] ), .A3(n909), .A4(
        \SB2_0_7/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[164] ) );
  XNOR2_X1 U4586 ( .A(n2053), .B(n194), .ZN(Ciphertext[15]) );
  NAND4_X1 U4587 ( .A1(\SB4_29/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_29/Component_Function_3/NAND4_in[0] ), .A3(n635), .A4(
        \SB4_29/Component_Function_3/NAND4_in[3] ), .ZN(n2053) );
  XNOR2_X1 U4588 ( .A(n2054), .B(n255), .ZN(Ciphertext[184]) );
  NAND4_X1 U4589 ( .A1(\SB4_1/Component_Function_4/NAND4_in[3] ), .A2(n2178), 
        .A3(\SB4_1/Component_Function_4/NAND4_in[2] ), .A4(n741), .ZN(n2054)
         );
  NAND4_X2 U4590 ( .A1(\SB2_0_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_10/Component_Function_3/NAND4_in[2] ), .A4(n1902), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[141] ) );
  NAND4_X1 U4591 ( .A1(\SB1_2_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_31/Component_Function_5/NAND4_in[0] ), .A4(n2055), .ZN(
        \RI3[2][5] ) );
  NAND3_X1 U4592 ( .A1(\SB2_1_9/i0[9] ), .A2(\SB2_1_9/i0_3 ), .A3(
        \SB2_1_9/i0[10] ), .ZN(\SB2_1_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4593 ( .A1(\SB1_3_21/i1[9] ), .A2(\SB1_3_21/i0_4 ), .A3(
        \SB1_3_21/i1_5 ), .ZN(\SB1_3_21/Component_Function_4/NAND4_in[3] ) );
  NAND4_X1 U4594 ( .A1(\SB3_16/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_5/NAND4_in[0] ), .A4(n2056), .ZN(
        \RI3[4][95] ) );
  NAND3_X1 U4595 ( .A1(\SB3_16/i1[9] ), .A2(\SB3_16/i0_3 ), .A3(\SB3_16/i0_4 ), 
        .ZN(n2056) );
  NAND3_X1 U4596 ( .A1(\SB1_1_9/i0_4 ), .A2(\SB1_1_9/i0[6] ), .A3(
        \SB1_1_9/i0[9] ), .ZN(\SB1_1_9/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U4597 ( .A1(n1754), .A2(\SB2_0_10/Component_Function_2/NAND4_in[1] ), .A3(\SB2_0_10/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_10/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[146] ) );
  NAND4_X4 U4598 ( .A1(n1793), .A2(\SB2_2_28/Component_Function_2/NAND4_in[0] ), .A3(n2064), .A4(\SB2_2_28/Component_Function_2/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[38] ) );
  NAND3_X1 U4599 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i1_5 ), .A3(
        \SB2_1_31/i0_4 ), .ZN(\SB2_1_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4600 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i0[6] ), .A3(
        \SB2_1_31/i0[10] ), .ZN(\SB2_1_31/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U4601 ( .A1(\SB1_3_19/i1[9] ), .A2(\SB1_3_19/i0_4 ), .A3(
        \SB1_3_19/i1_5 ), .ZN(\SB1_3_19/Component_Function_4/NAND4_in[3] ) );
  NAND4_X4 U4602 ( .A1(\SB2_2_23/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_23/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_23/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_23/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[58] ) );
  XNOR2_X1 U4603 ( .A(n1239), .B(n2057), .ZN(\RI1[2][35] ) );
  XNOR2_X1 U4604 ( .A(\MC_ARK_ARC_1_1/temp2[35] ), .B(
        \MC_ARK_ARC_1_1/temp4[35] ), .ZN(n2057) );
  BUF_X2 U4605 ( .A(\RI3[4][85] ), .Z(\SB4_17/i0[6] ) );
  NAND3_X1 U4606 ( .A1(\SB1_3_26/i0[10] ), .A2(\SB1_3_26/i1[9] ), .A3(
        \SB1_3_26/i1_5 ), .ZN(\SB1_3_26/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4607 ( .A1(\SB1_2_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_7/Component_Function_2/NAND4_in[2] ), .A4(n2058), .ZN(
        \RI3[2][164] ) );
  NAND3_X1 U4608 ( .A1(\SB1_2_7/i0_0 ), .A2(\SB1_2_7/i0_4 ), .A3(
        \SB1_2_7/i1_5 ), .ZN(n2058) );
  NAND3_X1 U4609 ( .A1(\SB2_3_4/i0[10] ), .A2(\SB2_3_4/i0_3 ), .A3(n2133), 
        .ZN(\SB2_3_4/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U4610 ( .A(n2059), .B(n218), .ZN(Ciphertext[80]) );
  NAND4_X1 U4611 ( .A1(\SB4_18/Component_Function_2/NAND4_in[2] ), .A2(n1335), 
        .A3(\SB4_18/Component_Function_2/NAND4_in[1] ), .A4(
        \SB4_18/Component_Function_2/NAND4_in[0] ), .ZN(n2059) );
  NAND3_X1 U4612 ( .A1(\SB1_3_15/i0[7] ), .A2(\SB1_3_15/i0_0 ), .A3(n1647), 
        .ZN(\SB1_3_15/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U4613 ( .A1(\SB3_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_18/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_5/NAND4_in[0] ), .A4(n2060), .ZN(
        \RI3[4][83] ) );
  NAND3_X1 U4614 ( .A1(\SB3_18/i0[6] ), .A2(\SB3_18/i0[9] ), .A3(\SB3_18/i0_4 ), .ZN(n2060) );
  XNOR2_X1 U4615 ( .A(\MC_ARK_ARC_1_3/temp6[79] ), .B(n2061), .ZN(\RI1[4][79] ) );
  XNOR2_X1 U4616 ( .A(\MC_ARK_ARC_1_3/temp2[79] ), .B(
        \MC_ARK_ARC_1_3/temp1[79] ), .ZN(n2061) );
  NAND4_X1 U4617 ( .A1(\SB1_3_4/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_4/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_4/Component_Function_5/NAND4_in[0] ), .A4(n2062), .ZN(
        \RI3[3][167] ) );
  NAND3_X1 U4618 ( .A1(\SB1_3_4/i1[9] ), .A2(\SB1_3_4/i0_3 ), .A3(
        \SB1_3_4/i0_4 ), .ZN(n2062) );
  NAND3_X1 U4619 ( .A1(\SB1_2_28/i3[0] ), .A2(\SB1_2_28/i0_0 ), .A3(
        \SB1_2_28/i1_7 ), .ZN(\SB1_2_28/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U4620 ( .A1(\SB2_3_2/i1[9] ), .A2(\SB2_3_2/i0_3 ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 U4621 ( .A1(\SB2_3_5/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_5/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_5/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_5/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[166] ) );
  NAND4_X1 U4622 ( .A1(\SB2_3_2/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_2/NAND4_in[0] ), .A4(n2063), .ZN(
        \RI5[3][2] ) );
  NAND3_X1 U4623 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i1_5 ), .A3(
        \SB2_3_2/i0_4 ), .ZN(n2063) );
  XNOR2_X1 U4624 ( .A(n2065), .B(n339), .ZN(Ciphertext[144]) );
  NAND4_X1 U4625 ( .A1(\SB4_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_7/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_7/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_7/Component_Function_0/NAND4_in[0] ), .ZN(n2065) );
  NAND3_X1 U4626 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0[10] ), .A3(
        \SB1_0_28/i0_4 ), .ZN(\SB1_0_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4627 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0_4 ), .A3(
        \SB2_1_15/i0_0 ), .ZN(\SB2_1_15/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U4628 ( .A1(n1576), .A2(\SB1_0_18/Component_Function_4/NAND4_in[2] ), .A3(\SB1_0_18/Component_Function_4/NAND4_in[1] ), .A4(n2066), .ZN(
        \RI3[0][88] ) );
  NAND3_X1 U4629 ( .A1(\SB1_0_18/i0[8] ), .A2(\SB1_0_18/i0[9] ), .A3(
        \SB1_0_18/i0_0 ), .ZN(n2066) );
  NAND3_X1 U4630 ( .A1(\SB3_10/i3[0] ), .A2(\SB3_10/i1_5 ), .A3(\SB3_10/i0[8] ), .ZN(\SB3_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4631 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i0_3 ), .A3(
        \SB1_2_10/i0_4 ), .ZN(\SB1_2_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4632 ( .A1(\SB2_3_26/i0[7] ), .A2(\SB2_3_26/i0[8] ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U4633 ( .A1(\SB3_6/i0[8] ), .A2(\SB3_6/i0[9] ), .A3(\SB3_6/i0_3 ), 
        .ZN(\SB3_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4634 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i0_0 ), .A3(
        \SB1_3_17/i0[6] ), .ZN(\SB1_3_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4635 ( .A1(\SB2_3_29/i0_3 ), .A2(\SB2_3_29/i0_4 ), .A3(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4636 ( .A1(\SB2_0_10/i0_3 ), .A2(\SB2_0_10/i0_0 ), .A3(
        \SB2_0_10/i0_4 ), .ZN(\SB2_0_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4637 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i1[9] ), .A3(
        \SB2_3_21/i0[6] ), .ZN(\SB2_3_21/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U4638 ( .A1(\SB4_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_8/Component_Function_3/NAND4_in[3] ), .A4(n2067), .ZN(
        \RI4[4][141] ) );
  NAND3_X1 U4639 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i1[9] ), .A3(\SB4_8/i1_7 ), 
        .ZN(n2067) );
  NAND3_X1 U4640 ( .A1(\SB2_0_22/i0[10] ), .A2(\SB2_0_22/i1[9] ), .A3(
        \SB2_0_22/i1_7 ), .ZN(\SB2_0_22/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U4641 ( .A1(\SB1_1_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_21/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_5/NAND4_in[0] ), .A4(n2068), .ZN(
        \RI3[1][65] ) );
  NAND3_X1 U4642 ( .A1(\SB1_1_21/i0[9] ), .A2(\SB1_1_21/i0_4 ), .A3(
        \SB1_1_21/i0[6] ), .ZN(n2068) );
  NAND4_X2 U4643 ( .A1(n1026), .A2(\SB2_1_29/Component_Function_3/NAND4_in[0] ), .A3(n1252), .A4(\SB2_1_29/Component_Function_3/NAND4_in[2] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[27] ) );
  NAND4_X2 U4644 ( .A1(\SB2_2_10/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_10/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[131] ) );
  NAND4_X2 U4645 ( .A1(\SB2_2_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_8/Component_Function_3/NAND4_in[0] ), .A3(n2069), .A4(n1169), 
        .ZN(\MC_ARK_ARC_1_2/buf_datainput[153] ) );
  NAND3_X1 U4646 ( .A1(\SB2_2_8/i0[10] ), .A2(\SB2_2_8/i1_7 ), .A3(
        \SB2_2_8/i1[9] ), .ZN(n2069) );
  NAND4_X1 U4647 ( .A1(\SB2_1_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_30/Component_Function_4/NAND4_in[1] ), .A4(n2070), .ZN(
        \RI5[1][16] ) );
  XNOR2_X1 U4648 ( .A(n2071), .B(n281), .ZN(Ciphertext[98]) );
  NAND4_X1 U4649 ( .A1(\SB4_15/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_15/Component_Function_2/NAND4_in[2] ), .A3(n1312), .A4(
        \SB4_15/Component_Function_2/NAND4_in[0] ), .ZN(n2071) );
  XNOR2_X1 U4650 ( .A(n2073), .B(n2072), .ZN(\RI1[2][104] ) );
  XNOR2_X1 U4651 ( .A(\MC_ARK_ARC_1_1/temp1[104] ), .B(
        \MC_ARK_ARC_1_1/temp4[104] ), .ZN(n2072) );
  XNOR2_X1 U4652 ( .A(\MC_ARK_ARC_1_1/temp3[104] ), .B(
        \MC_ARK_ARC_1_1/temp2[104] ), .ZN(n2073) );
  NAND4_X1 U4653 ( .A1(\SB2_1_28/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_28/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_28/Component_Function_2/NAND4_in[3] ), .A4(n2074), .ZN(
        \RI5[1][38] ) );
  NAND3_X1 U4654 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0[9] ), .A3(
        \SB2_1_28/i0[8] ), .ZN(n2074) );
  XNOR2_X1 U4655 ( .A(n2075), .B(n1732), .ZN(\RI1[1][41] ) );
  XNOR2_X1 U4656 ( .A(\MC_ARK_ARC_1_0/temp4[41] ), .B(
        \MC_ARK_ARC_1_0/temp1[41] ), .ZN(n2075) );
  NAND4_X2 U4657 ( .A1(\SB2_3_14/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_14/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_14/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_14/Component_Function_4/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[112] ) );
  XNOR2_X1 U4658 ( .A(n2076), .B(n283), .ZN(Ciphertext[29]) );
  NAND4_X1 U4659 ( .A1(\SB4_27/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_27/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_27/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_27/Component_Function_5/NAND4_in[0] ), .ZN(n2076) );
  NAND4_X1 U4660 ( .A1(\SB4_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_26/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_26/Component_Function_3/NAND4_in[3] ), .A4(n2077), .ZN(
        \RI4[4][33] ) );
  NAND3_X1 U4661 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i1[9] ), .A3(
        \SB4_26/i1_7 ), .ZN(n2077) );
  XNOR2_X1 U4662 ( .A(n2078), .B(n270), .ZN(Ciphertext[31]) );
  NAND4_X1 U4663 ( .A1(\SB4_26/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_26/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_26/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_26/Component_Function_1/NAND4_in[2] ), .ZN(n2078) );
  NAND3_X1 U4664 ( .A1(\SB1_1_11/i0[7] ), .A2(\SB1_1_11/i0_0 ), .A3(
        \SB1_1_11/i0_3 ), .ZN(\SB1_1_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4665 ( .A1(\SB2_3_19/i0_0 ), .A2(\SB2_3_19/i3[0] ), .A3(
        \SB2_3_19/i1_7 ), .ZN(\SB2_3_19/Component_Function_4/NAND4_in[1] ) );
  XNOR2_X1 U4666 ( .A(n2079), .B(n333), .ZN(Ciphertext[49]) );
  NAND4_X1 U4667 ( .A1(\SB4_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_23/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_23/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_23/Component_Function_1/NAND4_in[0] ), .ZN(n2079) );
  NAND4_X1 U4668 ( .A1(\SB2_1_20/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_20/Component_Function_0/NAND4_in[0] ), .A4(n2080), .ZN(
        \RI5[1][96] ) );
  NAND3_X1 U4669 ( .A1(\SB2_1_20/i0_3 ), .A2(\SB2_1_20/i0[7] ), .A3(
        \SB2_1_20/i0_0 ), .ZN(n2080) );
  NAND3_X1 U4670 ( .A1(\SB2_3_28/i0[10] ), .A2(\SB2_3_28/i1[9] ), .A3(
        \SB2_3_28/i1_5 ), .ZN(\SB2_3_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4671 ( .A1(\SB2_0_16/i0_4 ), .A2(\SB2_0_16/i1_5 ), .A3(
        \SB2_0_16/i0_0 ), .ZN(\SB2_0_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4672 ( .A1(\SB2_1_27/i0[9] ), .A2(\SB2_1_27/i0_3 ), .A3(
        \SB2_1_27/i0[8] ), .ZN(\SB2_1_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4673 ( .A1(\SB2_0_20/i0[9] ), .A2(\SB2_0_20/i0[10] ), .A3(
        \SB2_0_20/i0_3 ), .ZN(\SB2_0_20/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U4674 ( .A(n2081), .B(n242), .ZN(Ciphertext[145]) );
  NAND4_X1 U4675 ( .A1(n1101), .A2(\SB4_7/Component_Function_1/NAND4_in[1] ), 
        .A3(n1527), .A4(\SB4_7/Component_Function_1/NAND4_in[0] ), .ZN(n2081)
         );
  NAND3_X1 U4676 ( .A1(\SB1_3_31/i1[9] ), .A2(\SB1_3_31/i0[10] ), .A3(
        \SB1_3_31/i1_7 ), .ZN(\SB1_3_31/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U4677 ( .A1(\SB2_1_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_3/NAND4_in[2] ), .A4(n2082), .ZN(
        \RI5[1][51] ) );
  NAND3_X1 U4678 ( .A1(\SB2_1_25/i1_5 ), .A2(\SB2_1_25/i3[0] ), .A3(
        \SB2_1_25/i0[8] ), .ZN(n2082) );
  NAND4_X1 U4679 ( .A1(\SB1_3_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_4/NAND4_in[3] ), .A4(n2083), .ZN(
        \RI3[3][118] ) );
  NAND3_X1 U4680 ( .A1(\SB1_3_13/i0[10] ), .A2(\SB1_3_13/i0_3 ), .A3(
        \SB1_3_13/i0[9] ), .ZN(n2083) );
  NAND4_X1 U4681 ( .A1(\SB3_5/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_5/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_5/Component_Function_3/NAND4_in[2] ), .A4(n2084), .ZN(
        \RI3[4][171] ) );
  NAND3_X1 U4682 ( .A1(\SB3_5/i3[0] ), .A2(\SB3_5/i1_5 ), .A3(\SB3_5/i0[8] ), 
        .ZN(n2084) );
  XNOR2_X1 U4683 ( .A(n2085), .B(n257), .ZN(Ciphertext[74]) );
  NAND4_X1 U4684 ( .A1(\SB4_19/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_19/Component_Function_2/NAND4_in[2] ), .A3(n1614), .A4(
        \SB4_19/Component_Function_2/NAND4_in[0] ), .ZN(n2085) );
  NAND4_X1 U4685 ( .A1(\SB3_7/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_7/Component_Function_5/NAND4_in[0] ), .A4(n2086), .ZN(
        \RI3[4][149] ) );
  NAND3_X1 U4686 ( .A1(\SB3_7/i1[9] ), .A2(\SB3_7/i0_4 ), .A3(\SB3_7/i0_3 ), 
        .ZN(n2086) );
  NAND4_X1 U4687 ( .A1(\SB3_20/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_20/Component_Function_3/NAND4_in[2] ), .A3(
        \SB3_20/Component_Function_3/NAND4_in[0] ), .A4(n2087), .ZN(
        \RI3[4][81] ) );
  NAND3_X1 U4688 ( .A1(\SB3_20/i3[0] ), .A2(\SB3_20/i1_5 ), .A3(\SB3_20/i0[8] ), .ZN(n2087) );
  NAND4_X1 U4689 ( .A1(\SB3_12/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_12/Component_Function_2/NAND4_in[0] ), .A4(n2088), .ZN(
        \RI3[4][134] ) );
  NAND3_X1 U4690 ( .A1(\SB3_12/i0[9] ), .A2(\SB3_12/i0_3 ), .A3(\SB3_12/i0[8] ), .ZN(n2088) );
  NAND4_X1 U4691 ( .A1(\SB1_3_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_27/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_3_27/Component_Function_0/NAND4_in[1] ), .A4(n2089), .ZN(
        \RI3[3][54] ) );
  NAND3_X1 U4692 ( .A1(\SB1_3_27/i0[7] ), .A2(\SB1_3_27/i0_0 ), .A3(
        \SB1_3_27/i0_3 ), .ZN(n2089) );
  XNOR2_X1 U4693 ( .A(n2091), .B(n2090), .ZN(\RI1[1][44] ) );
  XNOR2_X1 U4694 ( .A(\MC_ARK_ARC_1_0/temp4[44] ), .B(
        \MC_ARK_ARC_1_0/temp1[44] ), .ZN(n2090) );
  XNOR2_X1 U4695 ( .A(\MC_ARK_ARC_1_0/temp2[44] ), .B(
        \MC_ARK_ARC_1_0/temp3[44] ), .ZN(n2091) );
  NAND4_X1 U4696 ( .A1(\SB2_0_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_23/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_23/Component_Function_4/NAND4_in[1] ), .A4(n2092), .ZN(
        \RI5[0][58] ) );
  NAND3_X1 U4697 ( .A1(\SB2_0_23/i0[9] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0[10] ), .ZN(n2092) );
  NAND3_X1 U4698 ( .A1(\SB2_1_13/i0[10] ), .A2(\SB2_1_13/i1[9] ), .A3(
        \SB2_1_13/i1_7 ), .ZN(\SB2_1_13/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U4699 ( .A1(\SB1_2_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_12/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_12/Component_Function_5/NAND4_in[0] ), .A4(n2093), .ZN(
        \RI3[2][119] ) );
  NAND3_X1 U4700 ( .A1(\SB1_2_12/i0[6] ), .A2(\SB1_2_12/i0[9] ), .A3(
        \SB1_2_12/i0_4 ), .ZN(n2093) );
  NAND4_X1 U4701 ( .A1(\SB2_2_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_22/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_22/Component_Function_4/NAND4_in[1] ), .A4(n2094), .ZN(
        \RI5[2][64] ) );
  NAND3_X1 U4702 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[10] ), .A3(
        \SB2_2_22/i0[9] ), .ZN(n2094) );
  INV_X1 U4703 ( .A(\RI3[0][53] ), .ZN(\SB2_0_23/i1_5 ) );
  NAND3_X1 U4704 ( .A1(\SB2_1_19/i0_0 ), .A2(\SB2_1_19/i3[0] ), .A3(
        \SB2_1_19/i1_7 ), .ZN(\SB2_1_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4705 ( .A1(\SB1_3_26/i1[9] ), .A2(\SB1_3_26/i0[10] ), .A3(
        \SB1_3_26/i1_7 ), .ZN(\SB1_3_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4706 ( .A1(\SB2_3_24/i0[10] ), .A2(\SB2_3_24/i1_5 ), .A3(
        \SB2_3_24/i1[9] ), .ZN(\SB2_3_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4707 ( .A1(\SB2_2_26/i0[10] ), .A2(\SB2_2_26/i1_5 ), .A3(
        \SB2_2_26/i1[9] ), .ZN(\SB2_2_26/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4708 ( .A1(\SB2_2_15/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_15/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_15/Component_Function_2/NAND4_in[1] ), .A4(n2095), .ZN(
        \RI5[2][116] ) );
  NAND3_X1 U4709 ( .A1(\SB2_2_15/i0_4 ), .A2(\SB2_2_15/i0_0 ), .A3(
        \SB2_2_15/i1_5 ), .ZN(n2095) );
  XNOR2_X1 U4710 ( .A(n2096), .B(n332), .ZN(Ciphertext[8]) );
  NAND3_X1 U4711 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0[7] ), .A3(
        \SB1_1_6/i0_0 ), .ZN(\SB1_1_6/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U4712 ( .A1(n1268), .A2(\SB2_1_1/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB2_1_1/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_1/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[8] ) );
  NAND3_X1 U4713 ( .A1(\SB2_1_16/i0[10] ), .A2(\SB2_1_16/i1[9] ), .A3(
        \SB2_1_16/i1_7 ), .ZN(\SB2_1_16/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X1 U4714 ( .A(Key[11]), .Z(n398) );
  NAND4_X1 U4715 ( .A1(\SB1_3_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_19/Component_Function_1/NAND4_in[3] ), .ZN(n2097) );
  NAND4_X1 U4716 ( .A1(\SB2_2_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_11/Component_Function_3/NAND4_in[2] ), .A4(n1048), .ZN(n2098)
         );
  NAND4_X1 U4717 ( .A1(\SB2_2_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_11/Component_Function_3/NAND4_in[2] ), .A4(n1048), .ZN(n2099)
         );
  NAND4_X1 U4718 ( .A1(\SB2_2_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_11/Component_Function_3/NAND4_in[2] ), .A4(n1048), .ZN(
        \RI5[2][135] ) );
  BUF_X1 U4719 ( .A(\RI1[4][2] ), .Z(\SB3_31/i1[9] ) );
  NAND4_X1 U4720 ( .A1(\SB3_23/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_23/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_23/Component_Function_5/NAND4_in[0] ), .A4(n980), .ZN(n2100) );
  BUF_X1 U4721 ( .A(\RI1[4][104] ), .Z(\SB3_14/i1[9] ) );
  NAND4_X1 U4722 ( .A1(n1584), .A2(\SB2_2_23/Component_Function_3/NAND4_in[1] ), .A3(\SB2_2_23/Component_Function_3/NAND4_in[2] ), .A4(n1014), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[63] ) );
  BUF_X1 U4723 ( .A(\RI1[4][110] ), .Z(\SB3_13/i1[9] ) );
  INV_X1 U4724 ( .A(\RI1[4][119] ), .ZN(\SB3_12/i0_3 ) );
  NAND4_X1 U4725 ( .A1(\SB2_3_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_23/Component_Function_4/NAND4_in[3] ), .ZN(n2102) );
  NAND4_X1 U4726 ( .A1(\SB2_3_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_23/Component_Function_4/NAND4_in[3] ), .ZN(n2103) );
  NAND4_X1 U4727 ( .A1(\SB2_3_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_23/Component_Function_4/NAND4_in[3] ), .ZN(\RI5[3][58] ) );
  NAND4_X1 U4728 ( .A1(\SB2_1_30/Component_Function_5/NAND4_in[2] ), .A2(n561), 
        .A3(\SB2_1_30/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_30/Component_Function_5/NAND4_in[0] ), .ZN(n2104) );
  NAND4_X1 U4729 ( .A1(\SB3_31/Component_Function_5/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_5/NAND4_in[3] ), .ZN(n2106) );
  NAND4_X1 U4730 ( .A1(\SB1_3_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_0/NAND4_in[3] ), .ZN(n2107) );
  NAND4_X1 U4731 ( .A1(n1322), .A2(\SB2_3_14/Component_Function_5/NAND4_in[1] ), .A3(\SB2_3_14/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_14/Component_Function_5/NAND4_in[0] ), .ZN(n2108) );
  NAND4_X1 U4732 ( .A1(n1322), .A2(\SB2_3_14/Component_Function_5/NAND4_in[1] ), .A3(\SB2_3_14/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_14/Component_Function_5/NAND4_in[0] ), .ZN(n2109) );
  NAND4_X1 U4733 ( .A1(n1322), .A2(\SB2_3_14/Component_Function_5/NAND4_in[1] ), .A3(\SB2_3_14/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_14/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[107] ) );
  NAND4_X1 U4734 ( .A1(\SB1_3_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_0/NAND4_in[3] ), .ZN(n2110) );
  NAND4_X2 U4735 ( .A1(\SB2_3_25/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_3_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_25/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_3_25/Component_Function_5/NAND4_in[3] ), .ZN(n2111) );
  INV_X1 U4736 ( .A(\RI1[4][113] ), .ZN(\SB3_13/i0_3 ) );
  CLKBUF_X1 U4737 ( .A(\RI1[1][46] ), .Z(\SB1_1_24/i0[7] ) );
  NAND4_X1 U4738 ( .A1(\SB2_3_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_21/Component_Function_5/NAND4_in[0] ), .ZN(n2112) );
  NAND4_X1 U4739 ( .A1(\SB2_3_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[65] ) );
  BUF_X1 U4740 ( .A(\RI3[4][125] ), .Z(n841) );
  NAND4_X1 U4741 ( .A1(\SB1_3_21/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_3_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_21/Component_Function_0/NAND4_in[0] ), .A4(n574), .ZN(n2114) );
  NAND4_X1 U4742 ( .A1(\SB1_3_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_1/Component_Function_1/NAND4_in[3] ), .ZN(n2115) );
  BUF_X1 U4743 ( .A(\RI1[4][38] ), .Z(\SB3_25/i1[9] ) );
  NAND4_X1 U4744 ( .A1(n1444), .A2(\SB2_0_6/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_6/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_6/Component_Function_5/NAND4_in[0] ), .ZN(n2116) );
  NAND4_X1 U4745 ( .A1(n1444), .A2(\SB2_0_6/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_6/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_6/Component_Function_5/NAND4_in[0] ), .ZN(n2117) );
  NAND4_X1 U4746 ( .A1(n1444), .A2(\SB2_0_6/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_0_6/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[155] ) );
  BUF_X1 U4747 ( .A(\RI1[1][147] ), .Z(\SB1_1_7/i0[8] ) );
  BUF_X1 U4748 ( .A(\RI5[3][158] ), .Z(n2119) );
  NAND4_X1 U4749 ( .A1(\SB2_3_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_6/Component_Function_5/NAND4_in[0] ), .ZN(n2120) );
  NAND4_X1 U4750 ( .A1(\SB2_3_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_6/Component_Function_5/NAND4_in[0] ), .ZN(n2121) );
  NAND4_X1 U4751 ( .A1(\SB2_3_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[155] ) );
  NAND4_X1 U4752 ( .A1(n633), .A2(\SB2_2_17/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB2_2_17/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_2_17/Component_Function_2/NAND4_in[3] ), .ZN(n2122) );
  NAND4_X1 U4753 ( .A1(n633), .A2(\SB2_2_17/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB2_2_17/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_2_17/Component_Function_2/NAND4_in[3] ), .ZN(n2123) );
  NAND4_X1 U4754 ( .A1(n633), .A2(\SB2_2_17/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB2_2_17/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_2_17/Component_Function_2/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[104] ) );
  NAND4_X2 U4755 ( .A1(\SB2_3_6/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_6/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_6/Component_Function_2/NAND4_in[1] ), .A4(n592), .ZN(
        \RI5[3][170] ) );
  NAND4_X1 U4756 ( .A1(\SB2_1_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_15/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_15/Component_Function_5/NAND4_in[0] ), .ZN(n2124) );
  NAND4_X1 U4757 ( .A1(\SB2_1_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_15/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_15/Component_Function_5/NAND4_in[0] ), .ZN(n2125) );
  NAND4_X1 U4758 ( .A1(\SB2_1_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_15/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_15/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[101] ) );
  BUF_X1 U4759 ( .A(\RI1[4][32] ), .Z(\SB3_26/i1[9] ) );
  NAND4_X4 U4760 ( .A1(\SB2_3_21/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_21/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_3_21/Component_Function_2/NAND4_in[3] ), .ZN(\RI5[3][80] ) );
  NAND4_X4 U4761 ( .A1(\SB2_3_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_19/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[77] ) );
  NAND4_X1 U4762 ( .A1(\SB2_2_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_15/Component_Function_5/NAND4_in[3] ), .ZN(n2126) );
  NAND4_X1 U4763 ( .A1(\SB2_2_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_15/Component_Function_5/NAND4_in[3] ), .ZN(n2127) );
  NAND4_X1 U4764 ( .A1(\SB2_3_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_26/Component_Function_2/NAND4_in[0] ), .ZN(n2128) );
  NAND4_X1 U4765 ( .A1(\SB2_3_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_26/Component_Function_2/NAND4_in[0] ), .ZN(n2129) );
  NAND4_X1 U4766 ( .A1(\SB2_2_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_15/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[101] ) );
  NAND4_X1 U4767 ( .A1(\SB2_3_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_26/Component_Function_2/NAND4_in[0] ), .ZN(\RI5[3][50] ) );
  NAND4_X1 U4768 ( .A1(\SB2_3_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_0/NAND4_in[3] ), .ZN(n2130) );
  NAND4_X1 U4769 ( .A1(\SB2_3_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_0/NAND4_in[3] ), .ZN(\RI5[3][84] ) );
  NAND4_X2 U4770 ( .A1(\SB3_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_30/Component_Function_4/NAND4_in[3] ), .A3(
        \SB3_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_30/Component_Function_4/NAND4_in[1] ), .ZN(n2131) );
  NAND4_X1 U4771 ( .A1(\SB1_0_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_0/NAND4_in[3] ), .ZN(n2132) );
  NAND4_X1 U4772 ( .A1(\SB1_3_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_9/Component_Function_0/NAND4_in[3] ), .ZN(n2133) );
  AND4_X1 U4773 ( .A1(\SB1_3_17/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_17/Component_Function_4/NAND4_in[0] ), .A3(n734), .A4(
        \SB1_3_17/Component_Function_4/NAND4_in[3] ), .ZN(n2134) );
  BUF_X1 U4774 ( .A(\RI3[4][47] ), .Z(n2135) );
  BUF_X1 U4775 ( .A(\RI3[4][47] ), .Z(\SB4_24/i0_3 ) );
  INV_X1 U4776 ( .A(n37), .ZN(n2136) );
  INV_X1 U4777 ( .A(n37), .ZN(\SB1_0_6/i0_3 ) );
  NAND4_X1 U4778 ( .A1(\SB2_0_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_8/Component_Function_2/NAND4_in[0] ), .ZN(n2137) );
  NAND4_X1 U4779 ( .A1(\SB2_0_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_8/Component_Function_2/NAND4_in[0] ), .ZN(n2138) );
  NAND4_X1 U4780 ( .A1(\SB2_0_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_8/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[158] ) );
  NAND4_X1 U4781 ( .A1(\SB2_2_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_9/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_9/Component_Function_3/NAND4_in[3] ), .ZN(n2139) );
  NAND4_X1 U4782 ( .A1(\SB2_2_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_9/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_9/Component_Function_3/NAND4_in[3] ), .ZN(n2140) );
  NAND4_X1 U4783 ( .A1(\SB2_2_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_9/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_9/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[2][147] ) );
  NAND4_X4 U4784 ( .A1(\SB2_2_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_2/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_2/Component_Function_3/NAND4_in[2] ), .A4(n1260), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[189] ) );
  INV_X1 U4785 ( .A(\RI1[1][125] ), .ZN(n2141) );
  INV_X1 U4786 ( .A(\RI1[1][125] ), .ZN(\SB1_1_11/i0_3 ) );
  CLKBUF_X1 U4787 ( .A(Key[71]), .Z(n397) );
  NAND4_X1 U4788 ( .A1(\SB1_3_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_1/NAND4_in[3] ), .ZN(n2143) );
  NAND4_X2 U4789 ( .A1(n1161), .A2(\SB2_2_6/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB2_2_6/Component_Function_2/NAND4_in[1] ), .A4(n1838), .ZN(n2144) );
  NAND4_X2 U4790 ( .A1(n1272), .A2(\SB2_3_9/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB2_3_9/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[137] ) );
  INV_X1 U4791 ( .A(\RI1[1][154] ), .ZN(\SB1_1_6/i0_4 ) );
  NAND4_X1 U4792 ( .A1(n1242), .A2(\SB2_3_16/Component_Function_5/NAND4_in[3] ), .A3(\SB2_3_16/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[95] ) );
  NAND4_X2 U4793 ( .A1(\SB2_2_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_3/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_3/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_3/Component_Function_5/NAND4_in[0] ), .ZN(n827) );
  INV_X1 U4794 ( .A(\RI1[1][124] ), .ZN(\SB1_1_11/i0_4 ) );
  NAND4_X1 U4795 ( .A1(\SB2_0_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_30/Component_Function_5/NAND4_in[1] ), .A3(n950), .A4(n1467), 
        .ZN(n2146) );
  NAND4_X1 U4796 ( .A1(\SB2_0_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_30/Component_Function_5/NAND4_in[1] ), .A3(n950), .A4(n1467), 
        .ZN(n2147) );
  NAND4_X1 U4797 ( .A1(\SB2_0_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_30/Component_Function_5/NAND4_in[1] ), .A3(n950), .A4(n1467), 
        .ZN(\MC_ARK_ARC_1_0/buf_datainput[11] ) );
  BUF_X1 U4798 ( .A(\RI3[4][113] ), .Z(n2148) );
  BUF_X1 U4799 ( .A(\RI3[4][113] ), .Z(\SB4_13/i0_3 ) );
  INV_X1 U4800 ( .A(\RI1[1][167] ), .ZN(n2149) );
  INV_X1 U4801 ( .A(\RI1[1][167] ), .ZN(\SB1_1_4/i0_3 ) );
  NAND4_X1 U4802 ( .A1(\SB2_0_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_3/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_3/Component_Function_5/NAND4_in[3] ), .ZN(n2150) );
  NAND4_X1 U4803 ( .A1(\SB2_0_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_3/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_3/Component_Function_5/NAND4_in[3] ), .ZN(n2151) );
  NAND4_X1 U4804 ( .A1(\SB2_1_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_6/Component_Function_5/NAND4_in[0] ), .ZN(n2152) );
  NAND4_X1 U4805 ( .A1(\SB2_1_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_6/Component_Function_5/NAND4_in[0] ), .ZN(n2153) );
  NAND4_X1 U4806 ( .A1(\SB2_0_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_3/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_3/Component_Function_5/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[173] ) );
  NAND4_X1 U4807 ( .A1(\SB2_1_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[155] ) );
  NAND4_X1 U4808 ( .A1(\SB4_30/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_30/Component_Function_0/NAND4_in[0] ), .A4(n2154), .ZN(n615) );
  NAND3_X1 U4809 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0[7] ), .A3(
        \SB4_30/i0[8] ), .ZN(n2154) );
  XNOR2_X1 U4810 ( .A(n2155), .B(n230), .ZN(Ciphertext[188]) );
  NAND4_X1 U4811 ( .A1(\SB4_0/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_0/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_0/Component_Function_2/NAND4_in[0] ), .A4(
        \SB4_0/Component_Function_2/NAND4_in[3] ), .ZN(n2155) );
  XNOR2_X1 U4812 ( .A(n2156), .B(n314), .ZN(Ciphertext[189]) );
  NAND4_X1 U4813 ( .A1(\SB2_1_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_11/Component_Function_2/NAND4_in[1] ), .A4(n2157), .ZN(
        \RI5[1][140] ) );
  NAND3_X1 U4814 ( .A1(\SB2_1_11/i0_4 ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB2_1_11/i0_0 ), .ZN(n2157) );
  NAND4_X1 U4815 ( .A1(\SB2_0_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_1/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_1/Component_Function_4/NAND4_in[1] ), .A4(n2158), .ZN(
        \RI5[0][190] ) );
  NAND3_X1 U4816 ( .A1(\SB2_0_1/i0_4 ), .A2(\SB2_0_1/i1[9] ), .A3(
        \SB2_0_1/i1_5 ), .ZN(n2158) );
  INV_X1 U4817 ( .A(\RI3[0][110] ), .ZN(\SB2_0_13/i1[9] ) );
  NAND4_X1 U4818 ( .A1(\SB1_0_16/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_16/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_0_16/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][110] ) );
  XNOR2_X1 U4819 ( .A(n2159), .B(n259), .ZN(Ciphertext[156]) );
  NAND4_X1 U4820 ( .A1(\SB4_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_5/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_5/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_5/Component_Function_0/NAND4_in[1] ), .ZN(n2159) );
  NAND4_X2 U4821 ( .A1(n2228), .A2(\SB2_1_19/Component_Function_4/NAND4_in[3] ), .A3(\SB2_1_19/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_19/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[82] ) );
  NAND3_X1 U4822 ( .A1(\SB1_3_23/i1[9] ), .A2(\SB1_3_23/i0[10] ), .A3(
        \SB1_3_23/i1_7 ), .ZN(\SB1_3_23/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U4823 ( .A1(\SB2_3_21/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_21/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_21/Component_Function_3/NAND4_in[2] ), .A4(n2160), .ZN(
        \RI5[3][75] ) );
  NAND3_X1 U4824 ( .A1(\SB2_3_21/i3[0] ), .A2(\SB2_3_21/i1_5 ), .A3(
        \SB2_3_21/i0[8] ), .ZN(n2160) );
  NAND3_X1 U4825 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i1[9] ), .A3(
        \SB2_1_10/i1_7 ), .ZN(\SB2_1_10/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U4826 ( .A1(\SB3_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_11/Component_Function_3/NAND4_in[2] ), .A3(
        \SB3_11/Component_Function_3/NAND4_in[0] ), .A4(n2161), .ZN(
        \RI3[4][135] ) );
  NAND3_X1 U4827 ( .A1(\SB3_11/i3[0] ), .A2(\SB3_11/i1_5 ), .A3(\SB3_11/i0[8] ), .ZN(n2161) );
  NAND4_X1 U4828 ( .A1(\SB1_1_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_2/NAND4_in[2] ), .A4(n2162), .ZN(
        \RI3[1][164] ) );
  NAND3_X1 U4829 ( .A1(\SB1_1_7/i0_0 ), .A2(\SB1_1_7/i1_5 ), .A3(
        \SB1_1_7/i0_4 ), .ZN(n2162) );
  NAND3_X1 U4830 ( .A1(\SB1_1_8/i0_0 ), .A2(\SB1_1_8/i0_4 ), .A3(
        \SB1_1_8/i1_5 ), .ZN(\SB1_1_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4831 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0_0 ), .A3(
        \SB2_3_17/i0[7] ), .ZN(\SB2_3_17/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U4832 ( .A1(\SB1_0_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_8/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_0_8/Component_Function_2/NAND4_in[1] ), .A4(n2163), .ZN(
        \RI3[0][158] ) );
  NAND3_X1 U4833 ( .A1(\SB1_0_8/i1_5 ), .A2(\SB1_0_8/i0_4 ), .A3(
        \SB1_0_8/i0_0 ), .ZN(n2163) );
  NAND3_X1 U4834 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i0[6] ), .A3(
        \SB2_1_31/i0[10] ), .ZN(\SB2_1_31/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X1 U4835 ( .A1(\SB2_1_17/i0[8] ), .A2(\SB2_1_17/i3[0] ), .A3(
        \SB2_1_17/i1_5 ), .ZN(n1194) );
  NAND4_X2 U4836 ( .A1(\SB2_0_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_24/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_24/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[57] ) );
  NAND4_X2 U4837 ( .A1(\SB2_0_30/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_30/Component_Function_2/NAND4_in[2] ), .A3(n701), .A4(
        \SB2_0_30/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[26] ) );
  XNOR2_X1 U4838 ( .A(n2164), .B(n370), .ZN(Ciphertext[153]) );
  NAND4_X1 U4839 ( .A1(\SB4_6/Component_Function_3/NAND4_in[2] ), .A2(
        \SB4_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_6/Component_Function_3/NAND4_in[0] ), .A4(
        \SB4_6/Component_Function_3/NAND4_in[3] ), .ZN(n2164) );
  XNOR2_X1 U4840 ( .A(n2166), .B(n2165), .ZN(\RI1[3][167] ) );
  XNOR2_X1 U4841 ( .A(\MC_ARK_ARC_1_2/temp3[167] ), .B(
        \MC_ARK_ARC_1_2/temp1[167] ), .ZN(n2165) );
  XNOR2_X1 U4842 ( .A(\MC_ARK_ARC_1_2/temp2[167] ), .B(
        \MC_ARK_ARC_1_2/temp4[167] ), .ZN(n2166) );
  NAND3_X1 U4843 ( .A1(\SB2_1_12/i0_3 ), .A2(\SB2_1_12/i0[10] ), .A3(
        \SB2_1_12/i0[9] ), .ZN(\SB2_1_12/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U4844 ( .A1(\SB1_3_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_4/NAND4_in[2] ), .A4(n2167), .ZN(
        \RI3[3][64] ) );
  NAND3_X1 U4845 ( .A1(\SB1_3_22/i1[9] ), .A2(\SB1_3_22/i0_4 ), .A3(
        \SB1_3_22/i1_5 ), .ZN(n2167) );
  XNOR2_X1 U4846 ( .A(n2168), .B(\MC_ARK_ARC_1_0/temp6[152] ), .ZN(
        \RI1[1][152] ) );
  XNOR2_X1 U4847 ( .A(\MC_ARK_ARC_1_0/temp1[152] ), .B(
        \MC_ARK_ARC_1_0/temp2[152] ), .ZN(n2168) );
  NAND3_X1 U4848 ( .A1(\SB2_0_9/i0_0 ), .A2(\SB2_0_9/i0_4 ), .A3(
        \SB2_0_9/i1_5 ), .ZN(n2169) );
  NAND4_X1 U4849 ( .A1(\SB2_0_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_13/Component_Function_2/NAND4_in[1] ), .A4(n2170), .ZN(
        \RI5[0][128] ) );
  NAND3_X1 U4850 ( .A1(\SB2_0_13/i0_0 ), .A2(\SB2_0_13/i0_4 ), .A3(
        \SB2_0_13/i1_5 ), .ZN(n2170) );
  NAND3_X1 U4851 ( .A1(\SB3_6/i0[10] ), .A2(\SB3_6/i0_0 ), .A3(\SB3_6/i0[6] ), 
        .ZN(\SB3_6/Component_Function_5/NAND4_in[1] ) );
  XNOR2_X1 U4852 ( .A(n2171), .B(n278), .ZN(Ciphertext[167]) );
  NAND4_X1 U4853 ( .A1(\SB4_4/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_4/Component_Function_5/NAND4_in[1] ), .A3(n1806), .A4(
        \SB4_4/Component_Function_5/NAND4_in[0] ), .ZN(n2171) );
  XNOR2_X1 U4854 ( .A(\MC_ARK_ARC_1_0/temp5[173] ), .B(n2172), .ZN(
        \RI1[1][173] ) );
  XNOR2_X1 U4855 ( .A(\MC_ARK_ARC_1_0/temp4[173] ), .B(
        \MC_ARK_ARC_1_0/temp3[173] ), .ZN(n2172) );
  XNOR2_X1 U4856 ( .A(n2173), .B(n365), .ZN(Ciphertext[99]) );
  NAND4_X1 U4857 ( .A1(\SB4_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_15/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_15/Component_Function_3/NAND4_in[3] ), .ZN(n2173) );
  NAND3_X1 U4858 ( .A1(\SB2_3_21/i0_0 ), .A2(\SB2_3_21/i1_5 ), .A3(
        \RI3[3][64] ), .ZN(\SB2_3_21/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U4859 ( .A1(\SB4_29/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_29/Component_Function_2/NAND4_in[1] ), .A3(n1770), .A4(n2174), 
        .ZN(n1905) );
  NAND3_X1 U4860 ( .A1(\SB4_29/i0_0 ), .A2(n2131), .A3(\SB4_29/i1_5 ), .ZN(
        n2174) );
  NAND3_X1 U4861 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i1_5 ), .A3(
        \SB2_1_0/i1[9] ), .ZN(\SB2_1_0/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4862 ( .A1(n1284), .A2(\SB2_2_26/Component_Function_2/NAND4_in[0] ), .A3(\SB2_2_26/Component_Function_2/NAND4_in[1] ), .A4(n2175), .ZN(
        \RI5[2][50] ) );
  NAND3_X1 U4863 ( .A1(\SB2_2_26/i0_4 ), .A2(\SB2_2_26/i0_0 ), .A3(
        \SB2_2_26/i1_5 ), .ZN(n2175) );
  NAND4_X1 U4864 ( .A1(\SB3_0/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_0/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_0/Component_Function_2/NAND4_in[0] ), .A4(n2176), .ZN(
        \RI3[4][14] ) );
  NAND3_X1 U4865 ( .A1(\SB3_0/i1_5 ), .A2(\SB3_0/i0_0 ), .A3(\SB3_0/i0_4 ), 
        .ZN(n2176) );
  NAND4_X1 U4866 ( .A1(\SB4_28/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_28/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_28/Component_Function_2/NAND4_in[0] ), .A4(n2177), .ZN(n1885) );
  NAND3_X1 U4867 ( .A1(\SB4_28/i0_4 ), .A2(\SB4_28/i0_0 ), .A3(\SB4_28/i1_5 ), 
        .ZN(n2177) );
  NAND3_X1 U4868 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0[9] ), .A3(
        \SB2_2_30/i0[8] ), .ZN(\SB2_2_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4869 ( .A1(\SB2_3_5/i0_0 ), .A2(\SB2_3_5/i1_5 ), .A3(
        \SB2_3_5/i0_4 ), .ZN(\SB2_3_5/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U4870 ( .A1(\SB1_3_6/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_3_6/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_5/i0_4 ) );
  NAND3_X1 U4871 ( .A1(\SB2_0_2/i0_0 ), .A2(\SB2_0_2/i1_5 ), .A3(
        \SB2_0_2/i0_4 ), .ZN(\SB2_0_2/Component_Function_2/NAND4_in[3] ) );
  NAND4_X4 U4872 ( .A1(\SB2_1_7/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_7/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_7/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_1_7/Component_Function_4/NAND4_in[1] ), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[154] ) );
  NAND3_X1 U4873 ( .A1(\SB1_0_5/i0_4 ), .A2(\SB1_0_5/i1_5 ), .A3(
        \SB1_0_5/i1[9] ), .ZN(\SB1_0_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4874 ( .A1(\SB1_2_21/i0_0 ), .A2(\SB1_2_21/i0_4 ), .A3(
        \SB1_2_21/i1_5 ), .ZN(n883) );
  NAND3_X1 U4875 ( .A1(\SB2_1_27/i0_3 ), .A2(\SB2_1_27/i0_4 ), .A3(
        \SB2_1_27/i1[9] ), .ZN(n1243) );
  NAND3_X1 U4876 ( .A1(\SB2_1_7/i0_0 ), .A2(\SB2_1_7/i3[0] ), .A3(
        \SB2_1_7/i1_7 ), .ZN(\SB2_1_7/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U4877 ( .A1(\SB2_2_23/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_23/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_2_23/Component_Function_2/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[68] ) );
  NAND3_X1 U4878 ( .A1(\SB1_0_9/i0[6] ), .A2(\SB1_0_9/i0[9] ), .A3(
        \SB1_0_9/i0_4 ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[3] ) );
  INV_X1 U4879 ( .A(\RI3[0][80] ), .ZN(\SB2_0_18/i1[9] ) );
  NAND4_X1 U4880 ( .A1(\SB1_0_21/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_0_21/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[0][80] ) );
  NAND3_X1 U4881 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0[8] ), .A3(\SB4_1/i0[9] ), 
        .ZN(n2178) );
  NAND3_X1 U4882 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0[10] ), .A3(
        \SB1_0_9/i0_4 ), .ZN(\SB1_0_9/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U4883 ( .A1(\SB2_0_14/Component_Function_3/NAND4_in[0] ), .A2(n2179), .A3(\SB2_0_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_14/Component_Function_3/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[117] ) );
  NAND3_X1 U4884 ( .A1(\SB2_0_14/i0_0 ), .A2(\SB2_0_14/i0_4 ), .A3(
        \SB2_0_14/i0_3 ), .ZN(n2179) );
  NAND3_X1 U4885 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i0_3 ), .A3(
        \SB1_3_10/i0[9] ), .ZN(\SB1_3_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4886 ( .A1(\SB4_2/i0_4 ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i1_5 ), 
        .ZN(\SB4_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4887 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i0[9] ), .A3(\SB3_7/i0_3 ), 
        .ZN(\SB3_7/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U4888 ( .A(n2180), .B(n340), .ZN(Ciphertext[185]) );
  NAND4_X1 U4889 ( .A1(\SB4_1/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_1/Component_Function_5/NAND4_in[2] ), .A3(n2187), .A4(
        \SB4_1/Component_Function_5/NAND4_in[0] ), .ZN(n2180) );
  INV_X2 U4890 ( .A(\RI1[1][107] ), .ZN(\SB1_1_14/i0_3 ) );
  XNOR2_X1 U4891 ( .A(\MC_ARK_ARC_1_0/temp6[107] ), .B(
        \MC_ARK_ARC_1_0/temp5[107] ), .ZN(\RI1[1][107] ) );
  NAND4_X2 U4892 ( .A1(\SB2_0_10/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_10/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_10/Component_Function_5/NAND4_in[1] ), .A4(n2181), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[131] ) );
  NAND2_X1 U4893 ( .A1(\SB2_0_10/i0_0 ), .A2(\SB2_0_10/i3[0] ), .ZN(n2181) );
  NAND3_X1 U4894 ( .A1(\SB2_3_4/i0[10] ), .A2(\SB2_3_4/i1_5 ), .A3(
        \SB2_3_4/i1[9] ), .ZN(\SB2_3_4/Component_Function_2/NAND4_in[0] ) );
  XNOR2_X1 U4895 ( .A(n2182), .B(n335), .ZN(Ciphertext[131]) );
  NAND4_X1 U4896 ( .A1(\SB4_10/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_10/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_10/Component_Function_5/NAND4_in[0] ), .ZN(n2182) );
  XNOR2_X1 U4897 ( .A(n2183), .B(n299), .ZN(Ciphertext[150]) );
  NAND4_X1 U4898 ( .A1(\SB4_6/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_6/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_6/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_6/Component_Function_0/NAND4_in[0] ), .ZN(n2183) );
  NAND4_X1 U4899 ( .A1(\SB2_2_29/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_29/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_29/Component_Function_4/NAND4_in[1] ), .A4(n2184), .ZN(
        \RI5[2][22] ) );
  NAND3_X1 U4900 ( .A1(\SB2_2_29/i0_4 ), .A2(\SB2_2_29/i1[9] ), .A3(
        \SB2_2_29/i1_5 ), .ZN(n2184) );
  NAND4_X2 U4901 ( .A1(\SB2_1_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_3/NAND4_in[1] ), .A3(n2185), .A4(
        \SB2_1_21/Component_Function_3/NAND4_in[3] ), .ZN(\RI5[1][75] ) );
  NAND3_X1 U4902 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i1[9] ), .A3(
        \SB2_1_21/i1_7 ), .ZN(n2185) );
  NAND4_X2 U4903 ( .A1(\SB2_3_27/Component_Function_5/NAND4_in[3] ), .A2(n690), 
        .A3(\SB2_3_27/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[29] ) );
  NAND4_X1 U4904 ( .A1(\SB2_3_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_17/Component_Function_5/NAND4_in[0] ), .A3(n1074), .A4(n2186), 
        .ZN(\RI5[3][89] ) );
  NAND3_X1 U4905 ( .A1(\SB2_3_17/i0[10] ), .A2(\SB2_3_17/i0_0 ), .A3(
        \SB2_3_17/i0[6] ), .ZN(n2186) );
  NAND3_X1 U4906 ( .A1(n828), .A2(\SB4_12/i0_4 ), .A3(\SB4_12/i1[9] ), .ZN(
        \SB4_12/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4907 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i1[9] ), .A3(\SB4_0/i1_5 ), 
        .ZN(\SB4_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4908 ( .A1(\SB3_19/i0_0 ), .A2(\SB3_19/i0[10] ), .A3(
        \SB3_19/i0[6] ), .ZN(\SB3_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4909 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i1[9] ), .ZN(n1276) );
  NAND3_X1 U4910 ( .A1(\SB2_3_14/i0_3 ), .A2(n1945), .A3(\SB2_3_14/i1[9] ), 
        .ZN(n1322) );
  NAND3_X1 U4911 ( .A1(\SB1_3_5/i0[6] ), .A2(\SB1_3_5/i0_0 ), .A3(
        \SB1_3_5/i0[10] ), .ZN(\SB1_3_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4912 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i1_5 ), .A3(
        \SB2_3_11/i1[9] ), .ZN(\SB2_3_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4913 ( .A1(\SB2_2_21/i0_4 ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB2_2_21/i0_0 ), .ZN(\SB2_2_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4914 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0[10] ), .A3(
        \SB1_0_23/i0[9] ), .ZN(\SB1_0_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4915 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0[10] ), .A3(\SB4_1/i0[6] ), 
        .ZN(n2187) );
  NAND4_X1 U4916 ( .A1(\SB2_1_30/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_30/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_30/Component_Function_2/NAND4_in[1] ), .A4(n2188), .ZN(
        \RI5[1][26] ) );
  NAND3_X1 U4917 ( .A1(\SB2_1_30/i0_4 ), .A2(\SB2_1_30/i0_0 ), .A3(
        \SB2_1_30/i1_5 ), .ZN(n2188) );
  NAND3_X1 U4918 ( .A1(\SB2_3_9/i0_0 ), .A2(\SB2_3_9/i3[0] ), .A3(
        \SB2_3_9/i1_7 ), .ZN(\SB2_3_9/Component_Function_4/NAND4_in[1] ) );
  NAND4_X1 U4919 ( .A1(\SB1_2_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_30/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_30/Component_Function_5/NAND4_in[0] ), .A4(n2189), .ZN(
        \RI3[2][11] ) );
  NAND3_X1 U4920 ( .A1(\SB1_2_30/i0_3 ), .A2(\SB1_2_30/i1[9] ), .A3(
        \SB1_2_30/i0_4 ), .ZN(n2189) );
  XNOR2_X1 U4921 ( .A(n2190), .B(n287), .ZN(Ciphertext[1]) );
  NAND4_X1 U4922 ( .A1(n1297), .A2(\SB4_31/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB4_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_31/Component_Function_1/NAND4_in[0] ), .ZN(n2190) );
  NAND4_X1 U4923 ( .A1(\SB3_0/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_0/Component_Function_4/NAND4_in[0] ), .A4(n2191), .ZN(\RI3[4][4] ) );
  NAND3_X1 U4924 ( .A1(\SB3_0/i1_5 ), .A2(\SB3_0/i1[9] ), .A3(\SB3_0/i0_4 ), 
        .ZN(n2191) );
  INV_X1 U4925 ( .A(\RI3[0][83] ), .ZN(\SB2_0_18/i1_5 ) );
  NAND4_X1 U4926 ( .A1(n1156), .A2(\SB1_0_18/Component_Function_5/NAND4_in[1] ), .A3(\SB1_0_18/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_18/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][83] ) );
  XNOR2_X1 U4927 ( .A(\MC_ARK_ARC_1_2/buf_datainput[155] ), .B(n802), .ZN(
        \MC_ARK_ARC_1_2/temp2[17] ) );
  NAND4_X2 U4928 ( .A1(\SB2_2_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_2/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_2/Component_Function_5/NAND4_in[1] ), .A4(n1028), .ZN(n802) );
  NAND3_X1 U4929 ( .A1(\SB2_0_16/i0[10] ), .A2(\SB2_0_16/i1[9] ), .A3(
        \SB2_0_16/i1_7 ), .ZN(\SB2_0_16/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U4930 ( .A(\RI1[1][95] ), .ZN(\SB1_1_16/i0_3 ) );
  XNOR2_X1 U4931 ( .A(n1356), .B(n1355), .ZN(\RI1[1][95] ) );
  NAND3_X1 U4932 ( .A1(n828), .A2(\SB4_12/i0[7] ), .A3(\SB4_12/i0_0 ), .ZN(
        \SB4_12/Component_Function_0/NAND4_in[3] ) );
  NAND4_X1 U4933 ( .A1(\SB3_4/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_4/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_4/Component_Function_2/NAND4_in[3] ), .A4(n2192), .ZN(
        \RI3[4][182] ) );
  NAND3_X1 U4934 ( .A1(\SB3_4/i0[8] ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0[9] ), 
        .ZN(n2192) );
  NAND3_X1 U4935 ( .A1(\SB2_1_16/i0_3 ), .A2(\SB2_1_16/i0[6] ), .A3(
        \SB2_1_16/i1[9] ), .ZN(\SB2_1_16/Component_Function_3/NAND4_in[0] ) );
  NAND4_X1 U4936 ( .A1(\SB1_1_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_16/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_1_16/Component_Function_5/NAND4_in[1] ), .A4(n2193), .ZN(
        \RI3[1][95] ) );
  NAND3_X1 U4937 ( .A1(\SB1_1_16/i0[9] ), .A2(\SB1_1_16/i0[6] ), .A3(
        \SB1_1_16/i0_4 ), .ZN(n2193) );
  NAND3_X1 U4938 ( .A1(\SB2_2_11/i0[10] ), .A2(\SB2_2_11/i0_0 ), .A3(
        \SB2_2_11/i0[6] ), .ZN(\SB2_2_11/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U4939 ( .A1(\SB2_0_15/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[126] ) );
  NAND4_X2 U4940 ( .A1(\SB1_0_16/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_16/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_0_16/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_0_15/i0_4 ) );
  NAND3_X1 U4941 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i1[9] ), .A3(
        \SB2_3_17/i0_4 ), .ZN(\SB2_3_17/Component_Function_5/NAND4_in[2] ) );
  XNOR2_X1 U4942 ( .A(n2194), .B(n244), .ZN(Ciphertext[35]) );
  NAND4_X1 U4943 ( .A1(\SB4_26/Component_Function_5/NAND4_in[2] ), .A2(n2215), 
        .A3(\SB4_26/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_26/Component_Function_5/NAND4_in[0] ), .ZN(n2194) );
  NAND4_X1 U4944 ( .A1(\SB1_2_2/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_2/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_2/Component_Function_0/NAND4_in[1] ), .A4(n2195), .ZN(
        \RI3[2][12] ) );
  NAND3_X1 U4945 ( .A1(n1648), .A2(\SB1_2_2/i0[10] ), .A3(\SB1_2_2/i0_4 ), 
        .ZN(n2195) );
  XNOR2_X1 U4946 ( .A(n2197), .B(n2196), .ZN(\RI1[1][167] ) );
  XNOR2_X1 U4947 ( .A(\MC_ARK_ARC_1_0/temp3[167] ), .B(
        \MC_ARK_ARC_1_0/temp4[167] ), .ZN(n2196) );
  XNOR2_X1 U4948 ( .A(\MC_ARK_ARC_1_0/temp1[167] ), .B(
        \MC_ARK_ARC_1_0/temp2[167] ), .ZN(n2197) );
  NAND3_X1 U4949 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0[10] ), .A3(
        \SB1_0_10/i0_4 ), .ZN(\SB1_0_10/Component_Function_0/NAND4_in[2] ) );
  XNOR2_X1 U4950 ( .A(n2198), .B(\MC_ARK_ARC_1_3/temp6[94] ), .ZN(\RI1[4][94] ) );
  XNOR2_X1 U4951 ( .A(\MC_ARK_ARC_1_3/temp2[94] ), .B(
        \MC_ARK_ARC_1_3/temp1[94] ), .ZN(n2198) );
  NAND4_X1 U4952 ( .A1(\SB1_3_5/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_5/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_5/Component_Function_2/NAND4_in[2] ), .A4(n2199), .ZN(
        \RI3[3][176] ) );
  NAND3_X1 U4953 ( .A1(\SB1_3_5/i0_4 ), .A2(\SB1_3_5/i0_0 ), .A3(
        \SB1_3_5/i1_5 ), .ZN(n2199) );
  NAND3_X1 U4954 ( .A1(\SB1_1_2/i0[8] ), .A2(\SB1_1_2/i0_0 ), .A3(
        \SB1_1_2/i0[9] ), .ZN(\SB1_1_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U4955 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i1[9] ), .A3(
        \SB1_2_2/i0_4 ), .ZN(n2230) );
  NAND4_X1 U4956 ( .A1(\SB1_1_18/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_1_18/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_18/Component_Function_1/NAND4_in[0] ), .A4(n2200), .ZN(
        \RI3[1][103] ) );
  NAND3_X1 U4957 ( .A1(\SB1_1_18/i1_7 ), .A2(\SB1_1_18/i0_3 ), .A3(
        \SB1_1_18/i0[8] ), .ZN(n2200) );
  NAND3_X1 U4958 ( .A1(\SB2_3_7/i0_0 ), .A2(\SB2_3_7/i3[0] ), .A3(
        \SB2_3_7/i1_7 ), .ZN(\SB2_3_7/Component_Function_4/NAND4_in[1] ) );
  INV_X2 U4959 ( .A(\RI1[2][185] ), .ZN(\SB1_2_1/i0_3 ) );
  XNOR2_X1 U4960 ( .A(n1813), .B(n1814), .ZN(\RI1[2][185] ) );
  NAND4_X2 U4961 ( .A1(\SB2_2_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_30/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_30/Component_Function_5/NAND4_in[1] ), .A4(n2201), .ZN(
        \MC_ARK_ARC_1_2/buf_datainput[11] ) );
  NAND2_X1 U4962 ( .A1(\SB2_2_30/i0_0 ), .A2(\SB2_2_30/i3[0] ), .ZN(n2201) );
  NAND4_X1 U4963 ( .A1(\SB2_1_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_29/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_1_29/Component_Function_4/NAND4_in[1] ), .A4(n2202), .ZN(
        \RI5[1][22] ) );
  NAND3_X1 U4964 ( .A1(\SB2_1_29/i0_4 ), .A2(\SB2_1_29/i1[9] ), .A3(
        \SB2_1_29/i1_5 ), .ZN(n2202) );
  NAND3_X1 U4965 ( .A1(\SB2_3_25/i0[10] ), .A2(\SB2_3_25/i1_5 ), .A3(
        \SB2_3_25/i1[9] ), .ZN(\SB2_3_25/Component_Function_2/NAND4_in[0] ) );
  NAND4_X1 U4966 ( .A1(\SB1_2_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_13/Component_Function_5/NAND4_in[0] ), .A4(n2203), .ZN(
        \RI3[2][113] ) );
  NAND3_X1 U4967 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i1[9] ), .A3(
        \SB1_2_13/i0_4 ), .ZN(n2203) );
  XNOR2_X1 U4968 ( .A(n2204), .B(n371), .ZN(Ciphertext[2]) );
  NAND4_X1 U4969 ( .A1(\SB4_31/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_31/Component_Function_2/NAND4_in[3] ), .A3(
        \SB4_31/Component_Function_2/NAND4_in[1] ), .A4(n1894), .ZN(n2204) );
  NAND3_X1 U4970 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0[9] ), .A3(
        \SB2_3_26/i0[10] ), .ZN(\SB2_3_26/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U4971 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i1[9] ), .A3(
        \SB2_3_4/i0_4 ), .ZN(n2205) );
  NAND3_X1 U4972 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0[10] ), .A3(
        \SB1_0_10/i0[9] ), .ZN(\SB1_0_10/Component_Function_4/NAND4_in[2] ) );
  XNOR2_X1 U4973 ( .A(\MC_ARK_ARC_1_1/temp5[105] ), .B(n2206), .ZN(
        \RI1[2][105] ) );
  XNOR2_X1 U4974 ( .A(\MC_ARK_ARC_1_1/temp3[105] ), .B(
        \MC_ARK_ARC_1_1/temp4[105] ), .ZN(n2206) );
  NAND4_X1 U4975 ( .A1(\SB1_1_17/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_17/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_17/Component_Function_5/NAND4_in[0] ), .A4(n2207), .ZN(
        \RI3[1][89] ) );
  NAND3_X1 U4976 ( .A1(\SB1_1_17/i1[9] ), .A2(\SB1_1_17/i0_4 ), .A3(
        \SB1_1_17/i0_3 ), .ZN(n2207) );
  NAND4_X1 U4977 ( .A1(\SB1_3_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_13/Component_Function_5/NAND4_in[0] ), .A4(n2208), .ZN(
        \RI3[3][113] ) );
  NAND3_X1 U4978 ( .A1(\SB1_3_13/i1[9] ), .A2(\SB1_3_13/i0_4 ), .A3(
        \SB1_3_13/i0_3 ), .ZN(n2208) );
  NAND3_X1 U4979 ( .A1(\SB2_1_26/i0[10] ), .A2(\SB2_1_26/i1_5 ), .A3(
        \SB2_1_26/i1[9] ), .ZN(n2209) );
  XNOR2_X1 U4980 ( .A(n2210), .B(n225), .ZN(Ciphertext[175]) );
  NAND4_X1 U4981 ( .A1(\SB4_2/Component_Function_1/NAND4_in[1] ), .A2(n1221), 
        .A3(\SB4_2/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_2/Component_Function_1/NAND4_in[2] ), .ZN(n2210) );
  INV_X2 U4982 ( .A(\RI1[1][47] ), .ZN(\SB1_1_24/i0_3 ) );
  XNOR2_X1 U4983 ( .A(n1697), .B(n1696), .ZN(\RI1[1][47] ) );
  NAND4_X1 U4984 ( .A1(\SB4_14/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_14/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_14/Component_Function_4/NAND4_in[1] ), .A4(n2211), .ZN(n1551) );
  NAND3_X1 U4985 ( .A1(\SB4_14/i1[9] ), .A2(n799), .A3(\SB4_14/i1_5 ), .ZN(
        n2211) );
  XNOR2_X1 U4986 ( .A(n2212), .B(n202), .ZN(Ciphertext[0]) );
  NAND4_X1 U4987 ( .A1(\SB4_31/Component_Function_0/NAND4_in[3] ), .A2(n2216), 
        .A3(n1108), .A4(\SB4_31/Component_Function_0/NAND4_in[0] ), .ZN(n2212)
         );
  XNOR2_X1 U4988 ( .A(\MC_ARK_ARC_1_2/temp5[92] ), .B(n2213), .ZN(\RI1[3][92] ) );
  XNOR2_X1 U4989 ( .A(\MC_ARK_ARC_1_2/temp3[92] ), .B(
        \MC_ARK_ARC_1_2/temp4[92] ), .ZN(n2213) );
  XNOR2_X1 U4990 ( .A(n2214), .B(n361), .ZN(Ciphertext[127]) );
  NAND4_X1 U4991 ( .A1(\SB4_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_10/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_10/Component_Function_1/NAND4_in[0] ), .A4(n1323), .ZN(n2214) );
  NAND3_X1 U4992 ( .A1(\SB1_3_0/i0[10] ), .A2(\SB1_3_0/i0_0 ), .A3(
        \SB1_3_0/i0[6] ), .ZN(\SB1_3_0/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U4993 ( .A1(\SB2_3_0/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_0/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_3_0/Component_Function_4/NAND4_in[3] ), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[4] ) );
  NAND3_X1 U4994 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i1_5 ), .A3(
        \SB2_1_24/i1[9] ), .ZN(\SB2_1_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4995 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[9] ), .A3(
        \SB3_30/i0[10] ), .ZN(\SB3_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4996 ( .A1(\SB1_2_6/i1[9] ), .A2(\SB1_2_6/i0_3 ), .A3(
        \SB1_2_6/i0_4 ), .ZN(\SB1_2_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4997 ( .A1(\SB4_26/i0_0 ), .A2(\SB4_26/i0[10] ), .A3(
        \SB4_26/i0[6] ), .ZN(n2215) );
  NAND3_X1 U4998 ( .A1(\SB4_31/i0_4 ), .A2(n1670), .A3(\SB4_31/i0[10] ), .ZN(
        n2216) );
  NAND3_X1 U4999 ( .A1(\SB2_0_7/i0_3 ), .A2(\SB2_0_7/i0[9] ), .A3(
        \SB2_0_7/i0[10] ), .ZN(n2217) );
  NAND3_X1 U5000 ( .A1(\SB1_0_14/i0[9] ), .A2(\SB1_0_14/i0[8] ), .A3(
        \SB1_0_14/i0_3 ), .ZN(\SB1_0_14/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U5001 ( .A1(\SB2_0_21/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_21/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_21/Component_Function_1/NAND4_in[0] ), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[85] ) );
  NAND4_X2 U5002 ( .A1(\SB2_1_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_3/NAND4_in[2] ), .A4(n2218), .ZN(
        \RI5[1][141] ) );
  NAND3_X1 U5003 ( .A1(\SB2_1_10/i3[0] ), .A2(\SB2_1_10/i0[8] ), .A3(
        \SB2_1_10/i1_5 ), .ZN(n2218) );
  NAND3_X1 U5004 ( .A1(\SB1_2_16/i0_0 ), .A2(\SB1_2_16/i0_4 ), .A3(
        \SB1_2_16/i1_5 ), .ZN(n1858) );
  NAND4_X1 U5005 ( .A1(\SB2_2_29/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_2_29/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_29/Component_Function_2/NAND4_in[2] ), .A4(n2219), .ZN(
        \RI5[2][32] ) );
  NAND3_X1 U5006 ( .A1(\SB2_2_29/i0_4 ), .A2(\SB2_2_29/i0_0 ), .A3(
        \SB2_2_29/i1_5 ), .ZN(n2219) );
  XNOR2_X1 U5007 ( .A(\MC_ARK_ARC_1_1/temp5[94] ), .B(n2220), .ZN(\RI1[2][94] ) );
  XNOR2_X1 U5008 ( .A(\MC_ARK_ARC_1_1/temp3[94] ), .B(
        \MC_ARK_ARC_1_1/temp4[94] ), .ZN(n2220) );
  NAND4_X1 U5009 ( .A1(\SB1_3_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_1/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_1/Component_Function_3/NAND4_in[3] ), .A4(n2221), .ZN(
        \RI3[3][3] ) );
  NAND3_X1 U5010 ( .A1(\SB1_3_1/i1[9] ), .A2(\SB1_3_1/i1_7 ), .A3(
        \SB1_3_1/i0[10] ), .ZN(n2221) );
  NAND4_X1 U5011 ( .A1(\SB1_2_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_12/Component_Function_0/NAND4_in[0] ), .A4(n2222), .ZN(
        \RI3[2][144] ) );
  NAND3_X1 U5012 ( .A1(\SB1_2_12/i0[7] ), .A2(\SB1_2_12/i0_0 ), .A3(
        \SB1_2_12/i0_3 ), .ZN(n2222) );
  NAND3_X1 U5013 ( .A1(\SB4_17/i0_0 ), .A2(\SB4_17/i3[0] ), .A3(\SB4_17/i1_7 ), 
        .ZN(n2223) );
  NAND4_X1 U5014 ( .A1(\SB1_2_15/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_15/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_15/Component_Function_2/NAND4_in[2] ), .A4(n2224), .ZN(
        \RI3[2][116] ) );
  NAND3_X1 U5015 ( .A1(\SB1_2_15/i0_0 ), .A2(\SB1_2_15/i0_4 ), .A3(
        \SB1_2_15/i1_5 ), .ZN(n2224) );
  NAND3_X1 U5016 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i1_5 ), .A3(
        \SB2_2_12/i1[9] ), .ZN(\SB2_2_12/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U5017 ( .A1(\SB2_0_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_29/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_29/Component_Function_5/NAND4_in[1] ), .A4(n2225), .ZN(
        \MC_ARK_ARC_1_0/buf_datainput[17] ) );
  NAND2_X1 U5018 ( .A1(\SB2_0_29/i0_0 ), .A2(\SB2_0_29/i3[0] ), .ZN(n2225) );
  XNOR2_X1 U5019 ( .A(n2227), .B(n2226), .ZN(\RI1[1][35] ) );
  XNOR2_X1 U5020 ( .A(\MC_ARK_ARC_1_0/temp4[35] ), .B(
        \MC_ARK_ARC_1_0/temp1[35] ), .ZN(n2226) );
  XNOR2_X1 U5021 ( .A(\MC_ARK_ARC_1_0/temp3[35] ), .B(
        \MC_ARK_ARC_1_0/temp2[35] ), .ZN(n2227) );
  NAND3_X1 U5022 ( .A1(\SB2_1_19/i0_3 ), .A2(\SB2_1_19/i0[9] ), .A3(
        \SB2_1_19/i0[10] ), .ZN(n2228) );
  NAND4_X1 U5023 ( .A1(\SB1_1_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_18/Component_Function_5/NAND4_in[0] ), .A4(n2229), .ZN(
        \RI3[1][83] ) );
  NAND3_X1 U5024 ( .A1(\SB1_1_18/i1[9] ), .A2(\SB1_1_18/i0_3 ), .A3(
        \SB1_1_18/i0_4 ), .ZN(n2229) );
  NAND4_X1 U5025 ( .A1(\SB1_2_2/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_2/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_2/Component_Function_5/NAND4_in[0] ), .A4(n2230), .ZN(
        \RI3[2][179] ) );
  XNOR2_X1 U5026 ( .A(n2231), .B(n410), .ZN(Ciphertext[30]) );
  NAND4_X1 U5027 ( .A1(\SB4_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_26/Component_Function_0/NAND4_in[3] ), .A3(n1545), .A4(
        \SB4_26/Component_Function_0/NAND4_in[0] ), .ZN(n2231) );
  NAND3_X1 U5028 ( .A1(\SB4_17/i0[9] ), .A2(\SB4_17/i0_0 ), .A3(\SB4_17/i0[8] ), .ZN(n2232) );
  NAND4_X1 U5029 ( .A1(\SB3_22/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_0/NAND4_in[0] ), .A4(n2233), .ZN(
        \RI3[4][84] ) );
  NAND3_X1 U5030 ( .A1(\SB3_22/i0[7] ), .A2(\SB3_22/i0_3 ), .A3(\SB3_22/i0_0 ), 
        .ZN(n2233) );
  NAND3_X1 U5031 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0[9] ), .A3(
        \SB1_0_6/i0[8] ), .ZN(\SB1_0_6/Component_Function_2/NAND4_in[2] ) );
  NAND4_X1 U5032 ( .A1(\SB1_3_26/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_26/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_26/Component_Function_2/NAND4_in[2] ), .A4(n2234), .ZN(
        \RI3[3][50] ) );
  NAND3_X1 U5033 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i0_4 ), .A3(
        \SB1_3_26/i1_5 ), .ZN(n2234) );
  NAND4_X1 U5034 ( .A1(\SB1_1_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_13/Component_Function_5/NAND4_in[0] ), .A4(n2235), .ZN(
        \RI3[1][113] ) );
  NAND3_X1 U5035 ( .A1(\SB1_1_13/i1[9] ), .A2(\SB1_1_13/i0_3 ), .A3(
        \SB1_1_13/i0_4 ), .ZN(n2235) );
  NAND4_X1 U5036 ( .A1(\SB1_1_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_5/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_1_5/Component_Function_5/NAND4_in[0] ), .A4(n2236), .ZN(
        \RI3[1][161] ) );
  NAND3_X1 U5037 ( .A1(\SB1_1_5/i1[9] ), .A2(\SB1_1_5/i0_3 ), .A3(
        \SB1_1_5/i0_4 ), .ZN(n2236) );
  INV_X1 U5038 ( .A(\RI3[0][116] ), .ZN(\SB2_0_12/i1[9] ) );
  NAND4_X1 U5039 ( .A1(\SB1_0_15/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_15/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_15/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_0_15/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][116] ) );
  NAND3_X1 U5040 ( .A1(\SB1_0_20/i0[7] ), .A2(\SB1_0_20/i0_3 ), .A3(
        \SB1_0_20/i0_0 ), .ZN(\SB1_0_20/Component_Function_0/NAND4_in[3] ) );
  XNOR2_X1 U5041 ( .A(n2237), .B(n210), .ZN(Ciphertext[136]) );
  NAND4_X1 U5042 ( .A1(n1572), .A2(\SB4_9/Component_Function_4/NAND4_in[0] ), 
        .A3(n1563), .A4(\SB4_9/Component_Function_4/NAND4_in[3] ), .ZN(n2237)
         );
  NAND4_X1 U5043 ( .A1(\SB1_3_26/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_26/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_26/Component_Function_5/NAND4_in[0] ), .A4(n2238), .ZN(
        \RI3[3][35] ) );
  NAND3_X1 U5044 ( .A1(\SB1_3_26/i1[9] ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0_4 ), .ZN(n2238) );
  NAND4_X1 U5045 ( .A1(\SB1_0_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_0_8/Component_Function_5/NAND4_in[0] ), .A4(n2239), .ZN(
        \RI3[0][143] ) );
  NAND3_X1 U5046 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0_4 ), .A3(
        \SB1_0_8/i1[9] ), .ZN(n2239) );
  NAND3_X1 U5047 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0[10] ), .A3(
        \SB1_0_0/i0_4 ), .ZN(\SB1_0_0/Component_Function_0/NAND4_in[2] ) );
  NAND4_X1 U5048 ( .A1(\SB1_3_14/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_14/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_14/Component_Function_5/NAND4_in[0] ), .A4(n2240), .ZN(
        \RI3[3][107] ) );
  NAND3_X1 U5049 ( .A1(\SB1_3_14/i1[9] ), .A2(\SB1_3_14/i0_3 ), .A3(
        \SB1_3_14/i0_4 ), .ZN(n2240) );
  NAND4_X1 U5050 ( .A1(\SB1_2_23/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_2_23/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_5/NAND4_in[0] ), .A4(n2241), .ZN(
        \RI3[2][53] ) );
  NAND3_X1 U5051 ( .A1(\SB1_2_23/i1[9] ), .A2(\SB1_2_23/i0_3 ), .A3(
        \SB1_2_23/i0_4 ), .ZN(n2241) );
  XNOR2_X1 U5052 ( .A(n2242), .B(n326), .ZN(Ciphertext[146]) );
  XNOR2_X1 U5053 ( .A(n2243), .B(\MC_ARK_ARC_1_3/temp6[123] ), .ZN(
        \RI1[4][123] ) );
  XNOR2_X1 U5054 ( .A(\MC_ARK_ARC_1_3/temp2[123] ), .B(
        \MC_ARK_ARC_1_3/temp1[123] ), .ZN(n2243) );
  NAND3_X1 U5055 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i0[10] ), .A3(
        \SB1_0_17/i0[9] ), .ZN(\SB1_0_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U5056 ( .A1(n877), .A2(\SB4_7/i0[7] ), .A3(\SB4_7/i0_0 ), .ZN(
        \SB4_7/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U5057 ( .A1(\SB2_1_3/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_3/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_3/Component_Function_2/NAND4_in[1] ), .A4(n613), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[188] ) );
  NAND3_X1 U5058 ( .A1(\SB4_3/i0[10] ), .A2(\SB4_3/i1_5 ), .A3(\SB4_3/i1[9] ), 
        .ZN(n2244) );
  NAND3_X1 U5059 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0[10] ), .A3(
        \SB1_0_12/i0_4 ), .ZN(\SB1_0_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U5060 ( .A1(\SB2_2_21/i0[10] ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB2_2_21/i1[9] ), .ZN(\SB2_2_21/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U5061 ( .A1(\SB1_3_23/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_4/NAND4_in[0] ), .A3(n1096), .A4(
        \SB1_3_23/Component_Function_4/NAND4_in[3] ), .ZN(\SB2_3_22/i0_4 ) );
  NAND4_X2 U5062 ( .A1(\SB2_1_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_7/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_7/Component_Function_2/NAND4_in[1] ), .A4(n1712), .ZN(n1625) );
  INV_X2 U5063 ( .A(\RI1[2][137] ), .ZN(n1657) );
  NAND4_X2 U5064 ( .A1(\SB2_2_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_12/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_12/Component_Function_5/NAND4_in[0] ), .ZN(n811) );
  NAND4_X2 U5065 ( .A1(\SB2_2_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[2][133] ) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFF_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CK(clk), .Q(reg_in[191]) );
  DFF_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CK(clk), .Q(reg_in[190]) );
  DFF_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CK(clk), .Q(reg_in[189]) );
  DFF_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CK(clk), .Q(reg_in[188]) );
  DFF_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CK(clk), .Q(reg_in[187]) );
  DFF_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CK(clk), .Q(reg_in[186]) );
  DFF_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CK(clk), .Q(reg_in[185]) );
  DFF_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CK(clk), .Q(reg_in[184]) );
  DFF_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CK(clk), .Q(reg_in[183]) );
  DFF_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CK(clk), .Q(reg_in[182]) );
  DFF_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CK(clk), .Q(reg_in[181]) );
  DFF_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CK(clk), .Q(reg_in[180]) );
  DFF_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CK(clk), .Q(reg_in[179]) );
  DFF_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CK(clk), .Q(reg_in[178]) );
  DFF_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CK(clk), .Q(reg_in[177]) );
  DFF_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CK(clk), .Q(reg_in[176]) );
  DFF_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CK(clk), .Q(reg_in[175]) );
  DFF_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CK(clk), .Q(reg_in[174]) );
  DFF_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CK(clk), .Q(reg_in[173]) );
  DFF_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CK(clk), .Q(reg_in[172]) );
  DFF_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CK(clk), .Q(reg_in[171]) );
  DFF_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CK(clk), .Q(reg_in[170]) );
  DFF_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CK(clk), .Q(reg_in[169]) );
  DFF_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CK(clk), .Q(reg_in[168]) );
  DFF_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CK(clk), .Q(reg_in[167]) );
  DFF_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CK(clk), .Q(reg_in[166]) );
  DFF_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CK(clk), .Q(reg_in[165]) );
  DFF_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CK(clk), .Q(reg_in[164]) );
  DFF_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CK(clk), .Q(reg_in[163]) );
  DFF_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CK(clk), .Q(reg_in[162]) );
  DFF_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CK(clk), .Q(reg_in[161]) );
  DFF_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CK(clk), .Q(reg_in[160]) );
  DFF_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CK(clk), .Q(reg_in[159]) );
  DFF_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CK(clk), .Q(reg_in[158]) );
  DFF_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CK(clk), .Q(reg_in[157]) );
  DFF_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CK(clk), .Q(reg_in[156]) );
  DFF_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CK(clk), .Q(reg_in[155]) );
  DFF_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CK(clk), .Q(reg_in[154]) );
  DFF_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CK(clk), .Q(reg_in[153]) );
  DFF_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CK(clk), .Q(reg_in[152]) );
  DFF_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CK(clk), .Q(reg_in[151]) );
  DFF_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CK(clk), .Q(reg_in[150]) );
  DFF_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CK(clk), .Q(reg_in[149]) );
  DFF_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CK(clk), .Q(reg_in[148]) );
  DFF_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CK(clk), .Q(reg_in[147]) );
  DFF_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CK(clk), .Q(reg_in[146]) );
  DFF_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CK(clk), .Q(reg_in[145]) );
  DFF_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CK(clk), .Q(reg_in[144]) );
  DFF_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CK(clk), .Q(reg_in[143]) );
  DFF_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CK(clk), .Q(reg_in[142]) );
  DFF_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CK(clk), .Q(reg_in[141]) );
  DFF_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CK(clk), .Q(reg_in[140]) );
  DFF_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CK(clk), .Q(reg_in[139]) );
  DFF_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CK(clk), .Q(reg_in[138]) );
  DFF_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CK(clk), .Q(reg_in[137]) );
  DFF_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CK(clk), .Q(reg_in[136]) );
  DFF_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CK(clk), .Q(reg_in[135]) );
  DFF_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CK(clk), .Q(reg_in[134]) );
  DFF_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CK(clk), .Q(reg_in[133]) );
  DFF_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CK(clk), .Q(reg_in[132]) );
  DFF_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CK(clk), .Q(reg_in[131]) );
  DFF_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CK(clk), .Q(reg_in[130]) );
  DFF_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CK(clk), .Q(reg_in[129]) );
  DFF_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CK(clk), .Q(reg_in[128]) );
  DFF_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CK(clk), .Q(reg_in[127]) );
  DFF_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CK(clk), .Q(reg_in[126]) );
  DFF_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CK(clk), .Q(reg_in[125]) );
  DFF_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CK(clk), .Q(reg_in[124]) );
  DFF_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CK(clk), .Q(reg_in[123]) );
  DFF_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CK(clk), .Q(reg_in[122]) );
  DFF_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CK(clk), .Q(reg_in[121]) );
  DFF_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CK(clk), .Q(reg_in[120]) );
  DFF_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CK(clk), .Q(reg_in[119]) );
  DFF_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CK(clk), .Q(reg_in[118]) );
  DFF_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CK(clk), .Q(reg_in[117]) );
  DFF_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CK(clk), .Q(reg_in[116]) );
  DFF_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CK(clk), .Q(reg_in[115]) );
  DFF_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CK(clk), .Q(reg_in[114]) );
  DFF_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CK(clk), .Q(reg_in[113]) );
  DFF_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CK(clk), .Q(reg_in[112]) );
  DFF_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CK(clk), .Q(reg_in[111]) );
  DFF_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CK(clk), .Q(reg_in[110]) );
  DFF_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CK(clk), .Q(reg_in[109]) );
  DFF_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CK(clk), .Q(reg_in[108]) );
  DFF_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CK(clk), .Q(reg_in[107]) );
  DFF_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CK(clk), .Q(reg_in[106]) );
  DFF_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CK(clk), .Q(reg_in[105]) );
  DFF_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CK(clk), .Q(reg_in[104]) );
  DFF_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CK(clk), .Q(reg_in[103]) );
  DFF_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CK(clk), .Q(reg_in[102]) );
  DFF_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CK(clk), .Q(reg_in[101]) );
  DFF_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CK(clk), .Q(reg_in[100]) );
  DFF_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CK(clk), .Q(reg_in[99]) );
  DFF_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CK(clk), .Q(reg_in[98]) );
  DFF_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CK(clk), .Q(reg_in[97]) );
  DFF_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CK(clk), .Q(reg_in[96]) );
  DFF_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CK(clk), .Q(reg_in[95]) );
  DFF_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CK(clk), .Q(reg_in[94]) );
  DFF_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CK(clk), .Q(reg_in[93]) );
  DFF_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CK(clk), .Q(reg_in[92]) );
  DFF_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CK(clk), .Q(reg_in[91]) );
  DFF_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CK(clk), .Q(reg_in[90]) );
  DFF_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CK(clk), .Q(reg_in[89]) );
  DFF_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CK(clk), .Q(reg_in[88]) );
  DFF_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CK(clk), .Q(reg_in[87]) );
  DFF_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CK(clk), .Q(reg_in[86]) );
  DFF_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CK(clk), .Q(reg_in[85]) );
  DFF_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CK(clk), .Q(reg_in[84]) );
  DFF_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CK(clk), .Q(reg_in[83]) );
  DFF_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CK(clk), .Q(reg_in[82]) );
  DFF_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CK(clk), .Q(reg_in[81]) );
  DFF_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CK(clk), .Q(reg_in[80]) );
  DFF_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CK(clk), .Q(reg_in[79]) );
  DFF_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CK(clk), .Q(reg_in[78]) );
  DFF_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CK(clk), .Q(reg_in[77]) );
  DFF_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CK(clk), .Q(reg_in[76]) );
  DFF_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CK(clk), .Q(reg_in[75]) );
  DFF_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CK(clk), .Q(reg_in[74]) );
  DFF_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CK(clk), .Q(reg_in[73]) );
  DFF_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CK(clk), .Q(reg_in[72]) );
  DFF_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CK(clk), .Q(reg_in[71]) );
  DFF_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CK(clk), .Q(reg_in[70]) );
  DFF_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CK(clk), .Q(reg_in[69]) );
  DFF_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CK(clk), .Q(reg_in[68]) );
  DFF_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CK(clk), .Q(reg_in[67]) );
  DFF_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CK(clk), .Q(reg_in[66]) );
  DFF_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CK(clk), .Q(reg_in[65]) );
  DFF_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CK(clk), .Q(reg_in[64]) );
  DFF_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CK(clk), .Q(reg_in[63]) );
  DFF_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CK(clk), .Q(reg_in[62]) );
  DFF_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CK(clk), .Q(reg_in[61]) );
  DFF_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CK(clk), .Q(reg_in[60]) );
  DFF_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CK(clk), .Q(reg_in[59]) );
  DFF_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CK(clk), .Q(reg_in[58]) );
  DFF_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CK(clk), .Q(reg_in[57]) );
  DFF_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CK(clk), .Q(reg_in[56]) );
  DFF_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CK(clk), .Q(reg_in[55]) );
  DFF_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CK(clk), .Q(reg_in[54]) );
  DFF_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CK(clk), .Q(reg_in[53]) );
  DFF_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CK(clk), .Q(reg_in[52]) );
  DFF_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CK(clk), .Q(reg_in[51]) );
  DFF_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CK(clk), .Q(reg_in[50]) );
  DFF_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CK(clk), .Q(reg_in[49]) );
  DFF_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CK(clk), .Q(reg_in[48]) );
  DFF_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CK(clk), .Q(reg_in[47]) );
  DFF_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CK(clk), .Q(reg_in[46]) );
  DFF_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CK(clk), .Q(reg_in[45]) );
  DFF_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CK(clk), .Q(reg_in[44]) );
  DFF_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CK(clk), .Q(reg_in[43]) );
  DFF_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CK(clk), .Q(reg_in[42]) );
  DFF_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CK(clk), .Q(reg_in[41]) );
  DFF_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CK(clk), .Q(reg_in[40]) );
  DFF_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CK(clk), .Q(reg_in[39]) );
  DFF_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CK(clk), .Q(reg_in[38]) );
  DFF_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CK(clk), .Q(reg_in[37]) );
  DFF_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CK(clk), .Q(reg_in[36]) );
  DFF_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CK(clk), .Q(reg_in[35]) );
  DFF_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CK(clk), .Q(reg_in[34]) );
  DFF_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CK(clk), .Q(reg_in[33]) );
  DFF_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CK(clk), .Q(reg_in[32]) );
  DFF_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CK(clk), .Q(reg_in[31]) );
  DFF_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CK(clk), .Q(reg_in[30]) );
  DFF_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CK(clk), .Q(reg_in[29]) );
  DFF_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CK(clk), .Q(reg_in[28]) );
  DFF_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CK(clk), .Q(reg_in[27]) );
  DFF_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CK(clk), .Q(reg_in[26]) );
  DFF_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CK(clk), .Q(reg_in[25]) );
  DFF_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CK(clk), .Q(reg_in[24]) );
  DFF_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CK(clk), .Q(reg_in[23]) );
  DFF_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CK(clk), .Q(reg_in[22]) );
  DFF_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CK(clk), .Q(reg_in[21]) );
  DFF_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CK(clk), .Q(reg_in[20]) );
  DFF_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CK(clk), .Q(reg_in[19]) );
  DFF_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CK(clk), .Q(reg_in[18]) );
  DFF_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CK(clk), .Q(reg_in[17]) );
  DFF_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CK(clk), .Q(reg_in[16]) );
  DFF_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CK(clk), .Q(reg_in[15]) );
  DFF_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CK(clk), .Q(reg_in[14]) );
  DFF_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CK(clk), .Q(reg_in[13]) );
  DFF_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CK(clk), .Q(reg_in[12]) );
  DFF_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CK(clk), .Q(reg_in[11]) );
  DFF_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CK(clk), .Q(reg_in[10]) );
  DFF_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CK(clk), .Q(reg_in[9]) );
  DFF_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CK(clk), .Q(reg_in[8]) );
  DFF_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CK(clk), .Q(reg_in[7]) );
  DFF_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CK(clk), .Q(reg_in[6]) );
  DFF_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CK(clk), .Q(reg_in[5]) );
  DFF_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CK(clk), .Q(reg_in[4]) );
  DFF_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CK(clk), .Q(reg_in[3]) );
  DFF_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CK(clk), .Q(reg_in[2]) );
  DFF_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CK(clk), .Q(reg_in[1]) );
  DFF_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CK(clk), .Q(reg_in[0]) );
  DFF_X1 \reg_key_reg[191]  ( .D(Key[191]), .CK(clk), .Q(reg_key[191]) );
  DFF_X1 \reg_key_reg[190]  ( .D(Key[190]), .CK(clk), .Q(reg_key[190]) );
  DFF_X1 \reg_key_reg[189]  ( .D(Key[189]), .CK(clk), .Q(reg_key[189]) );
  DFF_X1 \reg_key_reg[188]  ( .D(Key[188]), .CK(clk), .Q(reg_key[188]) );
  DFF_X1 \reg_key_reg[187]  ( .D(Key[187]), .CK(clk), .Q(reg_key[187]) );
  DFF_X1 \reg_key_reg[186]  ( .D(Key[186]), .CK(clk), .Q(reg_key[186]) );
  DFF_X1 \reg_key_reg[185]  ( .D(Key[185]), .CK(clk), .Q(reg_key[185]) );
  DFF_X1 \reg_key_reg[184]  ( .D(Key[184]), .CK(clk), .Q(reg_key[184]) );
  DFF_X1 \reg_key_reg[183]  ( .D(Key[183]), .CK(clk), .Q(reg_key[183]) );
  DFF_X1 \reg_key_reg[182]  ( .D(Key[182]), .CK(clk), .Q(reg_key[182]) );
  DFF_X1 \reg_key_reg[181]  ( .D(Key[181]), .CK(clk), .Q(reg_key[181]) );
  DFF_X1 \reg_key_reg[180]  ( .D(Key[180]), .CK(clk), .Q(reg_key[180]) );
  DFF_X1 \reg_key_reg[179]  ( .D(Key[179]), .CK(clk), .Q(reg_key[179]) );
  DFF_X1 \reg_key_reg[178]  ( .D(Key[178]), .CK(clk), .Q(reg_key[178]) );
  DFF_X1 \reg_key_reg[177]  ( .D(Key[177]), .CK(clk), .Q(reg_key[177]) );
  DFF_X1 \reg_key_reg[176]  ( .D(Key[176]), .CK(clk), .Q(reg_key[176]) );
  DFF_X1 \reg_key_reg[175]  ( .D(Key[175]), .CK(clk), .Q(reg_key[175]) );
  DFF_X1 \reg_key_reg[174]  ( .D(Key[174]), .CK(clk), .Q(reg_key[174]) );
  DFF_X1 \reg_key_reg[173]  ( .D(Key[173]), .CK(clk), .Q(reg_key[173]) );
  DFF_X1 \reg_key_reg[172]  ( .D(Key[172]), .CK(clk), .Q(reg_key[172]) );
  DFF_X1 \reg_key_reg[171]  ( .D(Key[171]), .CK(clk), .Q(reg_key[171]) );
  DFF_X1 \reg_key_reg[170]  ( .D(Key[170]), .CK(clk), .Q(reg_key[170]) );
  DFF_X1 \reg_key_reg[169]  ( .D(Key[169]), .CK(clk), .Q(reg_key[169]) );
  DFF_X1 \reg_key_reg[168]  ( .D(Key[168]), .CK(clk), .Q(reg_key[168]) );
  DFF_X1 \reg_key_reg[167]  ( .D(Key[167]), .CK(clk), .Q(reg_key[167]) );
  DFF_X1 \reg_key_reg[166]  ( .D(Key[166]), .CK(clk), .Q(reg_key[166]) );
  DFF_X1 \reg_key_reg[165]  ( .D(Key[165]), .CK(clk), .Q(reg_key[165]) );
  DFF_X1 \reg_key_reg[164]  ( .D(Key[164]), .CK(clk), .Q(reg_key[164]) );
  DFF_X1 \reg_key_reg[163]  ( .D(Key[163]), .CK(clk), .Q(reg_key[163]) );
  DFF_X1 \reg_key_reg[162]  ( .D(Key[162]), .CK(clk), .Q(reg_key[162]) );
  DFF_X1 \reg_key_reg[161]  ( .D(Key[161]), .CK(clk), .Q(reg_key[161]) );
  DFF_X1 \reg_key_reg[160]  ( .D(Key[160]), .CK(clk), .Q(reg_key[160]) );
  DFF_X1 \reg_key_reg[159]  ( .D(Key[159]), .CK(clk), .Q(reg_key[159]) );
  DFF_X1 \reg_key_reg[158]  ( .D(Key[158]), .CK(clk), .Q(reg_key[158]) );
  DFF_X1 \reg_key_reg[157]  ( .D(Key[157]), .CK(clk), .Q(reg_key[157]) );
  DFF_X1 \reg_key_reg[156]  ( .D(Key[156]), .CK(clk), .Q(reg_key[156]) );
  DFF_X1 \reg_key_reg[155]  ( .D(Key[155]), .CK(clk), .Q(reg_key[155]) );
  DFF_X1 \reg_key_reg[154]  ( .D(Key[154]), .CK(clk), .Q(reg_key[154]) );
  DFF_X1 \reg_key_reg[153]  ( .D(Key[153]), .CK(clk), .Q(reg_key[153]) );
  DFF_X1 \reg_key_reg[152]  ( .D(Key[152]), .CK(clk), .Q(reg_key[152]) );
  DFF_X1 \reg_key_reg[151]  ( .D(Key[151]), .CK(clk), .Q(reg_key[151]) );
  DFF_X1 \reg_key_reg[150]  ( .D(Key[150]), .CK(clk), .Q(reg_key[150]) );
  DFF_X1 \reg_key_reg[149]  ( .D(Key[149]), .CK(clk), .Q(reg_key[149]) );
  DFF_X1 \reg_key_reg[148]  ( .D(Key[148]), .CK(clk), .Q(reg_key[148]) );
  DFF_X1 \reg_key_reg[147]  ( .D(Key[147]), .CK(clk), .Q(reg_key[147]) );
  DFF_X1 \reg_key_reg[146]  ( .D(Key[146]), .CK(clk), .Q(reg_key[146]) );
  DFF_X1 \reg_key_reg[145]  ( .D(Key[145]), .CK(clk), .Q(reg_key[145]) );
  DFF_X1 \reg_key_reg[144]  ( .D(Key[144]), .CK(clk), .Q(reg_key[144]) );
  DFF_X1 \reg_key_reg[143]  ( .D(Key[143]), .CK(clk), .Q(reg_key[143]) );
  DFF_X1 \reg_key_reg[142]  ( .D(Key[142]), .CK(clk), .Q(reg_key[142]) );
  DFF_X1 \reg_key_reg[141]  ( .D(Key[141]), .CK(clk), .Q(reg_key[141]) );
  DFF_X1 \reg_key_reg[140]  ( .D(Key[140]), .CK(clk), .Q(reg_key[140]) );
  DFF_X1 \reg_key_reg[139]  ( .D(Key[139]), .CK(clk), .Q(reg_key[139]) );
  DFF_X1 \reg_key_reg[138]  ( .D(Key[138]), .CK(clk), .Q(reg_key[138]) );
  DFF_X1 \reg_key_reg[137]  ( .D(Key[137]), .CK(clk), .Q(reg_key[137]) );
  DFF_X1 \reg_key_reg[136]  ( .D(Key[136]), .CK(clk), .Q(reg_key[136]) );
  DFF_X1 \reg_key_reg[135]  ( .D(Key[135]), .CK(clk), .Q(reg_key[135]) );
  DFF_X1 \reg_key_reg[134]  ( .D(Key[134]), .CK(clk), .Q(reg_key[134]) );
  DFF_X1 \reg_key_reg[133]  ( .D(Key[133]), .CK(clk), .Q(reg_key[133]) );
  DFF_X1 \reg_key_reg[132]  ( .D(Key[132]), .CK(clk), .Q(reg_key[132]) );
  DFF_X1 \reg_key_reg[131]  ( .D(Key[131]), .CK(clk), .Q(reg_key[131]) );
  DFF_X1 \reg_key_reg[130]  ( .D(Key[130]), .CK(clk), .Q(reg_key[130]) );
  DFF_X1 \reg_key_reg[129]  ( .D(Key[129]), .CK(clk), .Q(reg_key[129]) );
  DFF_X1 \reg_key_reg[128]  ( .D(Key[128]), .CK(clk), .Q(reg_key[128]) );
  DFF_X1 \reg_key_reg[127]  ( .D(Key[127]), .CK(clk), .Q(reg_key[127]) );
  DFF_X1 \reg_key_reg[126]  ( .D(Key[126]), .CK(clk), .Q(reg_key[126]) );
  DFF_X1 \reg_key_reg[125]  ( .D(Key[125]), .CK(clk), .Q(reg_key[125]) );
  DFF_X1 \reg_key_reg[124]  ( .D(Key[124]), .CK(clk), .Q(reg_key[124]) );
  DFF_X1 \reg_key_reg[123]  ( .D(Key[123]), .CK(clk), .Q(reg_key[123]) );
  DFF_X1 \reg_key_reg[122]  ( .D(Key[122]), .CK(clk), .Q(reg_key[122]) );
  DFF_X1 \reg_key_reg[121]  ( .D(Key[121]), .CK(clk), .Q(reg_key[121]) );
  DFF_X1 \reg_key_reg[120]  ( .D(Key[120]), .CK(clk), .Q(reg_key[120]) );
  DFF_X1 \reg_key_reg[119]  ( .D(Key[119]), .CK(clk), .Q(reg_key[119]) );
  DFF_X1 \reg_key_reg[118]  ( .D(Key[118]), .CK(clk), .Q(reg_key[118]) );
  DFF_X1 \reg_key_reg[117]  ( .D(Key[117]), .CK(clk), .Q(reg_key[117]) );
  DFF_X1 \reg_key_reg[116]  ( .D(Key[116]), .CK(clk), .Q(reg_key[116]) );
  DFF_X1 \reg_key_reg[115]  ( .D(Key[115]), .CK(clk), .Q(reg_key[115]) );
  DFF_X1 \reg_key_reg[114]  ( .D(Key[114]), .CK(clk), .Q(reg_key[114]) );
  DFF_X1 \reg_key_reg[113]  ( .D(Key[113]), .CK(clk), .Q(reg_key[113]) );
  DFF_X1 \reg_key_reg[112]  ( .D(Key[112]), .CK(clk), .Q(reg_key[112]) );
  DFF_X1 \reg_key_reg[111]  ( .D(Key[111]), .CK(clk), .Q(reg_key[111]) );
  DFF_X1 \reg_key_reg[110]  ( .D(Key[110]), .CK(clk), .Q(reg_key[110]) );
  DFF_X1 \reg_key_reg[109]  ( .D(Key[109]), .CK(clk), .Q(reg_key[109]) );
  DFF_X1 \reg_key_reg[108]  ( .D(Key[108]), .CK(clk), .Q(reg_key[108]) );
  DFF_X1 \reg_key_reg[107]  ( .D(Key[107]), .CK(clk), .Q(reg_key[107]) );
  DFF_X1 \reg_key_reg[106]  ( .D(Key[106]), .CK(clk), .Q(reg_key[106]) );
  DFF_X1 \reg_key_reg[105]  ( .D(Key[105]), .CK(clk), .Q(reg_key[105]) );
  DFF_X1 \reg_key_reg[104]  ( .D(Key[104]), .CK(clk), .Q(reg_key[104]) );
  DFF_X1 \reg_key_reg[103]  ( .D(Key[103]), .CK(clk), .Q(reg_key[103]) );
  DFF_X1 \reg_key_reg[102]  ( .D(Key[102]), .CK(clk), .Q(reg_key[102]) );
  DFF_X1 \reg_key_reg[101]  ( .D(Key[101]), .CK(clk), .Q(reg_key[101]) );
  DFF_X1 \reg_key_reg[100]  ( .D(Key[100]), .CK(clk), .Q(reg_key[100]) );
  DFF_X1 \reg_key_reg[99]  ( .D(Key[99]), .CK(clk), .Q(reg_key[99]) );
  DFF_X1 \reg_key_reg[98]  ( .D(Key[98]), .CK(clk), .Q(reg_key[98]) );
  DFF_X1 \reg_key_reg[97]  ( .D(Key[97]), .CK(clk), .Q(reg_key[97]) );
  DFF_X1 \reg_key_reg[96]  ( .D(Key[96]), .CK(clk), .Q(reg_key[96]) );
  DFF_X1 \reg_key_reg[95]  ( .D(Key[95]), .CK(clk), .Q(reg_key[95]) );
  DFF_X1 \reg_key_reg[94]  ( .D(Key[94]), .CK(clk), .Q(reg_key[94]) );
  DFF_X1 \reg_key_reg[93]  ( .D(Key[93]), .CK(clk), .Q(reg_key[93]) );
  DFF_X1 \reg_key_reg[92]  ( .D(Key[92]), .CK(clk), .Q(reg_key[92]) );
  DFF_X1 \reg_key_reg[91]  ( .D(Key[91]), .CK(clk), .Q(reg_key[91]) );
  DFF_X1 \reg_key_reg[90]  ( .D(Key[90]), .CK(clk), .Q(reg_key[90]) );
  DFF_X1 \reg_key_reg[89]  ( .D(Key[89]), .CK(clk), .Q(reg_key[89]) );
  DFF_X1 \reg_key_reg[88]  ( .D(Key[88]), .CK(clk), .Q(reg_key[88]) );
  DFF_X1 \reg_key_reg[87]  ( .D(Key[87]), .CK(clk), .Q(reg_key[87]) );
  DFF_X1 \reg_key_reg[86]  ( .D(Key[86]), .CK(clk), .Q(reg_key[86]) );
  DFF_X1 \reg_key_reg[85]  ( .D(Key[85]), .CK(clk), .Q(reg_key[85]) );
  DFF_X1 \reg_key_reg[84]  ( .D(Key[84]), .CK(clk), .Q(reg_key[84]) );
  DFF_X1 \reg_key_reg[83]  ( .D(Key[83]), .CK(clk), .Q(reg_key[83]) );
  DFF_X1 \reg_key_reg[82]  ( .D(Key[82]), .CK(clk), .Q(reg_key[82]) );
  DFF_X1 \reg_key_reg[81]  ( .D(Key[81]), .CK(clk), .Q(reg_key[81]) );
  DFF_X1 \reg_key_reg[80]  ( .D(Key[80]), .CK(clk), .Q(reg_key[80]) );
  DFF_X1 \reg_key_reg[79]  ( .D(Key[79]), .CK(clk), .Q(reg_key[79]) );
  DFF_X1 \reg_key_reg[78]  ( .D(Key[78]), .CK(clk), .Q(reg_key[78]) );
  DFF_X1 \reg_key_reg[77]  ( .D(Key[77]), .CK(clk), .Q(reg_key[77]) );
  DFF_X1 \reg_key_reg[76]  ( .D(Key[76]), .CK(clk), .Q(reg_key[76]) );
  DFF_X1 \reg_key_reg[75]  ( .D(Key[75]), .CK(clk), .Q(reg_key[75]) );
  DFF_X1 \reg_key_reg[74]  ( .D(Key[74]), .CK(clk), .Q(reg_key[74]) );
  DFF_X1 \reg_key_reg[73]  ( .D(Key[73]), .CK(clk), .Q(reg_key[73]) );
  DFF_X1 \reg_key_reg[72]  ( .D(Key[72]), .CK(clk), .Q(reg_key[72]) );
  DFF_X1 \reg_key_reg[71]  ( .D(Key[71]), .CK(clk), .Q(reg_key[71]) );
  DFF_X1 \reg_key_reg[70]  ( .D(Key[70]), .CK(clk), .Q(reg_key[70]) );
  DFF_X1 \reg_key_reg[69]  ( .D(Key[69]), .CK(clk), .Q(reg_key[69]) );
  DFF_X1 \reg_key_reg[68]  ( .D(Key[68]), .CK(clk), .Q(reg_key[68]) );
  DFF_X1 \reg_key_reg[67]  ( .D(Key[67]), .CK(clk), .Q(reg_key[67]) );
  DFF_X1 \reg_key_reg[66]  ( .D(Key[66]), .CK(clk), .Q(reg_key[66]) );
  DFF_X1 \reg_key_reg[65]  ( .D(Key[65]), .CK(clk), .Q(reg_key[65]) );
  DFF_X1 \reg_key_reg[64]  ( .D(Key[64]), .CK(clk), .Q(reg_key[64]) );
  DFF_X1 \reg_key_reg[63]  ( .D(Key[63]), .CK(clk), .Q(reg_key[63]) );
  DFF_X1 \reg_key_reg[62]  ( .D(Key[62]), .CK(clk), .Q(reg_key[62]) );
  DFF_X1 \reg_key_reg[61]  ( .D(Key[61]), .CK(clk), .Q(reg_key[61]) );
  DFF_X1 \reg_key_reg[60]  ( .D(Key[60]), .CK(clk), .Q(reg_key[60]) );
  DFF_X1 \reg_key_reg[59]  ( .D(Key[59]), .CK(clk), .Q(reg_key[59]) );
  DFF_X1 \reg_key_reg[58]  ( .D(Key[58]), .CK(clk), .Q(reg_key[58]) );
  DFF_X1 \reg_key_reg[57]  ( .D(Key[57]), .CK(clk), .Q(reg_key[57]) );
  DFF_X1 \reg_key_reg[56]  ( .D(Key[56]), .CK(clk), .Q(reg_key[56]) );
  DFF_X1 \reg_key_reg[55]  ( .D(Key[55]), .CK(clk), .Q(reg_key[55]) );
  DFF_X1 \reg_key_reg[54]  ( .D(Key[54]), .CK(clk), .Q(reg_key[54]) );
  DFF_X1 \reg_key_reg[53]  ( .D(Key[53]), .CK(clk), .Q(reg_key[53]) );
  DFF_X1 \reg_key_reg[52]  ( .D(Key[52]), .CK(clk), .Q(reg_key[52]) );
  DFF_X1 \reg_key_reg[51]  ( .D(Key[51]), .CK(clk), .Q(reg_key[51]) );
  DFF_X1 \reg_key_reg[50]  ( .D(Key[50]), .CK(clk), .Q(reg_key[50]) );
  DFF_X1 \reg_key_reg[49]  ( .D(Key[49]), .CK(clk), .Q(reg_key[49]) );
  DFF_X1 \reg_key_reg[48]  ( .D(Key[48]), .CK(clk), .Q(reg_key[48]) );
  DFF_X1 \reg_key_reg[47]  ( .D(Key[47]), .CK(clk), .Q(reg_key[47]) );
  DFF_X1 \reg_key_reg[46]  ( .D(Key[46]), .CK(clk), .Q(reg_key[46]) );
  DFF_X1 \reg_key_reg[45]  ( .D(Key[45]), .CK(clk), .Q(reg_key[45]) );
  DFF_X1 \reg_key_reg[44]  ( .D(Key[44]), .CK(clk), .Q(reg_key[44]) );
  DFF_X1 \reg_key_reg[43]  ( .D(Key[43]), .CK(clk), .Q(reg_key[43]) );
  DFF_X1 \reg_key_reg[42]  ( .D(Key[42]), .CK(clk), .Q(reg_key[42]) );
  DFF_X1 \reg_key_reg[41]  ( .D(Key[41]), .CK(clk), .Q(reg_key[41]) );
  DFF_X1 \reg_key_reg[40]  ( .D(Key[40]), .CK(clk), .Q(reg_key[40]) );
  DFF_X1 \reg_key_reg[39]  ( .D(Key[39]), .CK(clk), .Q(reg_key[39]) );
  DFF_X1 \reg_key_reg[38]  ( .D(Key[38]), .CK(clk), .Q(reg_key[38]) );
  DFF_X1 \reg_key_reg[37]  ( .D(Key[37]), .CK(clk), .Q(reg_key[37]) );
  DFF_X1 \reg_key_reg[36]  ( .D(Key[36]), .CK(clk), .Q(reg_key[36]) );
  DFF_X1 \reg_key_reg[35]  ( .D(Key[35]), .CK(clk), .Q(reg_key[35]) );
  DFF_X1 \reg_key_reg[34]  ( .D(Key[34]), .CK(clk), .Q(reg_key[34]) );
  DFF_X1 \reg_key_reg[33]  ( .D(Key[33]), .CK(clk), .Q(reg_key[33]) );
  DFF_X1 \reg_key_reg[32]  ( .D(Key[32]), .CK(clk), .Q(reg_key[32]) );
  DFF_X1 \reg_key_reg[31]  ( .D(Key[31]), .CK(clk), .Q(reg_key[31]) );
  DFF_X1 \reg_key_reg[30]  ( .D(Key[30]), .CK(clk), .Q(reg_key[30]) );
  DFF_X1 \reg_key_reg[29]  ( .D(Key[29]), .CK(clk), .Q(reg_key[29]) );
  DFF_X1 \reg_key_reg[28]  ( .D(Key[28]), .CK(clk), .Q(reg_key[28]) );
  DFF_X1 \reg_key_reg[27]  ( .D(Key[27]), .CK(clk), .Q(reg_key[27]) );
  DFF_X1 \reg_key_reg[26]  ( .D(Key[26]), .CK(clk), .Q(reg_key[26]) );
  DFF_X1 \reg_key_reg[25]  ( .D(Key[25]), .CK(clk), .Q(reg_key[25]) );
  DFF_X1 \reg_key_reg[24]  ( .D(Key[24]), .CK(clk), .Q(reg_key[24]) );
  DFF_X1 \reg_key_reg[23]  ( .D(Key[23]), .CK(clk), .Q(reg_key[23]) );
  DFF_X1 \reg_key_reg[22]  ( .D(Key[22]), .CK(clk), .Q(reg_key[22]) );
  DFF_X1 \reg_key_reg[21]  ( .D(Key[21]), .CK(clk), .Q(reg_key[21]) );
  DFF_X1 \reg_key_reg[20]  ( .D(Key[20]), .CK(clk), .Q(reg_key[20]) );
  DFF_X1 \reg_key_reg[19]  ( .D(Key[19]), .CK(clk), .Q(reg_key[19]) );
  DFF_X1 \reg_key_reg[18]  ( .D(Key[18]), .CK(clk), .Q(reg_key[18]) );
  DFF_X1 \reg_key_reg[17]  ( .D(Key[17]), .CK(clk), .Q(reg_key[17]) );
  DFF_X1 \reg_key_reg[16]  ( .D(Key[16]), .CK(clk), .Q(reg_key[16]) );
  DFF_X1 \reg_key_reg[15]  ( .D(Key[15]), .CK(clk), .Q(reg_key[15]) );
  DFF_X1 \reg_key_reg[14]  ( .D(Key[14]), .CK(clk), .Q(reg_key[14]) );
  DFF_X1 \reg_key_reg[13]  ( .D(Key[13]), .CK(clk), .Q(reg_key[13]) );
  DFF_X1 \reg_key_reg[12]  ( .D(Key[12]), .CK(clk), .Q(reg_key[12]) );
  DFF_X1 \reg_key_reg[11]  ( .D(Key[11]), .CK(clk), .Q(reg_key[11]) );
  DFF_X1 \reg_key_reg[10]  ( .D(Key[10]), .CK(clk), .Q(reg_key[10]) );
  DFF_X1 \reg_key_reg[9]  ( .D(Key[9]), .CK(clk), .Q(reg_key[9]) );
  DFF_X1 \reg_key_reg[8]  ( .D(Key[8]), .CK(clk), .Q(reg_key[8]) );
  DFF_X1 \reg_key_reg[7]  ( .D(Key[7]), .CK(clk), .Q(reg_key[7]) );
  DFF_X1 \reg_key_reg[6]  ( .D(Key[6]), .CK(clk), .Q(reg_key[6]) );
  DFF_X1 \reg_key_reg[5]  ( .D(Key[5]), .CK(clk), .Q(reg_key[5]) );
  DFF_X1 \reg_key_reg[4]  ( .D(Key[4]), .CK(clk), .Q(reg_key[4]) );
  DFF_X1 \reg_key_reg[3]  ( .D(Key[3]), .CK(clk), .Q(reg_key[3]) );
  DFF_X1 \reg_key_reg[2]  ( .D(Key[2]), .CK(clk), .Q(reg_key[2]) );
  DFF_X1 \reg_key_reg[1]  ( .D(Key[1]), .CK(clk), .Q(reg_key[1]) );
  DFF_X1 \reg_key_reg[0]  ( .D(Key[0]), .CK(clk), .Q(reg_key[0]) );
  DFF_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CK(clk), .Q(
        Ciphertext[191]) );
  DFF_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CK(clk), .Q(
        Ciphertext[190]) );
  DFF_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CK(clk), .Q(
        Ciphertext[189]) );
  DFF_X1 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CK(clk), .Q(
        Ciphertext[188]) );
  DFF_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CK(clk), .Q(
        Ciphertext[187]) );
  DFF_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CK(clk), .Q(
        Ciphertext[186]) );
  DFF_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CK(clk), .Q(
        Ciphertext[185]) );
  DFF_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CK(clk), .Q(
        Ciphertext[184]) );
  DFF_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CK(clk), .Q(
        Ciphertext[183]) );
  DFF_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CK(clk), .Q(
        Ciphertext[182]) );
  DFF_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CK(clk), .Q(
        Ciphertext[181]) );
  DFF_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CK(clk), .Q(
        Ciphertext[180]) );
  DFF_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CK(clk), .Q(
        Ciphertext[179]) );
  DFF_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CK(clk), .Q(
        Ciphertext[178]) );
  DFF_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CK(clk), .Q(
        Ciphertext[177]) );
  DFF_X1 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CK(clk), .Q(
        Ciphertext[176]) );
  DFF_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CK(clk), .Q(
        Ciphertext[175]) );
  DFF_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CK(clk), .Q(
        Ciphertext[174]) );
  DFF_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CK(clk), .Q(
        Ciphertext[173]) );
  DFF_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CK(clk), .Q(
        Ciphertext[172]) );
  DFF_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CK(clk), .Q(
        Ciphertext[171]) );
  DFF_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CK(clk), .Q(
        Ciphertext[170]) );
  DFF_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CK(clk), .Q(
        Ciphertext[169]) );
  DFF_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CK(clk), .Q(
        Ciphertext[168]) );
  DFF_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CK(clk), .Q(
        Ciphertext[167]) );
  DFF_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CK(clk), .Q(
        Ciphertext[166]) );
  DFF_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CK(clk), .Q(
        Ciphertext[165]) );
  DFF_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CK(clk), .Q(
        Ciphertext[164]) );
  DFF_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CK(clk), .Q(
        Ciphertext[163]) );
  DFF_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CK(clk), .Q(
        Ciphertext[162]) );
  DFF_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CK(clk), .Q(
        Ciphertext[161]) );
  DFF_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CK(clk), .Q(
        Ciphertext[160]) );
  DFF_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CK(clk), .Q(
        Ciphertext[159]) );
  DFF_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CK(clk), .Q(
        Ciphertext[158]) );
  DFF_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CK(clk), .Q(
        Ciphertext[157]) );
  DFF_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CK(clk), .Q(
        Ciphertext[156]) );
  DFF_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CK(clk), .Q(
        Ciphertext[155]) );
  DFF_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CK(clk), .Q(
        Ciphertext[154]) );
  DFF_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CK(clk), .Q(
        Ciphertext[153]) );
  DFF_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CK(clk), .Q(
        Ciphertext[152]) );
  DFF_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CK(clk), .Q(
        Ciphertext[151]) );
  DFF_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CK(clk), .Q(
        Ciphertext[150]) );
  DFF_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CK(clk), .Q(
        Ciphertext[149]) );
  DFF_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CK(clk), .Q(
        Ciphertext[148]) );
  DFF_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CK(clk), .Q(
        Ciphertext[147]) );
  DFF_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CK(clk), .Q(
        Ciphertext[146]) );
  DFF_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CK(clk), .Q(
        Ciphertext[145]) );
  DFF_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CK(clk), .Q(
        Ciphertext[144]) );
  DFF_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CK(clk), .Q(
        Ciphertext[143]) );
  DFF_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CK(clk), .Q(
        Ciphertext[142]) );
  DFF_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CK(clk), .Q(
        Ciphertext[141]) );
  DFF_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CK(clk), .Q(
        Ciphertext[140]) );
  DFF_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CK(clk), .Q(
        Ciphertext[139]) );
  DFF_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CK(clk), .Q(
        Ciphertext[138]) );
  DFF_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CK(clk), .Q(
        Ciphertext[137]) );
  DFF_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CK(clk), .Q(
        Ciphertext[136]) );
  DFF_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CK(clk), .Q(
        Ciphertext[135]) );
  DFF_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CK(clk), .Q(
        Ciphertext[134]) );
  DFF_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CK(clk), .Q(
        Ciphertext[133]) );
  DFF_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CK(clk), .Q(
        Ciphertext[132]) );
  DFF_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CK(clk), .Q(
        Ciphertext[131]) );
  DFF_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CK(clk), .Q(
        Ciphertext[130]) );
  DFF_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CK(clk), .Q(
        Ciphertext[129]) );
  DFF_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CK(clk), .Q(
        Ciphertext[128]) );
  DFF_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CK(clk), .Q(
        Ciphertext[127]) );
  DFF_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CK(clk), .Q(
        Ciphertext[126]) );
  DFF_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CK(clk), .Q(
        Ciphertext[125]) );
  DFF_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CK(clk), .Q(
        Ciphertext[124]) );
  DFF_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CK(clk), .Q(
        Ciphertext[123]) );
  DFF_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CK(clk), .Q(
        Ciphertext[122]) );
  DFF_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CK(clk), .Q(
        Ciphertext[121]) );
  DFF_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CK(clk), .Q(
        Ciphertext[120]) );
  DFF_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CK(clk), .Q(
        Ciphertext[119]) );
  DFF_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CK(clk), .Q(
        Ciphertext[118]) );
  DFF_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CK(clk), .Q(
        Ciphertext[117]) );
  DFF_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CK(clk), .Q(
        Ciphertext[116]) );
  DFF_X1 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CK(clk), .Q(
        Ciphertext[115]) );
  DFF_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CK(clk), .Q(
        Ciphertext[114]) );
  DFF_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CK(clk), .Q(
        Ciphertext[113]) );
  DFF_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CK(clk), .Q(
        Ciphertext[112]) );
  DFF_X1 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CK(clk), .Q(
        Ciphertext[111]) );
  DFF_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CK(clk), .Q(
        Ciphertext[110]) );
  DFF_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CK(clk), .Q(
        Ciphertext[109]) );
  DFF_X1 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CK(clk), .Q(
        Ciphertext[108]) );
  DFF_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CK(clk), .Q(
        Ciphertext[107]) );
  DFF_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CK(clk), .Q(
        Ciphertext[106]) );
  DFF_X1 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CK(clk), .Q(
        Ciphertext[105]) );
  DFF_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CK(clk), .Q(
        Ciphertext[103]) );
  DFF_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CK(clk), .Q(
        Ciphertext[102]) );
  DFF_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CK(clk), .Q(
        Ciphertext[101]) );
  DFF_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CK(clk), .Q(
        Ciphertext[100]) );
  DFF_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CK(clk), .Q(Ciphertext[99])
         );
  DFF_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CK(clk), .Q(Ciphertext[98])
         );
  DFF_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CK(clk), .Q(Ciphertext[97])
         );
  DFF_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CK(clk), .Q(Ciphertext[96])
         );
  DFF_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CK(clk), .Q(Ciphertext[95])
         );
  DFF_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CK(clk), .Q(Ciphertext[94])
         );
  DFF_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CK(clk), .Q(Ciphertext[93])
         );
  DFF_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CK(clk), .Q(Ciphertext[92])
         );
  DFF_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CK(clk), .Q(Ciphertext[91])
         );
  DFF_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CK(clk), .Q(Ciphertext[90])
         );
  DFF_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CK(clk), .Q(Ciphertext[89])
         );
  DFF_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CK(clk), .Q(Ciphertext[88])
         );
  DFF_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CK(clk), .Q(Ciphertext[87])
         );
  DFF_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CK(clk), .Q(Ciphertext[86])
         );
  DFF_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CK(clk), .Q(Ciphertext[85])
         );
  DFF_X1 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CK(clk), .Q(Ciphertext[84])
         );
  DFF_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CK(clk), .Q(Ciphertext[83])
         );
  DFF_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CK(clk), .Q(Ciphertext[82])
         );
  DFF_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CK(clk), .Q(Ciphertext[81])
         );
  DFF_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CK(clk), .Q(Ciphertext[80])
         );
  DFF_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CK(clk), .Q(Ciphertext[79])
         );
  DFF_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CK(clk), .Q(Ciphertext[78])
         );
  DFF_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CK(clk), .Q(Ciphertext[77])
         );
  DFF_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CK(clk), .Q(Ciphertext[76])
         );
  DFF_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CK(clk), .Q(Ciphertext[75])
         );
  DFF_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CK(clk), .Q(Ciphertext[74])
         );
  DFF_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CK(clk), .Q(Ciphertext[73])
         );
  DFF_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CK(clk), .Q(Ciphertext[72])
         );
  DFF_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CK(clk), .Q(Ciphertext[71])
         );
  DFF_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CK(clk), .Q(Ciphertext[70])
         );
  DFF_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CK(clk), .Q(Ciphertext[69])
         );
  DFF_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CK(clk), .Q(Ciphertext[68])
         );
  DFF_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CK(clk), .Q(Ciphertext[67])
         );
  DFF_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CK(clk), .Q(Ciphertext[66])
         );
  DFF_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CK(clk), .Q(Ciphertext[65])
         );
  DFF_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CK(clk), .Q(Ciphertext[64])
         );
  DFF_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CK(clk), .Q(Ciphertext[63])
         );
  DFF_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CK(clk), .Q(Ciphertext[62])
         );
  DFF_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CK(clk), .Q(Ciphertext[61])
         );
  DFF_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CK(clk), .Q(Ciphertext[60])
         );
  DFF_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CK(clk), .Q(Ciphertext[59])
         );
  DFF_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CK(clk), .Q(Ciphertext[58])
         );
  DFF_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CK(clk), .Q(Ciphertext[57])
         );
  DFF_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CK(clk), .Q(Ciphertext[56])
         );
  DFF_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CK(clk), .Q(Ciphertext[55])
         );
  DFF_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CK(clk), .Q(Ciphertext[54])
         );
  DFF_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CK(clk), .Q(Ciphertext[53])
         );
  DFF_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CK(clk), .Q(Ciphertext[52])
         );
  DFF_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CK(clk), .Q(Ciphertext[51])
         );
  DFF_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CK(clk), .Q(Ciphertext[50])
         );
  DFF_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CK(clk), .Q(Ciphertext[49])
         );
  DFF_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CK(clk), .Q(Ciphertext[48])
         );
  DFF_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CK(clk), .Q(Ciphertext[47])
         );
  DFF_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CK(clk), .Q(Ciphertext[46])
         );
  DFF_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CK(clk), .Q(Ciphertext[45])
         );
  DFF_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CK(clk), .Q(Ciphertext[44])
         );
  DFF_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CK(clk), .Q(Ciphertext[43])
         );
  DFF_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CK(clk), .Q(Ciphertext[42])
         );
  DFF_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CK(clk), .Q(Ciphertext[40])
         );
  DFF_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CK(clk), .Q(Ciphertext[39])
         );
  DFF_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CK(clk), .Q(Ciphertext[38])
         );
  DFF_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CK(clk), .Q(Ciphertext[37])
         );
  DFF_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CK(clk), .Q(Ciphertext[36])
         );
  DFF_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CK(clk), .Q(Ciphertext[35])
         );
  DFF_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CK(clk), .Q(Ciphertext[34])
         );
  DFF_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CK(clk), .Q(Ciphertext[33])
         );
  DFF_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CK(clk), .Q(Ciphertext[32])
         );
  DFF_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CK(clk), .Q(Ciphertext[31])
         );
  DFF_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CK(clk), .Q(Ciphertext[30])
         );
  DFF_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CK(clk), .Q(Ciphertext[29])
         );
  DFF_X1 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CK(clk), .Q(Ciphertext[28])
         );
  DFF_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CK(clk), .Q(Ciphertext[27])
         );
  DFF_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CK(clk), .Q(Ciphertext[25])
         );
  DFF_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CK(clk), .Q(Ciphertext[24])
         );
  DFF_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CK(clk), .Q(Ciphertext[23])
         );
  DFF_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CK(clk), .Q(Ciphertext[22])
         );
  DFF_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CK(clk), .Q(Ciphertext[21])
         );
  DFF_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CK(clk), .Q(Ciphertext[20])
         );
  DFF_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CK(clk), .Q(Ciphertext[19])
         );
  DFF_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CK(clk), .Q(Ciphertext[18])
         );
  DFF_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CK(clk), .Q(Ciphertext[17])
         );
  DFF_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CK(clk), .Q(Ciphertext[15])
         );
  DFF_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CK(clk), .Q(Ciphertext[14])
         );
  DFF_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CK(clk), .Q(Ciphertext[13])
         );
  DFF_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CK(clk), .Q(Ciphertext[12])
         );
  DFF_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CK(clk), .Q(Ciphertext[11])
         );
  DFF_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CK(clk), .Q(Ciphertext[10])
         );
  DFF_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CK(clk), .Q(Ciphertext[9]) );
  DFF_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CK(clk), .Q(Ciphertext[8]) );
  DFF_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CK(clk), .Q(Ciphertext[7]) );
  DFF_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CK(clk), .Q(Ciphertext[6]) );
  DFF_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CK(clk), .Q(Ciphertext[5]) );
  DFF_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CK(clk), .Q(Ciphertext[4]) );
  DFF_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CK(clk), .Q(Ciphertext[3]) );
  DFF_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CK(clk), .Q(Ciphertext[2]) );
  DFF_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CK(clk), .Q(Ciphertext[1]) );
  DFF_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CK(clk), .Q(Ciphertext[0]) );
  SPEEDY_Rounds5_0 SPEEDY_instance ( .Plaintext(reg_in), .Key(reg_key), 
        .Ciphertext(reg_out) );
  DFFS_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CK(clk), .SN(1'b1), .Q(
        Ciphertext[16]) );
  DFF_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CK(clk), .Q(Ciphertext[26])
         );
  DFF_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CK(clk), .Q(Ciphertext[41])
         );
  DFF_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CK(clk), .Q(
        Ciphertext[104]) );
endmodule

