module SPEEDY_Rounds5_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   n1, n2, n3, n4, n6, n7, n8, n9, n11, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n40, n41, n44, n45, n46, n48, n49, n50, n52, n53, n55, n57,
         n60, n61, n63, n64, n65, n66, n67, n68, n70, n71, n73, n74, n75, n76,
         n78, n79, n80, n81, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93,
         n94, n95, n98, n99, n100, n102, n103, n104, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n117, n118, n119, n121, n122, n123,
         n125, n126, n128, n129, n130, n131, n132, n133, n134, n135, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n160, n163, n164, n169, n170, n176,
         n177, n178, n179, n180, n182, n190, n191, n192, n193, n195, n196,
         n197, n198, n199, n200, n201, n202, n204, n205, n207, n208, n209,
         n210, n212, n213, n214, n215, n216, n219, n220, n221, n222, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n273, n274, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n298, n299, n300, n301, n302, n303, n304, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n328, n329, n331,
         n332, n333, n334, n335, n336, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n382, n383, n385, n386, n387, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n409, n410, n411, n412, n415, n416, n417, n419, n420,
         n421, n422, n423, n424, n425, n427, n428, n429, n430, n431, n432,
         n434, n435, n436, n437, n439, n440, n443, n444, n445, n446, n447,
         n448, n449, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n469, n470, n471,
         n472, n473, n474, n475, n477, n478, n479, n480, n481, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n499, n502, n504, n505, n506, n507, n508, n509, n510, n512,
         n513, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n581,
         n582, n583, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n637, n638, n639,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n841, n842, n843, n844, n845, n846, n847,
         n848, n850, n851, n852, n854, n855, n856, n857, n859, n860, n861,
         n862, n864, n865, n868, n870, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n888, n889, n890,
         n891, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n946, n947, n948, n951, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1122,
         n1123, n1124, n1126, n1127, n1128, n1129, n1131, n1132, n1133, n1136,
         n1137, n1139, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1170, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1223, n1224, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1343, n1344,
         n1345, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1376, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1435, n1436, n1437, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1613, n1614, n1615, n1616, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1649, n1650, n1651,
         n1652, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1703, n1704,
         n1705, n1706, n1707, n1708, n1710, n1711, n1712, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1761, n1762, n1763, n1764, n1765, n1766, n1768, n1769,
         n1770, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1885, n1886, n1887, n1888, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2084, n2085,
         n2086, n2087, n2088, n2089, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2118,
         n2120, n2121, n2122, n2123, n2125, n2126, n2127, n2129, n2130, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2195, n2196, n2197, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2410, n2411, n2412, n2413, n2414, n2415,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2448,
         n2449, n2450, n2451, n2452, n2454, n2455, n2456, n2457, n2458, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2570, n2571, n2572, n2573, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2664, n2665, n2666, n2668, n2669, n2670, n2671, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2695, n2696, n2697,
         n2698, n2699, n2701, n2702, n2703, n2704, n2705, n2707, n2709, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2729, n2730, n2731, n2732,
         n2733, n2734, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2781, n2782, n2783, n2784, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2828, n2829,
         n2830, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2905, n2906, n2907, n2908, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2964, n2965, n2966,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3027, n3028, n3030,
         n3031, n3034, n3035, n3036, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3078, n3079, n3080, n3081, n3082, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3146, n3147, n3148, n3149, n3150, n3151,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3164, n3165, n3166, n3167, n3168, n3169, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3293, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3436,
         n3437, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3572,
         n3573, n3574, n3575, n3576, n3578, n3579, n3580, n3581, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3669, n3670, n3671, n3672, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3752, n3753, n3754, n3755, n3757, n3758, n3759, n3760, n3761,
         n3762, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3787, n3788, n3789, n3791, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3986, n3987, n3988, n3989, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4250, n4251, n4253, n4254, n4255, n4256, n4257, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4311, n4312, n4313,
         n4314, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4428,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4527, n4528, n4529, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4958, n4959, n4960, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5083,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5150, n5151, n5152, n5153, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5756, n5757, n5758, n5759, n5760, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5893, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5965, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7121, n7122, n7123, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7519, n7520, n7521, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7551, n7552, n7553, n7554, n7555, n7556, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7610, n7611, n7612,
         n7613, n7615, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7701, n7702, n7703, n7704, n7705, n7706, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7810, n7811, n7812,
         n7813, n7814, n7815, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n8000,
         n8001, n8002, n8003, n8004, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8230, n8232, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8577, n8578, n8579, n8580, n8581, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8676, n8677, n8678, n8679,
         n8680, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8754, n8755, n8756, n8757, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8939, n8940, n8941, n8942, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8993, n8994, n8995, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9204, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9255, n9256, n9257, n9258, n9260, n9261, n9262, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9834,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9891, n9892, n9893, n9894, n9895, n9898, n9899, n9900, n9901, n9902,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10625, n10626, n10627, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10964, n10965, n10966, n10967, n10968, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11191,
         n11192, n11193, n11194, n11195, n11196, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11512, n11513, n11514, n11515,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11553, n11554, n11555, n11556, n11557,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11791, n11792, n11793, n11794, n11795, n11796,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12147, n12148, n12149,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13004, n13005,
         n13006, n13007, n13008, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13778, n13779, n13780, n13781, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13797, n13798, n13799, n13800, n13801,
         n13802, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14047, n14049, n14050, n14051, n14052, n14053,
         n14054, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14171,
         n14172, n14173, n14174, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14203, n14204, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14287, n14288, n14289, n14290,
         n14291, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14367, n14368, n14369, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14501, n14502, n14504, n14505, n14506, n14507, n14508,
         n14509, n14511, n14512, n14513, n14514, n14515, n14516, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14596,
         n14597, n14598, n14599, n14600, n14601, n14603, n14604, n14606,
         n14607, n14608, n14609, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14648,
         n14649, n14651, n14652, n14653, n14654, n14655, n14656, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14673, n14674, n14675,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14726, n14727, n14728, n14729, n14730, n14731, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14826,
         n14827, n14828, n14829, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14911, n14913, n14914, n14915, n14916, n14917, n14918,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14997, n14998, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15453, n15454,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15485, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15640,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15733,
         n15734, n15735, n15736, n15737, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15793,
         n15794, n15796, n15797, n15798, n15800, n15801, n15802, n15803,
         n15804, n15805, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15919, n15920, n15921,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16159, n16160,
         n16161, n16163, n16164, n16165, n16166, n16167, n16168, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16251, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16579, n16580, n16581, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17135, n17136, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17238, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17656, n17658, n17659, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17705, n17706, n17707,
         n17708, n17709, n17710, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17793, n17794, n17795, n17796, n17797, n17799, n17800, n17802,
         n17803, n17804, n17805, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17822, n17823, n17824, n17825, n17826, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17860, n17861, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17872, n17873, n17874,
         n17875, n17876, n17878, n17879, n17881, n17882, n17883, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17925, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17943, n17944, n17945,
         n17946, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17985, n17986, n17987, n17988, n17989, n17991,
         n17992, n17993, n17994, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18054, n18055, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18168, n18169, n18170, n18171,
         n18172, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18240,
         n18241, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18311,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18364, n18365, n18366, n18367, n18368, n18369, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18389, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18448, n18449, n18450, n18451, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18575, n18576, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18644, n18645, n18646, n18647, n18648,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18735,
         n18736, n18737, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18749, n18750, n18751, n18752, n18753, n18754, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18822, n18823, n18825, n18826, n18827, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18901, n18902, n18903, n18904, n18905, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18946, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19100, n19101,
         n19102, n19103, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19288, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19324, n19325, n19326, n19327,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19418, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19472, n19474, n19475,
         n19476, n19485, n19488, n19490, n19492, n19496, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19557, n19558, n19559, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19672, n19673, n19674, n19675, n19676, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19697, n19698, n19699, n19700, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19713,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19794, n19796, n19797, n19798, n19799,
         n19802, n19803, n19804, n19805, n19806, n19807, n19809, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19871,
         n19872, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19927, n19928, n19929, n19930,
         n19931, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19962, n19963, n19964, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19977, n19978, n19979, n19980, n19983, n19984, n19985, n19986,
         n19988, n19989, n19990, n19992, n19993, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20076, n20077, n20079, n20080, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20117, n20119, n20120, n20121, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20239, n20240, n20241, n20242, n20243, n20244,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20281, n20282, n20283, n20284, n20285, n20286, n20288, n20290,
         n20291, n20292, n20293, n20294, n20295, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697;

  OR2_X1 U1 ( .A1(n19081), .A2(n19082), .ZN(n1) );
  OR2_X1 U2 ( .A1(n17858), .A2(n15), .ZN(n14) );
  AND2_X1 U8 ( .A1(n18948), .A2(n17812), .ZN(n20) );
  AND3_X1 U9 ( .A1(n3414), .A2(n3413), .A3(n15736), .ZN(n16988) );
  NAND2_X1 U11 ( .A1(n14372), .A2(n2720), .ZN(n16406) );
  OAI21_X1 U12 ( .B1(n15862), .B2(n15864), .A(n9), .ZN(n15173) );
  AND2_X1 U13 ( .A1(n15720), .A2(n15861), .ZN(n15328) );
  OR2_X1 U20 ( .A1(n13909), .A2(n14611), .ZN(n133) );
  OR2_X1 U21 ( .A1(n15121), .A2(n14520), .ZN(n14320) );
  BUF_X1 U22 ( .A(n12911), .Z(n14439) );
  OR2_X1 U28 ( .A1(n12606), .A2(n12237), .ZN(n12604) );
  OR2_X1 U29 ( .A1(n19833), .A2(n12479), .ZN(n6) );
  AND2_X1 U30 ( .A1(n12207), .A2(n12208), .ZN(n4) );
  BUF_X1 U32 ( .A(n10625), .Z(n11820) );
  INV_X1 U33 ( .A(n11598), .ZN(n11828) );
  AND2_X1 U34 ( .A1(n3630), .A2(n3629), .ZN(n122) );
  OR2_X1 U36 ( .A1(n10960), .A2(n20366), .ZN(n142) );
  INV_X1 U37 ( .A(n20366), .ZN(n143) );
  OR2_X1 U39 ( .A1(n11365), .A2(n10677), .ZN(n2765) );
  NOR2_X1 U41 ( .A1(n9570), .A2(n9569), .ZN(n9843) );
  OR2_X1 U43 ( .A1(n8547), .A2(n8546), .ZN(n10339) );
  OR2_X1 U45 ( .A1(n8946), .A2(n111), .ZN(n109) );
  AND3_X1 U47 ( .A1(n6957), .A2(n6956), .A3(n6955), .ZN(n9163) );
  INV_X1 U49 ( .A(n8127), .ZN(n9088) );
  OR2_X1 U53 ( .A1(n7507), .A2(n7508), .ZN(n1540) );
  XNOR2_X1 U54 ( .A(n6040), .B(n6732), .ZN(n8193) );
  XNOR2_X1 U55 ( .A(n7070), .B(n6947), .ZN(n6770) );
  CLKBUF_X1 U57 ( .A(Key[108]), .Z(n19027) );
  OAI21_X1 U59 ( .B1(n19790), .B2(n5929), .A(n41), .ZN(n5597) );
  OAI21_X1 U60 ( .B1(n6060), .B2(n6061), .A(n6059), .ZN(n6062) );
  OR2_X1 U61 ( .A1(n5349), .A2(n6150), .ZN(n6154) );
  INV_X1 U63 ( .A(n6042), .ZN(n135) );
  INV_X1 U64 ( .A(n5632), .ZN(n31) );
  INV_X1 U65 ( .A(n5215), .ZN(n32) );
  OR2_X1 U66 ( .A1(n4174), .A2(n4175), .ZN(n117) );
  AND2_X1 U69 ( .A1(n4819), .A2(n4820), .ZN(n5953) );
  NAND2_X1 U70 ( .A1(n2215), .A2(n2214), .ZN(n6017) );
  OR2_X1 U71 ( .A1(n5038), .A2(n303), .ZN(n1320) );
  AND2_X1 U72 ( .A1(n4524), .A2(n4342), .ZN(n87) );
  OR2_X1 U74 ( .A1(n176), .A2(n4685), .ZN(n4487) );
  AND2_X1 U76 ( .A1(n4313), .A2(n4601), .ZN(n29) );
  NAND2_X2 U78 ( .A1(n1186), .A2(n8561), .ZN(n10171) );
  OAI211_X1 U80 ( .C1(n11791), .C2(n14588), .A(n108), .B(n107), .ZN(n12658) );
  OAI21_X1 U83 ( .B1(n16679), .B2(n132), .A(n131), .ZN(n17675) );
  AND2_X1 U85 ( .A1(n19056), .A2(n19071), .ZN(n70) );
  OR2_X1 U88 ( .A1(n18935), .A2(n18936), .ZN(n7) );
  INV_X1 U90 ( .A(n19400), .ZN(n2) );
  OR2_X1 U92 ( .A1(n14010), .A2(n14406), .ZN(n35) );
  NOR3_X1 U93 ( .A1(n19292), .A2(n19283), .A3(n19282), .ZN(n19294) );
  OR2_X1 U94 ( .A1(n19290), .A2(n19304), .ZN(n138) );
  XNOR2_X1 U95 ( .A(n13834), .B(n13079), .ZN(n13389) );
  OAI22_X2 U96 ( .A1(n15472), .A2(n15471), .B1(n15470), .B2(n20503), .ZN(
        n17298) );
  INV_X1 U102 ( .A(n3516), .ZN(n139) );
  INV_X1 U103 ( .A(n701), .ZN(n14443) );
  XNOR2_X1 U106 ( .A(n6915), .B(n6916), .ZN(n8342) );
  AND2_X1 U107 ( .A1(n14601), .A2(n14250), .ZN(n14248) );
  OR2_X1 U110 ( .A1(n19402), .A2(n17650), .ZN(n81) );
  AND2_X1 U118 ( .A1(n19021), .A2(n19009), .ZN(n19004) );
  AND2_X1 U123 ( .A1(n6064), .A2(n5304), .ZN(n6061) );
  AOI21_X1 U125 ( .B1(n16638), .B2(n19353), .A(n16637), .ZN(n17935) );
  AND2_X1 U128 ( .A1(n17656), .A2(n19396), .ZN(n3) );
  INV_X1 U130 ( .A(n16306), .ZN(n17) );
  OR2_X1 U131 ( .A1(n19360), .A2(n17861), .ZN(n132) );
  NOR2_X1 U132 ( .A1(n15896), .A2(n15538), .ZN(n15890) );
  BUF_X1 U133 ( .A(n15896), .Z(n15402) );
  INV_X1 U134 ( .A(n14792), .ZN(n12627) );
  OR2_X1 U138 ( .A1(n15266), .A2(n15845), .ZN(n717) );
  NAND2_X2 U139 ( .A1(n14745), .A2(n14744), .ZN(n17294) );
  OAI21_X2 U143 ( .B1(n15231), .B2(n15449), .A(n15230), .ZN(n16861) );
  OR2_X1 U144 ( .A1(n8542), .A2(n9066), .ZN(n8860) );
  NAND2_X1 U146 ( .A1(n19080), .A2(n1), .ZN(n19084) );
  OAI21_X1 U147 ( .B1(n19511), .B2(n3), .A(n2), .ZN(n17658) );
  INV_X1 U149 ( .A(n17856), .ZN(n18) );
  OAI21_X1 U150 ( .B1(n1690), .B2(n8179), .A(n1851), .ZN(n8796) );
  NAND2_X1 U152 ( .A1(n12211), .A2(n4), .ZN(n12218) );
  OR2_X2 U156 ( .A1(n5538), .A2(n5537), .ZN(n5736) );
  AND2_X2 U158 ( .A1(n2750), .A2(n1002), .ZN(n2749) );
  NAND2_X1 U160 ( .A1(n11223), .A2(n6), .ZN(n12784) );
  NAND2_X1 U162 ( .A1(n3607), .A2(n3752), .ZN(n3658) );
  OR2_X1 U163 ( .A1(n352), .A2(n9563), .ZN(n2170) );
  NAND3_X1 U169 ( .A1(n18933), .A2(n18934), .A3(n7), .ZN(n2062) );
  NAND2_X1 U170 ( .A1(n8), .A2(n1912), .ZN(n8330) );
  NAND2_X1 U172 ( .A1(n4825), .A2(n4826), .ZN(n4831) );
  NAND2_X1 U174 ( .A1(n15862), .A2(n15327), .ZN(n9) );
  NAND2_X1 U176 ( .A1(n18923), .A2(n11), .ZN(n18925) );
  NAND2_X1 U177 ( .A1(n18920), .A2(n18921), .ZN(n11) );
  XNOR2_X2 U178 ( .A(n16910), .B(n16909), .ZN(n18221) );
  NAND2_X1 U182 ( .A1(n9527), .A2(n9530), .ZN(n9754) );
  NAND4_X2 U186 ( .A1(n5127), .A2(n5126), .A3(n5125), .A4(n1096), .ZN(n7179)
         );
  AND3_X2 U188 ( .A1(n1251), .A2(n1249), .A3(n1447), .ZN(n13577) );
  XNOR2_X2 U190 ( .A(n16100), .B(n16099), .ZN(n17891) );
  NAND2_X1 U194 ( .A1(n1487), .A2(n8832), .ZN(n2150) );
  INV_X1 U195 ( .A(n14285), .ZN(n15066) );
  OR2_X1 U199 ( .A1(n11664), .A2(n121), .ZN(n11666) );
  NOR2_X2 U200 ( .A1(n16), .A2(n14), .ZN(n19242) );
  NOR2_X1 U202 ( .A1(n18), .A2(n17), .ZN(n16) );
  NAND3_X1 U205 ( .A1(n5928), .A2(n6027), .A3(n5929), .ZN(n19) );
  INV_X2 U206 ( .A(n8129), .ZN(n9451) );
  MUX2_X2 U208 ( .A(n12086), .B(n12085), .S(n12416), .Z(n12906) );
  NAND2_X1 U209 ( .A1(n18047), .A2(n20), .ZN(n3544) );
  NAND2_X1 U210 ( .A1(n24), .A2(n21), .ZN(n7523) );
  NAND2_X1 U211 ( .A1(n23), .A2(n22), .ZN(n21) );
  INV_X1 U212 ( .A(n7922), .ZN(n22) );
  NAND2_X1 U213 ( .A1(n2176), .A2(n776), .ZN(n23) );
  NAND2_X1 U214 ( .A1(n7521), .A2(n7922), .ZN(n24) );
  NAND2_X1 U219 ( .A1(n15740), .A2(n26), .ZN(n25) );
  INV_X1 U220 ( .A(n15751), .ZN(n26) );
  NAND3_X1 U222 ( .A1(n12068), .A2(n12069), .A3(n1878), .ZN(n13710) );
  NAND2_X1 U227 ( .A1(n1938), .A2(n13892), .ZN(n1352) );
  INV_X1 U228 ( .A(n6117), .ZN(n6122) );
  NAND2_X1 U229 ( .A1(n5868), .A2(n6118), .ZN(n6117) );
  NAND2_X1 U230 ( .A1(n4354), .A2(n29), .ZN(n4314) );
  NAND2_X1 U233 ( .A1(n32), .A2(n31), .ZN(n30) );
  OAI21_X1 U235 ( .B1(n12032), .B2(n12033), .A(n12272), .ZN(n33) );
  NAND2_X1 U237 ( .A1(n703), .A2(n12185), .ZN(n1981) );
  AOI21_X1 U239 ( .B1(n11374), .B2(n11375), .A(n11373), .ZN(n12552) );
  OR2_X1 U241 ( .A1(n7965), .A2(n20490), .ZN(n8019) );
  AOI21_X1 U242 ( .B1(n34), .B2(n5530), .A(n5529), .ZN(n5536) );
  NAND2_X1 U243 ( .A1(n2940), .A2(n5569), .ZN(n34) );
  NAND2_X1 U248 ( .A1(n14007), .A2(n14236), .ZN(n36) );
  OR2_X1 U250 ( .A1(n11995), .A2(n11820), .ZN(n12327) );
  NAND3_X1 U251 ( .A1(n261), .A2(n9151), .A3(n2499), .ZN(n391) );
  OAI21_X1 U254 ( .B1(n3028), .B2(n19989), .A(n679), .ZN(n18862) );
  NAND3_X1 U258 ( .A1(n15794), .A2(n15791), .A3(n859), .ZN(n2309) );
  NAND2_X1 U265 ( .A1(n14211), .A2(n14213), .ZN(n14084) );
  OR2_X1 U267 ( .A1(n11921), .A2(n11920), .ZN(n40) );
  NAND2_X1 U269 ( .A1(n19790), .A2(n6025), .ZN(n41) );
  OAI21_X1 U270 ( .B1(n8814), .B2(n8812), .A(n8810), .ZN(n44) );
  INV_X1 U271 ( .A(n9119), .ZN(n45) );
  NOR2_X1 U272 ( .A1(n14441), .A2(n20262), .ZN(n140) );
  OAI22_X1 U273 ( .A1(n11126), .A2(n19949), .B1(n10814), .B2(n2729), .ZN(
        n11128) );
  OAI21_X1 U274 ( .B1(n48), .B2(n15150), .A(n46), .ZN(n14922) );
  NAND2_X1 U275 ( .A1(n15713), .A2(n19514), .ZN(n46) );
  NAND2_X1 U277 ( .A1(n49), .A2(n20178), .ZN(n48) );
  INV_X1 U278 ( .A(n15712), .ZN(n49) );
  NAND2_X1 U286 ( .A1(n1764), .A2(n5114), .ZN(n4068) );
  AOI22_X1 U288 ( .A1(n3703), .A2(n2749), .B1(n19606), .B2(n8544), .ZN(n88) );
  NAND2_X1 U290 ( .A1(n52), .A2(n50), .ZN(n18071) );
  NAND2_X1 U291 ( .A1(n18069), .A2(n17091), .ZN(n50) );
  NAND2_X1 U292 ( .A1(n18068), .A2(n2516), .ZN(n52) );
  NAND3_X2 U294 ( .A1(n11123), .A2(n11122), .A3(n2033), .ZN(n12463) );
  XNOR2_X1 U295 ( .A(n13222), .B(n13724), .ZN(n13761) );
  AOI21_X1 U298 ( .B1(n53), .B2(n19891), .A(n15256), .ZN(n15000) );
  NAND2_X1 U299 ( .A1(n2223), .A2(n19931), .ZN(n53) );
  NAND2_X1 U302 ( .A1(n15201), .A2(n3431), .ZN(n55) );
  NAND2_X1 U304 ( .A1(n15200), .A2(n15495), .ZN(n57) );
  NAND2_X1 U307 ( .A1(n1300), .A2(n1299), .ZN(n1298) );
  NAND2_X1 U311 ( .A1(n14101), .A2(n14102), .ZN(n14106) );
  INV_X1 U312 ( .A(n7462), .ZN(n7461) );
  NAND2_X1 U313 ( .A1(n8061), .A2(n8060), .ZN(n7462) );
  NAND2_X1 U314 ( .A1(n16662), .A2(n1173), .ZN(n60) );
  AOI21_X1 U316 ( .B1(n4345), .B2(n4344), .A(n4516), .ZN(n61) );
  AND2_X1 U318 ( .A1(n19998), .A2(n11500), .ZN(n11082) );
  XNOR2_X2 U319 ( .A(n10556), .B(n10555), .ZN(n11500) );
  NAND2_X1 U321 ( .A1(n12126), .A2(n1508), .ZN(n11703) );
  NAND2_X1 U323 ( .A1(n2241), .A2(n2242), .ZN(n63) );
  AND2_X1 U324 ( .A1(n11256), .A2(n11253), .ZN(n10774) );
  NAND2_X1 U326 ( .A1(n81), .A2(n16291), .ZN(n16497) );
  AND2_X2 U328 ( .A1(n65), .A2(n64), .ZN(n13791) );
  NAND2_X1 U329 ( .A1(n1439), .A2(n1440), .ZN(n64) );
  NAND2_X1 U330 ( .A1(n12292), .A2(n12291), .ZN(n65) );
  NAND2_X1 U334 ( .A1(n19294), .A2(n20515), .ZN(n18166) );
  OAI21_X1 U337 ( .B1(n18269), .B2(n17766), .A(n100), .ZN(n16869) );
  NAND3_X2 U345 ( .A1(n2543), .A2(n8199), .A3(n1361), .ZN(n9217) );
  NAND3_X1 U347 ( .A1(n15782), .A2(n15686), .A3(n15687), .ZN(n93) );
  NAND2_X1 U351 ( .A1(n13802), .A2(n14148), .ZN(n67) );
  NAND2_X1 U352 ( .A1(n6035), .A2(n6037), .ZN(n86) );
  NAND3_X1 U354 ( .A1(n2311), .A2(n2005), .A3(n15678), .ZN(n2003) );
  OR2_X2 U355 ( .A1(n4973), .A2(n4972), .ZN(n6036) );
  XNOR2_X1 U356 ( .A(n15218), .B(n15219), .ZN(n17245) );
  XNOR2_X1 U358 ( .A(n68), .B(n7303), .ZN(n5759) );
  XNOR2_X1 U359 ( .A(n6942), .B(n5754), .ZN(n68) );
  XNOR2_X1 U360 ( .A(n6872), .B(n106), .ZN(n6874) );
  NAND2_X1 U361 ( .A1(n495), .A2(n497), .ZN(n6872) );
  NAND2_X1 U362 ( .A1(n71), .A2(n70), .ZN(n2362) );
  NAND2_X1 U367 ( .A1(n153), .A2(n4706), .ZN(n4453) );
  XNOR2_X1 U369 ( .A(n12681), .B(n12682), .ZN(n13937) );
  NAND2_X1 U370 ( .A1(n10688), .A2(n11411), .ZN(n11006) );
  OR2_X1 U375 ( .A1(n8733), .A2(n8736), .ZN(n8333) );
  NAND3_X1 U377 ( .A1(n15507), .A2(n1758), .A3(n15188), .ZN(n14937) );
  NAND2_X1 U383 ( .A1(n4846), .A2(n4839), .ZN(n4661) );
  NAND2_X1 U384 ( .A1(n164), .A2(n4657), .ZN(n4846) );
  AND2_X1 U386 ( .A1(n11952), .A2(n11598), .ZN(n9613) );
  NAND2_X1 U389 ( .A1(n3873), .A2(n1920), .ZN(n5798) );
  NAND3_X1 U390 ( .A1(n3896), .A2(n74), .A3(n4467), .ZN(n3895) );
  NAND2_X1 U391 ( .A1(n4117), .A2(n4114), .ZN(n74) );
  NAND2_X1 U393 ( .A1(n4916), .A2(n76), .ZN(n75) );
  NAND2_X1 U394 ( .A1(n4952), .A2(n4953), .ZN(n76) );
  NAND2_X1 U396 ( .A1(n4955), .A2(n4954), .ZN(n78) );
  AND2_X2 U401 ( .A1(n10666), .A2(n10665), .ZN(n12110) );
  AND2_X2 U403 ( .A1(n80), .A2(n79), .ZN(n10570) );
  NAND2_X1 U404 ( .A1(n8452), .A2(n19880), .ZN(n79) );
  NAND2_X1 U405 ( .A1(n8453), .A2(n8454), .ZN(n80) );
  OR2_X1 U406 ( .A1(n3948), .A2(n4541), .ZN(n4538) );
  BUF_X1 U407 ( .A(n4220), .Z(n4845) );
  NAND3_X1 U417 ( .A1(n626), .A2(n2003), .A3(n625), .ZN(n17444) );
  AND3_X2 U419 ( .A1(n1291), .A2(n2715), .A3(n1287), .ZN(n16973) );
  NAND3_X1 U424 ( .A1(n8916), .A2(n19518), .A3(n8917), .ZN(n8918) );
  XNOR2_X2 U432 ( .A(n5854), .B(n5853), .ZN(n8040) );
  NAND2_X1 U434 ( .A1(n11469), .A2(n927), .ZN(n10884) );
  NAND3_X1 U437 ( .A1(n3431), .A2(n15607), .A3(n16128), .ZN(n417) );
  NAND2_X1 U443 ( .A1(n2626), .A2(n19748), .ZN(n2439) );
  NAND2_X1 U444 ( .A1(n1034), .A2(n1033), .ZN(n2626) );
  AND2_X2 U446 ( .A1(n16018), .A2(n16017), .ZN(n17347) );
  NAND3_X1 U448 ( .A1(n8259), .A2(n8159), .A3(n6831), .ZN(n6847) );
  NAND2_X1 U452 ( .A1(n9309), .A2(n1751), .ZN(n9229) );
  NAND3_X2 U454 ( .A1(n8207), .A2(n2885), .A3(n8206), .ZN(n9114) );
  NAND2_X1 U457 ( .A1(n595), .A2(n596), .ZN(n594) );
  NAND2_X1 U458 ( .A1(n84), .A2(n83), .ZN(n10787) );
  NAND2_X1 U459 ( .A1(n11879), .A2(n10259), .ZN(n83) );
  NAND2_X1 U460 ( .A1(n10786), .A2(n85), .ZN(n84) );
  INV_X1 U461 ( .A(n10259), .ZN(n85) );
  NAND2_X1 U462 ( .A1(n10808), .A2(n11884), .ZN(n10786) );
  NAND3_X1 U464 ( .A1(n15685), .A2(n15779), .A3(n20362), .ZN(n15689) );
  NAND2_X1 U465 ( .A1(n9338), .A2(n9070), .ZN(n8699) );
  BUF_X1 U469 ( .A(n4233), .Z(n4499) );
  NAND2_X1 U473 ( .A1(n86), .A2(n5531), .ZN(n1708) );
  XNOR2_X1 U474 ( .A(n13808), .B(n12614), .ZN(n12626) );
  XNOR2_X1 U475 ( .A(n13376), .B(n13518), .ZN(n13808) );
  OR2_X2 U478 ( .A1(n12039), .A2(n11172), .ZN(n12282) );
  NAND2_X1 U481 ( .A1(n3925), .A2(n87), .ZN(n4189) );
  NAND2_X1 U483 ( .A1(n4595), .A2(n4596), .ZN(n6477) );
  INV_X1 U487 ( .A(n7961), .ZN(n90) );
  INV_X1 U488 ( .A(n7773), .ZN(n91) );
  NAND3_X1 U489 ( .A1(n7961), .A2(n7917), .A3(n1231), .ZN(n92) );
  XNOR2_X2 U493 ( .A(Key[145]), .B(Plaintext[145]), .ZN(n5010) );
  AOI22_X2 U494 ( .A1(n9274), .A2(n3618), .B1(n8649), .B2(n8449), .ZN(n10114)
         );
  NAND3_X1 U496 ( .A1(n94), .A2(n14433), .A3(n2811), .ZN(n14488) );
  NAND3_X1 U497 ( .A1(n14485), .A2(n14486), .A3(n14487), .ZN(n94) );
  NAND2_X1 U498 ( .A1(n5425), .A2(n5668), .ZN(n5674) );
  NOR2_X2 U500 ( .A1(n14805), .A2(n14804), .ZN(n15812) );
  NAND2_X1 U502 ( .A1(n95), .A2(n11114), .ZN(n1813) );
  NOR2_X1 U503 ( .A1(n1812), .A2(n11452), .ZN(n95) );
  NAND2_X1 U511 ( .A1(n9363), .A2(n8958), .ZN(n8965) );
  BUF_X1 U515 ( .A(n10685), .Z(n11271) );
  NAND2_X1 U517 ( .A1(n98), .A2(n8083), .ZN(n7558) );
  OAI21_X1 U518 ( .B1(n8230), .B2(n20107), .A(n8085), .ZN(n98) );
  NAND2_X1 U519 ( .A1(n10677), .A2(n11231), .ZN(n11235) );
  NAND2_X1 U525 ( .A1(n18269), .A2(n18275), .ZN(n100) );
  NAND2_X1 U528 ( .A1(n8592), .A2(n9358), .ZN(n9530) );
  NAND3_X1 U529 ( .A1(n647), .A2(n11547), .A3(n258), .ZN(n10764) );
  NAND3_X1 U532 ( .A1(n15831), .A2(n15642), .A3(n2223), .ZN(n15646) );
  NAND2_X1 U534 ( .A1(n8565), .A2(n8884), .ZN(n8471) );
  NAND2_X1 U536 ( .A1(n443), .A2(n444), .ZN(n102) );
  NAND3_X1 U537 ( .A1(n2600), .A2(n2598), .A3(n12543), .ZN(n11798) );
  OAI211_X1 U551 ( .C1(n1714), .C2(n1729), .A(n103), .B(n1727), .ZN(
        Ciphertext[10]) );
  NAND2_X1 U552 ( .A1(n1714), .A2(n1728), .ZN(n103) );
  OR2_X1 U553 ( .A1(n11717), .A2(n12279), .ZN(n12278) );
  NAND2_X1 U558 ( .A1(n15600), .A2(n15275), .ZN(n15277) );
  AOI21_X1 U560 ( .B1(n11447), .B2(n11448), .A(n11446), .ZN(n104) );
  NAND2_X1 U565 ( .A1(n19375), .A2(n19380), .ZN(n17236) );
  NAND2_X2 U566 ( .A1(n435), .A2(n15570), .ZN(n17014) );
  NAND2_X1 U569 ( .A1(n14809), .A2(n14813), .ZN(n107) );
  NAND2_X1 U570 ( .A1(n474), .A2(n239), .ZN(n108) );
  NAND2_X1 U571 ( .A1(n110), .A2(n109), .ZN(n8491) );
  NAND2_X1 U572 ( .A1(n8940), .A2(n8644), .ZN(n8946) );
  NAND2_X1 U573 ( .A1(n8489), .A2(n111), .ZN(n110) );
  INV_X1 U574 ( .A(n8947), .ZN(n111) );
  BUF_X1 U575 ( .A(n16639), .Z(n17219) );
  OAI21_X2 U577 ( .B1(n11301), .B2(n11398), .A(n11300), .ZN(n12399) );
  OAI211_X2 U578 ( .C1(n17450), .C2(n17946), .A(n2290), .B(n2289), .ZN(n18697)
         );
  NAND3_X1 U581 ( .A1(n12335), .A2(n12339), .A3(n11992), .ZN(n11971) );
  XNOR2_X1 U582 ( .A(n13600), .B(n112), .ZN(n13257) );
  INV_X1 U583 ( .A(n13255), .ZN(n112) );
  NAND2_X1 U587 ( .A1(n5630), .A2(n5631), .ZN(n5634) );
  INV_X1 U588 ( .A(n17882), .ZN(n113) );
  NOR2_X1 U589 ( .A1(n5635), .A2(n5636), .ZN(n6301) );
  NAND2_X1 U593 ( .A1(n20258), .A2(n18238), .ZN(n114) );
  OR3_X1 U594 ( .A1(n15081), .A2(n15422), .A3(n15531), .ZN(n14257) );
  XNOR2_X1 U595 ( .A(n6667), .B(n6666), .ZN(n6671) );
  INV_X1 U597 ( .A(n5752), .ZN(n5750) );
  NAND2_X1 U598 ( .A1(n5744), .A2(n5743), .ZN(n5752) );
  NAND2_X1 U603 ( .A1(n12488), .A2(n12811), .ZN(n11693) );
  OR2_X1 U606 ( .A1(n11283), .A2(n10693), .ZN(n11286) );
  NAND2_X1 U607 ( .A1(n118), .A2(n117), .ZN(n5649) );
  NAND2_X1 U608 ( .A1(n4172), .A2(n4171), .ZN(n118) );
  NAND3_X1 U612 ( .A1(n11185), .A2(n2948), .A3(n2949), .ZN(n12141) );
  NAND2_X1 U613 ( .A1(n8126), .A2(n9453), .ZN(n8127) );
  NAND2_X1 U616 ( .A1(n8597), .A2(n8928), .ZN(n8598) );
  OAI22_X1 U618 ( .A1(n17396), .A2(n18264), .B1(n17762), .B2(n18750), .ZN(
        n17397) );
  AOI22_X2 U619 ( .A1(n1223), .A2(n228), .B1(n15815), .B2(n15036), .ZN(n17358)
         );
  OAI211_X1 U620 ( .C1(n11439), .C2(n11116), .A(n11034), .B(n119), .ZN(n3160)
         );
  OR2_X1 U621 ( .A1(n11115), .A2(n11440), .ZN(n119) );
  NAND2_X1 U631 ( .A1(n122), .A2(n11990), .ZN(n121) );
  OR2_X2 U632 ( .A1(n775), .A2(n3901), .ZN(n5428) );
  NAND2_X2 U634 ( .A1(n3998), .A2(n3997), .ZN(n6067) );
  NAND2_X1 U635 ( .A1(n201), .A2(n12500), .ZN(n2016) );
  AND2_X2 U636 ( .A1(n3981), .A2(n3320), .ZN(n3319) );
  OR2_X1 U638 ( .A1(n14796), .A2(n13891), .ZN(n14213) );
  MUX2_X2 U642 ( .A(n14383), .B(n14382), .S(n14381), .Z(n15838) );
  NAND2_X1 U643 ( .A1(n8768), .A2(n8477), .ZN(n1470) );
  NAND2_X1 U644 ( .A1(n1672), .A2(n1671), .ZN(n8768) );
  XNOR2_X2 U646 ( .A(n12496), .B(n12495), .ZN(n14789) );
  NAND2_X1 U648 ( .A1(n12759), .A2(n123), .ZN(n1828) );
  NOR2_X1 U649 ( .A1(n2523), .A2(n12754), .ZN(n123) );
  NAND2_X1 U651 ( .A1(n4555), .A2(n20229), .ZN(n4731) );
  NAND2_X1 U654 ( .A1(n2056), .A2(n12595), .ZN(n125) );
  XNOR2_X2 U655 ( .A(n2264), .B(n11682), .ZN(n14813) );
  OAI21_X1 U659 ( .B1(n12008), .B2(n12009), .A(n126), .ZN(n11662) );
  AND2_X1 U664 ( .A1(n11539), .A2(n11168), .ZN(n11537) );
  OR2_X1 U666 ( .A1(n18697), .A2(n18702), .ZN(n18706) );
  NAND2_X1 U667 ( .A1(n12412), .A2(n12390), .ZN(n3082) );
  NAND2_X1 U668 ( .A1(n128), .A2(n4206), .ZN(n4209) );
  NAND2_X1 U669 ( .A1(n5003), .A2(n4750), .ZN(n128) );
  NAND2_X1 U670 ( .A1(n20168), .A2(n17501), .ZN(n17503) );
  BUF_X2 U671 ( .A(n5250), .Z(n5323) );
  NAND2_X1 U673 ( .A1(n1976), .A2(n1977), .ZN(n129) );
  NAND2_X1 U678 ( .A1(n3734), .A2(n12261), .ZN(n1045) );
  AND3_X2 U686 ( .A1(n7555), .A2(n7554), .A3(n7553), .ZN(n8961) );
  OAI211_X2 U695 ( .C1(n10944), .C2(n12048), .A(n10942), .B(n130), .ZN(n13058)
         );
  NAND3_X1 U696 ( .A1(n10944), .A2(n10934), .A3(n11647), .ZN(n130) );
  NAND3_X1 U697 ( .A1(n1213), .A2(n12337), .A3(n12338), .ZN(n12342) );
  NAND2_X1 U698 ( .A1(n4108), .A2(n567), .ZN(n3290) );
  AND2_X2 U703 ( .A1(n14391), .A2(n1021), .ZN(n1288) );
  NAND3_X1 U704 ( .A1(n8892), .A2(n8893), .A3(n9010), .ZN(n8894) );
  OR2_X2 U706 ( .A1(n13926), .A2(n13925), .ZN(n14935) );
  NAND2_X1 U709 ( .A1(n11926), .A2(n11683), .ZN(n12579) );
  NAND3_X2 U710 ( .A1(n11004), .A2(n411), .A3(n11003), .ZN(n11926) );
  NAND3_X1 U712 ( .A1(n1266), .A2(n1265), .A3(n15314), .ZN(n1129) );
  OAI21_X2 U713 ( .B1(n15383), .B2(n3621), .A(n2862), .ZN(n16840) );
  MUX2_X2 U714 ( .A(n14030), .B(n14029), .S(n20120), .Z(n15491) );
  NOR2_X1 U715 ( .A1(n5251), .A2(n5323), .ZN(n5392) );
  NAND2_X2 U719 ( .A1(n10470), .A2(n10471), .ZN(n11995) );
  XNOR2_X2 U726 ( .A(n4040), .B(Key[120]), .ZN(n4708) );
  NAND2_X1 U729 ( .A1(n17670), .A2(n19360), .ZN(n131) );
  NAND3_X2 U732 ( .A1(n14144), .A2(n14145), .A3(n133), .ZN(n15509) );
  OR2_X2 U733 ( .A1(n14774), .A2(n14773), .ZN(n16964) );
  OAI21_X1 U735 ( .B1(n6041), .B2(n135), .A(n134), .ZN(n5889) );
  NAND2_X1 U736 ( .A1(n6041), .A2(n1214), .ZN(n134) );
  XNOR2_X1 U741 ( .A(n137), .B(n1259), .ZN(Ciphertext[171]) );
  NAND2_X2 U744 ( .A1(n9270), .A2(n1157), .ZN(n10360) );
  NAND2_X1 U752 ( .A1(n2596), .A2(n4137), .ZN(n4139) );
  NAND3_X1 U755 ( .A1(n2773), .A2(n140), .A3(n139), .ZN(n564) );
  OAI211_X1 U759 ( .C1(n19090), .C2(n19089), .A(n141), .B(n19088), .ZN(n19091)
         );
  NAND2_X1 U760 ( .A1(n19086), .A2(n19109), .ZN(n141) );
  BUF_X1 U766 ( .A(n14952), .Z(n15803) );
  OAI211_X1 U767 ( .C1(n143), .C2(n3515), .A(n142), .B(n11142), .ZN(n1669) );
  NAND2_X1 U768 ( .A1(n273), .A2(n8014), .ZN(n7992) );
  AOI21_X2 U769 ( .B1(n144), .B2(n307), .A(n1000), .ZN(n16961) );
  NOR2_X1 U770 ( .A1(n14983), .A2(n15522), .ZN(n144) );
  NOR2_X1 U774 ( .A1(n8879), .A2(n9249), .ZN(n1618) );
  OR2_X1 U779 ( .A1(n6090), .A2(n5176), .ZN(n806) );
  OR2_X1 U780 ( .A1(n6090), .A2(n6087), .ZN(n1468) );
  OR3_X1 U782 ( .A1(n5997), .A2(n5434), .A3(n5704), .ZN(n5814) );
  OR2_X1 U783 ( .A1(n19980), .A2(n6007), .ZN(n6014) );
  INV_X1 U784 ( .A(n7421), .ZN(n585) );
  OR2_X1 U786 ( .A1(n20257), .A2(n5941), .ZN(n1834) );
  AND2_X1 U787 ( .A1(n8542), .A2(n9065), .ZN(n8544) );
  INV_X1 U789 ( .A(n2749), .ZN(n545) );
  XNOR2_X1 U790 ( .A(n694), .B(n10027), .ZN(n10319) );
  NOR2_X1 U792 ( .A1(n15495), .A2(n747), .ZN(n3425) );
  OAI21_X1 U793 ( .B1(n15574), .B2(n15365), .A(n15796), .ZN(n15366) );
  OAI21_X1 U794 ( .B1(n18094), .B2(n19774), .A(n424), .ZN(n17166) );
  AND2_X1 U795 ( .A1(n19935), .A2(n18650), .ZN(n18645) );
  OR2_X1 U796 ( .A1(n19456), .A2(n19459), .ZN(n810) );
  AND2_X1 U797 ( .A1(n5955), .A2(n6107), .ZN(n145) );
  AND2_X1 U798 ( .A1(n5780), .A2(n5778), .ZN(n146) );
  AND2_X2 U799 ( .A1(n7636), .A2(n1404), .ZN(n8602) );
  NAND4_X2 U800 ( .A1(n7107), .A2(n7104), .A3(n7105), .A4(n7106), .ZN(n8851)
         );
  AND2_X1 U803 ( .A1(n951), .A2(n20443), .ZN(n147) );
  NAND2_X2 U805 ( .A1(n2152), .A2(n2153), .ZN(n15573) );
  OR2_X1 U806 ( .A1(n14916), .A2(n15863), .ZN(n148) );
  NAND2_X2 U807 ( .A1(n12933), .A2(n2535), .ZN(n15380) );
  OR2_X1 U808 ( .A1(n15093), .A2(n15636), .ZN(n149) );
  OR2_X1 U810 ( .A1(n19708), .A2(n19163), .ZN(n150) );
  OR2_X1 U812 ( .A1(n19031), .A2(n20074), .ZN(n151) );
  AND3_X1 U813 ( .A1(n19775), .A2(n16453), .A3(n16452), .ZN(n152) );
  XNOR2_X1 U821 ( .A(Key[122]), .B(Plaintext[122]), .ZN(n5031) );
  XNOR2_X1 U830 ( .A(Key[177]), .B(Plaintext[177]), .ZN(n4638) );
  MUX2_X2 U842 ( .A(n8346), .B(n8345), .S(n8344), .Z(n9135) );
  XNOR2_X2 U846 ( .A(n6893), .B(n6892), .ZN(n8347) );
  XNOR2_X1 U856 ( .A(Key[69]), .B(Plaintext[69]), .ZN(n4656) );
  XNOR2_X2 U858 ( .A(Key[162]), .B(Plaintext[162]), .ZN(n4539) );
  OAI21_X2 U867 ( .B1(n5210), .B2(n861), .A(n5209), .ZN(n6854) );
  INV_X2 U872 ( .A(n5106), .ZN(n5102) );
  AND2_X2 U874 ( .A1(n1131), .A2(n1393), .ZN(n7345) );
  AND2_X2 U879 ( .A1(n1445), .A2(n4900), .ZN(n5682) );
  XNOR2_X2 U888 ( .A(n13140), .B(n13471), .ZN(n14667) );
  XNOR2_X2 U894 ( .A(Key[87]), .B(Plaintext[87]), .ZN(n5073) );
  XNOR2_X2 U901 ( .A(n13170), .B(n13171), .ZN(n14666) );
  OAI21_X2 U905 ( .B1(n3193), .B2(n12878), .A(n12881), .ZN(n15167) );
  AOI22_X1 U911 ( .A1(n4655), .A2(n4654), .B1(n4863), .B2(n4653), .ZN(n6167)
         );
  XNOR2_X1 U932 ( .A(n6885), .B(n6884), .ZN(n8349) );
  BUF_X1 U934 ( .A(n4686), .Z(n177) );
  BUF_X1 U935 ( .A(n4686), .Z(n178) );
  XNOR2_X1 U936 ( .A(Key[57]), .B(Plaintext[57]), .ZN(n4686) );
  OAI21_X2 U937 ( .B1(n5708), .B2(n4113), .A(n622), .ZN(n7390) );
  OR2_X1 U950 ( .A1(n7967), .A2(n278), .ZN(n7976) );
  XNOR2_X2 U951 ( .A(n3953), .B(Key[187]), .ZN(n4614) );
  NAND2_X2 U952 ( .A1(n6197), .A2(n6198), .ZN(n7031) );
  NAND2_X2 U954 ( .A1(n1983), .A2(n1982), .ZN(n7134) );
  AOI22_X2 U956 ( .A1(n17980), .A2(n18752), .B1(n17979), .B2(n17978), .ZN(
        n18682) );
  OAI21_X2 U960 ( .B1(n8575), .B2(n9059), .A(n8574), .ZN(n10186) );
  AOI21_X2 U962 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n10240) );
  XNOR2_X2 U963 ( .A(n3880), .B(Key[0]), .ZN(n4169) );
  XNOR2_X2 U975 ( .A(n2745), .B(n2744), .ZN(n10677) );
  OAI22_X2 U977 ( .A1(n11969), .A2(n11631), .B1(n11629), .B2(n11630), .ZN(
        n12986) );
  OAI21_X2 U978 ( .B1(n6074), .B2(n6075), .A(n6073), .ZN(n7391) );
  BUF_X1 U984 ( .A(n11325), .Z(n190) );
  NOR2_X1 U987 ( .A1(n18454), .A2(n20139), .ZN(n18469) );
  OAI21_X1 U989 ( .B1(n17679), .B2(n20514), .A(n17678), .ZN(n1205) );
  OAI21_X1 U991 ( .B1(n222), .B2(n17876), .A(n600), .ZN(n19248) );
  OR2_X1 U993 ( .A1(n14838), .A2(n15018), .ZN(n322) );
  INV_X1 U994 ( .A(n16011), .ZN(n192) );
  INV_X1 U1002 ( .A(n12589), .ZN(n193) );
  CLKBUF_X1 U1005 ( .A(n10684), .Z(n12104) );
  NAND2_X1 U1006 ( .A1(n7284), .A2(n3210), .ZN(n8932) );
  NAND3_X1 U1009 ( .A1(n8151), .A2(n7864), .A3(n8261), .ZN(n7572) );
  NAND2_X1 U1010 ( .A1(n8175), .A2(n8179), .ZN(n7887) );
  CLKBUF_X1 U1012 ( .A(n7508), .Z(n7910) );
  NAND4_X1 U1014 ( .A1(n5353), .A2(n5352), .A3(n5351), .A4(n5350), .ZN(n7146)
         );
  CLKBUF_X1 U1017 ( .A(n4176), .Z(n4613) );
  CLKBUF_X1 U1019 ( .A(Key[14]), .Z(n16035) );
  CLKBUF_X1 U1020 ( .A(Key[118]), .Z(n2329) );
  CLKBUF_X1 U1021 ( .A(Key[104]), .Z(n2454) );
  CLKBUF_X1 U1022 ( .A(Key[147]), .Z(n2344) );
  CLKBUF_X1 U1023 ( .A(Key[141]), .Z(n2446) );
  CLKBUF_X1 U1024 ( .A(Key[128]), .Z(n2096) );
  CLKBUF_X1 U1025 ( .A(Key[45]), .Z(n17365) );
  CLKBUF_X1 U1027 ( .A(Key[32]), .Z(n1857) );
  CLKBUF_X1 U1028 ( .A(Key[68]), .Z(n18478) );
  CLKBUF_X1 U1029 ( .A(Key[29]), .Z(n18801) );
  CLKBUF_X1 U1031 ( .A(Key[157]), .Z(n1969) );
  CLKBUF_X1 U1032 ( .A(Key[145]), .Z(n2082) );
  CLKBUF_X1 U1033 ( .A(Key[101]), .Z(n18420) );
  CLKBUF_X1 U1034 ( .A(Key[67]), .Z(n18170) );
  CLKBUF_X1 U1035 ( .A(Key[171]), .Z(n17733) );
  AOI21_X1 U1036 ( .B1(n19267), .B2(n19276), .A(n658), .ZN(n19279) );
  NAND2_X1 U1038 ( .A1(n1557), .A2(n1556), .ZN(n19146) );
  MUX2_X1 U1043 ( .A(n16043), .B(n16042), .S(n19707), .Z(n19168) );
  INV_X1 U1044 ( .A(n19164), .ZN(n195) );
  AND2_X1 U1045 ( .A1(n3039), .A2(n17906), .ZN(n18358) );
  OAI211_X1 U1046 ( .C1(n220), .C2(n20127), .A(n17193), .B(n326), .ZN(n17820)
         );
  CLKBUF_X1 U1047 ( .A(n17225), .Z(n17510) );
  CLKBUF_X1 U1048 ( .A(n16251), .Z(n16629) );
  CLKBUF_X1 U1049 ( .A(n17394), .Z(n18754) );
  INV_X1 U1050 ( .A(n17676), .ZN(n1112) );
  XNOR2_X1 U1051 ( .A(n16935), .B(n16934), .ZN(n18948) );
  BUF_X1 U1055 ( .A(n16171), .Z(n17507) );
  XNOR2_X1 U1057 ( .A(n16433), .B(n16432), .ZN(n18092) );
  INV_X1 U1058 ( .A(n17876), .ZN(n196) );
  XNOR2_X1 U1061 ( .A(n15979), .B(n17143), .ZN(n16553) );
  INV_X1 U1065 ( .A(n15310), .ZN(n197) );
  INV_X1 U1066 ( .A(n15714), .ZN(n198) );
  INV_X1 U1067 ( .A(n14707), .ZN(n14273) );
  INV_X1 U1068 ( .A(n14547), .ZN(n199) );
  AND2_X1 U1069 ( .A1(n14562), .A2(n14566), .ZN(n14708) );
  INV_X1 U1072 ( .A(n14692), .ZN(n200) );
  XNOR2_X1 U1074 ( .A(n11789), .B(n11788), .ZN(n14199) );
  XNOR2_X1 U1076 ( .A(n12173), .B(n294), .ZN(n13636) );
  XNOR2_X1 U1077 ( .A(n12173), .B(n299), .ZN(n12850) );
  XNOR2_X1 U1078 ( .A(n12173), .B(n304), .ZN(n13049) );
  AND3_X1 U1082 ( .A1(n12164), .A2(n3476), .A3(n12163), .ZN(n12173) );
  OR2_X1 U1084 ( .A1(n1252), .A2(n193), .ZN(n1251) );
  INV_X1 U1085 ( .A(n248), .ZN(n685) );
  CLKBUF_X1 U1086 ( .A(n12275), .Z(n920) );
  NAND3_X1 U1093 ( .A1(n10847), .A2(n11202), .A3(n19920), .ZN(n10848) );
  AND3_X1 U1094 ( .A1(n11177), .A2(n11174), .A3(n9486), .ZN(n3219) );
  INV_X1 U1095 ( .A(n11330), .ZN(n202) );
  CLKBUF_X1 U1096 ( .A(n9548), .Z(n10952) );
  CLKBUF_X1 U1098 ( .A(n9351), .Z(n9486) );
  INV_X1 U1099 ( .A(n11216), .ZN(n204) );
  XNOR2_X1 U1100 ( .A(n9409), .B(n9410), .ZN(n10947) );
  INV_X1 U1101 ( .A(n11129), .ZN(n205) );
  XNOR2_X1 U1102 ( .A(n10030), .B(n298), .ZN(n9404) );
  XNOR2_X1 U1103 ( .A(n9646), .B(n296), .ZN(n8716) );
  XNOR2_X1 U1104 ( .A(n260), .B(n9646), .ZN(n9910) );
  XNOR2_X1 U1105 ( .A(n10030), .B(n300), .ZN(n9417) );
  NOR2_X1 U1107 ( .A1(n8847), .A2(n3201), .ZN(n9623) );
  INV_X1 U1113 ( .A(n8959), .ZN(n207) );
  OR2_X1 U1115 ( .A1(n1231), .A2(n277), .ZN(n377) );
  CLKBUF_X1 U1117 ( .A(n6734), .Z(n8373) );
  INV_X1 U1119 ( .A(n8016), .ZN(n208) );
  XNOR2_X1 U1120 ( .A(n1369), .B(n6630), .ZN(n8068) );
  XNOR2_X1 U1121 ( .A(n3570), .B(n3572), .ZN(n7479) );
  XNOR2_X1 U1122 ( .A(n5249), .B(n295), .ZN(n6386) );
  XNOR2_X1 U1123 ( .A(n5249), .B(n293), .ZN(n6620) );
  OR2_X1 U1125 ( .A1(n5947), .A2(n5946), .ZN(n7127) );
  NAND3_X1 U1126 ( .A1(n5187), .A2(n2978), .A3(n5186), .ZN(n7178) );
  AND2_X1 U1127 ( .A1(n355), .A2(n5848), .ZN(n354) );
  OAI211_X1 U1129 ( .C1(n5943), .C2(n6172), .A(n6175), .B(n5221), .ZN(n6873)
         );
  OR2_X1 U1131 ( .A1(n5816), .A2(n285), .ZN(n5820) );
  NAND2_X1 U1132 ( .A1(n827), .A2(n830), .ZN(n5435) );
  NOR3_X1 U1133 ( .A1(n6166), .A2(n170), .A3(n6171), .ZN(n569) );
  AND2_X1 U1135 ( .A1(n762), .A2(n3714), .ZN(n5747) );
  INV_X1 U1137 ( .A(n6067), .ZN(n209) );
  OR2_X1 U1139 ( .A1(n5079), .A2(n20002), .ZN(n4809) );
  INV_X1 U1141 ( .A(n4899), .ZN(n210) );
  CLKBUF_X1 U1142 ( .A(Key[85]), .Z(n18848) );
  CLKBUF_X1 U1143 ( .A(Key[46]), .Z(n632) );
  CLKBUF_X1 U1144 ( .A(Key[83]), .Z(n19336) );
  CLKBUF_X1 U1146 ( .A(Key[163]), .Z(n2347) );
  CLKBUF_X1 U1147 ( .A(Key[34]), .Z(n2376) );
  CLKBUF_X1 U1148 ( .A(Key[133]), .Z(n17170) );
  CLKBUF_X1 U1150 ( .A(Key[25]), .Z(n2218) );
  CLKBUF_X1 U1151 ( .A(Key[21]), .Z(n2375) );
  CLKBUF_X1 U1152 ( .A(Key[8]), .Z(n2298) );
  CLKBUF_X1 U1153 ( .A(Key[191]), .Z(n2123) );
  CLKBUF_X1 U1154 ( .A(Key[170]), .Z(n2284) );
  CLKBUF_X1 U1155 ( .A(Key[44]), .Z(n484) );
  CLKBUF_X1 U1156 ( .A(Key[18]), .Z(n19216) );
  CLKBUF_X1 U1157 ( .A(Key[96]), .Z(n2369) );
  CLKBUF_X1 U1158 ( .A(Key[58]), .Z(n1148) );
  CLKBUF_X1 U1159 ( .A(Key[182]), .Z(n1904) );
  CLKBUF_X1 U1160 ( .A(Key[90]), .Z(n18779) );
  CLKBUF_X1 U1161 ( .A(Key[11]), .Z(n2087) );
  CLKBUF_X1 U1162 ( .A(Key[111]), .Z(n16030) );
  CLKBUF_X1 U1163 ( .A(Key[168]), .Z(n2257) );
  CLKBUF_X1 U1164 ( .A(Key[15]), .Z(n16424) );
  CLKBUF_X1 U1165 ( .A(Key[161]), .Z(n2392) );
  CLKBUF_X1 U1166 ( .A(Key[125]), .Z(n19436) );
  CLKBUF_X1 U1167 ( .A(Key[89]), .Z(n1386) );
  CLKBUF_X1 U1168 ( .A(Key[86]), .Z(n2248) );
  CLKBUF_X1 U1169 ( .A(Key[0]), .Z(n2341) );
  CLKBUF_X1 U1170 ( .A(Key[64]), .Z(n457) );
  CLKBUF_X1 U1171 ( .A(Key[4]), .Z(n1996) );
  CLKBUF_X1 U1172 ( .A(Key[91]), .Z(n18006) );
  CLKBUF_X1 U1173 ( .A(Key[72]), .Z(n2122) );
  CLKBUF_X1 U1174 ( .A(Key[87]), .Z(n311) );
  CLKBUF_X1 U1175 ( .A(Key[116]), .Z(n16366) );
  CLKBUF_X1 U1176 ( .A(Key[150]), .Z(n642) );
  CLKBUF_X1 U1177 ( .A(Key[143]), .Z(n2448) );
  CLKBUF_X1 U1178 ( .A(Key[172]), .Z(n2323) );
  CLKBUF_X1 U1179 ( .A(Key[106]), .Z(n621) );
  CLKBUF_X1 U1180 ( .A(Key[37]), .Z(n2368) );
  CLKBUF_X1 U1181 ( .A(Key[130]), .Z(n573) );
  CLKBUF_X1 U1182 ( .A(Key[140]), .Z(n18090) );
  CLKBUF_X1 U1183 ( .A(Key[23]), .Z(n2410) );
  CLKBUF_X1 U1184 ( .A(Key[153]), .Z(n18070) );
  CLKBUF_X1 U1185 ( .A(Key[27]), .Z(n2395) );
  CLKBUF_X1 U1186 ( .A(Key[5]), .Z(n19018) );
  CLKBUF_X1 U1187 ( .A(Key[26]), .Z(n18433) );
  CLKBUF_X1 U1188 ( .A(Key[126]), .Z(n875) );
  CLKBUF_X1 U1190 ( .A(Key[71]), .Z(n18830) );
  CLKBUF_X1 U1191 ( .A(Key[92]), .Z(n15479) );
  CLKBUF_X1 U1193 ( .A(Key[40]), .Z(n347) );
  CLKBUF_X1 U1194 ( .A(Key[19]), .Z(n18208) );
  CLKBUF_X1 U1195 ( .A(Key[70]), .Z(n2067) );
  CLKBUF_X1 U1197 ( .A(Key[112]), .Z(n18304) );
  CLKBUF_X1 U1198 ( .A(Key[149]), .Z(n19243) );
  CLKBUF_X1 U1200 ( .A(Key[49]), .Z(n17587) );
  CLKBUF_X1 U1201 ( .A(Key[178]), .Z(n1869) );
  CLKBUF_X1 U1202 ( .A(Key[151]), .Z(n18716) );
  CLKBUF_X1 U1203 ( .A(Key[12]), .Z(n2280) );
  CLKBUF_X1 U1204 ( .A(Key[154]), .Z(n2424) );
  CLKBUF_X1 U1205 ( .A(Key[20]), .Z(n2222) );
  CLKBUF_X1 U1206 ( .A(Key[158]), .Z(n19321) );
  CLKBUF_X1 U1207 ( .A(Key[109]), .Z(n17466) );
  CLKBUF_X1 U1208 ( .A(Key[74]), .Z(n2356) );
  CLKBUF_X1 U1209 ( .A(Key[80]), .Z(n18988) );
  CLKBUF_X1 U1210 ( .A(Key[2]), .Z(n18203) );
  CLKBUF_X1 U1211 ( .A(Key[131]), .Z(n2385) );
  CLKBUF_X1 U1212 ( .A(Key[105]), .Z(n2208) );
  CLKBUF_X1 U1213 ( .A(Key[138]), .Z(n538) );
  CLKBUF_X1 U1214 ( .A(Key[152]), .Z(n2233) );
  CLKBUF_X1 U1216 ( .A(Key[166]), .Z(n2337) );
  CLKBUF_X1 U1217 ( .A(Key[134]), .Z(n641) );
  CLKBUF_X1 U1218 ( .A(Key[107]), .Z(n19205) );
  CLKBUF_X1 U1219 ( .A(Key[61]), .Z(n610) );
  CLKBUF_X1 U1220 ( .A(Key[115]), .Z(n16487) );
  CLKBUF_X1 U1221 ( .A(Key[135]), .Z(n19222) );
  CLKBUF_X1 U1222 ( .A(Key[77]), .Z(n17932) );
  CLKBUF_X1 U1225 ( .A(Key[122]), .Z(n18065) );
  CLKBUF_X1 U1226 ( .A(Key[16]), .Z(n404) );
  CLKBUF_X1 U1227 ( .A(Key[102]), .Z(n16242) );
  CLKBUF_X1 U1228 ( .A(Key[9]), .Z(n17089) );
  CLKBUF_X1 U1229 ( .A(Key[55]), .Z(n2310) );
  CLKBUF_X1 U1230 ( .A(Key[56]), .Z(n18338) );
  CLKBUF_X1 U1231 ( .A(Key[113]), .Z(n18863) );
  CLKBUF_X1 U1232 ( .A(Key[78]), .Z(n19467) );
  CLKBUF_X1 U1233 ( .A(Key[129]), .Z(n18439) );
  CLKBUF_X1 U1235 ( .A(Key[48]), .Z(n17804) );
  CLKBUF_X1 U1236 ( .A(Key[121]), .Z(n2296) );
  CLKBUF_X1 U1237 ( .A(Key[187]), .Z(n19158) );
  CLKBUF_X1 U1238 ( .A(Key[24]), .Z(n2164) );
  CLKBUF_X1 U1239 ( .A(Key[110]), .Z(n2307) );
  CLKBUF_X1 U1240 ( .A(Key[38]), .Z(n18887) );
  CLKBUF_X1 U1241 ( .A(Key[52]), .Z(n2203) );
  CLKBUF_X1 U1242 ( .A(Key[84]), .Z(n649) );
  CLKBUF_X1 U1243 ( .A(Key[76]), .Z(n18768) );
  CLKBUF_X1 U1244 ( .A(Key[169]), .Z(n18984) );
  CLKBUF_X1 U1245 ( .A(Key[148]), .Z(n2305) );
  CLKBUF_X1 U1246 ( .A(Key[114]), .Z(n2221) );
  CLKBUF_X1 U1248 ( .A(Key[47]), .Z(n19052) );
  CLKBUF_X1 U1249 ( .A(Key[73]), .Z(n2394) );
  CLKBUF_X1 U1250 ( .A(Key[17]), .Z(n18366) );
  CLKBUF_X1 U1251 ( .A(Key[62]), .Z(n18726) );
  CLKBUF_X1 U1252 ( .A(Key[127]), .Z(n2151) );
  CLKBUF_X1 U1253 ( .A(Key[188]), .Z(n18854) );
  CLKBUF_X1 U1254 ( .A(Key[146]), .Z(n17993) );
  CLKBUF_X1 U1255 ( .A(Key[155]), .Z(n17060) );
  CLKBUF_X1 U1256 ( .A(Key[10]), .Z(n18055) );
  CLKBUF_X1 U1257 ( .A(Key[181]), .Z(n2032) );
  CLKBUF_X1 U1258 ( .A(Key[162]), .Z(n18396) );
  CLKBUF_X1 U1259 ( .A(Key[120]), .Z(n16651) );
  CLKBUF_X1 U1261 ( .A(Key[43]), .Z(n2055) );
  CLKBUF_X1 U1262 ( .A(Key[66]), .Z(n2442) );
  CLKBUF_X1 U1263 ( .A(Key[31]), .Z(n2413) );
  CLKBUF_X1 U1264 ( .A(Key[35]), .Z(n18011) );
  CLKBUF_X1 U1265 ( .A(Key[3]), .Z(n2192) );
  INV_X1 U1267 ( .A(n19125), .ZN(n833) );
  MUX2_X1 U1269 ( .A(n17088), .B(n17087), .S(n19683), .Z(n17090) );
  OAI21_X1 U1270 ( .B1(n18201), .B2(n16446), .A(n2208), .ZN(n628) );
  OR2_X1 U1271 ( .A1(n17997), .A2(n18555), .ZN(n16459) );
  AND2_X1 U1272 ( .A1(n18646), .A2(n299), .ZN(n842) );
  OAI22_X1 U1274 ( .A1(n19692), .A2(n19163), .B1(n19948), .B2(n18306), .ZN(
        n19166) );
  CLKBUF_X1 U1275 ( .A(n18311), .Z(n19334) );
  NOR2_X1 U1277 ( .A1(n18465), .A2(n20110), .ZN(n18441) );
  OR2_X1 U1278 ( .A1(n18638), .A2(n18637), .ZN(n583) );
  AND2_X1 U1283 ( .A1(n930), .A2(n931), .ZN(n19460) );
  INV_X1 U1284 ( .A(n18009), .ZN(n18504) );
  AND2_X1 U1285 ( .A1(n19009), .A2(n19002), .ZN(n310) );
  AND3_X1 U1287 ( .A1(n16405), .A2(n1147), .A3(n1146), .ZN(n18559) );
  INV_X1 U1288 ( .A(n19190), .ZN(n19197) );
  INV_X1 U1292 ( .A(n19452), .ZN(n212) );
  INV_X1 U1293 ( .A(n18795), .ZN(n213) );
  AND3_X1 U1297 ( .A1(n1906), .A2(n1905), .A3(n982), .ZN(n19233) );
  INV_X1 U1298 ( .A(n18511), .ZN(n214) );
  OAI21_X1 U1306 ( .B1(n18268), .B2(n16869), .A(n16868), .ZN(n17054) );
  MUX2_X1 U1308 ( .A(n17151), .B(n17150), .S(n17957), .Z(n17152) );
  OAI21_X1 U1309 ( .B1(n612), .B2(n18262), .A(n611), .ZN(n17398) );
  INV_X1 U1311 ( .A(n1205), .ZN(n215) );
  NOR2_X1 U1312 ( .A1(n17164), .A2(n759), .ZN(n17165) );
  OR2_X1 U1313 ( .A1(n17864), .A2(n17595), .ZN(n601) );
  OR2_X1 U1314 ( .A1(n17762), .A2(n18264), .ZN(n18140) );
  OAI211_X1 U1316 ( .C1(n17161), .C2(n16792), .A(n16791), .B(n18542), .ZN(
        n17584) );
  INV_X1 U1317 ( .A(n18869), .ZN(n216) );
  OR2_X1 U1318 ( .A1(n196), .A2(n17879), .ZN(n17610) );
  NOR2_X1 U1319 ( .A1(n17495), .A2(n17492), .ZN(n17490) );
  INV_X1 U1320 ( .A(n17492), .ZN(n16801) );
  CLKBUF_X1 U1321 ( .A(n17458), .Z(n17559) );
  OR2_X1 U1322 ( .A1(n19846), .A2(n18948), .ZN(n17315) );
  MUX2_X1 U1324 ( .A(n17830), .B(n17829), .S(n20221), .Z(n17834) );
  AND2_X1 U1332 ( .A1(n18221), .A2(n18977), .ZN(n18224) );
  INV_X1 U1334 ( .A(n18956), .ZN(n219) );
  OR2_X1 U1335 ( .A1(n18273), .A2(n18033), .ZN(n17764) );
  INV_X1 U1337 ( .A(n19380), .ZN(n635) );
  XNOR2_X1 U1338 ( .A(n16060), .B(n16061), .ZN(n17879) );
  AOI21_X1 U1339 ( .B1(n18221), .B2(n20499), .A(n18976), .ZN(n320) );
  BUF_X1 U1340 ( .A(n17187), .Z(n18935) );
  INV_X1 U1341 ( .A(n17245), .ZN(n812) );
  XNOR2_X1 U1342 ( .A(n16520), .B(n16519), .ZN(n17861) );
  BUF_X1 U1344 ( .A(n16540), .Z(n19348) );
  INV_X1 U1345 ( .A(n18968), .ZN(n220) );
  INV_X1 U1348 ( .A(n18273), .ZN(n221) );
  XNOR2_X1 U1350 ( .A(n15949), .B(n15950), .ZN(n17825) );
  INV_X1 U1351 ( .A(n19823), .ZN(n815) );
  INV_X1 U1354 ( .A(n17881), .ZN(n222) );
  XNOR2_X1 U1356 ( .A(n16904), .B(n16903), .ZN(n18976) );
  INV_X1 U1359 ( .A(n18221), .ZN(n224) );
  INV_X1 U1360 ( .A(n20499), .ZN(n225) );
  XNOR2_X1 U1362 ( .A(n16585), .B(n16586), .ZN(n19396) );
  INV_X1 U1363 ( .A(n18092), .ZN(n226) );
  XNOR2_X1 U1364 ( .A(n15557), .B(n15556), .ZN(n16666) );
  INV_X1 U1365 ( .A(n17818), .ZN(n227) );
  XNOR2_X1 U1366 ( .A(n17102), .B(n334), .ZN(n16132) );
  INV_X1 U1367 ( .A(n15979), .ZN(n17005) );
  AND3_X1 U1369 ( .A1(n15035), .A2(n3314), .A3(n1898), .ZN(n16969) );
  AND3_X1 U1374 ( .A1(n1079), .A2(n1077), .A3(n1075), .ZN(n16240) );
  INV_X1 U1375 ( .A(n16045), .ZN(n335) );
  NAND2_X1 U1378 ( .A1(n565), .A2(n1154), .ZN(n16292) );
  NAND3_X1 U1379 ( .A1(n1645), .A2(n1644), .A3(n1650), .ZN(n16507) );
  NAND2_X1 U1381 ( .A1(n15796), .A2(n691), .ZN(n690) );
  OR2_X1 U1382 ( .A1(n15771), .A2(n15665), .ZN(n1443) );
  MUX2_X1 U1383 ( .A(n15058), .B(n15057), .S(n15409), .Z(n16269) );
  OR2_X1 U1385 ( .A1(n717), .A2(n15846), .ZN(n714) );
  OR2_X1 U1386 ( .A1(n15227), .A2(n15451), .ZN(n349) );
  OAI21_X1 U1387 ( .B1(n15307), .B2(n15306), .A(n361), .ZN(n2969) );
  MUX2_X1 U1388 ( .A(n15364), .B(n15045), .S(n1520), .Z(n14951) );
  INV_X1 U1389 ( .A(n717), .ZN(n15640) );
  AND2_X1 U1390 ( .A1(n13181), .A2(n2023), .ZN(n783) );
  NOR2_X1 U1391 ( .A1(n15857), .A2(n15720), .ZN(n15171) );
  NAND2_X1 U1392 ( .A1(n3496), .A2(n14586), .ZN(n15270) );
  AND2_X1 U1395 ( .A1(n16128), .A2(n15734), .ZN(n387) );
  INV_X1 U1398 ( .A(n14954), .ZN(n15808) );
  OR2_X1 U1399 ( .A1(n546), .A2(n15474), .ZN(n2113) );
  INV_X1 U1400 ( .A(n15060), .ZN(n15307) );
  NAND2_X1 U1401 ( .A1(n15812), .A2(n15813), .ZN(n3313) );
  CLKBUF_X1 U1403 ( .A(n14312), .Z(n15056) );
  AND2_X1 U1405 ( .A1(n15070), .A2(n15405), .ZN(n15617) );
  OR2_X1 U1406 ( .A1(n14754), .A2(n14757), .ZN(n15822) );
  AND2_X1 U1407 ( .A1(n2889), .A2(n14702), .ZN(n942) );
  INV_X1 U1408 ( .A(n15796), .ZN(n15364) );
  OAI21_X1 U1409 ( .B1(n914), .B2(n14489), .A(n14488), .ZN(n15132) );
  INV_X1 U1411 ( .A(n15311), .ZN(n361) );
  INV_X1 U1412 ( .A(n15028), .ZN(n3621) );
  INV_X1 U1413 ( .A(n15671), .ZN(n15666) );
  INV_X1 U1414 ( .A(n15812), .ZN(n228) );
  AND3_X1 U1415 ( .A1(n1743), .A2(n1741), .A3(n1739), .ZN(n15673) );
  AOI21_X1 U1417 ( .B1(n14538), .B2(n2676), .A(n14537), .ZN(n14997) );
  NOR2_X1 U1420 ( .A1(n14670), .A2(n14671), .ZN(n859) );
  INV_X1 U1421 ( .A(n15657), .ZN(n229) );
  INV_X1 U1422 ( .A(n15846), .ZN(n230) );
  INV_X1 U1429 ( .A(n15491), .ZN(n15755) );
  OAI22_X1 U1431 ( .A1(n13953), .A2(n13952), .B1(n2642), .B2(n14134), .ZN(
        n16011) );
  INV_X1 U1432 ( .A(n15490), .ZN(n15588) );
  INV_X1 U1433 ( .A(n20183), .ZN(n232) );
  OR2_X1 U1435 ( .A1(n15815), .A2(n15813), .ZN(n15035) );
  INV_X1 U1436 ( .A(n15813), .ZN(n233) );
  OR3_X1 U1437 ( .A1(n14198), .A2(n14197), .A3(n14590), .ZN(n2789) );
  INV_X1 U1438 ( .A(n15667), .ZN(n234) );
  OR2_X1 U1439 ( .A1(n13957), .A2(n14705), .ZN(n402) );
  MUX2_X1 U1441 ( .A(n14669), .B(n14668), .S(n14667), .Z(n14670) );
  XNOR2_X1 U1442 ( .A(n13680), .B(n13681), .ZN(n14718) );
  MUX2_X1 U1443 ( .A(n13948), .B(n13947), .S(n200), .Z(n13949) );
  BUF_X1 U1445 ( .A(n13901), .Z(n14782) );
  BUF_X1 U1446 ( .A(n14727), .Z(n14408) );
  INV_X1 U1447 ( .A(n14548), .ZN(n14654) );
  INV_X1 U1448 ( .A(n13940), .ZN(n2039) );
  XNOR2_X1 U1450 ( .A(n3236), .B(n12015), .ZN(n14203) );
  AND2_X1 U1452 ( .A1(n13865), .A2(n14441), .ZN(n2983) );
  XNOR2_X1 U1457 ( .A(n13187), .B(n13188), .ZN(n14548) );
  INV_X1 U1459 ( .A(n14818), .ZN(n3444) );
  INV_X1 U1460 ( .A(n14820), .ZN(n235) );
  CLKBUF_X1 U1462 ( .A(n13872), .Z(n14524) );
  INV_X1 U1463 ( .A(n14724), .ZN(n236) );
  AND2_X1 U1464 ( .A1(n951), .A2(n14648), .ZN(n779) );
  XNOR2_X1 U1465 ( .A(n13034), .B(n2240), .ZN(n13868) );
  INV_X1 U1467 ( .A(n14522), .ZN(n237) );
  INV_X1 U1469 ( .A(n14442), .ZN(n238) );
  INV_X1 U1471 ( .A(n14199), .ZN(n239) );
  XNOR2_X1 U1472 ( .A(n13669), .B(n13670), .ZN(n14714) );
  XNOR2_X1 U1473 ( .A(n13286), .B(n13285), .ZN(n14563) );
  XNOR2_X1 U1475 ( .A(n13801), .B(n13800), .ZN(n14239) );
  INV_X1 U1476 ( .A(n14228), .ZN(n240) );
  INV_X1 U1477 ( .A(n20266), .ZN(n241) );
  XNOR2_X1 U1478 ( .A(n13242), .B(n627), .ZN(n13246) );
  XNOR2_X1 U1479 ( .A(n13028), .B(n979), .ZN(n1089) );
  INV_X1 U1480 ( .A(n12977), .ZN(n13757) );
  INV_X1 U1481 ( .A(n13231), .ZN(n13706) );
  XNOR2_X1 U1482 ( .A(n13136), .B(n13088), .ZN(n13382) );
  XNOR2_X1 U1483 ( .A(n13193), .B(n18478), .ZN(n12999) );
  XNOR2_X1 U1485 ( .A(n13755), .B(n13687), .ZN(n627) );
  XNOR2_X1 U1490 ( .A(n12173), .B(n357), .ZN(n13086) );
  XNOR2_X1 U1493 ( .A(n13703), .B(n13059), .ZN(n12826) );
  AND4_X1 U1494 ( .A1(n3530), .A2(n11139), .A3(n11137), .A4(n11138), .ZN(
        n13330) );
  INV_X1 U1496 ( .A(n12709), .ZN(n13827) );
  AND2_X1 U1497 ( .A1(n553), .A2(n552), .ZN(n551) );
  OR2_X1 U1501 ( .A1(n12557), .A2(n12558), .ZN(n13017) );
  OAI21_X1 U1505 ( .B1(n12815), .B2(n12814), .A(n12813), .ZN(n13287) );
  NAND3_X1 U1506 ( .A1(n2432), .A2(n12140), .A3(n2431), .ZN(n13446) );
  XNOR2_X1 U1507 ( .A(n13511), .B(n19205), .ZN(n3365) );
  INV_X1 U1509 ( .A(n12770), .ZN(n13745) );
  OAI211_X1 U1511 ( .C1(n12359), .C2(n12506), .A(n12012), .B(n12011), .ZN(
        n13673) );
  OAI211_X1 U1513 ( .C1(n741), .C2(n11730), .A(n3816), .B(n740), .ZN(n12770)
         );
  OR2_X1 U1514 ( .A1(n1366), .A2(n685), .ZN(n684) );
  AOI22_X1 U1515 ( .A1(n10822), .A2(n12206), .B1(n2713), .B2(n12211), .ZN(
        n2711) );
  OAI21_X1 U1516 ( .B1(n11983), .B2(n12619), .A(n11982), .ZN(n13634) );
  OR2_X1 U1519 ( .A1(n11832), .A2(n11833), .ZN(n1471) );
  INV_X1 U1520 ( .A(n11793), .ZN(n850) );
  OR2_X1 U1523 ( .A1(n20457), .A2(n12642), .ZN(n491) );
  AND2_X1 U1524 ( .A1(n13145), .A2(n13147), .ZN(n356) );
  AND2_X1 U1526 ( .A1(n12589), .A2(n12202), .ZN(n563) );
  OR2_X1 U1527 ( .A1(n11658), .A2(n11951), .ZN(n488) );
  NOR2_X1 U1528 ( .A1(n12639), .A2(n12455), .ZN(n12637) );
  OAI21_X1 U1529 ( .B1(n698), .B2(n12131), .A(n12130), .ZN(n697) );
  NOR2_X1 U1531 ( .A1(n12084), .A2(n12416), .ZN(n369) );
  INV_X1 U1532 ( .A(n12174), .ZN(n415) );
  OR2_X1 U1534 ( .A1(n11670), .A2(n12180), .ZN(n11672) );
  OR2_X1 U1535 ( .A1(n12514), .A2(n11997), .ZN(n521) );
  AND3_X1 U1536 ( .A1(n10848), .A2(n2060), .A3(n2061), .ZN(n12201) );
  INV_X1 U1537 ( .A(n12250), .ZN(n242) );
  OAI211_X1 U1538 ( .C1(n12437), .C2(n12442), .A(n11942), .B(n12443), .ZN(
        n10686) );
  OR2_X1 U1539 ( .A1(n11845), .A2(n20427), .ZN(n588) );
  OR2_X1 U1543 ( .A1(n11478), .A2(n3481), .ZN(n313) );
  INV_X1 U1544 ( .A(n12532), .ZN(n243) );
  OR2_X1 U1545 ( .A1(n12636), .A2(n12449), .ZN(n11948) );
  OR3_X1 U1546 ( .A1(n12576), .A2(n11683), .A3(n11926), .ZN(n3816) );
  INV_X1 U1549 ( .A(n953), .ZN(n3586) );
  AND2_X1 U1551 ( .A1(n3639), .A2(n3638), .ZN(n12257) );
  INV_X1 U1552 ( .A(n12255), .ZN(n244) );
  INV_X1 U1553 ( .A(n12759), .ZN(n245) );
  INV_X1 U1554 ( .A(n11618), .ZN(n246) );
  INV_X1 U1556 ( .A(n948), .ZN(n247) );
  OR2_X1 U1558 ( .A1(n10930), .A2(n10926), .ZN(n1892) );
  CLKBUF_X1 U1560 ( .A(n11061), .Z(n12016) );
  INV_X1 U1561 ( .A(n12417), .ZN(n12084) );
  INV_X1 U1562 ( .A(n12263), .ZN(n248) );
  NAND3_X1 U1564 ( .A1(n11576), .A2(n11575), .A3(n3151), .ZN(n12273) );
  INV_X1 U1566 ( .A(n12349), .ZN(n249) );
  OAI21_X1 U1569 ( .B1(n11407), .B2(n19506), .A(n2810), .ZN(n12544) );
  INV_X1 U1570 ( .A(n12554), .ZN(n250) );
  INV_X1 U1571 ( .A(n12442), .ZN(n251) );
  INV_X1 U1575 ( .A(n12180), .ZN(n252) );
  INV_X1 U1576 ( .A(n12399), .ZN(n253) );
  INV_X1 U1577 ( .A(n12408), .ZN(n254) );
  OR2_X1 U1579 ( .A1(n1279), .A2(n1280), .ZN(n766) );
  AND2_X1 U1580 ( .A1(n2043), .A2(n10861), .ZN(n874) );
  AND2_X1 U1582 ( .A1(n727), .A2(n725), .ZN(n724) );
  INV_X1 U1583 ( .A(n12126), .ZN(n255) );
  NOR2_X1 U1585 ( .A1(n9413), .A2(n11281), .ZN(n606) );
  INV_X1 U1586 ( .A(n11673), .ZN(n256) );
  INV_X1 U1587 ( .A(n12415), .ZN(n257) );
  OAI21_X1 U1589 ( .B1(n11340), .B2(n10198), .A(n10197), .ZN(n11992) );
  OAI211_X1 U1590 ( .C1(n11458), .C2(n1814), .A(n11457), .B(n1813), .ZN(n12290) );
  CLKBUF_X1 U1592 ( .A(n10785), .Z(n10814) );
  OR2_X1 U1593 ( .A1(n11200), .A2(n11493), .ZN(n798) );
  MUX2_X1 U1594 ( .A(n11525), .B(n11524), .S(n11523), .Z(n11741) );
  OR2_X1 U1595 ( .A1(n10845), .A2(n10726), .ZN(n11203) );
  INV_X1 U1597 ( .A(n12107), .ZN(n765) );
  OR2_X1 U1598 ( .A1(n11264), .A2(n11339), .ZN(n753) );
  INV_X1 U1599 ( .A(n11574), .ZN(n723) );
  OR2_X1 U1601 ( .A1(n11006), .A2(n11005), .ZN(n411) );
  OR2_X1 U1602 ( .A1(n11079), .A2(n3482), .ZN(n11080) );
  OAI21_X1 U1603 ( .B1(n732), .B2(n11539), .A(n731), .ZN(n10738) );
  NOR2_X1 U1604 ( .A1(n11168), .A2(n11538), .ZN(n732) );
  AND2_X1 U1605 ( .A1(n12103), .A2(n11381), .ZN(n12107) );
  INV_X1 U1607 ( .A(n11538), .ZN(n11171) );
  MUX2_X1 U1608 ( .A(n10758), .B(n10757), .S(n10756), .Z(n10759) );
  INV_X1 U1609 ( .A(n11275), .ZN(n764) );
  OR2_X1 U1610 ( .A1(n20517), .A2(n11866), .ZN(n1403) );
  BUF_X1 U1611 ( .A(n9616), .Z(n10701) );
  INV_X1 U1612 ( .A(n11087), .ZN(n11114) );
  OR2_X1 U1613 ( .A1(n11538), .A2(n10640), .ZN(n11540) );
  OR2_X1 U1614 ( .A1(n9830), .A2(n10673), .ZN(n756) );
  NAND2_X1 U1615 ( .A1(n11133), .A2(n19959), .ZN(n3295) );
  OR2_X1 U1616 ( .A1(n11476), .A2(n11475), .ZN(n10893) );
  NOR2_X1 U1617 ( .A1(n3588), .A2(n11294), .ZN(n11405) );
  OR2_X1 U1620 ( .A1(n11489), .A2(n11493), .ZN(n11198) );
  OR2_X1 U1622 ( .A1(n11437), .A2(n11440), .ZN(n11916) );
  XNOR2_X1 U1625 ( .A(n9428), .B(n9944), .ZN(n11277) );
  CLKBUF_X1 U1627 ( .A(n10726), .Z(n11201) );
  XNOR2_X1 U1628 ( .A(n10269), .B(n10268), .ZN(n11325) );
  INV_X1 U1631 ( .A(n11535), .ZN(n731) );
  OR2_X1 U1632 ( .A1(n11302), .A2(n19750), .ZN(n11387) );
  INV_X1 U1634 ( .A(n11550), .ZN(n258) );
  XNOR2_X1 U1635 ( .A(n9816), .B(n9815), .ZN(n9830) );
  XNOR2_X1 U1636 ( .A(n2938), .B(n9997), .ZN(n11513) );
  INV_X1 U1637 ( .A(n11510), .ZN(n259) );
  CLKBUF_X1 U1638 ( .A(n11113), .Z(n11456) );
  CLKBUF_X1 U1640 ( .A(n9551), .Z(n11010) );
  XNOR2_X1 U1643 ( .A(n8900), .B(n8899), .ZN(n11539) );
  XNOR2_X1 U1644 ( .A(n10162), .B(n10161), .ZN(n11428) );
  XNOR2_X1 U1646 ( .A(n9829), .B(n9828), .ZN(n11339) );
  XNOR2_X1 U1647 ( .A(n10408), .B(n10407), .ZN(n10829) );
  XNOR2_X1 U1653 ( .A(n802), .B(n801), .ZN(n9603) );
  INV_X1 U1655 ( .A(n9462), .ZN(n790) );
  XNOR2_X1 U1656 ( .A(n9602), .B(n9983), .ZN(n802) );
  CLKBUF_X1 U1657 ( .A(n9537), .Z(n10483) );
  XNOR2_X1 U1658 ( .A(n9646), .B(n768), .ZN(n10238) );
  XNOR2_X1 U1659 ( .A(n10281), .B(n9862), .ZN(n10563) );
  INV_X1 U1660 ( .A(n10185), .ZN(n10441) );
  XNOR2_X1 U1661 ( .A(n9623), .B(n9624), .ZN(n10343) );
  XNOR2_X1 U1662 ( .A(n9646), .B(n767), .ZN(n9388) );
  INV_X1 U1665 ( .A(n9414), .ZN(n10143) );
  BUF_X1 U1666 ( .A(n9856), .Z(n10205) );
  XNOR2_X1 U1667 ( .A(n10237), .B(n1228), .ZN(n1227) );
  NAND4_X1 U1670 ( .A1(n3200), .A2(n8935), .A3(n3199), .A4(n3799), .ZN(n9624)
         );
  NAND3_X1 U1672 ( .A1(n7900), .A2(n7901), .A3(n7899), .ZN(n10528) );
  OAI211_X1 U1674 ( .C1(n9218), .C2(n8670), .A(n8669), .B(n8668), .ZN(n10332)
         );
  XNOR2_X1 U1675 ( .A(n9414), .B(n17024), .ZN(n801) );
  OAI211_X1 U1676 ( .C1(n6215), .C2(n9238), .A(n6214), .B(n6213), .ZN(n9819)
         );
  NAND2_X1 U1681 ( .A1(n7658), .A2(n2336), .ZN(n9430) );
  AND3_X1 U1682 ( .A1(n8851), .A2(n590), .A3(n589), .ZN(n7175) );
  AND2_X1 U1683 ( .A1(n9160), .A2(n436), .ZN(n1257) );
  OAI211_X1 U1685 ( .C1(n9152), .C2(n1544), .A(n1543), .B(n1542), .ZN(n10061)
         );
  AND2_X1 U1688 ( .A1(n8475), .A2(n8976), .ZN(n577) );
  OR2_X1 U1692 ( .A1(n9566), .A2(n9346), .ZN(n2171) );
  INV_X1 U1693 ( .A(n10157), .ZN(n260) );
  OR2_X1 U1694 ( .A1(n9059), .A2(n9031), .ZN(n3072) );
  OR2_X1 U1695 ( .A1(n9298), .A2(n7424), .ZN(n7440) );
  NOR2_X1 U1696 ( .A1(n8987), .A2(n9172), .ZN(n8763) );
  OR2_X1 U1697 ( .A1(n1765), .A2(n9031), .ZN(n1766) );
  OR2_X1 U1698 ( .A1(n8498), .A2(n8499), .ZN(n704) );
  OR2_X1 U1699 ( .A1(n8965), .A2(n207), .ZN(n838) );
  OR2_X1 U1702 ( .A1(n8960), .A2(n8959), .ZN(n7559) );
  OR2_X1 U1703 ( .A1(n8338), .A2(n8790), .ZN(n8439) );
  INV_X1 U1706 ( .A(n9300), .ZN(n9297) );
  OR2_X1 U1707 ( .A1(n978), .A2(n19490), .ZN(n464) );
  INV_X1 U1709 ( .A(n2097), .ZN(n9238) );
  AND2_X1 U1711 ( .A1(n778), .A2(n777), .ZN(n7996) );
  AND2_X1 U1712 ( .A1(n8499), .A2(n8733), .ZN(n7665) );
  INV_X1 U1714 ( .A(n8923), .ZN(n3645) );
  INV_X1 U1715 ( .A(n8786), .ZN(n261) );
  NOR2_X1 U1716 ( .A1(n8125), .A2(n8124), .ZN(n8995) );
  NAND2_X1 U1719 ( .A1(n737), .A2(n7509), .ZN(n9049) );
  OAI211_X1 U1720 ( .C1(n7505), .C2(n7931), .A(n7506), .B(n1402), .ZN(n9287)
         );
  AND2_X1 U1721 ( .A1(n9114), .A2(n9113), .ZN(n9219) );
  INV_X1 U1722 ( .A(n9333), .ZN(n262) );
  OR2_X1 U1723 ( .A1(n9168), .A2(n8569), .ZN(n777) );
  INV_X1 U1726 ( .A(n9210), .ZN(n263) );
  NAND3_X1 U1727 ( .A1(n2156), .A2(n2155), .A3(n6894), .ZN(n9228) );
  INV_X1 U1728 ( .A(n655), .ZN(n9233) );
  INV_X1 U1729 ( .A(n8569), .ZN(n264) );
  OAI21_X1 U1730 ( .B1(n8137), .B2(n8138), .A(n8136), .ZN(n352) );
  OAI21_X1 U1732 ( .B1(n6701), .B2(n8261), .A(n6700), .ZN(n9305) );
  INV_X1 U1733 ( .A(n8985), .ZN(n265) );
  INV_X1 U1736 ( .A(n9162), .ZN(n437) );
  INV_X1 U1741 ( .A(n9189), .ZN(n266) );
  INV_X1 U1742 ( .A(n6587), .ZN(n267) );
  INV_X1 U1745 ( .A(n9242), .ZN(n268) );
  INV_X1 U1747 ( .A(n8568), .ZN(n269) );
  INV_X1 U1748 ( .A(n9018), .ZN(n270) );
  INV_X1 U1751 ( .A(n770), .ZN(n8434) );
  INV_X1 U1753 ( .A(n9166), .ZN(n8705) );
  AND3_X1 U1756 ( .A1(n493), .A2(n6284), .A3(n6283), .ZN(n8470) );
  OR2_X1 U1757 ( .A1(n7807), .A2(n462), .ZN(n461) );
  OR2_X1 U1758 ( .A1(n8236), .A2(n6539), .ZN(n770) );
  OR2_X1 U1760 ( .A1(n7499), .A2(n163), .ZN(n3377) );
  CLKBUF_X1 U1761 ( .A(n7717), .Z(n7723) );
  AND3_X1 U1764 ( .A1(n7760), .A2(n6903), .A3(n3089), .ZN(n9162) );
  AOI21_X1 U1767 ( .B1(n1198), .B2(n7541), .A(n1197), .ZN(n8823) );
  AND3_X1 U1769 ( .A1(n2934), .A2(n8368), .A3(n8367), .ZN(n8420) );
  AND2_X1 U1770 ( .A1(n7513), .A2(n7514), .ZN(n738) );
  AOI211_X1 U1771 ( .C1(n7912), .C2(n7745), .A(n6908), .B(n7911), .ZN(n6909)
         );
  INV_X1 U1772 ( .A(n7602), .ZN(n7793) );
  OR2_X1 U1773 ( .A1(n7417), .A2(n8068), .ZN(n428) );
  INV_X1 U1774 ( .A(n8091), .ZN(n718) );
  OR2_X1 U1775 ( .A1(n6539), .A2(n19826), .ZN(n358) );
  NAND3_X1 U1776 ( .A1(n8183), .A2(n7464), .A3(n7463), .ZN(n9023) );
  BUF_X1 U1777 ( .A(n7389), .Z(n7807) );
  AND2_X1 U1778 ( .A1(n20195), .A2(n7936), .ZN(n6244) );
  AND2_X1 U1779 ( .A1(n8010), .A2(n1560), .ZN(n427) );
  INV_X1 U1780 ( .A(n1726), .ZN(n505) );
  INV_X1 U1783 ( .A(n8003), .ZN(n324) );
  OR2_X1 U1785 ( .A1(n7903), .A2(n7530), .ZN(n494) );
  OR2_X1 U1786 ( .A1(n7918), .A2(n7917), .ZN(n376) );
  AND2_X1 U1787 ( .A1(n8212), .A2(n8095), .ZN(n8091) );
  NOR2_X1 U1788 ( .A1(n7801), .A2(n208), .ZN(n629) );
  AND2_X1 U1789 ( .A1(n8300), .A2(n5941), .ZN(n7787) );
  INV_X1 U1790 ( .A(n7967), .ZN(n776) );
  XNOR2_X1 U1794 ( .A(n1074), .B(n1073), .ZN(n8251) );
  XNOR2_X1 U1796 ( .A(n6823), .B(n6822), .ZN(n8159) );
  BUF_X1 U1799 ( .A(n6312), .Z(n7982) );
  OR2_X1 U1800 ( .A1(n7833), .A2(n8910), .ZN(n7773) );
  INV_X1 U1801 ( .A(n7991), .ZN(n273) );
  INV_X1 U1802 ( .A(n7908), .ZN(n274) );
  XNOR2_X1 U1806 ( .A(n639), .B(n6691), .ZN(n895) );
  INV_X1 U1807 ( .A(n8325), .ZN(n276) );
  XNOR2_X1 U1808 ( .A(n6372), .B(n6371), .ZN(n7709) );
  XNOR2_X1 U1809 ( .A(n6583), .B(n6582), .ZN(n8111) );
  XNOR2_X1 U1810 ( .A(n6291), .B(n6292), .ZN(n7978) );
  INV_X1 U1811 ( .A(n7631), .ZN(n2703) );
  INV_X1 U1812 ( .A(n2977), .ZN(n277) );
  XNOR2_X1 U1813 ( .A(n2622), .B(n5898), .ZN(n5941) );
  INV_X1 U1814 ( .A(n7971), .ZN(n278) );
  XNOR2_X1 U1815 ( .A(n7075), .B(n7076), .ZN(n1560) );
  INV_X1 U1817 ( .A(n7855), .ZN(n279) );
  INV_X1 U1819 ( .A(n7754), .ZN(n280) );
  INV_X1 U1820 ( .A(n7475), .ZN(n281) );
  XNOR2_X1 U1821 ( .A(n7236), .B(n7235), .ZN(n8016) );
  INV_X1 U1823 ( .A(n6830), .ZN(n282) );
  AND2_X1 U1826 ( .A1(n6217), .A2(n6221), .ZN(n7360) );
  INV_X1 U1827 ( .A(n6690), .ZN(n639) );
  XNOR2_X1 U1828 ( .A(n459), .B(n6032), .ZN(n6040) );
  XNOR2_X1 U1829 ( .A(n7178), .B(n7273), .ZN(n6838) );
  XNOR2_X1 U1830 ( .A(n6024), .B(n7333), .ZN(n459) );
  INV_X1 U1833 ( .A(n3068), .ZN(n7305) );
  INV_X1 U1834 ( .A(n7143), .ZN(n353) );
  OAI21_X1 U1836 ( .B1(n6148), .B2(n6147), .A(n6146), .ZN(n7206) );
  XNOR2_X1 U1838 ( .A(n354), .B(n7274), .ZN(n6593) );
  OAI211_X1 U1840 ( .C1(n5620), .C2(n6143), .A(n5619), .B(n5618), .ZN(n6713)
         );
  AND2_X1 U1844 ( .A1(n6207), .A2(n6208), .ZN(n6221) );
  INV_X1 U1846 ( .A(n354), .ZN(n6793) );
  XNOR2_X1 U1847 ( .A(n3663), .B(n7146), .ZN(n6506) );
  NAND2_X1 U1853 ( .A1(n2524), .A2(n480), .ZN(n6719) );
  OR2_X1 U1854 ( .A1(n5359), .A2(n5358), .ZN(n7142) );
  OAI21_X1 U1859 ( .B1(n6192), .B2(n5234), .A(n5233), .ZN(n6919) );
  INV_X1 U1862 ( .A(n6220), .ZN(n3674) );
  AOI22_X1 U1864 ( .A1(n5348), .A2(n5720), .B1(n3664), .B2(n5347), .ZN(n5984)
         );
  MUX2_X1 U1865 ( .A(n4689), .B(n4688), .S(n6172), .Z(n4690) );
  MUX2_X1 U1869 ( .A(n5446), .B(n5445), .S(n5645), .Z(n7257) );
  OR2_X1 U1870 ( .A1(n6003), .A2(n6000), .ZN(n3602) );
  NOR2_X1 U1873 ( .A1(n6173), .A2(n5842), .ZN(n568) );
  OR2_X1 U1875 ( .A1(n5868), .A2(n6119), .ZN(n2092) );
  AOI21_X1 U1877 ( .B1(n2407), .B2(n5790), .A(n5428), .ZN(n2879) );
  OR2_X1 U1878 ( .A1(n6379), .A2(n5847), .ZN(n5848) );
  INV_X1 U1879 ( .A(n5953), .ZN(n283) );
  OR2_X1 U1880 ( .A1(n5622), .A2(n5623), .ZN(n6134) );
  OR2_X1 U1881 ( .A1(n5745), .A2(n5742), .ZN(n1883) );
  OAI21_X1 U1883 ( .B1(n5322), .B2(n5395), .A(n1838), .ZN(n533) );
  AND2_X1 U1884 ( .A1(n5930), .A2(n6027), .ZN(n5596) );
  AND2_X1 U1885 ( .A1(n5201), .A2(n5745), .ZN(n455) );
  OR3_X1 U1886 ( .A1(n5823), .A2(n6017), .A3(n6016), .ZN(n5829) );
  AND2_X1 U1888 ( .A1(n618), .A2(n617), .ZN(n5742) );
  NOR2_X1 U1890 ( .A1(n1685), .A2(n3606), .ZN(n5718) );
  OR2_X1 U1891 ( .A1(n5393), .A2(n5395), .ZN(n5369) );
  BUF_X1 U1892 ( .A(n5483), .Z(n5716) );
  INV_X1 U1893 ( .A(n3701), .ZN(n5748) );
  OR2_X1 U1894 ( .A1(n5328), .A2(n6049), .ZN(n3919) );
  INV_X1 U1895 ( .A(n6124), .ZN(n6120) );
  AND2_X1 U1896 ( .A1(n4282), .A2(n4281), .ZN(n508) );
  INV_X1 U1898 ( .A(n5952), .ZN(n284) );
  INV_X1 U1902 ( .A(n733), .ZN(n5571) );
  INV_X1 U1905 ( .A(n5985), .ZN(n285) );
  NAND4_X1 U1906 ( .A1(n760), .A2(n761), .A3(n3714), .A4(n762), .ZN(n3701) );
  NAND2_X1 U1907 ( .A1(n2572), .A2(n2573), .ZN(n5611) );
  INV_X1 U1908 ( .A(n5802), .ZN(n5378) );
  INV_X1 U1909 ( .A(n6068), .ZN(n473) );
  NAND2_X1 U1910 ( .A1(n4301), .A2(n4300), .ZN(n5363) );
  NAND2_X1 U1911 ( .A1(n4120), .A2(n4121), .ZN(n5971) );
  OAI21_X1 U1912 ( .B1(n4124), .B2(n4985), .A(n4123), .ZN(n5699) );
  INV_X1 U1917 ( .A(n5251), .ZN(n5398) );
  INV_X1 U1918 ( .A(n5172), .ZN(n5957) );
  NOR2_X1 U1919 ( .A1(n5531), .A2(n6036), .ZN(n5566) );
  INV_X1 U1921 ( .A(n5747), .ZN(n286) );
  OAI21_X1 U1926 ( .B1(n4364), .B2(n604), .A(n603), .ZN(n4375) );
  OR2_X1 U1927 ( .A1(n4034), .A2(n4033), .ZN(n1214) );
  OAI211_X1 U1930 ( .C1(n4980), .C2(n4979), .A(n4978), .B(n3517), .ZN(n5563)
         );
  OAI211_X1 U1931 ( .C1(n4964), .C2(n210), .A(n3232), .B(n3229), .ZN(n5531) );
  MUX2_X1 U1932 ( .A(n4949), .B(n4948), .S(n4947), .Z(n5532) );
  OAI21_X1 U1933 ( .B1(n4506), .B2(n4567), .A(n4505), .ZN(n5766) );
  OR2_X1 U1936 ( .A1(n821), .A2(n4652), .ZN(n4873) );
  OAI211_X1 U1937 ( .C1(n4607), .C2(n4153), .A(n1253), .B(n680), .ZN(n733) );
  INV_X1 U1938 ( .A(n6205), .ZN(n287) );
  OR2_X1 U1940 ( .A1(n665), .A2(n4569), .ZN(n643) );
  INV_X1 U1941 ( .A(n19475), .ZN(n288) );
  INV_X1 U1942 ( .A(n5072), .ZN(n828) );
  OR2_X1 U1943 ( .A1(n4681), .A2(n4387), .ZN(n523) );
  AND2_X1 U1944 ( .A1(n4337), .A2(n20487), .ZN(n4535) );
  OR2_X1 U1945 ( .A1(n3624), .A2(n20487), .ZN(n393) );
  OR2_X1 U1947 ( .A1(n3854), .A2(n4674), .ZN(n306) );
  OR2_X1 U1948 ( .A1(n4732), .A2(n3683), .ZN(n3682) );
  AND2_X1 U1949 ( .A1(n4365), .A2(n4013), .ZN(n1535) );
  BUF_X1 U1950 ( .A(n4021), .Z(n4976) );
  OR2_X1 U1951 ( .A1(n896), .A2(n20357), .ZN(n453) );
  OR2_X1 U1953 ( .A1(n5100), .A2(n5101), .ZN(n4049) );
  OR2_X1 U1954 ( .A1(n4652), .A2(n20357), .ZN(n4863) );
  CLKBUF_X1 U1955 ( .A(n3995), .Z(n4387) );
  OR2_X1 U1956 ( .A1(n4548), .A2(n4152), .ZN(n4153) );
  CLKBUF_X1 U1957 ( .A(n4232), .Z(n4902) );
  CLKBUF_X1 U1959 ( .A(n4445), .Z(n4585) );
  OR2_X1 U1961 ( .A1(n4271), .A2(n4268), .ZN(n556) );
  INV_X1 U1962 ( .A(n2233), .ZN(n357) );
  INV_X1 U1963 ( .A(n20355), .ZN(n289) );
  INV_X1 U1964 ( .A(n5079), .ZN(n378) );
  AND2_X1 U1966 ( .A1(n5022), .A2(n19788), .ZN(n315) );
  INV_X1 U1967 ( .A(n4365), .ZN(n290) );
  INV_X1 U1968 ( .A(n4663), .ZN(n291) );
  CLKBUF_X1 U1969 ( .A(n4602), .Z(n4361) );
  OR2_X1 U1970 ( .A1(n4638), .A2(n4528), .ZN(n4636) );
  BUF_X1 U1971 ( .A(n4439), .Z(n5042) );
  CLKBUF_X1 U1972 ( .A(n4187), .Z(n4522) );
  OR2_X1 U1973 ( .A1(n4110), .A2(n4277), .ZN(n672) );
  XNOR2_X1 U1974 ( .A(n1581), .B(Key[76]), .ZN(n4214) );
  OR2_X1 U1975 ( .A1(n20143), .A2(n4285), .ZN(n4630) );
  CLKBUF_X1 U1976 ( .A(n4048), .Z(n5105) );
  AND2_X1 U1977 ( .A1(n4623), .A2(n4626), .ZN(n531) );
  BUF_X1 U1979 ( .A(n4575), .Z(n4372) );
  CLKBUF_X1 U1980 ( .A(Key[183]), .Z(n18997) );
  CLKBUF_X1 U1982 ( .A(Key[190]), .Z(n2035) );
  CLKBUF_X1 U1983 ( .A(Key[176]), .Z(n2382) );
  INV_X1 U1984 ( .A(n4894), .ZN(n292) );
  CLKBUF_X1 U1985 ( .A(Key[136]), .Z(n2417) );
  INV_X1 U1987 ( .A(n2082), .ZN(n293) );
  INV_X1 U1988 ( .A(n1857), .ZN(n294) );
  INV_X1 U1989 ( .A(n2218), .ZN(n295) );
  XNOR2_X1 U1990 ( .A(Key[81]), .B(Plaintext[81]), .ZN(n5117) );
  CLKBUF_X1 U1991 ( .A(Key[50]), .Z(n19457) );
  INV_X1 U1992 ( .A(n18801), .ZN(n296) );
  CLKBUF_X1 U1993 ( .A(Key[1]), .Z(n17787) );
  CLKBUF_X1 U1995 ( .A(Key[22]), .Z(n2275) );
  CLKBUF_X1 U1996 ( .A(Key[165]), .Z(n2381) );
  CLKBUF_X1 U2000 ( .A(Key[95]), .Z(n17989) );
  CLKBUF_X1 U2001 ( .A(Key[81]), .Z(n17024) );
  CLKBUF_X1 U2002 ( .A(Key[53]), .Z(n18146) );
  CLKBUF_X1 U2003 ( .A(Key[99]), .Z(n18308) );
  CLKBUF_X1 U2004 ( .A(Key[97]), .Z(n19410) );
  CLKBUF_X1 U2005 ( .A(Key[177]), .Z(n17686) );
  INV_X1 U2006 ( .A(n17544), .ZN(n298) );
  CLKBUF_X1 U2007 ( .A(Key[184]), .Z(n2401) );
  CLKBUF_X1 U2008 ( .A(Key[132]), .Z(n18809) );
  CLKBUF_X1 U2009 ( .A(Key[79]), .Z(n19180) );
  CLKBUF_X1 U2010 ( .A(Key[139]), .Z(n2383) );
  CLKBUF_X1 U2011 ( .A(Key[160]), .Z(n18819) );
  CLKBUF_X1 U2012 ( .A(Key[13]), .Z(n2455) );
  CLKBUF_X1 U2013 ( .A(Key[65]), .Z(n1840) );
  XNOR2_X1 U2015 ( .A(Key[72]), .B(Plaintext[72]), .ZN(n4829) );
  CLKBUF_X1 U2016 ( .A(Key[59]), .Z(n18078) );
  INV_X1 U2017 ( .A(n2096), .ZN(n299) );
  CLKBUF_X1 U2018 ( .A(Key[174]), .Z(n2108) );
  CLKBUF_X1 U2019 ( .A(Key[180]), .Z(n17637) );
  INV_X1 U2020 ( .A(n17733), .ZN(n300) );
  INV_X1 U2022 ( .A(n4541), .ZN(n301) );
  CLKBUF_X1 U2023 ( .A(Key[164]), .Z(n2384) );
  INV_X1 U2024 ( .A(n1969), .ZN(n302) );
  CLKBUF_X1 U2025 ( .A(Key[189]), .Z(n2420) );
  XNOR2_X1 U2026 ( .A(Key[166]), .B(Plaintext[166]), .ZN(n4349) );
  INV_X1 U2031 ( .A(n4107), .ZN(n303) );
  CLKBUF_X1 U2032 ( .A(Key[42]), .Z(n2216) );
  INV_X1 U2033 ( .A(n16035), .ZN(n304) );
  CLKBUF_X1 U2034 ( .A(Key[7]), .Z(n2423) );
  CLKBUF_X1 U2035 ( .A(Key[28]), .Z(n1911) );
  CLKBUF_X1 U2036 ( .A(Key[98]), .Z(n17791) );
  NAND2_X1 U2038 ( .A1(n4828), .A2(n19688), .ZN(n4674) );
  NOR2_X1 U2039 ( .A1(n14984), .A2(n15180), .ZN(n307) );
  NAND3_X1 U2040 ( .A1(n1822), .A2(n262), .A3(n8121), .ZN(n8122) );
  NOR3_X1 U2041 ( .A1(n12223), .A2(n308), .A3(n10925), .ZN(n12225) );
  INV_X1 U2042 ( .A(n12220), .ZN(n308) );
  AND2_X1 U2043 ( .A1(n8937), .A2(n8729), .ZN(n8942) );
  NAND2_X1 U2044 ( .A1(n8097), .A2(n309), .ZN(n8103) );
  OAI21_X1 U2045 ( .B1(n8210), .B2(n8091), .A(n7631), .ZN(n309) );
  NAND2_X1 U2046 ( .A1(n19724), .A2(n310), .ZN(n18992) );
  OAI21_X1 U2049 ( .B1(n19751), .B2(n19753), .A(n312), .ZN(n17630) );
  NAND2_X1 U2050 ( .A1(n18703), .A2(n18697), .ZN(n312) );
  NAND3_X1 U2052 ( .A1(n3711), .A2(n11218), .A3(n3482), .ZN(n11220) );
  NAND2_X1 U2053 ( .A1(n1142), .A2(n1144), .ZN(n1236) );
  NAND2_X1 U2054 ( .A1(n314), .A2(n1235), .ZN(n11597) );
  NAND2_X1 U2055 ( .A1(n1234), .A2(n245), .ZN(n314) );
  NAND2_X1 U2057 ( .A1(n4581), .A2(n315), .ZN(n4583) );
  INV_X1 U2060 ( .A(n8941), .ZN(n317) );
  NAND2_X1 U2061 ( .A1(n8942), .A2(n8941), .ZN(n318) );
  NAND2_X1 U2063 ( .A1(n321), .A2(n320), .ZN(n319) );
  NAND2_X1 U2064 ( .A1(n20129), .A2(n225), .ZN(n321) );
  OR2_X1 U2066 ( .A1(n5444), .A2(n5641), .ZN(n5640) );
  NAND3_X1 U2067 ( .A1(n3109), .A2(n4610), .A3(n4615), .ZN(n3108) );
  NAND3_X1 U2068 ( .A1(n7601), .A2(n7602), .A3(n8286), .ZN(n2315) );
  OAI21_X2 U2069 ( .B1(n14840), .B2(n14839), .A(n322), .ZN(n16614) );
  OAI21_X1 U2070 ( .B1(n8004), .B2(n324), .A(n323), .ZN(n8009) );
  NAND2_X1 U2071 ( .A1(n281), .A2(n8004), .ZN(n323) );
  NOR2_X1 U2072 ( .A1(n325), .A2(n147), .ZN(n2152) );
  NOR2_X1 U2073 ( .A1(n14652), .A2(n14651), .ZN(n325) );
  NAND2_X1 U2074 ( .A1(n17818), .A2(n18962), .ZN(n326) );
  NAND3_X1 U2075 ( .A1(n4789), .A2(n5092), .A3(n4782), .ZN(n4070) );
  NAND2_X1 U2076 ( .A1(n2460), .A2(n4405), .ZN(n4789) );
  NAND3_X1 U2078 ( .A1(n4604), .A2(n4603), .A3(n4354), .ZN(n4606) );
  NAND2_X1 U2079 ( .A1(n329), .A2(n2281), .ZN(n478) );
  NAND2_X1 U2080 ( .A1(n13955), .A2(n14566), .ZN(n329) );
  NAND2_X1 U2081 ( .A1(n10995), .A2(n10996), .ZN(n10997) );
  NAND2_X1 U2082 ( .A1(n4495), .A2(n4496), .ZN(n4500) );
  NAND3_X1 U2083 ( .A1(n20368), .A2(n6013), .A3(n5921), .ZN(n5516) );
  OAI211_X1 U2084 ( .C1(n245), .C2(n12754), .A(n331), .B(n12389), .ZN(n609) );
  NAND2_X1 U2085 ( .A1(n12410), .A2(n254), .ZN(n331) );
  NAND2_X1 U2086 ( .A1(n12399), .A2(n953), .ZN(n11912) );
  NAND2_X1 U2089 ( .A1(n11336), .A2(n11265), .ZN(n332) );
  NAND2_X1 U2090 ( .A1(n11335), .A2(n11337), .ZN(n333) );
  OAI22_X1 U2091 ( .A1(n252), .A2(n256), .B1(n11673), .B2(n20427), .ZN(n703)
         );
  NAND2_X1 U2092 ( .A1(n7600), .A2(n8033), .ZN(n7602) );
  NAND2_X1 U2094 ( .A1(n4696), .A2(n4795), .ZN(n4029) );
  NAND2_X1 U2096 ( .A1(n7864), .A2(n8153), .ZN(n6698) );
  OAI211_X1 U2097 ( .C1(n9314), .C2(n9313), .A(n9312), .B(n9311), .ZN(n9856)
         );
  XNOR2_X1 U2098 ( .A(n17406), .B(n335), .ZN(n334) );
  NAND3_X1 U2101 ( .A1(n336), .A2(n15467), .A3(n15466), .ZN(n15472) );
  NAND2_X1 U2102 ( .A1(n20502), .A2(n15465), .ZN(n336) );
  OAI21_X1 U2103 ( .B1(n3725), .B2(n15257), .A(n1349), .ZN(n15261) );
  NAND3_X1 U2105 ( .A1(n5465), .A2(n5464), .A3(n5633), .ZN(n5469) );
  NAND2_X1 U2106 ( .A1(n5632), .A2(n5364), .ZN(n5465) );
  NAND2_X1 U2111 ( .A1(n12662), .A2(n12661), .ZN(n338) );
  INV_X1 U2112 ( .A(n339), .ZN(n17499) );
  NOR2_X1 U2114 ( .A1(n20648), .A2(n17504), .ZN(n339) );
  NAND2_X1 U2115 ( .A1(n7766), .A2(n7919), .ZN(n7536) );
  NAND2_X1 U2118 ( .A1(n358), .A2(n7425), .ZN(n7427) );
  NAND2_X1 U2120 ( .A1(n14045), .A2(n14826), .ZN(n340) );
  NAND2_X1 U2121 ( .A1(n14833), .A2(n19859), .ZN(n341) );
  NAND2_X1 U2122 ( .A1(n1955), .A2(n15339), .ZN(n2069) );
  NAND2_X1 U2124 ( .A1(n5435), .A2(n5704), .ZN(n6003) );
  NAND3_X1 U2125 ( .A1(n19916), .A2(n17687), .A3(n18042), .ZN(n17813) );
  NAND3_X1 U2126 ( .A1(n15895), .A2(n19838), .A3(n15896), .ZN(n15897) );
  NAND2_X1 U2127 ( .A1(n5037), .A2(n153), .ZN(n713) );
  XNOR2_X1 U2128 ( .A(n9987), .B(n9947), .ZN(n10417) );
  OAI21_X1 U2129 ( .B1(n18223), .B2(n18977), .A(n342), .ZN(n16911) );
  NAND2_X1 U2130 ( .A1(n224), .A2(n18977), .ZN(n342) );
  OAI21_X1 U2131 ( .B1(n684), .B2(n11726), .A(n683), .ZN(n682) );
  NAND2_X1 U2132 ( .A1(n1177), .A2(n14954), .ZN(n14743) );
  NAND2_X1 U2134 ( .A1(n12250), .A2(n12573), .ZN(n541) );
  NAND2_X1 U2137 ( .A1(n6100), .A2(n283), .ZN(n343) );
  NAND2_X1 U2138 ( .A1(n5663), .A2(n5952), .ZN(n6100) );
  NAND2_X1 U2141 ( .A1(n11364), .A2(n2765), .ZN(n344) );
  OR2_X1 U2142 ( .A1(n8386), .A2(n8132), .ZN(n2441) );
  XNOR2_X1 U2143 ( .A(n10593), .B(n10592), .ZN(n3051) );
  INV_X1 U2144 ( .A(n5428), .ZN(n5797) );
  NAND2_X1 U2145 ( .A1(n5338), .A2(n6124), .ZN(n1382) );
  AND2_X2 U2146 ( .A1(n1051), .A2(n1050), .ZN(n6124) );
  NAND2_X1 U2147 ( .A1(n19476), .A2(n6379), .ZN(n5844) );
  NAND3_X1 U2149 ( .A1(n6056), .A2(n20670), .A3(n5785), .ZN(n5305) );
  NAND2_X1 U2151 ( .A1(n346), .A2(n2618), .ZN(n2617) );
  NAND2_X1 U2152 ( .A1(n9174), .A2(n9175), .ZN(n346) );
  NAND3_X1 U2153 ( .A1(n820), .A2(n8202), .A3(n8201), .ZN(n8207) );
  NAND3_X1 U2154 ( .A1(n3532), .A2(n14600), .A3(n20181), .ZN(n1824) );
  NAND3_X1 U2155 ( .A1(n3410), .A2(n5931), .A3(n5930), .ZN(n5932) );
  NAND2_X1 U2157 ( .A1(n14866), .A2(n15684), .ZN(n15226) );
  NAND2_X1 U2159 ( .A1(n9874), .A2(n11230), .ZN(n348) );
  NAND2_X1 U2161 ( .A1(n1987), .A2(n1183), .ZN(n350) );
  NAND3_X1 U2163 ( .A1(n6844), .A2(n279), .A3(n7852), .ZN(n6845) );
  NOR2_X1 U2164 ( .A1(n351), .A2(n18504), .ZN(n1660) );
  AOI21_X1 U2165 ( .B1(n18518), .B2(n18511), .A(n18512), .ZN(n351) );
  AOI22_X1 U2166 ( .A1(n11835), .A2(n12506), .B1(n12507), .B2(n12505), .ZN(
        n11840) );
  NOR2_X1 U2167 ( .A1(n390), .A2(n12642), .ZN(n389) );
  NAND2_X1 U2168 ( .A1(n352), .A2(n9564), .ZN(n9193) );
  NAND2_X1 U2169 ( .A1(n9338), .A2(n352), .ZN(n8155) );
  XNOR2_X1 U2171 ( .A(n353), .B(n6793), .ZN(n7089) );
  XNOR2_X1 U2172 ( .A(n354), .B(n7088), .ZN(n6722) );
  NAND2_X1 U2173 ( .A1(n5850), .A2(n5849), .ZN(n355) );
  NAND2_X1 U2174 ( .A1(n356), .A2(n244), .ZN(n12018) );
  NAND2_X1 U2175 ( .A1(n242), .A2(n356), .ZN(n542) );
  INV_X1 U2176 ( .A(n358), .ZN(n7859) );
  NAND2_X1 U2178 ( .A1(n359), .A2(n9559), .ZN(n3489) );
  NAND2_X1 U2179 ( .A1(n2734), .A2(n10996), .ZN(n359) );
  INV_X1 U2180 ( .A(n1640), .ZN(n360) );
  NAND2_X1 U2181 ( .A1(n15397), .A2(n361), .ZN(n15064) );
  AND3_X2 U2182 ( .A1(n3267), .A2(n3266), .A3(n3268), .ZN(n15311) );
  OAI21_X1 U2183 ( .B1(n8439), .B2(n2499), .A(n364), .ZN(n362) );
  AOI21_X1 U2184 ( .B1(n365), .B2(n8337), .A(n9144), .ZN(n363) );
  NAND2_X1 U2185 ( .A1(n9145), .A2(n2499), .ZN(n364) );
  NAND2_X1 U2186 ( .A1(n8338), .A2(n8786), .ZN(n365) );
  NAND2_X1 U2187 ( .A1(n8338), .A2(n2499), .ZN(n8337) );
  NAND2_X1 U2188 ( .A1(n6105), .A2(n6109), .ZN(n368) );
  NAND2_X1 U2189 ( .A1(n1623), .A2(n368), .ZN(n1620) );
  NOR2_X1 U2193 ( .A1(n5957), .A2(n368), .ZN(n367) );
  NAND2_X1 U2195 ( .A1(n12502), .A2(n12004), .ZN(n12345) );
  NAND2_X1 U2197 ( .A1(n19999), .A2(n11521), .ZN(n370) );
  NAND3_X1 U2199 ( .A1(n372), .A2(n1446), .A3(n10930), .ZN(n371) );
  NAND2_X1 U2200 ( .A1(n10889), .A2(n11550), .ZN(n10930) );
  NAND2_X1 U2201 ( .A1(n10068), .A2(n11544), .ZN(n372) );
  NAND2_X1 U2202 ( .A1(n374), .A2(n646), .ZN(n373) );
  NAND2_X1 U2203 ( .A1(n648), .A2(n647), .ZN(n374) );
  INV_X1 U2204 ( .A(n4349), .ZN(n4199) );
  NAND2_X1 U2205 ( .A1(n4349), .A2(n4541), .ZN(n4536) );
  XNOR2_X2 U2206 ( .A(Key[167]), .B(Plaintext[167]), .ZN(n4541) );
  NAND2_X1 U2207 ( .A1(n15766), .A2(n15474), .ZN(n12664) );
  NAND3_X1 U2208 ( .A1(n15766), .A2(n15474), .A3(n15769), .ZN(n375) );
  NAND3_X1 U2209 ( .A1(n7916), .A2(n377), .A3(n376), .ZN(n9143) );
  NAND2_X1 U2210 ( .A1(n8910), .A2(n7956), .ZN(n1231) );
  NAND2_X1 U2211 ( .A1(n20431), .A2(n378), .ZN(n4083) );
  OAI21_X1 U2212 ( .B1(n378), .B2(n5074), .A(n4809), .ZN(n4084) );
  NAND2_X1 U2213 ( .A1(n4810), .A2(n378), .ZN(n1047) );
  NAND2_X2 U2214 ( .A1(n379), .A2(n14033), .ZN(n15760) );
  NAND2_X1 U2215 ( .A1(n14301), .A2(n14512), .ZN(n379) );
  NAND2_X1 U2216 ( .A1(n13986), .A2(n2972), .ZN(n14301) );
  NAND4_X2 U2217 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n7128)
         );
  NAND2_X1 U2220 ( .A1(n10784), .A2(n11435), .ZN(n382) );
  NAND2_X1 U2221 ( .A1(n5664), .A2(n5949), .ZN(n5458) );
  NOR3_X1 U2222 ( .A1(n9296), .A2(n9300), .A3(n9295), .ZN(n2225) );
  OAI21_X1 U2224 ( .B1(n8297), .B2(n20485), .A(n383), .ZN(n7582) );
  NAND2_X1 U2225 ( .A1(n7581), .A2(n8297), .ZN(n383) );
  AOI22_X1 U2227 ( .A1(n19166), .A2(n19165), .B1(n386), .B2(n19948), .ZN(
        n19167) );
  NAND2_X1 U2228 ( .A1(n19161), .A2(n150), .ZN(n386) );
  OR2_X2 U2229 ( .A1(n1967), .A2(n7423), .ZN(n9018) );
  NAND2_X1 U2230 ( .A1(n439), .A2(n387), .ZN(n15735) );
  INV_X1 U2233 ( .A(n12639), .ZN(n390) );
  NAND2_X1 U2234 ( .A1(n8682), .A2(n9149), .ZN(n392) );
  NAND2_X1 U2237 ( .A1(n1525), .A2(n15148), .ZN(n15149) );
  OAI21_X1 U2238 ( .B1(n9211), .B2(n263), .A(n394), .ZN(n8448) );
  NAND2_X1 U2239 ( .A1(n9211), .A2(n8444), .ZN(n394) );
  XNOR2_X1 U2241 ( .A(n395), .B(n9787), .ZN(n9789) );
  XNOR2_X1 U2242 ( .A(n9788), .B(n10387), .ZN(n395) );
  AOI21_X1 U2243 ( .B1(n17982), .B2(n18238), .A(n396), .ZN(n3208) );
  INV_X1 U2244 ( .A(n17981), .ZN(n396) );
  OAI22_X1 U2246 ( .A1(n19385), .A2(n17221), .B1(n17218), .B2(n19383), .ZN(
        n19387) );
  NAND3_X1 U2247 ( .A1(n4739), .A2(n5059), .A3(n5060), .ZN(n4102) );
  OR2_X2 U2248 ( .A1(n4103), .A2(n4104), .ZN(n5985) );
  OR2_X1 U2250 ( .A1(n8296), .A2(n8299), .ZN(n397) );
  NOR2_X1 U2251 ( .A1(n20000), .A2(n9107), .ZN(n8555) );
  AOI21_X2 U2252 ( .B1(n12506), .B2(n9887), .A(n398), .ZN(n13746) );
  OAI22_X1 U2253 ( .A1(n9885), .A2(n12506), .B1(n9886), .B2(n12008), .ZN(n398)
         );
  OAI21_X2 U2254 ( .B1(n8130), .B2(n8129), .A(n399), .ZN(n9999) );
  OAI211_X1 U2255 ( .C1(n8127), .C2(n8128), .A(n1651), .B(n8889), .ZN(n399) );
  NOR2_X2 U2256 ( .A1(n8724), .A2(n8725), .ZN(n10273) );
  MUX2_X1 U2257 ( .A(n7724), .B(n8161), .S(n8160), .Z(n8164) );
  NAND2_X1 U2258 ( .A1(n7855), .A2(n8157), .ZN(n8160) );
  NOR2_X1 U2259 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  NAND2_X1 U2260 ( .A1(n3959), .A2(n3960), .ZN(n5583) );
  NAND2_X1 U2262 ( .A1(n15373), .A2(n548), .ZN(n16996) );
  XNOR2_X1 U2263 ( .A(n400), .B(n18985), .ZN(Ciphertext[108]) );
  NAND2_X1 U2264 ( .A1(n2050), .A2(n18983), .ZN(n400) );
  OAI211_X1 U2265 ( .C1(n6439), .C2(n8128), .A(n401), .B(n9090), .ZN(n6440) );
  NAND3_X1 U2268 ( .A1(n1118), .A2(n17913), .A3(n17914), .ZN(n403) );
  OAI21_X1 U2270 ( .B1(n650), .B2(n11423), .A(n2440), .ZN(n12524) );
  XNOR2_X1 U2271 ( .A(n403), .B(n302), .ZN(Ciphertext[24]) );
  OR2_X1 U2272 ( .A1(n4306), .A2(n4305), .ZN(n4004) );
  XNOR2_X1 U2273 ( .A(n405), .B(n17783), .ZN(Ciphertext[87]) );
  NAND3_X1 U2274 ( .A1(n2219), .A2(n2177), .A3(n17782), .ZN(n405) );
  NAND2_X1 U2277 ( .A1(n3770), .A2(n410), .ZN(n409) );
  OR2_X1 U2278 ( .A1(n4233), .A2(n4856), .ZN(n410) );
  NAND3_X1 U2279 ( .A1(n412), .A2(n4153), .A3(n4607), .ZN(n4154) );
  NAND2_X1 U2280 ( .A1(n4546), .A2(n4603), .ZN(n412) );
  NOR2_X1 U2281 ( .A1(n5581), .A2(n733), .ZN(n5000) );
  OAI21_X1 U2285 ( .B1(n415), .B2(n249), .A(n12002), .ZN(n2260) );
  NAND3_X1 U2287 ( .A1(n1687), .A2(n2465), .A3(n5145), .ZN(n6674) );
  NAND2_X1 U2288 ( .A1(n416), .A2(n7963), .ZN(n7966) );
  NAND2_X1 U2289 ( .A1(n208), .A2(n7801), .ZN(n416) );
  OAI21_X1 U2290 ( .B1(n14131), .B2(n15606), .A(n417), .ZN(n14139) );
  OR2_X1 U2293 ( .A1(n10673), .A2(n10194), .ZN(n11341) );
  NAND3_X2 U2294 ( .A1(n419), .A2(n3107), .A3(n3106), .ZN(n10229) );
  NAND3_X1 U2296 ( .A1(n14728), .A2(n14731), .A3(n14224), .ZN(n420) );
  OAI211_X1 U2297 ( .C1(n12347), .C2(n201), .A(n421), .B(n12346), .ZN(n12348)
         );
  NAND2_X1 U2298 ( .A1(n12345), .A2(n201), .ZN(n421) );
  OR3_X1 U2299 ( .A1(n3366), .A2(n14666), .A3(n14663), .ZN(n14037) );
  NAND2_X1 U2300 ( .A1(n806), .A2(n5495), .ZN(n805) );
  AND3_X2 U2301 ( .A1(n422), .A2(n1307), .A3(n1306), .ZN(n13275) );
  NAND2_X1 U2302 ( .A1(n10366), .A2(n11451), .ZN(n422) );
  NAND2_X1 U2303 ( .A1(n9028), .A2(n9031), .ZN(n9034) );
  NAND2_X1 U2304 ( .A1(n2504), .A2(n8545), .ZN(n544) );
  OAI21_X1 U2305 ( .B1(n8263), .B2(n8262), .A(n423), .ZN(n8265) );
  NAND2_X1 U2306 ( .A1(n8263), .A2(n895), .ZN(n423) );
  NAND3_X1 U2307 ( .A1(n10705), .A2(n10708), .A3(n10953), .ZN(n2045) );
  NAND2_X1 U2308 ( .A1(n20470), .A2(n10952), .ZN(n10705) );
  NAND2_X1 U2309 ( .A1(n18101), .A2(n19774), .ZN(n424) );
  NAND2_X1 U2310 ( .A1(n14998), .A2(n15835), .ZN(n15001) );
  OAI211_X2 U2311 ( .C1(n12515), .C2(n1305), .A(n2491), .B(n1304), .ZN(n13136)
         );
  XNOR2_X2 U2312 ( .A(n425), .B(Key[93]), .ZN(n5093) );
  INV_X1 U2313 ( .A(Plaintext[93]), .ZN(n425) );
  NAND2_X1 U2319 ( .A1(n7418), .A2(n19901), .ZN(n429) );
  NAND2_X1 U2320 ( .A1(n9243), .A2(n430), .ZN(n8715) );
  NAND2_X1 U2321 ( .A1(n431), .A2(n1777), .ZN(n430) );
  OR2_X1 U2323 ( .A1(n7584), .A2(n2548), .ZN(n7588) );
  OR2_X1 U2324 ( .A1(n4667), .A2(n19688), .ZN(n4672) );
  AND2_X1 U2325 ( .A1(n18094), .A2(n18096), .ZN(n759) );
  NAND3_X1 U2326 ( .A1(n4026), .A2(n4027), .A3(n20464), .ZN(n432) );
  NAND2_X1 U2327 ( .A1(n4029), .A2(n4698), .ZN(n434) );
  NAND2_X1 U2328 ( .A1(n15564), .A2(n232), .ZN(n435) );
  AOI22_X1 U2329 ( .A1(n14741), .A2(n14740), .B1(n14739), .B2(n14738), .ZN(
        n14952) );
  NAND2_X1 U2330 ( .A1(n9163), .A2(n437), .ZN(n436) );
  INV_X1 U2331 ( .A(n12430), .ZN(n3649) );
  XNOR2_X1 U2332 ( .A(n6415), .B(n6414), .ZN(n7750) );
  OR2_X1 U2333 ( .A1(n8353), .A2(n8352), .ZN(n823) );
  OAI211_X1 U2335 ( .C1(n1334), .C2(n803), .A(n1333), .B(n3454), .ZN(n9748) );
  NAND2_X1 U2336 ( .A1(n747), .A2(n16126), .ZN(n439) );
  INV_X1 U2337 ( .A(n14410), .ZN(n14132) );
  AND2_X1 U2338 ( .A1(n236), .A2(n14410), .ZN(n14223) );
  OAI211_X1 U2340 ( .C1(n18472), .C2(n18471), .A(n18470), .B(n440), .ZN(n18474) );
  NAND3_X1 U2341 ( .A1(n18466), .A2(n20110), .A3(n20148), .ZN(n440) );
  OR2_X1 U2342 ( .A1(n20451), .A2(n14410), .ZN(n14134) );
  NAND3_X1 U2343 ( .A1(n11275), .A2(n10684), .A3(n11271), .ZN(n11249) );
  AND2_X1 U2346 ( .A1(n11428), .A2(n11106), .ZN(n10769) );
  NAND2_X1 U2347 ( .A1(n17817), .A2(n227), .ZN(n443) );
  NAND2_X1 U2348 ( .A1(n18966), .A2(n18968), .ZN(n17817) );
  NAND2_X1 U2349 ( .A1(n18965), .A2(n20127), .ZN(n444) );
  NAND2_X1 U2352 ( .A1(n5316), .A2(n3533), .ZN(n446) );
  NAND2_X2 U2353 ( .A1(n447), .A2(n7004), .ZN(n9046) );
  NAND3_X1 U2355 ( .A1(n16010), .A2(n15333), .A3(n13968), .ZN(n527) );
  OAI21_X1 U2356 ( .B1(n5078), .B2(n5077), .A(n448), .ZN(n5503) );
  NAND2_X1 U2357 ( .A1(n2162), .A2(n11418), .ZN(n2161) );
  NAND3_X1 U2358 ( .A1(n12685), .A2(n1091), .A3(n12686), .ZN(n1092) );
  OR3_X1 U2359 ( .A1(n7754), .A2(n7530), .A3(n7903), .ZN(n644) );
  NAND2_X1 U2360 ( .A1(n7998), .A2(n1425), .ZN(n449) );
  NAND2_X1 U2363 ( .A1(n8256), .A2(n8258), .ZN(n7726) );
  NAND2_X1 U2365 ( .A1(n3133), .A2(n3134), .ZN(n2680) );
  INV_X1 U2366 ( .A(n15094), .ZN(n451) );
  AND2_X2 U2367 ( .A1(n451), .A2(n149), .ZN(n17035) );
  NAND3_X1 U2369 ( .A1(n4867), .A2(n2072), .A3(n453), .ZN(n452) );
  NAND2_X1 U2370 ( .A1(n11712), .A2(n454), .ZN(n13138) );
  OR2_X1 U2371 ( .A1(n11713), .A2(n12155), .ZN(n454) );
  OAI21_X1 U2372 ( .B1(n10789), .B2(n10788), .A(n10787), .ZN(n12636) );
  NAND2_X1 U2374 ( .A1(n4632), .A2(n455), .ZN(n5179) );
  OR2_X1 U2375 ( .A1(n8411), .A2(n655), .ZN(n9183) );
  NOR2_X1 U2376 ( .A1(n3468), .A2(n5985), .ZN(n5438) );
  XNOR2_X1 U2377 ( .A(n10600), .B(n9860), .ZN(n550) );
  XNOR2_X2 U2378 ( .A(n7214), .B(n7215), .ZN(n8004) );
  NAND2_X1 U2379 ( .A1(n4652), .A2(n4867), .ZN(n3562) );
  NAND3_X1 U2382 ( .A1(n11962), .A2(n2140), .A3(n2139), .ZN(n458) );
  INV_X1 U2385 ( .A(n8289), .ZN(n462) );
  NAND2_X1 U2386 ( .A1(n7468), .A2(n7807), .ZN(n463) );
  NAND2_X1 U2387 ( .A1(n1658), .A2(n464), .ZN(n9011) );
  OAI211_X2 U2389 ( .C1(n7819), .C2(n7818), .A(n7817), .B(n465), .ZN(n8895) );
  NAND3_X1 U2390 ( .A1(n466), .A2(n8379), .A3(n8378), .ZN(n8445) );
  NAND3_X1 U2391 ( .A1(n8371), .A2(n8369), .A3(n8370), .ZN(n466) );
  NOR2_X2 U2393 ( .A1(n7490), .A2(n467), .ZN(n9122) );
  AOI21_X1 U2394 ( .B1(n7489), .B2(n7488), .A(n22), .ZN(n467) );
  XNOR2_X1 U2395 ( .A(n20018), .B(n13527), .ZN(n12367) );
  OAI21_X1 U2397 ( .B1(n5345), .B2(n6139), .A(n469), .ZN(n6724) );
  NAND2_X1 U2398 ( .A1(n5343), .A2(n5344), .ZN(n469) );
  XNOR2_X1 U2399 ( .A(n470), .B(n790), .ZN(n8777) );
  XNOR2_X1 U2400 ( .A(n8776), .B(n10030), .ZN(n470) );
  NAND2_X1 U2401 ( .A1(n5593), .A2(n5590), .ZN(n5591) );
  NAND2_X1 U2402 ( .A1(n8950), .A2(n8603), .ZN(n9367) );
  NAND2_X1 U2403 ( .A1(n2070), .A2(n1882), .ZN(n3981) );
  NAND2_X1 U2405 ( .A1(n472), .A2(n471), .ZN(n4001) );
  NAND2_X1 U2406 ( .A1(n3993), .A2(n6068), .ZN(n471) );
  NAND2_X1 U2407 ( .A1(n3992), .A2(n473), .ZN(n472) );
  NAND2_X1 U2408 ( .A1(n12473), .A2(n12142), .ZN(n12393) );
  AOI21_X2 U2409 ( .B1(n8351), .B2(n7549), .A(n2778), .ZN(n8960) );
  AOI22_X1 U2410 ( .A1(n9369), .A2(n904), .B1(n9370), .B2(n9371), .ZN(n9373)
         );
  NOR2_X1 U2412 ( .A1(n14590), .A2(n19781), .ZN(n474) );
  AOI22_X1 U2414 ( .A1(n3250), .A2(n8141), .B1(n8270), .B2(n8350), .ZN(n475)
         );
  NAND2_X1 U2415 ( .A1(n12591), .A2(n12589), .ZN(n12596) );
  NAND2_X1 U2416 ( .A1(n15395), .A2(n14990), .ZN(n3247) );
  OR2_X1 U2417 ( .A1(n12658), .A2(n15657), .ZN(n546) );
  NAND2_X1 U2422 ( .A1(n7529), .A2(n274), .ZN(n477) );
  NOR2_X1 U2423 ( .A1(n13318), .A2(n478), .ZN(n15672) );
  NOR2_X1 U2426 ( .A1(n479), .A2(n17748), .ZN(n780) );
  AND2_X1 U2427 ( .A1(n18028), .A2(n17749), .ZN(n479) );
  OAI22_X1 U2428 ( .A1(n10688), .A2(n19851), .B1(n9547), .B2(n11277), .ZN(
        n11276) );
  OAI211_X1 U2429 ( .C1(n5745), .C2(n5741), .A(n20509), .B(n481), .ZN(n480) );
  NAND2_X1 U2430 ( .A1(n5741), .A2(n286), .ZN(n481) );
  XNOR2_X1 U2431 ( .A(n19844), .B(n16429), .ZN(n14163) );
  NAND2_X1 U2435 ( .A1(n2541), .A2(n14277), .ZN(n1409) );
  OAI21_X1 U2441 ( .B1(n2320), .B2(n12147), .A(n12149), .ZN(n485) );
  NAND2_X1 U2443 ( .A1(n486), .A2(n4334), .ZN(n6165) );
  NAND2_X1 U2444 ( .A1(n4333), .A2(n5632), .ZN(n486) );
  NAND2_X1 U2445 ( .A1(n15550), .A2(n15056), .ZN(n14979) );
  NAND2_X1 U2448 ( .A1(n11660), .A2(n11951), .ZN(n487) );
  NAND2_X1 U2449 ( .A1(n19248), .A2(n3345), .ZN(n17667) );
  NOR2_X2 U2450 ( .A1(n13998), .A2(n13999), .ZN(n15701) );
  NAND2_X1 U2451 ( .A1(n8263), .A2(n8262), .ZN(n8106) );
  NAND2_X1 U2453 ( .A1(n490), .A2(n489), .ZN(n18861) );
  NAND2_X1 U2454 ( .A1(n18860), .A2(n216), .ZN(n489) );
  NAND2_X1 U2455 ( .A1(n18859), .A2(n18869), .ZN(n490) );
  NAND2_X1 U2457 ( .A1(n492), .A2(n491), .ZN(n11947) );
  NAND2_X1 U2458 ( .A1(n11946), .A2(n20457), .ZN(n492) );
  NAND2_X1 U2459 ( .A1(n6272), .A2(n494), .ZN(n493) );
  NAND3_X1 U2461 ( .A1(n1812), .A2(n11452), .A3(n11455), .ZN(n10733) );
  XNOR2_X2 U2462 ( .A(n16759), .B(n16758), .ZN(n18954) );
  NAND3_X1 U2464 ( .A1(n14675), .A2(n13981), .A3(n14674), .ZN(n687) );
  OAI22_X1 U2465 ( .A1(n15475), .A2(n15244), .B1(n15656), .B2(n15243), .ZN(
        n14859) );
  NAND2_X1 U2466 ( .A1(n15658), .A2(n15474), .ZN(n15244) );
  INV_X1 U2467 ( .A(n496), .ZN(n495) );
  OAI21_X1 U2468 ( .B1(n5713), .B2(n5985), .A(n5712), .ZN(n496) );
  NAND2_X1 U2469 ( .A1(n5710), .A2(n5986), .ZN(n497) );
  NAND2_X1 U2470 ( .A1(n12606), .A2(n3305), .ZN(n11628) );
  NAND3_X2 U2471 ( .A1(n1893), .A2(n1892), .A3(n10892), .ZN(n12606) );
  INV_X1 U2475 ( .A(n8070), .ZN(n8204) );
  NAND2_X1 U2476 ( .A1(n4633), .A2(n20487), .ZN(n4156) );
  NOR2_X1 U2477 ( .A1(n12528), .A2(n12525), .ZN(n12526) );
  NAND2_X1 U2478 ( .A1(n182), .A2(n12523), .ZN(n12525) );
  AND2_X1 U2479 ( .A1(n1907), .A2(n17886), .ZN(n17600) );
  XNOR2_X1 U2480 ( .A(n13711), .B(n13659), .ZN(n12079) );
  AND2_X1 U2483 ( .A1(n11154), .A2(n1580), .ZN(n532) );
  NOR3_X1 U2486 ( .A1(n10979), .A2(n19506), .A3(n10982), .ZN(n10984) );
  XNOR2_X1 U2487 ( .A(n16568), .B(n17433), .ZN(n17135) );
  INV_X1 U2490 ( .A(n11168), .ZN(n11533) );
  NAND2_X1 U2491 ( .A1(n11337), .A2(n11267), .ZN(n755) );
  XNOR2_X1 U2492 ( .A(n657), .B(n18177), .ZN(n6832) );
  NAND2_X1 U2493 ( .A1(n4405), .A2(n5093), .ZN(n5096) );
  NAND2_X1 U2494 ( .A1(n2234), .A2(n2235), .ZN(n11922) );
  AND2_X1 U2497 ( .A1(n9559), .A2(n19779), .ZN(n11287) );
  NAND2_X1 U2498 ( .A1(n4901), .A2(n4492), .ZN(n4494) );
  NAND2_X1 U2499 ( .A1(n504), .A2(n502), .ZN(n1725) );
  NAND2_X1 U2501 ( .A1(n7536), .A2(n505), .ZN(n504) );
  NAND3_X1 U2503 ( .A1(n9368), .A2(n8953), .A3(n8952), .ZN(n506) );
  OAI22_X1 U2505 ( .A1(n3598), .A2(n3167), .B1(n5107), .B2(n507), .ZN(n3166)
         );
  NAND2_X1 U2506 ( .A1(n5099), .A2(n4048), .ZN(n507) );
  NAND2_X1 U2507 ( .A1(n1338), .A2(n11574), .ZN(n11576) );
  NAND2_X1 U2508 ( .A1(n5326), .A2(n508), .ZN(n4284) );
  NAND2_X1 U2509 ( .A1(n510), .A2(n509), .ZN(n12275) );
  NAND2_X1 U2511 ( .A1(n11551), .A2(n11550), .ZN(n510) );
  NAND2_X1 U2512 ( .A1(n12030), .A2(n12304), .ZN(n512) );
  NAND2_X1 U2513 ( .A1(n12031), .A2(n11782), .ZN(n513) );
  NAND2_X1 U2516 ( .A1(n14506), .A2(n14305), .ZN(n13507) );
  NAND2_X1 U2518 ( .A1(n19113), .A2(n19112), .ZN(n19120) );
  OAI21_X1 U2520 ( .B1(n5951), .B2(n5950), .A(n5949), .ZN(n515) );
  OR3_X1 U2522 ( .A1(n5796), .A2(n5795), .A3(n5300), .ZN(n5794) );
  NAND2_X1 U2523 ( .A1(n551), .A2(n516), .ZN(n13231) );
  NAND2_X1 U2524 ( .A1(n11624), .A2(n12441), .ZN(n516) );
  NAND2_X1 U2526 ( .A1(n5407), .A2(n517), .ZN(n6404) );
  OR2_X1 U2527 ( .A1(n5409), .A2(n5408), .ZN(n517) );
  OAI21_X1 U2528 ( .B1(n239), .B2(n19781), .A(n518), .ZN(n14200) );
  NAND2_X1 U2529 ( .A1(n19781), .A2(n14811), .ZN(n518) );
  NAND3_X2 U2531 ( .A1(n2452), .A2(n537), .A3(n536), .ZN(n10247) );
  NAND2_X1 U2533 ( .A1(n2373), .A2(n921), .ZN(n519) );
  NAND2_X1 U2534 ( .A1(n520), .A2(n828), .ZN(n827) );
  NAND2_X1 U2535 ( .A1(n575), .A2(n829), .ZN(n520) );
  NAND2_X1 U2536 ( .A1(n522), .A2(n521), .ZN(n10630) );
  NAND2_X1 U2537 ( .A1(n12325), .A2(n12514), .ZN(n522) );
  INV_X1 U2539 ( .A(n15333), .ZN(n1817) );
  NAND2_X1 U2540 ( .A1(n15879), .A2(n15153), .ZN(n15333) );
  OR2_X2 U2542 ( .A1(n9554), .A2(n9553), .ZN(n11598) );
  NOR2_X1 U2543 ( .A1(n12974), .A2(n3820), .ZN(n12975) );
  NAND2_X1 U2545 ( .A1(n7797), .A2(n7466), .ZN(n7963) );
  NAND2_X1 U2547 ( .A1(n1090), .A2(n14837), .ZN(n14840) );
  OAI211_X2 U2548 ( .C1(n10317), .C2(n10316), .A(n525), .B(n524), .ZN(n13352)
         );
  NAND2_X1 U2549 ( .A1(n10313), .A2(n12336), .ZN(n524) );
  NAND2_X1 U2550 ( .A1(n10315), .A2(n10314), .ZN(n525) );
  XNOR2_X1 U2551 ( .A(n526), .B(n2145), .ZN(n11113) );
  XNOR2_X1 U2552 ( .A(n10371), .B(n10370), .ZN(n526) );
  INV_X1 U2553 ( .A(n4714), .ZN(n5097) );
  OAI22_X1 U2554 ( .A1(n3804), .A2(n5891), .B1(n20670), .B2(n3249), .ZN(n5893)
         );
  NAND2_X1 U2555 ( .A1(n2217), .A2(n3662), .ZN(n1989) );
  NAND2_X1 U2558 ( .A1(n527), .A2(n15154), .ZN(n15155) );
  XNOR2_X2 U2560 ( .A(n9736), .B(n9737), .ZN(n11395) );
  OR2_X1 U2561 ( .A1(n5093), .A2(n4405), .ZN(n4782) );
  NOR2_X1 U2562 ( .A1(n12366), .A2(n12365), .ZN(n915) );
  OAI22_X1 U2564 ( .A1(n8944), .A2(n8945), .B1(n8947), .B2(n8946), .ZN(n528)
         );
  NAND2_X1 U2565 ( .A1(n5093), .A2(n5098), .ZN(n4714) );
  AOI21_X2 U2566 ( .B1(n15001), .B2(n15831), .A(n15000), .ZN(n16706) );
  INV_X1 U2567 ( .A(n14626), .ZN(n14192) );
  XNOR2_X1 U2568 ( .A(n11901), .B(n11900), .ZN(n14626) );
  OAI21_X1 U2569 ( .B1(n4349), .B2(n301), .A(n4540), .ZN(n3932) );
  NAND2_X1 U2570 ( .A1(n17977), .A2(n17758), .ZN(n17762) );
  NAND3_X1 U2572 ( .A1(n637), .A2(n9054), .A3(n9306), .ZN(n529) );
  AOI21_X1 U2574 ( .B1(n3056), .B2(n13682), .A(n13963), .ZN(n530) );
  NAND2_X1 U2575 ( .A1(n5394), .A2(n5395), .ZN(n5326) );
  NAND2_X1 U2576 ( .A1(n4167), .A2(n531), .ZN(n4017) );
  OR3_X1 U2577 ( .A1(n17480), .A2(n20354), .A3(n17479), .ZN(n17485) );
  AOI21_X2 U2578 ( .B1(n1971), .B2(n3382), .A(n532), .ZN(n12280) );
  NAND2_X1 U2579 ( .A1(n534), .A2(n533), .ZN(n5253) );
  NAND2_X1 U2580 ( .A1(n5252), .A2(n5323), .ZN(n534) );
  NAND2_X1 U2581 ( .A1(n3457), .A2(n15245), .ZN(n12663) );
  NAND2_X1 U2582 ( .A1(n8290), .A2(n20189), .ZN(n7370) );
  OAI21_X1 U2583 ( .B1(n5792), .B2(n1026), .A(n535), .ZN(n5157) );
  NAND2_X1 U2584 ( .A1(n5792), .A2(n5156), .ZN(n535) );
  NAND2_X1 U2585 ( .A1(n8800), .A2(n8799), .ZN(n536) );
  NAND2_X1 U2586 ( .A1(n908), .A2(n8798), .ZN(n537) );
  NAND2_X1 U2587 ( .A1(n539), .A2(n16364), .ZN(n18556) );
  OAI21_X1 U2588 ( .B1(n17966), .B2(n16363), .A(n18112), .ZN(n539) );
  NOR2_X1 U2589 ( .A1(n8468), .A2(n8467), .ZN(n9647) );
  OAI211_X1 U2590 ( .C1(n3373), .C2(n20424), .A(n2402), .B(n14020), .ZN(n688)
         );
  XNOR2_X1 U2591 ( .A(n540), .B(n12679), .ZN(n12681) );
  XNOR2_X1 U2592 ( .A(n12680), .B(n13018), .ZN(n540) );
  NAND2_X1 U2593 ( .A1(n10896), .A2(n10745), .ZN(n10059) );
  NAND2_X1 U2596 ( .A1(n12534), .A2(n12162), .ZN(n11804) );
  NOR2_X1 U2597 ( .A1(n8547), .A2(n8546), .ZN(n872) );
  NAND2_X1 U2598 ( .A1(n544), .A2(n543), .ZN(n8546) );
  NAND2_X1 U2599 ( .A1(n8544), .A2(n2749), .ZN(n543) );
  INV_X1 U2600 ( .A(n11133), .ZN(n650) );
  NAND2_X1 U2602 ( .A1(n4622), .A2(n4285), .ZN(n4167) );
  NOR2_X2 U2603 ( .A1(n14560), .A2(n14561), .ZN(n15644) );
  AND2_X2 U2606 ( .A1(n1132), .A2(n1133), .ZN(n12359) );
  NAND3_X1 U2607 ( .A1(n749), .A2(n748), .A3(n4610), .ZN(n762) );
  NAND2_X1 U2608 ( .A1(n20146), .A2(n9204), .ZN(n771) );
  INV_X1 U2610 ( .A(Plaintext[188]), .ZN(n547) );
  NAND2_X1 U2611 ( .A1(n549), .A2(n232), .ZN(n548) );
  INV_X1 U2612 ( .A(n15374), .ZN(n549) );
  NAND2_X1 U2614 ( .A1(n11623), .A2(n12442), .ZN(n552) );
  NAND2_X1 U2615 ( .A1(n11622), .A2(n1522), .ZN(n553) );
  AOI21_X1 U2616 ( .B1(n11540), .B2(n11541), .A(n11539), .ZN(n11542) );
  NAND2_X1 U2618 ( .A1(n5708), .A2(n5815), .ZN(n5816) );
  NAND2_X1 U2619 ( .A1(n557), .A2(n554), .ZN(n4273) );
  NAND2_X1 U2620 ( .A1(n555), .A2(n4765), .ZN(n554) );
  NAND2_X1 U2621 ( .A1(n4764), .A2(n556), .ZN(n555) );
  NAND2_X1 U2622 ( .A1(n4270), .A2(n19788), .ZN(n557) );
  XOR2_X1 U2623 ( .A(n7087), .B(n7316), .Z(n826) );
  NOR2_X1 U2625 ( .A1(n3247), .A2(n15306), .ZN(n15062) );
  NAND2_X1 U2626 ( .A1(n17882), .A2(n17881), .ZN(n558) );
  NAND2_X1 U2627 ( .A1(n17883), .A2(n222), .ZN(n559) );
  NAND3_X1 U2628 ( .A1(n593), .A2(n4437), .A3(n4438), .ZN(n1919) );
  NAND2_X1 U2629 ( .A1(n562), .A2(n560), .ZN(n17698) );
  NAND2_X1 U2630 ( .A1(n17694), .A2(n17819), .ZN(n560) );
  NAND2_X1 U2631 ( .A1(n17693), .A2(n935), .ZN(n562) );
  NAND3_X1 U2633 ( .A1(n564), .A2(n773), .A3(n3087), .ZN(n15059) );
  OAI211_X1 U2635 ( .C1(n15462), .C2(n1458), .A(n15351), .B(n15352), .ZN(n565)
         );
  OR2_X1 U2637 ( .A1(n2867), .A2(n2869), .ZN(n566) );
  NAND2_X1 U2638 ( .A1(n4707), .A2(n4706), .ZN(n567) );
  NAND2_X1 U2640 ( .A1(n1535), .A2(n619), .ZN(n1534) );
  NOR2_X1 U2641 ( .A1(n569), .A2(n568), .ZN(n5843) );
  NAND2_X1 U2642 ( .A1(n572), .A2(n570), .ZN(n12597) );
  NAND2_X1 U2643 ( .A1(n571), .A2(n12595), .ZN(n570) );
  NAND2_X1 U2644 ( .A1(n12593), .A2(n20430), .ZN(n571) );
  NAND2_X1 U2645 ( .A1(n12596), .A2(n11637), .ZN(n572) );
  NAND2_X1 U2646 ( .A1(n8851), .A2(n9038), .ZN(n1979) );
  OAI211_X1 U2648 ( .C1(n2600), .C2(n11977), .A(n574), .B(n250), .ZN(n11414)
         );
  NAND2_X1 U2649 ( .A1(n2600), .A2(n12545), .ZN(n574) );
  XNOR2_X1 U2650 ( .A(n638), .B(n6732), .ZN(n3484) );
  OR2_X1 U2651 ( .A1(n291), .A2(n5073), .ZN(n575) );
  NAND2_X1 U2653 ( .A1(n9098), .A2(n10646), .ZN(n576) );
  NAND2_X1 U2654 ( .A1(n1959), .A2(n20149), .ZN(n578) );
  XNOR2_X1 U2658 ( .A(n581), .B(n295), .ZN(Ciphertext[60]) );
  NAND3_X1 U2659 ( .A1(n582), .A2(n18641), .A3(n18640), .ZN(n581) );
  NAND2_X1 U2661 ( .A1(n19745), .A2(n583), .ZN(n18639) );
  NAND2_X1 U2663 ( .A1(n5760), .A2(n7421), .ZN(n586) );
  NAND2_X1 U2664 ( .A1(n18441), .A2(n18466), .ZN(n18446) );
  XNOR2_X2 U2665 ( .A(n587), .B(n13076), .ZN(n14514) );
  XNOR2_X1 U2666 ( .A(n2200), .B(n13077), .ZN(n587) );
  NAND3_X1 U2667 ( .A1(n243), .A2(n12537), .A3(n12534), .ZN(n2328) );
  NAND2_X1 U2669 ( .A1(n608), .A2(n20516), .ZN(n607) );
  NAND2_X1 U2670 ( .A1(n8852), .A2(n9038), .ZN(n589) );
  NAND2_X1 U2671 ( .A1(n8849), .A2(n591), .ZN(n590) );
  INV_X1 U2672 ( .A(n9038), .ZN(n591) );
  NAND2_X1 U2673 ( .A1(n592), .A2(n8492), .ZN(n7701) );
  NAND3_X1 U2675 ( .A1(n5429), .A2(n1776), .A3(n5790), .ZN(n2956) );
  NAND2_X1 U2676 ( .A1(n9009), .A2(n9007), .ZN(n1671) );
  OAI21_X1 U2677 ( .B1(n4807), .B2(n4802), .A(n4801), .ZN(n593) );
  XNOR2_X1 U2678 ( .A(n594), .B(n17365), .ZN(Ciphertext[8]) );
  NAND2_X1 U2680 ( .A1(n3455), .A2(n3456), .ZN(n596) );
  NAND2_X1 U2681 ( .A1(n1106), .A2(n3388), .ZN(n18394) );
  OAI21_X2 U2682 ( .B1(n11679), .B2(n12500), .A(n1149), .ZN(n12979) );
  AOI22_X1 U2683 ( .A1(n20111), .A2(n18384), .B1(n20611), .B2(n18376), .ZN(
        n18393) );
  NAND3_X1 U2684 ( .A1(n4609), .A2(n4613), .A3(n4177), .ZN(n3109) );
  NAND2_X1 U2685 ( .A1(n14005), .A2(n2304), .ZN(n14119) );
  AND2_X2 U2686 ( .A1(n751), .A2(n752), .ZN(n15696) );
  NAND2_X1 U2687 ( .A1(n5444), .A2(n5641), .ZN(n4179) );
  NAND3_X2 U2688 ( .A1(n3110), .A2(n3108), .A3(n4178), .ZN(n5444) );
  INV_X1 U2689 ( .A(n598), .ZN(n597) );
  NAND2_X1 U2691 ( .A1(n800), .A2(n9363), .ZN(n599) );
  NOR2_X1 U2692 ( .A1(n20005), .A2(n20133), .ZN(n750) );
  NAND2_X1 U2693 ( .A1(n17876), .A2(n16308), .ZN(n600) );
  OR2_X1 U2694 ( .A1(n10808), .A2(n10259), .ZN(n10809) );
  NAND2_X1 U2695 ( .A1(n4750), .A2(n4204), .ZN(n4558) );
  AOI22_X1 U2697 ( .A1(n11266), .A2(n11265), .B1(n11335), .B2(n11267), .ZN(
        n602) );
  OAI211_X2 U2698 ( .C1(n14521), .C2(n14520), .A(n15126), .B(n15125), .ZN(
        n15018) );
  NAND2_X1 U2699 ( .A1(n14518), .A2(n14519), .ZN(n15126) );
  NAND2_X1 U2701 ( .A1(n4366), .A2(n290), .ZN(n603) );
  NAND2_X1 U2702 ( .A1(n605), .A2(n4365), .ZN(n604) );
  NAND2_X1 U2703 ( .A1(n4011), .A2(n4614), .ZN(n605) );
  NAND2_X1 U2704 ( .A1(n11671), .A2(n11672), .ZN(n11676) );
  NAND2_X1 U2706 ( .A1(n8330), .A2(n8331), .ZN(n9861) );
  NAND2_X1 U2707 ( .A1(n2238), .A2(n7643), .ZN(n8603) );
  NOR2_X1 U2709 ( .A1(n15896), .A2(n15536), .ZN(n15539) );
  AOI22_X1 U2710 ( .A1(n11735), .A2(n242), .B1(n13149), .B2(n20153), .ZN(
        n11736) );
  NAND2_X1 U2711 ( .A1(n10803), .A2(n191), .ZN(n10804) );
  NAND2_X1 U2712 ( .A1(n18645), .A2(n18656), .ZN(n18282) );
  INV_X1 U2713 ( .A(n4615), .ZN(n748) );
  INV_X1 U2715 ( .A(n11159), .ZN(n608) );
  INV_X1 U2717 ( .A(n4931), .ZN(n4977) );
  OAI21_X1 U2718 ( .B1(n3877), .B2(n3876), .A(n4931), .ZN(n3878) );
  NAND2_X1 U2719 ( .A1(n4979), .A2(n4297), .ZN(n4931) );
  NAND2_X1 U2721 ( .A1(n17395), .A2(n18257), .ZN(n611) );
  OR2_X1 U2722 ( .A1(n18260), .A2(n18257), .ZN(n612) );
  NAND2_X1 U2725 ( .A1(n613), .A2(n4010), .ZN(n3955) );
  NAND2_X1 U2726 ( .A1(n4364), .A2(n4614), .ZN(n613) );
  NAND2_X1 U2728 ( .A1(n2682), .A2(n14599), .ZN(n3532) );
  INV_X1 U2729 ( .A(n9602), .ZN(n10289) );
  NAND2_X1 U2730 ( .A1(n7624), .A2(n7625), .ZN(n8741) );
  NAND4_X1 U2731 ( .A1(n4636), .A2(n4634), .A3(n4637), .A4(n4635), .ZN(n614)
         );
  NAND2_X1 U2732 ( .A1(n5319), .A2(n5406), .ZN(n615) );
  NAND2_X1 U2733 ( .A1(n13924), .A2(n3599), .ZN(n3254) );
  NAND2_X1 U2736 ( .A1(n6042), .A2(n1214), .ZN(n5308) );
  AND2_X2 U2737 ( .A1(n687), .A2(n688), .ZN(n15796) );
  NAND2_X1 U2738 ( .A1(n4616), .A2(n748), .ZN(n617) );
  NAND2_X1 U2739 ( .A1(n3715), .A2(n619), .ZN(n618) );
  INV_X1 U2740 ( .A(n3717), .ZN(n619) );
  MUX2_X1 U2742 ( .A(n4112), .B(n5711), .S(n5709), .Z(n622) );
  AOI21_X1 U2743 ( .B1(n1270), .B2(n3832), .A(n20105), .ZN(n623) );
  NAND2_X1 U2744 ( .A1(n624), .A2(n9346), .ZN(n2168) );
  NAND2_X1 U2745 ( .A1(n2170), .A2(n2169), .ZN(n624) );
  NAND2_X1 U2746 ( .A1(n4237), .A2(n4238), .ZN(n2215) );
  NAND2_X1 U2748 ( .A1(n15680), .A2(n15679), .ZN(n625) );
  NAND2_X1 U2749 ( .A1(n15681), .A2(n15682), .ZN(n626) );
  NOR2_X1 U2750 ( .A1(n152), .A2(n628), .ZN(n16460) );
  NAND2_X1 U2751 ( .A1(n630), .A2(n629), .ZN(n3681) );
  INV_X1 U2752 ( .A(n8017), .ZN(n630) );
  NAND2_X1 U2753 ( .A1(n631), .A2(n14800), .ZN(n14211) );
  XNOR2_X2 U2754 ( .A(n12249), .B(n12248), .ZN(n14800) );
  INV_X1 U2755 ( .A(n3440), .ZN(n631) );
  NAND3_X1 U2756 ( .A1(n252), .A2(n12179), .A3(n20427), .ZN(n1980) );
  XNOR2_X1 U2757 ( .A(n735), .B(n9478), .ZN(n9551) );
  NAND3_X1 U2758 ( .A1(n19742), .A2(n1089), .A3(n14501), .ZN(n13053) );
  NAND2_X1 U2759 ( .A1(n4807), .A2(n633), .ZN(n4699) );
  AND2_X1 U2760 ( .A1(n5087), .A2(n20202), .ZN(n633) );
  NAND2_X1 U2763 ( .A1(n16579), .A2(n635), .ZN(n634) );
  NAND2_X1 U2765 ( .A1(n1751), .A2(n9313), .ZN(n637) );
  XNOR2_X1 U2766 ( .A(n6731), .B(n6730), .ZN(n638) );
  NAND2_X1 U2767 ( .A1(n14731), .A2(n14729), .ZN(n14137) );
  NAND2_X1 U2768 ( .A1(n3086), .A2(n5602), .ZN(n5485) );
  AND2_X2 U2773 ( .A1(n5245), .A2(n5244), .ZN(n5249) );
  NAND2_X1 U2774 ( .A1(n7904), .A2(n7754), .ZN(n3272) );
  NAND2_X1 U2775 ( .A1(n7903), .A2(n20166), .ZN(n7904) );
  OAI211_X2 U2776 ( .C1(n7758), .C2(n7757), .A(n7756), .B(n644), .ZN(n8657) );
  NAND2_X1 U2780 ( .A1(n10069), .A2(n11548), .ZN(n646) );
  INV_X1 U2781 ( .A(n11548), .ZN(n647) );
  NAND2_X1 U2782 ( .A1(n11544), .A2(n10760), .ZN(n648) );
  AND2_X1 U2783 ( .A1(n205), .A2(n11133), .ZN(n10830) );
  NAND2_X1 U2784 ( .A1(n11052), .A2(n650), .ZN(n11053) );
  NAND2_X1 U2785 ( .A1(n11130), .A2(n650), .ZN(n2106) );
  NAND2_X1 U2788 ( .A1(n16685), .A2(n651), .ZN(n654) );
  AOI22_X2 U2792 ( .A1(n16686), .A2(n654), .B1(n19399), .B2(n16687), .ZN(
        n19463) );
  NAND2_X1 U2793 ( .A1(n654), .A2(n17654), .ZN(n17659) );
  OR2_X2 U2794 ( .A1(n5137), .A2(n5136), .ZN(n655) );
  NOR2_X1 U2795 ( .A1(n655), .A2(n9234), .ZN(n8633) );
  NAND2_X1 U2796 ( .A1(n19716), .A2(n655), .ZN(n9236) );
  NAND3_X1 U2797 ( .A1(n8411), .A2(n9234), .A3(n655), .ZN(n6214) );
  NAND2_X1 U2798 ( .A1(n8630), .A2(n655), .ZN(n8632) );
  NAND2_X1 U2800 ( .A1(n656), .A2(n912), .ZN(n2249) );
  MUX2_X1 U2801 ( .A(n14327), .B(n14352), .S(n14818), .Z(n656) );
  XNOR2_X1 U2802 ( .A(n20224), .B(n657), .ZN(n6554) );
  XNOR2_X1 U2803 ( .A(n657), .B(n18792), .ZN(n6848) );
  XNOR2_X1 U2804 ( .A(n7206), .B(n657), .ZN(n6962) );
  XNOR2_X1 U2805 ( .A(n6743), .B(n657), .ZN(n7303) );
  INV_X1 U2806 ( .A(n2816), .ZN(n660) );
  NOR2_X1 U2807 ( .A1(n2816), .A2(n215), .ZN(n658) );
  NAND3_X1 U2808 ( .A1(n19278), .A2(n19269), .A3(n660), .ZN(n19256) );
  MUX2_X1 U2809 ( .A(n19246), .B(n19269), .S(n2816), .Z(n17682) );
  NAND2_X1 U2810 ( .A1(n19274), .A2(n2816), .ZN(n659) );
  AOI21_X1 U2811 ( .B1(n19275), .B2(n660), .A(n20448), .ZN(n19277) );
  OR2_X1 U2812 ( .A1(n5021), .A2(n4277), .ZN(n662) );
  NAND2_X1 U2813 ( .A1(n4554), .A2(n663), .ZN(n661) );
  NAND2_X1 U2814 ( .A1(n5803), .A2(n5378), .ZN(n5733) );
  AND2_X1 U2815 ( .A1(n4734), .A2(n4555), .ZN(n663) );
  MUX2_X1 U2816 ( .A(n666), .B(n4568), .S(n1391), .Z(n664) );
  INV_X1 U2817 ( .A(n666), .ZN(n665) );
  NAND2_X1 U2818 ( .A1(n4563), .A2(n4754), .ZN(n666) );
  NAND2_X1 U2820 ( .A1(n7725), .A2(n7851), .ZN(n667) );
  NAND2_X1 U2822 ( .A1(n669), .A2(n8972), .ZN(n3354) );
  OAI21_X1 U2823 ( .B1(n8971), .B2(n9255), .A(n8976), .ZN(n669) );
  NAND2_X1 U2824 ( .A1(n671), .A2(n670), .ZN(n8976) );
  INV_X1 U2825 ( .A(n9250), .ZN(n671) );
  NAND2_X1 U2826 ( .A1(n4731), .A2(n672), .ZN(n4276) );
  NAND2_X1 U2827 ( .A1(n4110), .A2(n5012), .ZN(n5013) );
  NAND3_X1 U2828 ( .A1(n5016), .A2(n4110), .A3(n4734), .ZN(n4735) );
  NAND3_X1 U2829 ( .A1(n5020), .A2(n5019), .A3(n673), .ZN(n6027) );
  OR2_X1 U2830 ( .A1(n5021), .A2(n4110), .ZN(n673) );
  XNOR2_X1 U2831 ( .A(n674), .B(n18308), .ZN(Ciphertext[98]) );
  NAND2_X1 U2832 ( .A1(n677), .A2(n675), .ZN(n674) );
  NAND2_X1 U2833 ( .A1(n676), .A2(n19988), .ZN(n675) );
  MUX2_X1 U2834 ( .A(n20259), .B(n18857), .S(n20418), .Z(n676) );
  NAND2_X1 U2836 ( .A1(n678), .A2(n20535), .ZN(n677) );
  OAI21_X1 U2839 ( .B1(n5404), .B2(n5571), .A(n5408), .ZN(n5147) );
  NAND3_X1 U2840 ( .A1(n4607), .A2(n1908), .A3(n4312), .ZN(n680) );
  NAND2_X1 U2842 ( .A1(n14658), .A2(n19748), .ZN(n681) );
  XNOR2_X1 U2843 ( .A(n13185), .B(n13248), .ZN(n13186) );
  NAND2_X1 U2844 ( .A1(n11725), .A2(n685), .ZN(n683) );
  NAND2_X1 U2845 ( .A1(n686), .A2(n924), .ZN(n2143) );
  NAND2_X1 U2846 ( .A1(n12537), .A2(n686), .ZN(n11488) );
  INV_X1 U2847 ( .A(n12534), .ZN(n686) );
  INV_X1 U2849 ( .A(n17315), .ZN(n689) );
  NOR2_X1 U2850 ( .A1(n690), .A2(n15573), .ZN(n692) );
  INV_X1 U2851 ( .A(n15577), .ZN(n691) );
  NAND2_X1 U2852 ( .A1(n15791), .A2(n15796), .ZN(n693) );
  XNOR2_X1 U2854 ( .A(n694), .B(n17851), .ZN(n10418) );
  XNOR2_X1 U2855 ( .A(n694), .B(n9462), .ZN(n9656) );
  XNOR2_X1 U2856 ( .A(n9799), .B(n694), .ZN(n8427) );
  XNOR2_X1 U2857 ( .A(n694), .B(n9754), .ZN(n9465) );
  NAND2_X1 U2859 ( .A1(n699), .A2(n12126), .ZN(n12134) );
  NAND2_X1 U2860 ( .A1(n696), .A2(n699), .ZN(n695) );
  NAND2_X1 U2863 ( .A1(n2983), .A2(n238), .ZN(n3172) );
  NAND2_X1 U2864 ( .A1(n20262), .A2(n2983), .ZN(n700) );
  NAND3_X1 U2866 ( .A1(n9278), .A2(n9275), .A3(n8991), .ZN(n702) );
  INV_X1 U2867 ( .A(n11650), .ZN(n11674) );
  OAI21_X1 U2868 ( .B1(n3645), .B2(n8736), .A(n19518), .ZN(n708) );
  INV_X1 U2869 ( .A(n8921), .ZN(n705) );
  NAND2_X1 U2870 ( .A1(n8497), .A2(n707), .ZN(n706) );
  NOR2_X1 U2871 ( .A1(n19518), .A2(n8923), .ZN(n707) );
  NAND2_X1 U2872 ( .A1(n8324), .A2(n276), .ZN(n709) );
  NAND2_X1 U2873 ( .A1(n711), .A2(n710), .ZN(n9103) );
  NAND2_X1 U2874 ( .A1(n8323), .A2(n1425), .ZN(n710) );
  NAND2_X1 U2875 ( .A1(n3611), .A2(n19856), .ZN(n711) );
  NAND2_X1 U2876 ( .A1(n3161), .A2(n3160), .ZN(n712) );
  OAI22_X1 U2878 ( .A1(n12383), .A2(n12138), .B1(n11917), .B2(n712), .ZN(
        n11918) );
  NAND2_X1 U2881 ( .A1(n2146), .A2(n15266), .ZN(n716) );
  NAND3_X1 U2882 ( .A1(n717), .A2(n15636), .A3(n716), .ZN(n715) );
  NAND3_X1 U2883 ( .A1(n8214), .A2(n8213), .A3(n718), .ZN(n9113) );
  INV_X1 U2884 ( .A(n17886), .ZN(n719) );
  NAND2_X1 U2885 ( .A1(n719), .A2(n17887), .ZN(n3214) );
  NAND2_X1 U2886 ( .A1(n720), .A2(n12004), .ZN(n1861) );
  NAND2_X1 U2887 ( .A1(n12498), .A2(n12500), .ZN(n720) );
  NAND2_X1 U2890 ( .A1(n10007), .A2(n11575), .ZN(n722) );
  NAND2_X1 U2892 ( .A1(n10740), .A2(n11572), .ZN(n727) );
  NAND2_X1 U2894 ( .A1(n729), .A2(n3642), .ZN(n728) );
  NAND2_X1 U2895 ( .A1(n730), .A2(n14675), .ZN(n729) );
  NAND2_X1 U2896 ( .A1(n19530), .A2(n14542), .ZN(n730) );
  XNOR2_X2 U2897 ( .A(n8757), .B(n8756), .ZN(n11538) );
  NAND2_X1 U2898 ( .A1(n733), .A2(n5148), .ZN(n3960) );
  AOI21_X1 U2899 ( .B1(n5404), .B2(n733), .A(n5582), .ZN(n5409) );
  MUX2_X1 U2900 ( .A(n5404), .B(n733), .S(n5148), .Z(n3961) );
  XNOR2_X1 U2902 ( .A(n10494), .B(n9477), .ZN(n735) );
  XNOR2_X1 U2903 ( .A(n734), .B(n10126), .ZN(n10494) );
  INV_X1 U2904 ( .A(n9824), .ZN(n734) );
  MUX2_X1 U2906 ( .A(n9576), .B(n9291), .S(n9049), .Z(n736) );
  NAND2_X1 U2907 ( .A1(n1541), .A2(n1538), .ZN(n737) );
  NAND2_X1 U2910 ( .A1(n11730), .A2(n11683), .ZN(n740) );
  NAND2_X1 U2911 ( .A1(n742), .A2(n11926), .ZN(n741) );
  NAND2_X1 U2912 ( .A1(n11923), .A2(n11922), .ZN(n742) );
  OAI211_X1 U2913 ( .C1(n9576), .C2(n9287), .A(n743), .B(n9291), .ZN(n744) );
  NAND2_X1 U2914 ( .A1(n9576), .A2(n19715), .ZN(n743) );
  NAND2_X1 U2916 ( .A1(n9579), .A2(n746), .ZN(n745) );
  OR2_X1 U2917 ( .A1(n19519), .A2(n9576), .ZN(n746) );
  NAND2_X1 U2918 ( .A1(n747), .A2(n15607), .ZN(n14975) );
  MUX2_X1 U2919 ( .A(n15608), .B(n16126), .S(n16129), .Z(n14977) );
  NAND2_X1 U2920 ( .A1(n20007), .A2(n747), .ZN(n15737) );
  NAND2_X1 U2921 ( .A1(n15494), .A2(n747), .ZN(n3432) );
  NAND2_X1 U2922 ( .A1(n3415), .A2(n747), .ZN(n3414) );
  NAND2_X1 U2924 ( .A1(n749), .A2(n4610), .ZN(n4616) );
  NAND2_X1 U2925 ( .A1(n4365), .A2(n4013), .ZN(n4610) );
  NAND2_X1 U2926 ( .A1(n290), .A2(n4613), .ZN(n749) );
  NAND2_X1 U2927 ( .A1(n750), .A2(n20449), .ZN(n1998) );
  NAND2_X1 U2928 ( .A1(n14119), .A2(n19503), .ZN(n751) );
  NAND2_X1 U2929 ( .A1(n14006), .A2(n14232), .ZN(n752) );
  NAND2_X1 U2930 ( .A1(n754), .A2(n753), .ZN(n11809) );
  NAND2_X1 U2931 ( .A1(n1282), .A2(n9832), .ZN(n754) );
  NAND2_X1 U2933 ( .A1(n758), .A2(n757), .ZN(n16441) );
  NAND2_X1 U2934 ( .A1(n16434), .A2(n160), .ZN(n757) );
  NAND2_X1 U2935 ( .A1(n759), .A2(n226), .ZN(n758) );
  NAND2_X1 U2936 ( .A1(n4649), .A2(n4648), .ZN(n760) );
  MUX2_X1 U2937 ( .A(n4644), .B(n4643), .S(n4642), .Z(n761) );
  NAND2_X1 U2938 ( .A1(n12107), .A2(n764), .ZN(n974) );
  INV_X1 U2939 ( .A(n1840), .ZN(n767) );
  INV_X1 U2940 ( .A(n2317), .ZN(n768) );
  NAND2_X1 U2942 ( .A1(n18953), .A2(n17831), .ZN(n17830) );
  OR2_X1 U2943 ( .A1(n7560), .A2(n8249), .ZN(n769) );
  NAND2_X1 U2944 ( .A1(n3540), .A2(n3541), .ZN(n8435) );
  AND3_X2 U2945 ( .A1(n3540), .A2(n3541), .A3(n770), .ZN(n9780) );
  NAND2_X1 U2946 ( .A1(n3542), .A2(n9780), .ZN(n772) );
  NAND2_X1 U2947 ( .A1(n2983), .A2(n2773), .ZN(n773) );
  NAND2_X1 U2948 ( .A1(n15059), .A2(n15309), .ZN(n15060) );
  NOR2_X1 U2950 ( .A1(n14431), .A2(n14481), .ZN(n774) );
  AOI21_X1 U2951 ( .B1(n3900), .B2(n3899), .A(n19822), .ZN(n775) );
  MUX2_X1 U2952 ( .A(n5791), .B(n5300), .S(n5428), .Z(n5158) );
  NAND2_X1 U2953 ( .A1(n776), .A2(n7922), .ZN(n7923) );
  AOI21_X1 U2956 ( .B1(n8705), .B2(n9168), .A(n9167), .ZN(n778) );
  NAND2_X1 U2957 ( .A1(n237), .A2(n779), .ZN(n3244) );
  NAND2_X1 U2958 ( .A1(n18332), .A2(n213), .ZN(n18334) );
  INV_X1 U2959 ( .A(n781), .ZN(n784) );
  AOI21_X1 U2960 ( .B1(n13182), .B2(n13181), .A(n2023), .ZN(n781) );
  NAND2_X1 U2962 ( .A1(n784), .A2(n782), .ZN(n13183) );
  NAND2_X1 U2963 ( .A1(n13182), .A2(n783), .ZN(n782) );
  XNOR2_X1 U2964 ( .A(n785), .B(n18587), .ZN(n16573) );
  XNOR2_X1 U2965 ( .A(n785), .B(n2376), .ZN(n16046) );
  XNOR2_X1 U2966 ( .A(n785), .B(n3162), .ZN(n16386) );
  XNOR2_X1 U2967 ( .A(n16095), .B(n785), .ZN(n16828) );
  OR2_X1 U2968 ( .A1(n7855), .A2(n282), .ZN(n8259) );
  NAND2_X1 U2969 ( .A1(n786), .A2(n8157), .ZN(n7725) );
  NAND2_X1 U2970 ( .A1(n7855), .A2(n282), .ZN(n786) );
  NAND3_X1 U2971 ( .A1(n279), .A2(n7724), .A3(n8157), .ZN(n7554) );
  NAND2_X1 U2975 ( .A1(n15535), .A2(n15898), .ZN(n789) );
  NAND2_X1 U2976 ( .A1(n19838), .A2(n15401), .ZN(n15535) );
  XNOR2_X1 U2977 ( .A(n10030), .B(n791), .ZN(n10383) );
  INV_X1 U2978 ( .A(Key[63]), .ZN(n791) );
  NAND3_X1 U2979 ( .A1(n14023), .A2(n20266), .A3(n19748), .ZN(n1977) );
  NAND2_X1 U2982 ( .A1(n792), .A2(n20405), .ZN(n2796) );
  XNOR2_X1 U2983 ( .A(n794), .B(n793), .ZN(Ciphertext[124]) );
  INV_X1 U2984 ( .A(n1386), .ZN(n793) );
  NAND2_X1 U2985 ( .A1(n797), .A2(n795), .ZN(n794) );
  AOI22_X1 U2986 ( .A1(n796), .A2(n19069), .B1(n19653), .B2(n19070), .ZN(n795)
         );
  INV_X1 U2987 ( .A(n19071), .ZN(n796) );
  NAND2_X1 U2988 ( .A1(n19072), .A2(n19071), .ZN(n797) );
  NAND2_X1 U2989 ( .A1(n19074), .A2(n19059), .ZN(n19071) );
  NAND3_X2 U2990 ( .A1(n11199), .A2(n799), .A3(n798), .ZN(n12478) );
  NAND3_X1 U2991 ( .A1(n19913), .A2(n19719), .A3(n11198), .ZN(n799) );
  XNOR2_X2 U2992 ( .A(n10622), .B(n3049), .ZN(n11493) );
  INV_X1 U2993 ( .A(n7559), .ZN(n800) );
  XNOR2_X1 U2994 ( .A(n5249), .B(n302), .ZN(n7027) );
  NAND2_X1 U2996 ( .A1(n803), .A2(n9135), .ZN(n2726) );
  NAND2_X1 U2997 ( .A1(n9137), .A2(n803), .ZN(n9215) );
  AOI22_X1 U2998 ( .A1(n9135), .A2(n8446), .B1(n9134), .B2(n803), .ZN(n8447)
         );
  NOR2_X1 U2999 ( .A1(n953), .A2(n12488), .ZN(n11910) );
  NAND2_X1 U3000 ( .A1(n5908), .A2(n890), .ZN(n5495) );
  NAND2_X1 U3001 ( .A1(n805), .A2(n5494), .ZN(n804) );
  NAND2_X1 U3003 ( .A1(n19462), .A2(n19463), .ZN(n809) );
  XNOR2_X1 U3004 ( .A(n807), .B(n16688), .ZN(Ciphertext[189]) );
  NAND3_X1 U3005 ( .A1(n810), .A2(n808), .A3(n16682), .ZN(n807) );
  OAI211_X1 U3006 ( .C1(n19463), .C2(n17091), .A(n809), .B(n20140), .ZN(n808)
         );
  NAND2_X1 U3007 ( .A1(n301), .A2(n4539), .ZN(n4544) );
  NAND2_X1 U3008 ( .A1(n4349), .A2(n301), .ZN(n3760) );
  MUX2_X1 U3009 ( .A(n4347), .B(n4348), .S(n4541), .Z(n4352) );
  NAND3_X1 U3013 ( .A1(n17483), .A2(n17243), .A3(n812), .ZN(n811) );
  NAND3_X1 U3014 ( .A1(n815), .A2(n17479), .A3(n17480), .ZN(n814) );
  NAND2_X1 U3015 ( .A1(n817), .A2(n1718), .ZN(n816) );
  OAI21_X1 U3016 ( .B1(n17243), .B2(n17479), .A(n818), .ZN(n817) );
  NAND2_X1 U3017 ( .A1(n17479), .A2(n20353), .ZN(n818) );
  NAND2_X1 U3019 ( .A1(n2470), .A2(n10756), .ZN(n11531) );
  NAND2_X1 U3020 ( .A1(n819), .A2(n8200), .ZN(n820) );
  INV_X1 U3021 ( .A(n8070), .ZN(n819) );
  XNOR2_X2 U3022 ( .A(n5639), .B(n5638), .ZN(n8070) );
  NAND2_X1 U3023 ( .A1(n289), .A2(n20459), .ZN(n821) );
  NAND2_X1 U3024 ( .A1(n1312), .A2(n1311), .ZN(n822) );
  MUX2_X1 U3025 ( .A(n263), .B(n9135), .S(n9209), .Z(n1334) );
  NAND2_X1 U3026 ( .A1(n8351), .A2(n8350), .ZN(n824) );
  XNOR2_X1 U3027 ( .A(n825), .B(n6593), .ZN(n5854) );
  INV_X1 U3028 ( .A(n3590), .ZN(n825) );
  XNOR2_X1 U3029 ( .A(n3590), .B(n826), .ZN(n6638) );
  NAND2_X1 U3030 ( .A1(n5073), .A2(n4664), .ZN(n829) );
  NAND3_X1 U3031 ( .A1(n4814), .A2(n5072), .A3(n4409), .ZN(n830) );
  NAND2_X1 U3032 ( .A1(n4410), .A2(n5073), .ZN(n4409) );
  XNOR2_X1 U3033 ( .A(n831), .B(n18339), .ZN(Ciphertext[133]) );
  NAND2_X1 U3034 ( .A1(n834), .A2(n832), .ZN(n831) );
  NAND2_X1 U3035 ( .A1(n835), .A2(n833), .ZN(n832) );
  OAI22_X1 U3036 ( .A1(n835), .A2(n19130), .B1(n20508), .B2(n19148), .ZN(n834)
         );
  NAND2_X1 U3037 ( .A1(n20508), .A2(n19135), .ZN(n19130) );
  AND2_X1 U3038 ( .A1(n18337), .A2(n19134), .ZN(n835) );
  NAND2_X1 U3039 ( .A1(n8322), .A2(n2548), .ZN(n836) );
  AOI21_X1 U3040 ( .B1(n7585), .B2(n8325), .A(n8001), .ZN(n837) );
  NAND2_X1 U3041 ( .A1(n8532), .A2(n8577), .ZN(n839) );
  NAND3_X1 U3042 ( .A1(n846), .A2(n843), .A3(n841), .ZN(Ciphertext[61]) );
  NAND2_X1 U3043 ( .A1(n18647), .A2(n842), .ZN(n841) );
  NAND2_X1 U3044 ( .A1(n845), .A2(n844), .ZN(n843) );
  AOI21_X1 U3045 ( .B1(n18647), .B2(n18646), .A(n299), .ZN(n844) );
  NAND2_X1 U3046 ( .A1(n848), .A2(n18659), .ZN(n845) );
  NAND2_X1 U3047 ( .A1(n848), .A2(n847), .ZN(n846) );
  AND2_X1 U3048 ( .A1(n18659), .A2(n299), .ZN(n847) );
  INV_X1 U3049 ( .A(n18645), .ZN(n848) );
  OAI21_X1 U3050 ( .B1(n850), .B2(n11794), .A(n11792), .ZN(n852) );
  NAND3_X1 U3053 ( .A1(n1511), .A2(n907), .A3(n12523), .ZN(n851) );
  INV_X1 U3054 ( .A(n12165), .ZN(n1511) );
  INV_X1 U3055 ( .A(n16025), .ZN(n854) );
  NAND2_X1 U3056 ( .A1(n2732), .A2(n1339), .ZN(n855) );
  OAI211_X1 U3057 ( .C1(n8984), .C2(n8983), .A(n8982), .B(n3797), .ZN(n856) );
  OR2_X1 U3058 ( .A1(n11128), .A2(n2029), .ZN(n857) );
  OAI211_X1 U3059 ( .C1(n1597), .C2(n2462), .A(n1595), .B(n1594), .ZN(n861) );
  OAI211_X1 U3060 ( .C1(n1597), .C2(n2462), .A(n1595), .B(n1594), .ZN(n862) );
  OAI211_X1 U3062 ( .C1(n1597), .C2(n2462), .A(n1595), .B(n1594), .ZN(n5920)
         );
  NAND2_X1 U3065 ( .A1(n2300), .A2(n2299), .ZN(n865) );
  OAI21_X1 U3068 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(n15843) );
  XNOR2_X1 U3069 ( .A(n5690), .B(n6534), .ZN(n5727) );
  AOI21_X1 U3070 ( .B1(n16726), .B2(n20127), .A(n16725), .ZN(n19143) );
  XNOR2_X1 U3072 ( .A(Key[126]), .B(Plaintext[126]), .ZN(n873) );
  INV_X1 U3073 ( .A(n12041), .ZN(n876) );
  OAI211_X1 U3074 ( .C1(n9260), .C2(n19516), .A(n9258), .B(n9257), .ZN(n878)
         );
  OAI211_X1 U3075 ( .C1(n15850), .C2(n15851), .A(n15849), .B(n15848), .ZN(n879) );
  OAI211_X1 U3076 ( .C1(n15850), .C2(n15851), .A(n15849), .B(n15848), .ZN(n880) );
  XNOR2_X1 U3077 ( .A(n11593), .B(n11592), .ZN(n14779) );
  OAI211_X1 U3078 ( .C1(n9260), .C2(n19516), .A(n9258), .B(n9257), .ZN(n9878)
         );
  OR2_X1 U3080 ( .A1(n18382), .A2(n18384), .ZN(n881) );
  NAND2_X1 U3081 ( .A1(n881), .A2(n18394), .ZN(n2274) );
  OAI21_X1 U3082 ( .B1(n11016), .B2(n1579), .A(n10956), .ZN(n882) );
  OAI211_X1 U3083 ( .C1(n5242), .C2(n5714), .A(n4376), .B(n2207), .ZN(n883) );
  OAI21_X1 U3084 ( .B1(n11016), .B2(n1579), .A(n10956), .ZN(n12127) );
  OAI211_X1 U3085 ( .C1(n5242), .C2(n5714), .A(n4376), .B(n2207), .ZN(n7325)
         );
  OAI211_X2 U3086 ( .C1(n14576), .C2(n14570), .A(n14272), .B(n14271), .ZN(
        n15400) );
  INV_X1 U3087 ( .A(n7457), .ZN(n8053) );
  OR2_X1 U3088 ( .A1(n8361), .A2(n7709), .ZN(n884) );
  NAND2_X1 U3089 ( .A1(n884), .A2(n1994), .ZN(n7512) );
  NAND2_X1 U3090 ( .A1(n7875), .A2(n7874), .ZN(n885) );
  XNOR2_X1 U3092 ( .A(n10609), .B(n10610), .ZN(n888) );
  XOR2_X1 U3093 ( .A(n17031), .B(n17030), .Z(n889) );
  XOR2_X1 U3095 ( .A(n6856), .B(n6857), .Z(n6862) );
  NAND2_X1 U3096 ( .A1(n4838), .A2(n4837), .ZN(n890) );
  INV_X1 U3097 ( .A(n9018), .ZN(n891) );
  INV_X1 U3098 ( .A(n17729), .ZN(n893) );
  AND2_X1 U3099 ( .A1(n19755), .A2(n10873), .ZN(n894) );
  XNOR2_X1 U3100 ( .A(Key[63]), .B(Plaintext[63]), .ZN(n896) );
  XNOR2_X1 U3103 ( .A(Key[63]), .B(Plaintext[63]), .ZN(n4866) );
  NAND2_X1 U3105 ( .A1(n14877), .A2(n14878), .ZN(n897) );
  XNOR2_X1 U3106 ( .A(n9964), .B(n9963), .ZN(n898) );
  NAND2_X1 U3107 ( .A1(n14877), .A2(n14878), .ZN(n16336) );
  XNOR2_X1 U3108 ( .A(n9964), .B(n9963), .ZN(n11182) );
  BUF_X1 U3110 ( .A(n15957), .Z(n902) );
  OAI22_X1 U3111 ( .A1(n15707), .A2(n15706), .B1(n2625), .B2(n16009), .ZN(
        n15957) );
  NAND2_X1 U3112 ( .A1(n5976), .A2(n5977), .ZN(n903) );
  INV_X1 U3113 ( .A(n905), .ZN(n904) );
  NAND2_X1 U3114 ( .A1(n5976), .A2(n5977), .ZN(n7372) );
  NAND2_X1 U3115 ( .A1(n3850), .A2(n3849), .ZN(n906) );
  INV_X1 U3116 ( .A(n11493), .ZN(n3521) );
  OAI21_X1 U3118 ( .B1(n11463), .B2(n11886), .A(n11462), .ZN(n907) );
  INV_X1 U3119 ( .A(n8795), .ZN(n908) );
  XNOR2_X1 U3120 ( .A(n16347), .B(n17411), .ZN(n16921) );
  INV_X1 U3121 ( .A(n9748), .ZN(n9977) );
  NOR2_X1 U3123 ( .A1(n15819), .A2(n2114), .ZN(n911) );
  XNOR2_X1 U3124 ( .A(n10602), .B(n10601), .ZN(n913) );
  XNOR2_X1 U3126 ( .A(n12830), .B(n12829), .ZN(n14820) );
  XNOR2_X1 U3129 ( .A(n12071), .B(n12070), .ZN(n13206) );
  XNOR2_X1 U3130 ( .A(n13720), .B(n13719), .ZN(n14228) );
  AND2_X1 U3131 ( .A1(n20263), .A2(n14482), .ZN(n914) );
  OR2_X1 U3132 ( .A1(n12359), .A2(n12509), .ZN(n916) );
  NOR2_X1 U3133 ( .A1(n12366), .A2(n12365), .ZN(n13781) );
  NAND3_X1 U3134 ( .A1(n8170), .A2(n8169), .A3(n8168), .ZN(n917) );
  NAND3_X1 U3135 ( .A1(n8170), .A2(n8169), .A3(n8168), .ZN(n918) );
  XOR2_X1 U3136 ( .A(n13286), .B(n13285), .Z(n919) );
  INV_X1 U3138 ( .A(n14159), .ZN(n921) );
  XNOR2_X1 U3139 ( .A(n6638), .B(n6637), .ZN(n923) );
  XNOR2_X1 U3140 ( .A(n6638), .B(n6637), .ZN(n8066) );
  OR2_X1 U3141 ( .A1(n17937), .A2(n18349), .ZN(n925) );
  NAND2_X1 U3142 ( .A1(n925), .A2(n17908), .ZN(n17910) );
  XNOR2_X1 U3143 ( .A(n9440), .B(n9439), .ZN(n926) );
  XNOR2_X1 U3144 ( .A(n9956), .B(n926), .ZN(n927) );
  OAI211_X1 U3145 ( .C1(n9142), .C2(n9213), .A(n9141), .B(n9140), .ZN(n928) );
  XNOR2_X1 U3147 ( .A(n9956), .B(n926), .ZN(n11566) );
  OAI211_X1 U3148 ( .C1(n9142), .C2(n9213), .A(n9141), .B(n9140), .ZN(n10358)
         );
  AOI21_X1 U3149 ( .B1(n19387), .B2(n15731), .A(n15730), .ZN(n18412) );
  XNOR2_X1 U3150 ( .A(n10621), .B(n10321), .ZN(n9951) );
  XNOR2_X2 U3151 ( .A(n6807), .B(n6806), .ZN(n7855) );
  XNOR2_X1 U3152 ( .A(n10247), .B(n10008), .ZN(n929) );
  NAND2_X1 U3153 ( .A1(n17863), .A2(n16681), .ZN(n930) );
  NAND2_X1 U3154 ( .A1(n16680), .A2(n16679), .ZN(n931) );
  XNOR2_X1 U3155 ( .A(n13453), .B(n13369), .ZN(n933) );
  XNOR2_X1 U3156 ( .A(n7378), .B(n7379), .ZN(n934) );
  INV_X1 U3158 ( .A(n17729), .ZN(n18485) );
  OAI211_X2 U3159 ( .C1(n2781), .C2(n8614), .A(n8613), .B(n8612), .ZN(n9879)
         );
  XNOR2_X1 U3160 ( .A(n16700), .B(n16699), .ZN(n935) );
  XNOR2_X1 U3161 ( .A(n16084), .B(n16335), .ZN(n936) );
  OR2_X1 U3162 ( .A1(n17698), .A2(n17697), .ZN(n938) );
  OR2_X1 U3163 ( .A1(n14818), .A2(n14091), .ZN(n939) );
  OAI21_X1 U3165 ( .B1(n11618), .B2(n11897), .A(n11896), .ZN(n940) );
  OAI211_X1 U3167 ( .C1(n5874), .C2(n5873), .A(n5872), .B(n5871), .ZN(n943) );
  OAI211_X1 U3171 ( .C1(n5874), .C2(n5873), .A(n5872), .B(n5871), .ZN(n6249)
         );
  OAI21_X2 U3172 ( .B1(n4416), .B2(n4415), .A(n4414), .ZN(n6123) );
  AND2_X1 U3174 ( .A1(n5573), .A2(n5574), .ZN(n946) );
  OAI211_X2 U3176 ( .C1(n14137), .C2(n14408), .A(n14136), .B(n14135), .ZN(
        n16129) );
  INV_X1 U3179 ( .A(Plaintext[142]), .ZN(n2990) );
  XNOR2_X1 U3181 ( .A(n5727), .B(n5726), .ZN(n8200) );
  XNOR2_X1 U3182 ( .A(n6512), .B(n6811), .ZN(n7334) );
  XNOR2_X1 U3183 ( .A(n5759), .B(n1863), .ZN(n2886) );
  XNOR2_X1 U3184 ( .A(n6509), .B(n3321), .ZN(n8247) );
  OR2_X1 U3185 ( .A1(n6904), .A2(n7753), .ZN(n3271) );
  INV_X1 U3187 ( .A(n2886), .ZN(n7421) );
  AND2_X1 U3188 ( .A1(n8178), .A2(n8179), .ZN(n7416) );
  INV_X1 U3189 ( .A(n8247), .ZN(n8245) );
  INV_X1 U3190 ( .A(n8113), .ZN(n7844) );
  OR2_X1 U3191 ( .A1(n7722), .A2(n8352), .ZN(n2155) );
  AND2_X1 U3192 ( .A1(n7833), .A2(n8910), .ZN(n7918) );
  OR2_X1 U3193 ( .A1(n7507), .A2(n7748), .ZN(n1548) );
  XNOR2_X1 U3195 ( .A(n10461), .B(n10061), .ZN(n10356) );
  XNOR2_X1 U3196 ( .A(n1031), .B(n1029), .ZN(n9432) );
  XNOR2_X1 U3197 ( .A(n10621), .B(n3050), .ZN(n3049) );
  XNOR2_X1 U3198 ( .A(n10620), .B(n1605), .ZN(n3050) );
  INV_X1 U3199 ( .A(n10960), .ZN(n11143) );
  OR2_X1 U3200 ( .A1(n11124), .A2(n85), .ZN(n2033) );
  OR2_X1 U3201 ( .A1(n11540), .A2(n11168), .ZN(n3279) );
  AND2_X1 U3202 ( .A1(n12289), .A2(n12288), .ZN(n1440) );
  INV_X1 U3203 ( .A(n13697), .ZN(n12769) );
  INV_X1 U3204 ( .A(n11640), .ZN(n13792) );
  OAI211_X1 U3205 ( .C1(n11647), .C2(n11646), .A(n12227), .B(n11692), .ZN(
        n11648) );
  XNOR2_X1 U3206 ( .A(n13503), .B(n13502), .ZN(n14490) );
  XNOR2_X1 U3207 ( .A(n13139), .B(n3498), .ZN(n13471) );
  XNOR2_X1 U3208 ( .A(n12872), .B(n12871), .ZN(n13927) );
  AND2_X1 U3209 ( .A1(n13927), .A2(n14451), .ZN(n13559) );
  INV_X1 U3210 ( .A(n14493), .ZN(n1936) );
  NOR2_X1 U3211 ( .A1(n15424), .A2(n14238), .ZN(n14243) );
  XNOR2_X1 U3212 ( .A(n3543), .B(Key[53]), .ZN(n4233) );
  INV_X1 U3213 ( .A(n4950), .ZN(n3265) );
  XNOR2_X1 U3214 ( .A(Plaintext[45]), .B(Key[45]), .ZN(n4969) );
  AND2_X1 U3215 ( .A1(n5055), .A2(n4100), .ZN(n5053) );
  INV_X1 U3216 ( .A(n4887), .ZN(n4947) );
  INV_X1 U3217 ( .A(Plaintext[64]), .ZN(n1088) );
  INV_X1 U3218 ( .A(n6410), .ZN(n7025) );
  OR2_X1 U3219 ( .A1(n5763), .A2(n5736), .ZN(n2239) );
  OR2_X1 U3220 ( .A1(n5805), .A2(n6192), .ZN(n4593) );
  XNOR2_X1 U3221 ( .A(n7054), .B(n7053), .ZN(n2977) );
  NOR2_X1 U3222 ( .A1(n4062), .A2(n956), .ZN(n1131) );
  INV_X1 U3223 ( .A(n6510), .ZN(n8248) );
  OR2_X1 U3224 ( .A1(n7982), .A2(n7981), .ZN(n7767) );
  INV_X1 U3225 ( .A(n1507), .ZN(n1574) );
  AND2_X1 U3226 ( .A1(n7312), .A2(n7311), .ZN(n8323) );
  AND2_X1 U3227 ( .A1(n3395), .A2(n3394), .ZN(n1841) );
  INV_X1 U3228 ( .A(n7311), .ZN(n7590) );
  AND2_X1 U3229 ( .A1(n7958), .A2(n2977), .ZN(n2976) );
  AOI21_X1 U3230 ( .B1(n8013), .B2(n8012), .A(n7826), .ZN(n3625) );
  OR2_X1 U3231 ( .A1(n8035), .A2(n8286), .ZN(n2165) );
  NOR2_X1 U3233 ( .A1(n7909), .A2(n274), .ZN(n1785) );
  XNOR2_X1 U3234 ( .A(n6717), .B(n6720), .ZN(n2824) );
  INV_X1 U3235 ( .A(n7675), .ZN(n1994) );
  OR2_X1 U3236 ( .A1(n7622), .A2(n8177), .ZN(n3523) );
  OR2_X1 U3237 ( .A1(n7003), .A2(n7755), .ZN(n7004) );
  NOR2_X1 U3238 ( .A1(n8002), .A2(n3076), .ZN(n3075) );
  XNOR2_X1 U3242 ( .A(n10151), .B(n10491), .ZN(n10549) );
  INV_X1 U3243 ( .A(n10980), .ZN(n11291) );
  AND2_X1 U3244 ( .A1(n10980), .A2(n11294), .ZN(n11406) );
  XNOR2_X1 U3245 ( .A(n1284), .B(n1283), .ZN(n1285) );
  INV_X1 U3246 ( .A(n10808), .ZN(n11883) );
  INV_X1 U3247 ( .A(n1040), .ZN(n1317) );
  OR2_X1 U3248 ( .A1(n3789), .A2(n11177), .ZN(n10966) );
  XNOR2_X1 U3249 ( .A(n2202), .B(n7664), .ZN(n10945) );
  XNOR2_X1 U3250 ( .A(n10510), .B(n1479), .ZN(n11302) );
  XNOR2_X1 U3251 ( .A(n9771), .B(n18379), .ZN(n9772) );
  INV_X1 U3252 ( .A(n12463), .ZN(n11915) );
  OR2_X1 U3254 ( .A1(n11217), .A2(n11475), .ZN(n3768) );
  OR2_X1 U3255 ( .A1(n11289), .A2(n10950), .ZN(n3023) );
  INV_X1 U3257 ( .A(n12252), .ZN(n3637) );
  OR2_X1 U3258 ( .A1(n11078), .A2(n11474), .ZN(n2464) );
  OR2_X1 U3260 ( .A1(n11006), .A2(n19851), .ZN(n3175) );
  NAND2_X1 U3261 ( .A1(n1663), .A2(n1664), .ZN(n12255) );
  INV_X1 U3262 ( .A(n11243), .ZN(n1599) );
  OAI21_X1 U3263 ( .B1(n1748), .B2(n11140), .A(n1747), .ZN(n11146) );
  INV_X1 U3264 ( .A(n12600), .ZN(n12072) );
  INV_X1 U3265 ( .A(n14623), .ZN(n14001) );
  XNOR2_X1 U3266 ( .A(n13204), .B(n977), .ZN(n12654) );
  XNOR2_X1 U3268 ( .A(n13481), .B(n13081), .ZN(n13199) );
  INV_X1 U3269 ( .A(n12479), .ZN(n2553) );
  XNOR2_X1 U3270 ( .A(n13204), .B(n13205), .ZN(n13209) );
  OR2_X1 U3271 ( .A1(n1208), .A2(n14020), .ZN(n1207) );
  XNOR2_X1 U3272 ( .A(n13807), .B(n13251), .ZN(n2832) );
  XNOR2_X1 U3273 ( .A(n3742), .B(n3743), .ZN(n14120) );
  XNOR2_X1 U3274 ( .A(n13773), .B(n13770), .ZN(n2623) );
  INV_X1 U3275 ( .A(n15313), .ZN(n14146) );
  BUF_X1 U3276 ( .A(n14103), .Z(n14788) );
  OR2_X1 U3278 ( .A1(n14127), .A2(n19921), .ZN(n13950) );
  INV_X1 U3279 ( .A(n14599), .ZN(n1264) );
  XNOR2_X1 U3280 ( .A(n12972), .B(n12971), .ZN(n14032) );
  OR2_X1 U3281 ( .A1(n14442), .A2(n14168), .ZN(n2773) );
  NAND2_X1 U3284 ( .A1(n15488), .A2(n15487), .ZN(n15758) );
  OR2_X1 U3285 ( .A1(n2808), .A2(n14196), .ZN(n3006) );
  INV_X1 U3286 ( .A(n15421), .ZN(n2974) );
  AND2_X1 U3287 ( .A1(n19752), .A2(n15921), .ZN(n1119) );
  OR2_X1 U3288 ( .A1(n3174), .A2(n12919), .ZN(n2088) );
  OR2_X1 U3289 ( .A1(n13866), .A2(n15121), .ZN(n1789) );
  OR2_X1 U3290 ( .A1(n1795), .A2(n13559), .ZN(n1794) );
  AND2_X1 U3291 ( .A1(n14172), .A2(n14171), .ZN(n13883) );
  OR2_X1 U3292 ( .A1(n14750), .A2(n14747), .ZN(n3267) );
  OR2_X1 U3293 ( .A1(n14981), .A2(n15553), .ZN(n3042) );
  OR2_X1 U3294 ( .A1(n4824), .A2(n5258), .ZN(n4825) );
  XNOR2_X1 U3295 ( .A(n3874), .B(Key[23]), .ZN(n4021) );
  OR2_X1 U3297 ( .A1(n177), .A2(n3995), .ZN(n4682) );
  OR2_X1 U3298 ( .A1(n4391), .A2(n4685), .ZN(n4854) );
  OR2_X1 U3299 ( .A1(n5079), .A2(n4719), .ZN(n1163) );
  OR2_X1 U3300 ( .A1(n5080), .A2(n5075), .ZN(n5078) );
  INV_X1 U3302 ( .A(n4532), .ZN(n3551) );
  INV_X1 U3303 ( .A(n5226), .ZN(n6202) );
  INV_X1 U3304 ( .A(n4793), .ZN(n3167) );
  OR2_X1 U3305 ( .A1(n4056), .A2(n4060), .ZN(n4741) );
  INV_X1 U3306 ( .A(n4796), .ZN(n2670) );
  OR2_X1 U3307 ( .A1(n4088), .A2(n5046), .ZN(n5044) );
  INV_X1 U3308 ( .A(n4198), .ZN(n1391) );
  OR2_X1 U3309 ( .A1(n4504), .A2(n4565), .ZN(n4753) );
  XNOR2_X1 U3310 ( .A(n3204), .B(Key[124]), .ZN(n4706) );
  OR2_X1 U3311 ( .A1(n4618), .A2(n4982), .ZN(n1803) );
  OR2_X1 U3312 ( .A1(n4114), .A2(n4940), .ZN(n2389) );
  INV_X1 U3313 ( .A(n4271), .ZN(n5025) );
  INV_X1 U3314 ( .A(n4440), .ZN(n5040) );
  INV_X1 U3316 ( .A(n6168), .ZN(n1867) );
  INV_X1 U3317 ( .A(n292), .ZN(n3231) );
  OR2_X1 U3318 ( .A1(n4613), .A2(n4614), .ZN(n3716) );
  OR2_X1 U3319 ( .A1(n4674), .A2(n4673), .ZN(n3191) );
  OR2_X1 U3320 ( .A1(n4969), .A2(n4968), .ZN(n4971) );
  OR2_X1 U3321 ( .A1(n5054), .A2(n5055), .ZN(n2266) );
  OR2_X1 U3322 ( .A1(n6003), .A2(n6002), .ZN(n1454) );
  OR2_X1 U3323 ( .A1(n6138), .A2(n3188), .ZN(n4461) );
  AND2_X1 U3324 ( .A1(n5996), .A2(n5998), .ZN(n3604) );
  OR2_X1 U3325 ( .A1(n4114), .A2(n4118), .ZN(n3896) );
  MUX2_X1 U3326 ( .A(n4481), .B(n4480), .S(n4479), .Z(n3043) );
  OR2_X2 U3327 ( .A1(n4666), .A2(n4665), .ZN(n6172) );
  OR2_X1 U3329 ( .A1(n7445), .A2(n19686), .ZN(n3662) );
  OR2_X1 U3331 ( .A1(n5733), .A2(n6194), .ZN(n2866) );
  INV_X1 U3332 ( .A(n7500), .ZN(n8358) );
  INV_X1 U3333 ( .A(n7739), .ZN(n8357) );
  AND2_X1 U3335 ( .A1(n8112), .A2(n8241), .ZN(n1271) );
  OR2_X1 U3336 ( .A1(n9021), .A2(n8672), .ZN(n8838) );
  OR2_X1 U3337 ( .A1(n9023), .A2(n8510), .ZN(n1631) );
  INV_X1 U3338 ( .A(n2499), .ZN(n2501) );
  AND2_X1 U3339 ( .A1(n8947), .A2(n8945), .ZN(n8731) );
  INV_X1 U3340 ( .A(n7748), .ZN(n7911) );
  INV_X1 U3341 ( .A(n7749), .ZN(n7745) );
  OAI211_X1 U3343 ( .C1(n8011), .C2(n7830), .A(n8013), .B(n273), .ZN(n7831) );
  INV_X1 U3344 ( .A(n9121), .ZN(n9124) );
  NOR2_X1 U3345 ( .A1(n8815), .A2(n8813), .ZN(n9123) );
  AND2_X1 U3346 ( .A1(n7745), .A2(n7507), .ZN(n7694) );
  AND2_X1 U3347 ( .A1(n7749), .A2(n3446), .ZN(n7691) );
  OAI21_X1 U3348 ( .B1(n3445), .B2(n1308), .A(n3368), .ZN(n8125) );
  AOI21_X1 U3349 ( .B1(n7769), .B2(n3376), .A(n3375), .ZN(n8772) );
  INV_X1 U3350 ( .A(n3271), .ZN(n7758) );
  INV_X1 U3351 ( .A(n9113), .ZN(n1602) );
  AND2_X1 U3352 ( .A1(n6617), .A2(n1962), .ZN(n1961) );
  OR2_X1 U3353 ( .A1(n8786), .A2(n2499), .ZN(n2498) );
  OR2_X1 U3354 ( .A1(n9236), .A2(n9235), .ZN(n9237) );
  OAI21_X1 U3355 ( .B1(n8439), .B2(n261), .A(n8789), .ZN(n1737) );
  AOI21_X1 U3356 ( .B1(n8332), .B2(n7533), .A(n8499), .ZN(n2747) );
  AOI21_X1 U3357 ( .B1(n19518), .B2(n8920), .A(n8923), .ZN(n2746) );
  INV_X1 U3359 ( .A(n9067), .ZN(n2503) );
  AOI21_X1 U3360 ( .B1(n9134), .B2(n9213), .A(n1324), .ZN(n1323) );
  XNOR2_X1 U3361 ( .A(n10280), .B(n10087), .ZN(n10397) );
  OR2_X1 U3362 ( .A1(n9069), .A2(n2749), .ZN(n8075) );
  OAI211_X1 U3363 ( .C1(n9840), .C2(n2749), .A(n9839), .B(n9838), .ZN(n9841)
         );
  XNOR2_X1 U3364 ( .A(n3628), .B(n10091), .ZN(n1040) );
  OR2_X1 U3365 ( .A1(n7661), .A2(n8596), .ZN(n2478) );
  OR2_X1 U3366 ( .A1(n8924), .A2(n8749), .ZN(n2479) );
  AND2_X1 U3367 ( .A1(n9167), .A2(n9171), .ZN(n7989) );
  NAND2_X1 U3368 ( .A1(n2300), .A2(n2299), .ZN(n10542) );
  OR2_X1 U3369 ( .A1(n9064), .A2(n8829), .ZN(n2299) );
  NAND2_X1 U3370 ( .A1(n8922), .A2(n2301), .ZN(n10039) );
  AND2_X1 U3371 ( .A1(n8411), .A2(n9233), .ZN(n2650) );
  OAI21_X1 U3372 ( .B1(n9238), .B2(n8411), .A(n2653), .ZN(n2651) );
  AND2_X1 U3373 ( .A1(n11883), .A2(n3441), .ZN(n11887) );
  OR2_X1 U3374 ( .A1(n8941), .A2(n8945), .ZN(n2400) );
  OR2_X1 U3375 ( .A1(n3400), .A2(n12634), .ZN(n1387) );
  OR2_X1 U3376 ( .A1(n9147), .A2(n9145), .ZN(n1542) );
  INV_X1 U3377 ( .A(n10046), .ZN(n2689) );
  OR2_X1 U3378 ( .A1(n8701), .A2(n9070), .ZN(n8169) );
  INV_X1 U3379 ( .A(n9919), .ZN(n11476) );
  INV_X1 U3381 ( .A(n11359), .ZN(n3458) );
  OR2_X1 U3382 ( .A1(n12129), .A2(n1508), .ZN(n1546) );
  INV_X1 U3383 ( .A(n10683), .ZN(n3601) );
  INV_X1 U3384 ( .A(n11500), .ZN(n3234) );
  AND2_X1 U3385 ( .A1(n19897), .A2(n20233), .ZN(n2536) );
  INV_X1 U3386 ( .A(n3260), .ZN(n12147) );
  OR2_X1 U3387 ( .A1(n11293), .A2(n11294), .ZN(n3585) );
  MUX2_X1 U3388 ( .A(n11520), .B(n11519), .S(n12533), .Z(n13293) );
  NAND3_X1 U3389 ( .A1(n12632), .A2(n1689), .A3(n1240), .ZN(n13596) );
  INV_X1 U3390 ( .A(n12002), .ZN(n12355) );
  AOI21_X1 U3391 ( .B1(n1396), .B2(n1397), .A(n12338), .ZN(n11669) );
  NOR2_X1 U3393 ( .A1(n3781), .A2(n11699), .ZN(n3780) );
  NOR2_X1 U3396 ( .A1(n11642), .A2(n11586), .ZN(n11590) );
  XNOR2_X1 U3397 ( .A(n13293), .B(n13344), .ZN(n13569) );
  OR2_X1 U3398 ( .A1(n11018), .A2(n12576), .ZN(n2345) );
  INV_X1 U3399 ( .A(n11730), .ZN(n11017) );
  AOI22_X1 U3400 ( .A1(n11938), .A2(n12443), .B1(n11937), .B2(n1522), .ZN(
        n11941) );
  OR2_X1 U3401 ( .A1(n11943), .A2(n11942), .ZN(n1400) );
  XNOR2_X1 U3402 ( .A(n1260), .B(n13330), .ZN(n13332) );
  OAI21_X1 U3403 ( .B1(n1578), .B2(n11953), .A(n11659), .ZN(n3024) );
  AND3_X1 U3404 ( .A1(n1633), .A2(n12002), .A3(n11032), .ZN(n1634) );
  OR2_X1 U3405 ( .A1(n1636), .A2(n9380), .ZN(n1635) );
  AOI22_X1 U3406 ( .A1(n11775), .A2(n12281), .B1(n11776), .B2(n12282), .ZN(
        n11780) );
  XNOR2_X1 U3407 ( .A(n13201), .B(n13202), .ZN(n14021) );
  AND2_X1 U3408 ( .A1(n12684), .A2(n12429), .ZN(n3647) );
  AND2_X1 U3409 ( .A1(n12525), .A2(n12528), .ZN(n12172) );
  OR2_X1 U3410 ( .A1(n12231), .A2(n11646), .ZN(n12233) );
  AND2_X1 U3411 ( .A1(n11033), .A2(n11032), .ZN(n3536) );
  XNOR2_X1 U3412 ( .A(n13319), .B(n13596), .ZN(n13842) );
  OR2_X1 U3414 ( .A1(n3156), .A2(n19728), .ZN(n3154) );
  OR2_X1 U3415 ( .A1(n14032), .A2(n14642), .ZN(n2972) );
  INV_X1 U3416 ( .A(n15120), .ZN(n1802) );
  NOR2_X1 U3417 ( .A1(n14487), .A2(n14172), .ZN(n14481) );
  INV_X1 U3418 ( .A(n13872), .ZN(n14651) );
  NOR2_X1 U3419 ( .A1(n14516), .A2(n14321), .ZN(n14519) );
  XNOR2_X1 U3421 ( .A(n13061), .B(n13062), .ZN(n15119) );
  XNOR2_X1 U3423 ( .A(n2947), .B(n13549), .ZN(n13553) );
  OR2_X1 U3424 ( .A1(n13908), .A2(n14203), .ZN(n13909) );
  INV_X1 U3425 ( .A(n13927), .ZN(n14447) );
  NOR2_X1 U3426 ( .A1(n192), .A2(n19740), .ZN(n15335) );
  AND2_X1 U3427 ( .A1(n15445), .A2(n15678), .ZN(n2437) );
  OAI21_X1 U3428 ( .B1(n15076), .B2(n15077), .A(n15906), .ZN(n1412) );
  OR2_X1 U3429 ( .A1(n3019), .A2(n3778), .ZN(n3576) );
  NOR2_X1 U3430 ( .A1(n15081), .A2(n15430), .ZN(n15433) );
  AND2_X1 U3431 ( .A1(n14371), .A2(n2721), .ZN(n2720) );
  AND3_X1 U3432 ( .A1(n1181), .A2(n1925), .A3(n20094), .ZN(n15877) );
  NAND3_X1 U3433 ( .A1(n15189), .A2(n14935), .A3(n13933), .ZN(n1757) );
  OR2_X1 U3435 ( .A1(n3688), .A2(n15768), .ZN(n3686) );
  OR2_X1 U3436 ( .A1(n14938), .A2(n20449), .ZN(n3136) );
  NOR2_X1 U3437 ( .A1(n18948), .A2(n18946), .ZN(n3546) );
  OR2_X1 U3438 ( .A1(n15703), .A2(n15702), .ZN(n1877) );
  AND2_X1 U3439 ( .A1(n2364), .A2(n2363), .ZN(n2862) );
  AOI21_X1 U3440 ( .B1(n15439), .B2(n15775), .A(n1639), .ZN(n15440) );
  XNOR2_X1 U3441 ( .A(n16335), .B(n16084), .ZN(n16696) );
  INV_X1 U3444 ( .A(n17098), .ZN(n15970) );
  XNOR2_X1 U3445 ( .A(n16597), .B(n16598), .ZN(n19389) );
  AND2_X1 U3446 ( .A1(n19501), .A2(n18382), .ZN(n2794) );
  INV_X1 U3447 ( .A(n17221), .ZN(n3389) );
  INV_X1 U3448 ( .A(n16251), .ZN(n17211) );
  NOR2_X1 U3449 ( .A1(n17211), .A2(n19975), .ZN(n17214) );
  AND2_X1 U3450 ( .A1(n17210), .A2(n17208), .ZN(n2841) );
  XNOR2_X1 U3451 ( .A(n3736), .B(n16240), .ZN(n3735) );
  XNOR2_X1 U3452 ( .A(n16921), .B(n17291), .ZN(n3574) );
  XNOR2_X1 U3453 ( .A(n16361), .B(n16362), .ZN(n18112) );
  NOR2_X1 U3454 ( .A1(n17080), .A2(n17824), .ZN(n3293) );
  XNOR2_X1 U3455 ( .A(n16033), .B(n17371), .ZN(n17181) );
  XNOR2_X1 U3456 ( .A(n16040), .B(n16041), .ZN(n16781) );
  NOR2_X1 U3457 ( .A1(n4011), .A2(n1537), .ZN(n1536) );
  INV_X1 U3458 ( .A(n20002), .ZN(n3451) );
  OR2_X1 U3459 ( .A1(n4960), .A2(n292), .ZN(n4898) );
  INV_X1 U3461 ( .A(n5075), .ZN(n4457) );
  OR2_X1 U3462 ( .A1(n4539), .A2(n4350), .ZN(n4348) );
  AND2_X1 U3463 ( .A1(n3607), .A2(n3752), .ZN(n3606) );
  INV_X1 U3465 ( .A(n5088), .ZN(n5090) );
  OAI211_X1 U3466 ( .C1(n5069), .C2(n2971), .A(n5073), .B(n291), .ZN(n5505) );
  OR2_X1 U3467 ( .A1(n4438), .A2(n4804), .ZN(n2115) );
  INV_X1 U3468 ( .A(n5866), .ZN(n2158) );
  OR2_X1 U3470 ( .A1(n5674), .A2(n5424), .ZN(n4212) );
  AND2_X1 U3471 ( .A1(n6113), .A2(n6107), .ZN(n5658) );
  OR2_X1 U3472 ( .A1(n5104), .A2(n5102), .ZN(n1420) );
  AOI22_X1 U3473 ( .A1(n4885), .A2(n4946), .B1(n4467), .B2(n4002), .ZN(n5250)
         );
  OR2_X1 U3474 ( .A1(n3760), .A2(n4540), .ZN(n3759) );
  INV_X1 U3475 ( .A(n287), .ZN(n3071) );
  INV_X1 U3476 ( .A(n5401), .ZN(n4282) );
  INV_X1 U3477 ( .A(n6183), .ZN(n3196) );
  OR2_X1 U3478 ( .A1(n5114), .A2(n1915), .ZN(n3650) );
  OR2_X1 U3479 ( .A1(n5798), .A2(n1776), .ZN(n5156) );
  OR2_X1 U3480 ( .A1(n4722), .A2(n5076), .ZN(n1569) );
  INV_X1 U3481 ( .A(n5927), .ZN(n6026) );
  OR2_X1 U3482 ( .A1(n5200), .A2(n5492), .ZN(n6092) );
  OR2_X1 U3483 ( .A1(n5697), .A2(n5699), .ZN(n5528) );
  OAI21_X1 U3484 ( .B1(n5929), .B2(n5030), .A(n3371), .ZN(n5521) );
  OAI211_X1 U3485 ( .C1(n6206), .C2(n287), .A(n3044), .B(n6204), .ZN(n3672) );
  AND2_X1 U3486 ( .A1(n6207), .A2(n6208), .ZN(n1890) );
  OR2_X1 U3487 ( .A1(n4449), .A2(n5107), .ZN(n3453) );
  OR2_X1 U3488 ( .A1(n5188), .A2(n5675), .ZN(n2978) );
  AOI21_X1 U3489 ( .B1(n5969), .B2(n5973), .A(n971), .ZN(n5977) );
  OR2_X1 U3490 ( .A1(n5044), .A2(n5045), .ZN(n4444) );
  OR2_X1 U3491 ( .A1(n4048), .A2(n5100), .ZN(n4076) );
  NAND2_X1 U3492 ( .A1(n2870), .A2(n2873), .ZN(n5845) );
  XNOR2_X1 U3493 ( .A(n3513), .B(n6786), .ZN(n7098) );
  INV_X1 U3494 ( .A(n6687), .ZN(n3513) );
  OR2_X1 U3495 ( .A1(n5495), .A2(n5494), .ZN(n2099) );
  OR2_X1 U3496 ( .A1(n5683), .A2(n5682), .ZN(n5477) );
  NAND2_X1 U3497 ( .A1(n2640), .A2(n3351), .ZN(n2639) );
  OR2_X1 U3498 ( .A1(n5855), .A2(n6159), .ZN(n4403) );
  NOR2_X1 U3499 ( .A1(n6193), .A2(n6192), .ZN(n2869) );
  INV_X1 U3500 ( .A(n6016), .ZN(n5826) );
  OR2_X1 U3501 ( .A1(n4239), .A2(n4383), .ZN(n2214) );
  OAI21_X1 U3502 ( .B1(n7622), .B2(n8068), .A(n19901), .ZN(n2386) );
  INV_X1 U3503 ( .A(n8184), .ZN(n2649) );
  OR2_X1 U3504 ( .A1(n5474), .A2(n5475), .ZN(n1885) );
  INV_X1 U3505 ( .A(n6072), .ZN(n3999) );
  OR2_X1 U3506 ( .A1(n5216), .A2(n5360), .ZN(n1947) );
  XNOR2_X1 U3508 ( .A(n1081), .B(n6985), .ZN(n7377) );
  XNOR2_X1 U3509 ( .A(n6776), .B(n6641), .ZN(n7238) );
  OAI211_X1 U3510 ( .C1(n5993), .C2(n5818), .A(n3469), .B(n3467), .ZN(n6947)
         );
  OR2_X1 U3511 ( .A1(n3319), .A2(n6068), .ZN(n1982) );
  AND2_X1 U3512 ( .A1(n1958), .A2(n1274), .ZN(n1957) );
  AND2_X1 U3513 ( .A1(n6206), .A2(n287), .ZN(n5838) );
  OR2_X1 U3515 ( .A1(n5752), .A2(n5753), .ZN(n2294) );
  OR2_X1 U3516 ( .A1(n5320), .A2(n3319), .ZN(n6071) );
  INV_X1 U3517 ( .A(n8720), .ZN(n2756) );
  AND2_X1 U3518 ( .A1(n20154), .A2(n1560), .ZN(n7408) );
  OR2_X1 U3519 ( .A1(n7096), .A2(n20154), .ZN(n7407) );
  AND3_X1 U3520 ( .A1(n7642), .A2(n7641), .A3(n7640), .ZN(n2238) );
  INV_X1 U3521 ( .A(n8347), .ZN(n8271) );
  OR2_X1 U3522 ( .A1(n6618), .A2(n8095), .ZN(n1962) );
  INV_X1 U3523 ( .A(n9623), .ZN(n10231) );
  INV_X1 U3525 ( .A(n9006), .ZN(n8622) );
  OR2_X1 U3526 ( .A1(n9007), .A2(n9008), .ZN(n1484) );
  OR2_X1 U3528 ( .A1(n9346), .A2(n8156), .ZN(n8700) );
  OR2_X1 U3529 ( .A1(n2727), .A2(n9210), .ZN(n1326) );
  OR2_X1 U3530 ( .A1(n9252), .A2(n9251), .ZN(n1616) );
  INV_X1 U3531 ( .A(n8748), .ZN(n8747) );
  INV_X1 U3533 ( .A(n9287), .ZN(n8577) );
  OR2_X1 U3534 ( .A1(n8727), .A2(n8961), .ZN(n2850) );
  INV_X1 U3535 ( .A(n7668), .ZN(n8336) );
  AOI21_X1 U3536 ( .B1(n8728), .B2(n2955), .A(n8731), .ZN(n9382) );
  AND2_X1 U3537 ( .A1(n9121), .A2(n1233), .ZN(n8553) );
  AND2_X1 U3539 ( .A1(n9333), .A2(n9331), .ZN(n9075) );
  OR2_X1 U3540 ( .A1(n9122), .A2(n8552), .ZN(n9127) );
  OR2_X1 U3541 ( .A1(n9173), .A2(n9176), .ZN(n2618) );
  OAI211_X1 U3542 ( .C1(n9451), .C2(n6442), .A(n6441), .B(n6440), .ZN(n9957)
         );
  NAND2_X1 U3543 ( .A1(n2690), .A2(n8651), .ZN(n10351) );
  OR2_X1 U3544 ( .A1(n8660), .A2(n8995), .ZN(n3552) );
  XNOR2_X1 U3545 ( .A(n10171), .B(n19853), .ZN(n1283) );
  XNOR2_X1 U3546 ( .A(n9977), .B(n9596), .ZN(n1284) );
  XNOR2_X1 U3547 ( .A(n10472), .B(n875), .ZN(n9596) );
  XNOR2_X1 U3548 ( .A(n9646), .B(n9991), .ZN(n10348) );
  XNOR2_X1 U3549 ( .A(n9940), .B(n9939), .ZN(n10882) );
  INV_X1 U3550 ( .A(n9054), .ZN(n1761) );
  NAND2_X1 U3551 ( .A1(n8888), .A2(n1030), .ZN(n9429) );
  OR2_X1 U3552 ( .A1(n8889), .A2(n9451), .ZN(n1030) );
  INV_X1 U3553 ( .A(n11378), .ZN(n2611) );
  BUF_X1 U3554 ( .A(n10856), .Z(n11331) );
  OR2_X1 U3555 ( .A1(n8795), .A2(n9217), .ZN(n8670) );
  AOI21_X1 U3556 ( .B1(n1830), .B2(n8995), .A(n1829), .ZN(n8442) );
  AND2_X1 U3557 ( .A1(n8998), .A2(n8997), .ZN(n1829) );
  OR2_X1 U3559 ( .A1(n8420), .A2(n8445), .ZN(n8444) );
  OR2_X1 U3560 ( .A1(n9264), .A2(n9271), .ZN(n1321) );
  INV_X1 U3561 ( .A(n9583), .ZN(n9582) );
  XNOR2_X1 U3562 ( .A(n10617), .B(n3812), .ZN(n11489) );
  OR2_X1 U3563 ( .A1(n7897), .A2(n8649), .ZN(n7900) );
  OR2_X1 U3564 ( .A1(n8818), .A2(n8817), .ZN(n1964) );
  OR2_X1 U3565 ( .A1(n8785), .A2(n9149), .ZN(n8788) );
  INV_X1 U3566 ( .A(n9600), .ZN(n8769) );
  INV_X1 U3567 ( .A(n10163), .ZN(n8450) );
  INV_X1 U3568 ( .A(n9697), .ZN(n9587) );
  INV_X1 U3569 ( .A(n9430), .ZN(n9967) );
  INV_X1 U3570 ( .A(n9429), .ZN(n10304) );
  OAI211_X1 U3571 ( .C1(n8814), .C2(n8815), .A(n8813), .B(n2752), .ZN(n8456)
         );
  NOR2_X1 U3572 ( .A1(n9546), .A2(n11412), .ZN(n3617) );
  OAI21_X1 U3574 ( .B1(n2611), .B2(n11331), .A(n11375), .ZN(n2610) );
  XNOR2_X1 U3575 ( .A(n2570), .B(n9608), .ZN(n3588) );
  OR2_X1 U3576 ( .A1(n11460), .A2(n11880), .ZN(n10246) );
  NOR2_X1 U3577 ( .A1(n11093), .A2(n11446), .ZN(n11204) );
  AOI21_X1 U3578 ( .B1(n11233), .B2(n11366), .A(n1600), .ZN(n11252) );
  INV_X1 U3579 ( .A(n3482), .ZN(n3481) );
  AND2_X1 U3580 ( .A1(n11489), .A2(n11493), .ZN(n2135) );
  NOR2_X1 U3581 ( .A1(n11952), .A2(n11598), .ZN(n11658) );
  OR2_X1 U3582 ( .A1(n10998), .A2(n10999), .ZN(n2234) );
  INV_X1 U3584 ( .A(n12207), .ZN(n3692) );
  OR2_X1 U3585 ( .A1(n11401), .A2(n2724), .ZN(n1460) );
  INV_X1 U3586 ( .A(n11683), .ZN(n12577) );
  INV_X1 U3590 ( .A(n11942), .ZN(n12439) );
  AND2_X1 U3591 ( .A1(n11942), .A2(n12110), .ZN(n11938) );
  INV_X1 U3592 ( .A(n12606), .ZN(n12603) );
  OR2_X1 U3593 ( .A1(n11323), .A2(n11324), .ZN(n10806) );
  BUF_X1 U3595 ( .A(n13451), .Z(n12859) );
  NOR2_X1 U3596 ( .A1(n20363), .A2(n924), .ZN(n3811) );
  OR2_X1 U3598 ( .A1(n12416), .A2(n11602), .ZN(n2760) );
  AND2_X1 U3599 ( .A1(n246), .A2(n180), .ZN(n3405) );
  INV_X1 U3600 ( .A(n12429), .ZN(n12685) );
  OAI21_X1 U3601 ( .B1(n1547), .B2(n11642), .A(n1546), .ZN(n11705) );
  XNOR2_X1 U3602 ( .A(n13596), .B(n13715), .ZN(n13204) );
  INV_X1 U3603 ( .A(n12041), .ZN(n12283) );
  INV_X1 U3605 ( .A(n924), .ZN(n3164) );
  XNOR2_X1 U3606 ( .A(n13103), .B(n13383), .ZN(n13631) );
  NOR2_X1 U3607 ( .A1(n11194), .A2(n3234), .ZN(n11195) );
  OAI21_X1 U3608 ( .B1(n11618), .B2(n11897), .A(n11896), .ZN(n13686) );
  AND2_X1 U3609 ( .A1(n248), .A2(n12568), .ZN(n11893) );
  OR2_X1 U3610 ( .A1(n11173), .A2(n10912), .ZN(n3360) );
  AOI21_X1 U3611 ( .B1(n11210), .B2(n11480), .A(n2536), .ZN(n11215) );
  XNOR2_X1 U3613 ( .A(n12745), .B(n13634), .ZN(n12996) );
  XNOR2_X1 U3614 ( .A(n13677), .B(n13833), .ZN(n13433) );
  XNOR2_X1 U3616 ( .A(n12713), .B(n13330), .ZN(n2947) );
  OR2_X1 U3617 ( .A1(n14790), .A2(n14787), .ZN(n14102) );
  OR2_X1 U3618 ( .A1(n14775), .A2(n14781), .ZN(n13905) );
  OR2_X1 U3619 ( .A1(n13270), .A2(n13275), .ZN(n1304) );
  OR2_X1 U3620 ( .A1(n11627), .A2(n12237), .ZN(n3754) );
  OR2_X1 U3621 ( .A1(n11628), .A2(n12237), .ZN(n2910) );
  INV_X1 U3622 ( .A(n13335), .ZN(n2312) );
  OR2_X1 U3623 ( .A1(n14556), .A2(n14554), .ZN(n2125) );
  OAI211_X1 U3624 ( .C1(n11030), .C2(n12355), .A(n3278), .B(n1637), .ZN(n3276)
         );
  INV_X1 U3625 ( .A(n2748), .ZN(n14275) );
  INV_X1 U3626 ( .A(n19781), .ZN(n1295) );
  XNOR2_X1 U3627 ( .A(n2657), .B(n12913), .ZN(n3236) );
  AND2_X1 U3628 ( .A1(n12321), .A2(n2838), .ZN(n14850) );
  NOR2_X1 U3629 ( .A1(n14623), .A2(n19875), .ZN(n15316) );
  INV_X1 U3630 ( .A(n19906), .ZN(n14612) );
  INV_X1 U3631 ( .A(n14268), .ZN(n14740) );
  INV_X1 U3632 ( .A(n14693), .ZN(n1104) );
  NOR2_X1 U3633 ( .A1(n14935), .A2(n15504), .ZN(n3778) );
  NOR2_X1 U3634 ( .A1(n14641), .A2(n14637), .ZN(n14635) );
  INV_X1 U3635 ( .A(n14148), .ZN(n14237) );
  OR2_X1 U3636 ( .A1(n14497), .A2(n1089), .ZN(n1876) );
  AND2_X1 U3637 ( .A1(n2748), .A2(n14566), .ZN(n14276) );
  AND2_X1 U3638 ( .A1(n14673), .A2(n13981), .ZN(n14263) );
  INV_X1 U3639 ( .A(n14746), .ZN(n3158) );
  AND2_X1 U3640 ( .A1(n15906), .A2(n2723), .ZN(n2722) );
  INV_X1 U3641 ( .A(n19986), .ZN(n13913) );
  OR2_X1 U3642 ( .A1(n14828), .A2(n14826), .ZN(n13914) );
  AND2_X1 U3643 ( .A1(n13904), .A2(n3697), .ZN(n3696) );
  OR2_X1 U3645 ( .A1(n14728), .A2(n986), .ZN(n1642) );
  OR2_X1 U3646 ( .A1(n14644), .A2(n12973), .ZN(n13986) );
  NOR2_X1 U3647 ( .A1(n15378), .A2(n14874), .ZN(n14875) );
  XNOR2_X1 U3648 ( .A(n1809), .B(n12672), .ZN(n14420) );
  XNOR2_X1 U3649 ( .A(n12678), .B(n12677), .ZN(n14052) );
  OR2_X1 U3650 ( .A1(n20147), .A2(n15409), .ZN(n2129) );
  OR2_X1 U3651 ( .A1(n15544), .A2(n15070), .ZN(n2800) );
  INV_X1 U3652 ( .A(n15608), .ZN(n3427) );
  OR2_X1 U3653 ( .A1(n15615), .A2(n15071), .ZN(n15407) );
  INV_X1 U3654 ( .A(n17128), .ZN(n3273) );
  OAI211_X1 U3655 ( .C1(n14691), .C2(n19895), .A(n14693), .B(n2094), .ZN(n2186) );
  INV_X1 U3656 ( .A(n15625), .ZN(n15836) );
  OR2_X1 U3657 ( .A1(n15914), .A2(n15915), .ZN(n1152) );
  INV_X1 U3658 ( .A(n15409), .ZN(n15413) );
  AND2_X1 U3659 ( .A1(n14514), .A2(n14323), .ZN(n3149) );
  INV_X1 U3660 ( .A(n15353), .ZN(n1155) );
  OR2_X1 U3661 ( .A1(n198), .A2(n20178), .ZN(n15715) );
  OR2_X1 U3662 ( .A1(n15870), .A2(n15709), .ZN(n15711) );
  OAI21_X1 U3663 ( .B1(n2674), .B2(n2677), .A(n2673), .ZN(n15712) );
  INV_X1 U3664 ( .A(n2678), .ZN(n2674) );
  NOR2_X1 U3665 ( .A1(n18105), .A2(n17954), .ZN(n2661) );
  OR2_X1 U3666 ( .A1(n14016), .A2(n14015), .ZN(n2110) );
  INV_X1 U3667 ( .A(n17946), .ZN(n3475) );
  NOR2_X1 U3668 ( .A1(n15030), .A2(n15380), .ZN(n2988) );
  NOR2_X1 U3669 ( .A1(n16373), .A2(n2385), .ZN(n16051) );
  AND2_X1 U3670 ( .A1(n16373), .A2(n2385), .ZN(n16052) );
  INV_X1 U3671 ( .A(n2216), .ZN(n3102) );
  OR2_X1 U3673 ( .A1(n19891), .A2(n15828), .ZN(n14581) );
  OR2_X1 U3675 ( .A1(n17511), .A2(n16633), .ZN(n2335) );
  OAI21_X1 U3676 ( .B1(n20240), .B2(n19352), .A(n2668), .ZN(n16638) );
  AND2_X1 U3677 ( .A1(n20436), .A2(n17238), .ZN(n3485) );
  OR2_X1 U3678 ( .A1(n19647), .A2(n20436), .ZN(n3486) );
  OAI21_X1 U3681 ( .B1(n17492), .B2(n17491), .A(n17155), .ZN(n17158) );
  INV_X1 U3682 ( .A(n18131), .ZN(n17777) );
  AND2_X1 U3683 ( .A1(n20101), .A2(n19744), .ZN(n17449) );
  BUF_X1 U3684 ( .A(n18138), .Z(n18264) );
  XNOR2_X1 U3685 ( .A(n1529), .B(n1528), .ZN(n17981) );
  XNOR2_X1 U3686 ( .A(n17297), .B(n17301), .ZN(n1528) );
  XNOR2_X1 U3687 ( .A(n1417), .B(n17290), .ZN(n3207) );
  NOR2_X1 U3688 ( .A1(n225), .A2(n18016), .ZN(n18979) );
  XNOR2_X1 U3689 ( .A(n16138), .B(n16137), .ZN(n16731) );
  INV_X1 U3692 ( .A(n3287), .ZN(n3150) );
  XNOR2_X1 U3693 ( .A(n2994), .B(n16825), .ZN(n2991) );
  XNOR2_X1 U3694 ( .A(n17355), .B(n3749), .ZN(n2993) );
  AND2_X1 U3695 ( .A1(n17069), .A2(n19707), .ZN(n17184) );
  INV_X1 U3696 ( .A(n17887), .ZN(n1907) );
  AND2_X1 U3697 ( .A1(n17536), .A2(n17537), .ZN(n3535) );
  INV_X1 U3698 ( .A(n16465), .ZN(n1115) );
  OR2_X1 U3699 ( .A1(n17211), .A2(n20092), .ZN(n1395) );
  OR2_X1 U3700 ( .A1(n20111), .A2(n18392), .ZN(n3455) );
  NAND2_X1 U3701 ( .A1(n20111), .A2(n2793), .ZN(n1733) );
  INV_X1 U3703 ( .A(n18078), .ZN(n1728) );
  INV_X1 U3704 ( .A(n19352), .ZN(n2669) );
  NAND2_X1 U3705 ( .A1(n16468), .A2(n17507), .ZN(n3080) );
  OAI21_X1 U3706 ( .B1(n17214), .B2(n2841), .A(n20135), .ZN(n1844) );
  NOR2_X1 U3707 ( .A1(n16249), .A2(n16248), .ZN(n18501) );
  AND2_X1 U3712 ( .A1(n17789), .A2(n1668), .ZN(n19157) );
  OAI21_X1 U3713 ( .B1(n17596), .B2(n16657), .A(n16656), .ZN(n19452) );
  OR2_X1 U3714 ( .A1(n3078), .A2(n4952), .ZN(n4910) );
  NOR2_X1 U3715 ( .A1(n5018), .A2(n4555), .ZN(n3683) );
  INV_X1 U3716 ( .A(n5520), .ZN(n3410) );
  AND2_X1 U3717 ( .A1(n19789), .A2(n6027), .ZN(n5030) );
  OR2_X1 U3718 ( .A1(n4355), .A2(n4601), .ZN(n3095) );
  INV_X1 U3719 ( .A(n6101), .ZN(n5664) );
  OR2_X1 U3721 ( .A1(n4482), .A2(n4965), .ZN(n4481) );
  INV_X1 U3724 ( .A(n4960), .ZN(n3657) );
  INV_X1 U3725 ( .A(n5023), .ZN(n4765) );
  OR2_X1 U3726 ( .A1(n1232), .A2(n5073), .ZN(n3838) );
  NOR2_X1 U3727 ( .A1(n6171), .A2(n6168), .ZN(n2434) );
  AND2_X1 U3728 ( .A1(n6172), .A2(n6171), .ZN(n2435) );
  INV_X1 U3729 ( .A(n6172), .ZN(n2629) );
  OR2_X1 U3730 ( .A1(n4840), .A2(n4656), .ZN(n3980) );
  AND2_X1 U3731 ( .A1(n6202), .A2(n6201), .ZN(n1891) );
  OR2_X1 U3732 ( .A1(n5363), .A2(n5364), .ZN(n5464) );
  INV_X1 U3733 ( .A(n5631), .ZN(n5467) );
  INV_X1 U3734 ( .A(n6118), .ZN(n3483) );
  OR2_X1 U3735 ( .A1(n5387), .A2(n6124), .ZN(n2093) );
  INV_X1 U3736 ( .A(n6050), .ZN(n5138) );
  INV_X1 U3737 ( .A(n5471), .ZN(n5475) );
  INV_X1 U3738 ( .A(n5569), .ZN(n6033) );
  AND2_X1 U3739 ( .A1(n5676), .A2(n5279), .ZN(n3128) );
  INV_X1 U3740 ( .A(n5628), .ZN(n5632) );
  INV_X1 U3741 ( .A(n5930), .ZN(n3434) );
  INV_X1 U3743 ( .A(n5930), .ZN(n5929) );
  OR2_X1 U3744 ( .A1(n5899), .A2(n3098), .ZN(n3096) );
  INV_X1 U3745 ( .A(n5201), .ZN(n1695) );
  AND2_X1 U3746 ( .A1(n3802), .A2(n5218), .ZN(n1465) );
  OR2_X1 U3747 ( .A1(n4745), .A2(n5005), .ZN(n4748) );
  OAI21_X1 U3748 ( .B1(n6166), .B2(n1867), .A(n6172), .ZN(n1866) );
  OR2_X1 U3749 ( .A1(n4737), .A2(n4736), .ZN(n3008) );
  NOR2_X1 U3750 ( .A1(n3606), .A2(n3605), .ZN(n3608) );
  OR2_X1 U3751 ( .A1(n5570), .A2(n5569), .ZN(n2377) );
  INV_X1 U3752 ( .A(n3188), .ZN(n6148) );
  NOR2_X1 U3754 ( .A1(n6138), .A2(n5859), .ZN(n5864) );
  OR2_X1 U3755 ( .A1(n4507), .A2(n4370), .ZN(n3907) );
  AND2_X1 U3757 ( .A1(n4305), .A2(n2490), .ZN(n4124) );
  OR2_X1 U3758 ( .A1(n4087), .A2(n19562), .ZN(n2136) );
  OR2_X1 U3759 ( .A1(n5279), .A2(n2719), .ZN(n2718) );
  INV_X1 U3760 ( .A(n5444), .ZN(n5647) );
  INV_X1 U3761 ( .A(n2557), .ZN(n6742) );
  AND2_X1 U3762 ( .A1(n6067), .A2(n6068), .ZN(n2286) );
  AND2_X1 U3763 ( .A1(n5803), .A2(n6189), .ZN(n1986) );
  INV_X1 U3765 ( .A(n6022), .ZN(n5447) );
  AND2_X1 U3766 ( .A1(n3418), .A2(n9300), .ZN(n2985) );
  OR2_X1 U3767 ( .A1(n7974), .A2(n7972), .ZN(n2176) );
  OR2_X1 U3768 ( .A1(n5397), .A2(n5251), .ZN(n5399) );
  OR2_X1 U3770 ( .A1(n5826), .A2(n1096), .ZN(n1095) );
  OR2_X1 U3771 ( .A1(n6175), .A2(n170), .ZN(n6177) );
  INV_X1 U3772 ( .A(n8284), .ZN(n3660) );
  OR2_X1 U3773 ( .A1(n5235), .A2(n1746), .ZN(n1745) );
  NOR2_X1 U3774 ( .A1(n5793), .A2(n5429), .ZN(n2880) );
  OR2_X1 U3775 ( .A1(n7990), .A2(n7096), .ZN(n8013) );
  OR2_X1 U3776 ( .A1(n8014), .A2(n7096), .ZN(n7828) );
  OR2_X1 U3777 ( .A1(n8070), .A2(n7420), .ZN(n2379) );
  OR2_X1 U3778 ( .A1(n6023), .A2(n6022), .ZN(n1483) );
  INV_X1 U3779 ( .A(n6046), .ZN(n5777) );
  AND2_X1 U3780 ( .A1(n8271), .A2(n8272), .ZN(n1608) );
  NAND3_X1 U3781 ( .A1(n1568), .A2(n5384), .A3(n1570), .ZN(n7065) );
  OR2_X1 U3782 ( .A1(n5385), .A2(n19475), .ZN(n1570) );
  OR2_X1 U3784 ( .A1(n5870), .A2(n6124), .ZN(n2175) );
  OR2_X1 U3785 ( .A1(n7930), .A2(n2030), .ZN(n1402) );
  XNOR2_X1 U3786 ( .A(n5337), .B(n6630), .ZN(n7600) );
  INV_X1 U3787 ( .A(n8132), .ZN(n7497) );
  INV_X1 U3788 ( .A(n8220), .ZN(n3655) );
  XNOR2_X1 U3789 ( .A(n3068), .B(n7304), .ZN(n3067) );
  INV_X1 U3792 ( .A(n8114), .ZN(n1143) );
  AND2_X1 U3793 ( .A1(n8060), .A2(n8062), .ZN(n4730) );
  AND2_X1 U3794 ( .A1(n8344), .A2(n8341), .ZN(n3122) );
  AND2_X1 U3795 ( .A1(n8239), .A2(n8238), .ZN(n2987) );
  OR2_X1 U3796 ( .A1(n7432), .A2(n2687), .ZN(n7433) );
  AND2_X1 U3797 ( .A1(n7416), .A2(n8068), .ZN(n8793) );
  INV_X1 U3798 ( .A(n8603), .ZN(n8952) );
  INV_X1 U3799 ( .A(n7898), .ZN(n1405) );
  OR2_X1 U3800 ( .A1(n7618), .A2(n8204), .ZN(n1410) );
  AOI21_X1 U3801 ( .B1(n266), .B2(n9241), .A(n6587), .ZN(n2476) );
  INV_X1 U3802 ( .A(n9129), .ZN(n8805) );
  INV_X1 U3803 ( .A(n7445), .ZN(n8281) );
  INV_X1 U3804 ( .A(n8068), .ZN(n8181) );
  INV_X1 U3806 ( .A(n8354), .ZN(n7695) );
  AND2_X1 U3807 ( .A1(n6750), .A2(n8142), .ZN(n1197) );
  OAI21_X1 U3808 ( .B1(n8264), .B2(n8262), .A(n3765), .ZN(n6701) );
  OAI21_X1 U3809 ( .B1(n7556), .B2(n1791), .A(n7558), .ZN(n8500) );
  OR2_X1 U3810 ( .A1(n7678), .A2(n8363), .ZN(n3491) );
  OAI21_X1 U3811 ( .B1(n8264), .B2(n8261), .A(n8263), .ZN(n3597) );
  AND2_X1 U3812 ( .A1(n8420), .A2(n9210), .ZN(n8803) );
  OR2_X1 U3813 ( .A1(n8111), .A2(n8098), .ZN(n7436) );
  INV_X1 U3814 ( .A(n8248), .ZN(n3312) );
  OR2_X1 U3815 ( .A1(n8250), .A2(n8248), .ZN(n3311) );
  OAI22_X1 U3816 ( .A1(n1810), .A2(n8294), .B1(n7469), .B2(n8031), .ZN(n8811)
         );
  AND2_X1 U3817 ( .A1(n7469), .A2(n7471), .ZN(n1810) );
  INV_X1 U3818 ( .A(n1560), .ZN(n8015) );
  AND2_X1 U3819 ( .A1(n7466), .A2(n7811), .ZN(n7467) );
  AND2_X1 U3820 ( .A1(n9210), .A2(n9135), .ZN(n1324) );
  INV_X1 U3821 ( .A(n1567), .ZN(n8515) );
  AND2_X1 U3822 ( .A1(n8140), .A2(n8347), .ZN(n3250) );
  NOR2_X1 U3823 ( .A1(n8140), .A2(n8352), .ZN(n8270) );
  INV_X1 U3824 ( .A(n9357), .ZN(n1204) );
  OR2_X1 U3825 ( .A1(n9359), .A2(n9528), .ZN(n1201) );
  OR2_X1 U3826 ( .A1(n9215), .A2(n9214), .ZN(n1333) );
  NOR2_X1 U3827 ( .A1(n9176), .A2(n8761), .ZN(n8693) );
  XNOR2_X1 U3828 ( .A(n9934), .B(n6461), .ZN(n9935) );
  INV_X1 U3829 ( .A(n9105), .ZN(n8779) );
  NOR2_X1 U3830 ( .A1(n8077), .A2(n3795), .ZN(n3794) );
  INV_X1 U3831 ( .A(n9266), .ZN(n1587) );
  OR2_X1 U3833 ( .A1(n8998), .A2(n8772), .ZN(n1831) );
  AND2_X1 U3834 ( .A1(n7408), .A2(n7826), .ZN(n2405) );
  AND2_X1 U3835 ( .A1(n8272), .A2(n8349), .ZN(n1607) );
  INV_X1 U3836 ( .A(n6656), .ZN(n9190) );
  INV_X1 U3838 ( .A(n9453), .ZN(n8565) );
  OR2_X1 U3839 ( .A1(n7863), .A2(n1502), .ZN(n1499) );
  OR2_X1 U3840 ( .A1(n8146), .A2(n8145), .ZN(n8147) );
  OR2_X1 U3841 ( .A1(n8708), .A2(n1037), .ZN(n9182) );
  INV_X1 U3842 ( .A(n1032), .ZN(n10016) );
  BUF_X1 U3843 ( .A(n8550), .Z(n8818) );
  AND2_X1 U3844 ( .A1(n9262), .A2(n9266), .ZN(n8771) );
  INV_X1 U3847 ( .A(n1037), .ZN(n2653) );
  AND2_X1 U3848 ( .A1(n8708), .A2(n1037), .ZN(n8630) );
  INV_X1 U3850 ( .A(n7562), .ZN(n7564) );
  OR2_X1 U3851 ( .A1(n9300), .A2(n9018), .ZN(n9019) );
  INV_X1 U3852 ( .A(n8846), .ZN(n9298) );
  INV_X1 U3853 ( .A(n9624), .ZN(n9978) );
  AND2_X1 U3854 ( .A1(n9836), .A2(n2749), .ZN(n8467) );
  AND2_X1 U3855 ( .A1(n9305), .A2(n9228), .ZN(n1752) );
  INV_X1 U3856 ( .A(n20011), .ZN(n1754) );
  INV_X1 U3857 ( .A(n8500), .ZN(n9363) );
  INV_X1 U3858 ( .A(n8961), .ZN(n8726) );
  OR2_X1 U3859 ( .A1(n7659), .A2(n9038), .ZN(n2336) );
  INV_X1 U3861 ( .A(n8729), .ZN(n8939) );
  AND2_X1 U3862 ( .A1(n20146), .A2(n9129), .ZN(n9202) );
  INV_X1 U3863 ( .A(n9201), .ZN(n8665) );
  AND2_X1 U3864 ( .A1(n9130), .A2(n9201), .ZN(n9782) );
  INV_X1 U3865 ( .A(n8812), .ZN(n8552) );
  OR2_X1 U3866 ( .A1(n7477), .A2(n7476), .ZN(n3609) );
  OR2_X1 U3867 ( .A1(n8815), .A2(n8812), .ZN(n2752) );
  OR2_X1 U3868 ( .A1(n3518), .A2(n7752), .ZN(n1401) );
  INV_X1 U3869 ( .A(n8124), .ZN(n3520) );
  INV_X1 U3872 ( .A(n10805), .ZN(n10802) );
  MUX2_X1 U3873 ( .A(n9455), .B(n9454), .S(n9453), .Z(n9868) );
  AND2_X1 U3874 ( .A1(n10649), .A2(n10945), .ZN(n11156) );
  OR2_X1 U3875 ( .A1(n10960), .A2(n10701), .ZN(n9614) );
  XNOR2_X1 U3876 ( .A(n9429), .B(n9430), .ZN(n1029) );
  OR2_X1 U3877 ( .A1(n10971), .A2(n11162), .ZN(n3487) );
  NOR2_X1 U3878 ( .A1(n2498), .A2(n9145), .ZN(n7942) );
  OR2_X1 U3879 ( .A1(n11430), .A2(n11428), .ZN(n1970) );
  XNOR2_X1 U3880 ( .A(n10496), .B(n10495), .ZN(n10783) );
  INV_X1 U3881 ( .A(n11440), .ZN(n2272) );
  INV_X1 U3882 ( .A(n9960), .ZN(n2506) );
  XNOR2_X1 U3883 ( .A(n9778), .B(n1032), .ZN(n9860) );
  XNOR2_X1 U3884 ( .A(n9389), .B(n9390), .ZN(n10946) );
  OR2_X1 U3885 ( .A1(n9381), .A2(n9382), .ZN(n9383) );
  NOR2_X1 U3886 ( .A1(n247), .A2(n12209), .ZN(n2713) );
  OR2_X1 U3887 ( .A1(n204), .A2(n3507), .ZN(n3712) );
  INV_X1 U3888 ( .A(n11383), .ZN(n1330) );
  INV_X1 U3889 ( .A(n12212), .ZN(n12067) );
  AND2_X1 U3890 ( .A1(n12208), .A2(n247), .ZN(n1879) );
  OAI21_X1 U3891 ( .B1(n11463), .B2(n11886), .A(n11462), .ZN(n12168) );
  OR2_X1 U3893 ( .A1(n11460), .A2(n11120), .ZN(n11124) );
  OR2_X1 U3894 ( .A1(n11256), .A2(n191), .ZN(n10805) );
  INV_X1 U3895 ( .A(n10783), .ZN(n11438) );
  NOR2_X1 U3896 ( .A1(n12084), .A2(n12422), .ZN(n2761) );
  AND2_X1 U3897 ( .A1(n12639), .A2(n12449), .ZN(n12638) );
  XNOR2_X1 U3898 ( .A(n9850), .B(n9849), .ZN(n11365) );
  XNOR2_X1 U3899 ( .A(n9853), .B(n9855), .ZN(n2744) );
  INV_X1 U3900 ( .A(n11322), .ZN(n1124) );
  INV_X1 U3902 ( .A(n12636), .ZN(n2256) );
  NOR2_X1 U3903 ( .A1(n11562), .A2(n11561), .ZN(n11563) );
  OR2_X1 U3904 ( .A1(n12274), .A2(n12273), .ZN(n11748) );
  INV_X1 U3905 ( .A(n2605), .ZN(n2604) );
  OAI21_X1 U3906 ( .B1(n2606), .B2(n2610), .A(n10858), .ZN(n2605) );
  BUF_X1 U3907 ( .A(n11709), .Z(n12153) );
  INV_X1 U3908 ( .A(n12211), .ZN(n12206) );
  INV_X1 U3909 ( .A(n11011), .ZN(n3382) );
  INV_X1 U3910 ( .A(n11513), .ZN(n11509) );
  AND4_X1 U3912 ( .A1(n3488), .A2(n3489), .A3(n10949), .A4(n3487), .ZN(n11761)
         );
  INV_X1 U3913 ( .A(n11539), .ZN(n11532) );
  INV_X1 U3914 ( .A(n12282), .ZN(n11582) );
  XNOR2_X1 U3915 ( .A(n6657), .B(n6658), .ZN(n1523) );
  OR2_X1 U3917 ( .A1(n2610), .A2(n2606), .ZN(n2607) );
  OR2_X1 U3918 ( .A1(n11889), .A2(n11890), .ZN(n3732) );
  OR2_X1 U3919 ( .A1(n11042), .A2(n11041), .ZN(n10192) );
  OR2_X1 U3920 ( .A1(n12041), .A2(n12280), .ZN(n1299) );
  AND2_X1 U3921 ( .A1(n1387), .A2(n3676), .ZN(n1414) );
  INV_X1 U3922 ( .A(n3617), .ZN(n3614) );
  INV_X1 U3923 ( .A(n10756), .ZN(n11523) );
  INV_X1 U3924 ( .A(n10742), .ZN(n11572) );
  AND2_X1 U3925 ( .A1(n11365), .A2(n11230), .ZN(n10679) );
  INV_X1 U3926 ( .A(n10677), .ZN(n11366) );
  NOR2_X1 U3927 ( .A1(n10851), .A2(n11231), .ZN(n11364) );
  INV_X1 U3928 ( .A(n19878), .ZN(n3361) );
  INV_X1 U3929 ( .A(n2598), .ZN(n2160) );
  NAND2_X1 U3930 ( .A1(n2043), .A2(n10861), .ZN(n12240) );
  AND2_X1 U3931 ( .A1(n12554), .A2(n12542), .ZN(n11795) );
  INV_X1 U3932 ( .A(n12440), .ZN(n11939) );
  AOI21_X1 U3933 ( .B1(n10871), .B2(n20235), .A(n10870), .ZN(n12617) );
  INV_X1 U3934 ( .A(n12269), .ZN(n12020) );
  OR2_X1 U3935 ( .A1(n2707), .A2(n12002), .ZN(n3241) );
  AND2_X1 U3936 ( .A1(n12250), .A2(n11733), .ZN(n1139) );
  INV_X1 U3937 ( .A(n11717), .ZN(n11776) );
  AOI21_X1 U3939 ( .B1(n10310), .B2(n11254), .A(n11327), .ZN(n10312) );
  AND2_X1 U3940 ( .A1(n3733), .A2(n12261), .ZN(n1366) );
  OR2_X1 U3941 ( .A1(n12374), .A2(n12373), .ZN(n12375) );
  OR2_X1 U3942 ( .A1(n10737), .A2(n19915), .ZN(n10739) );
  OR2_X1 U3943 ( .A1(n11599), .A2(n1578), .ZN(n3633) );
  INV_X1 U3944 ( .A(n12273), .ZN(n12298) );
  INV_X1 U3945 ( .A(n12274), .ZN(n11781) );
  AND2_X1 U3946 ( .A1(n12648), .A2(n12686), .ZN(n12646) );
  NOR2_X1 U3947 ( .A1(n3601), .A2(n1330), .ZN(n12105) );
  OR2_X1 U3948 ( .A1(n10900), .A2(n11210), .ZN(n2898) );
  OR2_X1 U3950 ( .A1(n10961), .A2(n10960), .ZN(n1673) );
  AND2_X1 U3951 ( .A1(n11761), .A2(n11586), .ZN(n1735) );
  OAI211_X1 U3952 ( .C1(n10829), .C2(n11131), .A(n11418), .B(n11051), .ZN(
        n10413) );
  OR2_X1 U3953 ( .A1(n10372), .A2(n11456), .ZN(n1307) );
  OR2_X1 U3954 ( .A1(n12002), .A2(n12354), .ZN(n3278) );
  AND2_X1 U3955 ( .A1(n11399), .A2(n2724), .ZN(n9747) );
  OR2_X1 U3958 ( .A1(n10924), .A2(n11526), .ZN(n2522) );
  INV_X1 U3959 ( .A(n1260), .ZN(n13790) );
  INV_X1 U3960 ( .A(n11646), .ZN(n1952) );
  OR2_X1 U3961 ( .A1(n11603), .A2(n12417), .ZN(n12083) );
  NOR2_X1 U3962 ( .A1(n12103), .A2(n11380), .ZN(n1280) );
  OAI21_X1 U3963 ( .B1(n10674), .B2(n10673), .A(n10672), .ZN(n12437) );
  INV_X1 U3964 ( .A(n13199), .ZN(n2657) );
  OR2_X1 U3965 ( .A1(n631), .A2(n14800), .ZN(n12321) );
  XNOR2_X1 U3966 ( .A(n20155), .B(n6461), .ZN(n2518) );
  INV_X1 U3967 ( .A(n14420), .ZN(n1808) );
  AND2_X1 U3968 ( .A1(n12295), .A2(n20363), .ZN(n2220) );
  INV_X1 U3969 ( .A(n13735), .ZN(n2764) );
  OR2_X1 U3970 ( .A1(n1819), .A2(n14269), .ZN(n14270) );
  INV_X1 U3971 ( .A(n18517), .ZN(n2954) );
  XNOR2_X1 U3972 ( .A(n13795), .B(n2323), .ZN(n3237) );
  INV_X1 U3973 ( .A(n3405), .ZN(n3396) );
  XNOR2_X1 U3974 ( .A(n1260), .B(n2035), .ZN(n11653) );
  OR2_X1 U3975 ( .A1(n11803), .A2(n19626), .ZN(n3168) );
  OR2_X1 U3976 ( .A1(n11804), .A2(n20363), .ZN(n11805) );
  OR2_X1 U3977 ( .A1(n12145), .A2(n19833), .ZN(n2147) );
  INV_X1 U3978 ( .A(n13344), .ZN(n12937) );
  INV_X1 U3979 ( .A(n13330), .ZN(n12955) );
  AND2_X1 U3980 ( .A1(n13971), .A2(n20380), .ZN(n2563) );
  AND2_X1 U3981 ( .A1(n14326), .A2(n14327), .ZN(n14353) );
  INV_X1 U3982 ( .A(n14449), .ZN(n1364) );
  OAI21_X1 U3983 ( .B1(n19907), .B2(n14148), .A(n2979), .ZN(n15424) );
  INV_X1 U3984 ( .A(n240), .ZN(n2891) );
  NOR2_X1 U3985 ( .A1(n14599), .A2(n1262), .ZN(n1261) );
  NAND2_X1 U3986 ( .A1(n2439), .A2(n13951), .ZN(n15153) );
  OAI21_X1 U3987 ( .B1(n1699), .B2(n1593), .A(n14023), .ZN(n13951) );
  BUF_X1 U3988 ( .A(n14153), .Z(n14598) );
  OR2_X1 U3989 ( .A1(n14656), .A2(n14021), .ZN(n3280) );
  NOR2_X1 U3990 ( .A1(n241), .A2(n1593), .ZN(n1740) );
  INV_X1 U3991 ( .A(n14023), .ZN(n1744) );
  OR2_X1 U3992 ( .A1(n13118), .A2(n13980), .ZN(n14674) );
  AND2_X1 U3994 ( .A1(n15256), .A2(n15828), .ZN(n3722) );
  OAI21_X1 U3995 ( .B1(n14035), .B2(n2937), .A(n13164), .ZN(n14038) );
  INV_X1 U3996 ( .A(n14481), .ZN(n2811) );
  INV_X1 U3997 ( .A(n15905), .ZN(n15008) );
  AND2_X1 U3998 ( .A1(n2696), .A2(n2695), .ZN(n2167) );
  XNOR2_X1 U3999 ( .A(n12714), .B(n2947), .ZN(n1755) );
  INV_X1 U4000 ( .A(n3252), .ZN(n3299) );
  OR2_X1 U4001 ( .A1(n14554), .A2(n14679), .ZN(n14283) );
  NAND2_X1 U4002 ( .A1(n14235), .A2(n14596), .ZN(n15430) );
  XNOR2_X1 U4003 ( .A(n13314), .B(n13315), .ZN(n2748) );
  AND2_X1 U4004 ( .A1(n20471), .A2(n14021), .ZN(n1699) );
  AND2_X1 U4005 ( .A1(n20266), .A2(n14656), .ZN(n1698) );
  INV_X1 U4006 ( .A(n15906), .ZN(n15078) );
  OR2_X1 U4007 ( .A1(n14217), .A2(n3697), .ZN(n3538) );
  OR2_X1 U4008 ( .A1(n14141), .A2(n14593), .ZN(n2809) );
  OAI211_X1 U4010 ( .C1(n20262), .C2(n14167), .A(n3088), .B(n238), .ZN(n3087)
         );
  OAI21_X1 U4011 ( .B1(n14447), .B2(n14455), .A(n1363), .ZN(n1362) );
  OR2_X1 U4012 ( .A1(n12911), .A2(n1724), .ZN(n1723) );
  OR2_X1 U4013 ( .A1(n13979), .A2(n14678), .ZN(n2353) );
  INV_X1 U4014 ( .A(n13868), .ZN(n14498) );
  OR2_X1 U4015 ( .A1(n14265), .A2(n13981), .ZN(n1573) );
  NOR2_X1 U4016 ( .A1(n15327), .A2(n2655), .ZN(n15722) );
  INV_X1 U4017 ( .A(n2655), .ZN(n15863) );
  INV_X1 U4018 ( .A(n15007), .ZN(n2578) );
  INV_X1 U4019 ( .A(n2723), .ZN(n15910) );
  INV_X1 U4020 ( .A(n15397), .ZN(n2500) );
  OAI21_X1 U4021 ( .B1(n14186), .B2(n14185), .A(n14184), .ZN(n15308) );
  INV_X1 U4022 ( .A(n1288), .ZN(n1286) );
  INV_X1 U4023 ( .A(n14935), .ZN(n15506) );
  AND2_X1 U4024 ( .A1(n15845), .A2(n15266), .ZN(n15091) );
  INV_X1 U4025 ( .A(n19007), .ZN(n1782) );
  NOR2_X1 U4026 ( .A1(n20480), .A2(n14381), .ZN(n3705) );
  AOI22_X1 U4027 ( .A1(n15007), .A2(n15906), .B1(n15907), .B2(n15905), .ZN(
        n15419) );
  INV_X1 U4030 ( .A(n15628), .ZN(n15839) );
  INV_X1 U4031 ( .A(n15573), .ZN(n1520) );
  INV_X1 U4032 ( .A(n15697), .ZN(n15386) );
  INV_X1 U4033 ( .A(n15702), .ZN(n15385) );
  INV_X1 U4034 ( .A(n15243), .ZN(n3689) );
  AND2_X1 U4035 ( .A1(n15767), .A2(n15657), .ZN(n3690) );
  INV_X1 U4036 ( .A(n15698), .ZN(n3138) );
  AND2_X1 U4037 ( .A1(n15495), .A2(n15606), .ZN(n3430) );
  INV_X1 U4038 ( .A(n15442), .ZN(n15446) );
  OAI21_X1 U4039 ( .B1(n15316), .B2(n15315), .A(n2731), .ZN(n1226) );
  NAND2_X1 U4040 ( .A1(n20506), .A2(n17078), .ZN(n1166) );
  NOR2_X1 U4041 ( .A1(n14224), .A2(n14729), .ZN(n2642) );
  INV_X1 U4042 ( .A(n19739), .ZN(n16010) );
  OR2_X1 U4043 ( .A1(n12664), .A2(n15767), .ZN(n1383) );
  OR2_X1 U4045 ( .A1(n13950), .A2(n14693), .ZN(n2952) );
  OR2_X1 U4046 ( .A1(n14387), .A2(n14695), .ZN(n2716) );
  AND2_X1 U4047 ( .A1(n19884), .A2(n1638), .ZN(n1639) );
  AND2_X1 U4048 ( .A1(n15574), .A2(n15365), .ZN(n15045) );
  INV_X1 U4049 ( .A(n19828), .ZN(n15642) );
  INV_X1 U4050 ( .A(n14119), .ZN(n14123) );
  OR2_X1 U4051 ( .A1(n14312), .A2(n14903), .ZN(n14978) );
  INV_X1 U4052 ( .A(n15682), .ZN(n2005) );
  INV_X1 U4054 ( .A(n15587), .ZN(n15990) );
  AND2_X1 U4055 ( .A1(n15282), .A2(n15284), .ZN(n1656) );
  AOI21_X1 U4056 ( .B1(n12876), .B2(n14339), .A(n19485), .ZN(n3193) );
  OR2_X1 U4058 ( .A1(n14866), .A2(n15684), .ZN(n13180) );
  OR2_X1 U4059 ( .A1(n13868), .A2(n1089), .ZN(n2276) );
  NOR2_X1 U4060 ( .A1(n15413), .A2(n15551), .ZN(n15412) );
  OR2_X1 U4061 ( .A1(n15864), .A2(n15861), .ZN(n1974) );
  NOR2_X1 U4062 ( .A1(n13906), .A2(n3696), .ZN(n3695) );
  INV_X1 U4064 ( .A(n15308), .ZN(n15306) );
  INV_X1 U4065 ( .A(n15110), .ZN(n2644) );
  OR2_X1 U4067 ( .A1(n17494), .A2(n17493), .ZN(n2422) );
  OR2_X1 U4068 ( .A1(n15407), .A2(n2803), .ZN(n2802) );
  INV_X1 U4069 ( .A(n642), .ZN(n3209) );
  XNOR2_X1 U4070 ( .A(n17289), .B(n17291), .ZN(n1417) );
  OR2_X1 U4071 ( .A1(n18927), .A2(n18928), .ZN(n1068) );
  OAI21_X1 U4073 ( .B1(n196), .B2(n16308), .A(n20162), .ZN(n3343) );
  XNOR2_X1 U4075 ( .A(n16045), .B(n16269), .ZN(n16906) );
  OR2_X1 U4077 ( .A1(n15052), .A2(n15237), .ZN(n13566) );
  XNOR2_X1 U4078 ( .A(n16330), .B(n880), .ZN(n3448) );
  XNOR2_X1 U4079 ( .A(n16374), .B(n16507), .ZN(n15726) );
  XNOR2_X1 U4080 ( .A(n14376), .B(n14375), .ZN(n17511) );
  OR2_X1 U4081 ( .A1(n17149), .A2(n17956), .ZN(n2662) );
  OR2_X1 U4082 ( .A1(n18092), .A2(n20109), .ZN(n17569) );
  OR3_X1 U4083 ( .A1(n17973), .A2(n19771), .A3(n2836), .ZN(n2835) );
  INV_X1 U4084 ( .A(n18130), .ZN(n18126) );
  OR2_X1 U4085 ( .A1(n19787), .A2(n18753), .ZN(n18263) );
  NAND4_X1 U4087 ( .A1(n3548), .A2(n3544), .A3(n3545), .A4(n3547), .ZN(n18890)
         );
  OR2_X1 U4088 ( .A1(n17812), .A2(n16959), .ZN(n3547) );
  NOR2_X1 U4089 ( .A1(n16153), .A2(n17715), .ZN(n16730) );
  OR2_X1 U4092 ( .A1(n20221), .A2(n2907), .ZN(n2906) );
  OR2_X1 U4093 ( .A1(n17891), .A2(n16261), .ZN(n3216) );
  OR2_X1 U4094 ( .A1(n17898), .A2(n17896), .ZN(n1924) );
  XNOR2_X1 U4095 ( .A(n1436), .B(n16509), .ZN(n19363) );
  OR2_X1 U4096 ( .A1(n18335), .A2(n18332), .ZN(n2219) );
  OR2_X1 U4097 ( .A1(n18404), .A2(n18425), .ZN(n1875) );
  NOR2_X1 U4098 ( .A1(n18414), .A2(n15529), .ZN(n2018) );
  AND2_X1 U4099 ( .A1(n2544), .A2(n2545), .ZN(n2546) );
  OR2_X1 U4100 ( .A1(n18423), .A2(n18412), .ZN(n2544) );
  AOI21_X1 U4101 ( .B1(n3045), .B2(n18436), .A(n18444), .ZN(n18445) );
  AND2_X1 U4102 ( .A1(n17642), .A2(n17641), .ZN(n2852) );
  AND2_X1 U4103 ( .A1(n18500), .A2(n18485), .ZN(n17639) );
  AND2_X1 U4104 ( .A1(n18497), .A2(n18498), .ZN(n1174) );
  INV_X1 U4106 ( .A(n18546), .ZN(n18552) );
  INV_X1 U4107 ( .A(n17584), .ZN(n17923) );
  AND2_X1 U4108 ( .A1(n18559), .A2(n18555), .ZN(n1862) );
  AND2_X1 U4109 ( .A1(n19509), .A2(n18600), .ZN(n1080) );
  OR2_X1 U4110 ( .A1(n19757), .A2(n18600), .ZN(n18603) );
  AND2_X1 U4111 ( .A1(n3436), .A2(n3437), .ZN(n1799) );
  INV_X1 U4112 ( .A(n18688), .ZN(n17985) );
  INV_X1 U4113 ( .A(n18671), .ZN(n17964) );
  OR2_X1 U4114 ( .A1(n18667), .A2(n18671), .ZN(n1532) );
  AND2_X1 U4115 ( .A1(n18698), .A2(n18701), .ZN(n17631) );
  OR2_X1 U4116 ( .A1(n19766), .A2(n18834), .ZN(n18814) );
  NOR2_X1 U4118 ( .A1(n18882), .A2(n18921), .ZN(n18918) );
  NOR2_X1 U4121 ( .A1(n19151), .A2(n20508), .ZN(n17807) );
  INV_X1 U4123 ( .A(n18306), .ZN(n2918) );
  OAI21_X1 U4124 ( .B1(n2918), .B2(n19165), .A(n17790), .ZN(n17793) );
  OR2_X1 U4125 ( .A1(n195), .A2(n18306), .ZN(n17789) );
  NOR2_X1 U4126 ( .A1(n20460), .A2(n19168), .ZN(n19171) );
  OR2_X1 U4127 ( .A1(n17201), .A2(n16153), .ZN(n2236) );
  INV_X1 U4128 ( .A(n17184), .ZN(n1248) );
  OR2_X1 U4129 ( .A1(n19241), .A2(n19242), .ZN(n3338) );
  INV_X1 U4130 ( .A(n17665), .ZN(n2819) );
  INV_X1 U4131 ( .A(n1205), .ZN(n19274) );
  OR2_X1 U4132 ( .A1(n20515), .A2(n18164), .ZN(n2227) );
  INV_X1 U4133 ( .A(n17542), .ZN(n2996) );
  OR2_X1 U4134 ( .A1(n19404), .A2(n16306), .ZN(n2965) );
  OR2_X1 U4135 ( .A1(n19463), .A2(n20152), .ZN(n1145) );
  OR2_X1 U4136 ( .A1(n19453), .A2(n19452), .ZN(n19456) );
  NOR2_X1 U4137 ( .A1(n212), .A2(n19459), .ZN(n2515) );
  INV_X1 U4138 ( .A(n17091), .ZN(n2516) );
  OR2_X1 U4139 ( .A1(n2514), .A2(n17095), .ZN(n2509) );
  OR2_X1 U4140 ( .A1(n17907), .A2(n18365), .ZN(n16649) );
  NAND4_X1 U4142 ( .A1(n1732), .A2(n18376), .A3(n1733), .A4(n1728), .ZN(n1727)
         );
  AND2_X1 U4143 ( .A1(n18409), .A2(n18407), .ZN(n16492) );
  OR2_X1 U4145 ( .A1(n17739), .A2(n2084), .ZN(n17740) );
  OR2_X1 U4146 ( .A1(n18583), .A2(n18596), .ZN(n3411) );
  OAI211_X1 U4147 ( .C1(n19917), .C2(n19988), .A(n3028), .B(n18857), .ZN(
        n18852) );
  INV_X1 U4148 ( .A(n610), .ZN(n2361) );
  INV_X1 U4149 ( .A(n17535), .ZN(n2193) );
  OR2_X1 U4151 ( .A1(n18164), .A2(n19298), .ZN(n1775) );
  INV_X1 U4153 ( .A(n13918), .ZN(n3516) );
  INV_X1 U4154 ( .A(n14250), .ZN(n2682) );
  INV_X1 U4155 ( .A(n8212), .ZN(n8209) );
  INV_X1 U4157 ( .A(n8262), .ZN(n3766) );
  XNOR2_X1 U4158 ( .A(n3062), .B(n13583), .ZN(n14396) );
  AND2_X1 U4159 ( .A1(n4052), .A2(n135), .ZN(n956) );
  INV_X1 U4160 ( .A(n5250), .ZN(n1838) );
  XNOR2_X1 U4161 ( .A(n962), .B(n7252), .ZN(n7801) );
  AND2_X1 U4163 ( .A1(n5968), .A2(n5967), .ZN(n957) );
  AND2_X1 U4164 ( .A1(n11446), .A2(n11201), .ZN(n958) );
  OR2_X1 U4165 ( .A1(n19885), .A2(n17559), .ZN(n959) );
  OR2_X1 U4166 ( .A1(n16462), .A2(n17483), .ZN(n960) );
  INV_X1 U4167 ( .A(n5684), .ZN(n3529) );
  INV_X1 U4168 ( .A(n18600), .ZN(n3693) );
  INV_X1 U4169 ( .A(n9047), .ZN(n3395) );
  INV_X1 U4170 ( .A(n11244), .ZN(n2861) );
  INV_X1 U4171 ( .A(n11297), .ZN(n2724) );
  XOR2_X1 U4172 ( .A(n10252), .B(n10249), .Z(n961) );
  INV_X1 U4173 ( .A(n4013), .ZN(n1537) );
  XNOR2_X1 U4174 ( .A(n10338), .B(n10337), .ZN(n11458) );
  INV_X1 U4175 ( .A(n14566), .ZN(n2282) );
  INV_X1 U4176 ( .A(n14781), .ZN(n3697) );
  XOR2_X1 U4177 ( .A(n7247), .B(n7246), .Z(n962) );
  XOR2_X1 U4178 ( .A(n17139), .B(n17138), .Z(n963) );
  XNOR2_X1 U4179 ( .A(n9631), .B(n9630), .ZN(n11381) );
  INV_X1 U4181 ( .A(n11990), .ZN(n1213) );
  INV_X1 U4184 ( .A(n12004), .ZN(n1859) );
  INV_X1 U4185 ( .A(n8179), .ZN(n1850) );
  INV_X1 U4186 ( .A(n12262), .ZN(n3734) );
  XNOR2_X1 U4187 ( .A(n1756), .B(n1755), .ZN(n14465) );
  INV_X1 U4188 ( .A(n3319), .ZN(n6069) );
  INV_X1 U4189 ( .A(n15443), .ZN(n1494) );
  OR2_X1 U4190 ( .A1(n5003), .A2(n4745), .ZN(n964) );
  OR2_X1 U4192 ( .A1(n10814), .A2(n10113), .ZN(n965) );
  OR2_X1 U4193 ( .A1(n9209), .A2(n9135), .ZN(n966) );
  OAI211_X1 U4194 ( .C1(n11396), .C2(n11395), .A(n1460), .B(n11400), .ZN(
        n12554) );
  OR2_X1 U4195 ( .A1(n12282), .A2(n11721), .ZN(n967) );
  INV_X1 U4196 ( .A(n11142), .ZN(n1749) );
  OR2_X1 U4197 ( .A1(n3373), .A2(n14020), .ZN(n968) );
  OR3_X1 U4198 ( .A1(n9178), .A2(n9177), .A3(n9176), .ZN(n969) );
  INV_X1 U4199 ( .A(n15844), .ZN(n2146) );
  OR2_X1 U4200 ( .A1(n8309), .A2(n20057), .ZN(n970) );
  INV_X1 U4202 ( .A(n4892), .ZN(n4377) );
  INV_X1 U4203 ( .A(n12617), .ZN(n1591) );
  AND2_X1 U4204 ( .A1(n5968), .A2(n5971), .ZN(n971) );
  XNOR2_X1 U4205 ( .A(n6437), .B(n6436), .ZN(n7507) );
  INV_X1 U4206 ( .A(n7750), .ZN(n7912) );
  OR2_X1 U4207 ( .A1(n9158), .A2(n8696), .ZN(n972) );
  OR2_X1 U4208 ( .A1(n4226), .A2(n4853), .ZN(n973) );
  XNOR2_X1 U4209 ( .A(n9970), .B(n9969), .ZN(n11466) );
  INV_X1 U4210 ( .A(n5563), .ZN(n2940) );
  INV_X1 U4211 ( .A(n8445), .ZN(n2727) );
  NAND3_X1 U4212 ( .A1(n17504), .A2(n19898), .A3(n19815), .ZN(n975) );
  INV_X1 U4213 ( .A(n15627), .ZN(n2472) );
  INV_X1 U4215 ( .A(n14584), .ZN(n1351) );
  XNOR2_X1 U4216 ( .A(n12367), .B(n12368), .ZN(n14584) );
  OR3_X1 U4217 ( .A1(n12016), .A2(n12262), .A3(n12264), .ZN(n976) );
  INV_X1 U4218 ( .A(n5115), .ZN(n1915) );
  INV_X1 U4219 ( .A(n17831), .ZN(n2907) );
  INV_X1 U4220 ( .A(n12437), .ZN(n1099) );
  INV_X1 U4221 ( .A(n9135), .ZN(n9213) );
  INV_X1 U4222 ( .A(n14666), .ZN(n2676) );
  XNOR2_X1 U4223 ( .A(n1524), .B(n1523), .ZN(n11158) );
  XNOR2_X1 U4224 ( .A(n13740), .B(n13739), .ZN(n14229) );
  XOR2_X1 U4225 ( .A(n13260), .B(n17089), .Z(n977) );
  INV_X1 U4226 ( .A(n5112), .ZN(n2042) );
  AND2_X1 U4227 ( .A1(n9008), .A2(n9007), .ZN(n978) );
  OAI211_X1 U4228 ( .C1(n18930), .C2(n18929), .A(n1067), .B(n1066), .ZN(n19013) );
  INV_X1 U4229 ( .A(n19013), .ZN(n2058) );
  XNOR2_X1 U4230 ( .A(n6601), .B(n6600), .ZN(n8211) );
  INV_X1 U4231 ( .A(n5328), .ZN(n6054) );
  XNOR2_X1 U4232 ( .A(n9377), .B(n9376), .ZN(n10962) );
  XOR2_X1 U4233 ( .A(n13026), .B(n13025), .Z(n979) );
  OAI22_X1 U4234 ( .A1(n11050), .A2(n11887), .B1(n11049), .B2(n11886), .ZN(
        n12263) );
  XOR2_X1 U4235 ( .A(n6946), .B(n2208), .Z(n980) );
  AND2_X1 U4236 ( .A1(n11659), .A2(n11829), .ZN(n981) );
  OR3_X1 U4238 ( .A1(n17891), .A2(n16261), .A3(n17890), .ZN(n982) );
  XNOR2_X1 U4239 ( .A(n13575), .B(n3823), .ZN(n14154) );
  INV_X1 U4240 ( .A(n14154), .ZN(n2926) );
  AND3_X1 U4241 ( .A1(n4698), .A2(n5048), .A3(n4697), .ZN(n983) );
  INV_X1 U4242 ( .A(n12684), .ZN(n2805) );
  AND2_X1 U4243 ( .A1(n20513), .A2(n14601), .ZN(n984) );
  INV_X1 U4244 ( .A(n14000), .ZN(n14624) );
  XNOR2_X1 U4246 ( .A(n6298), .B(n6297), .ZN(n6312) );
  INV_X1 U4247 ( .A(n6312), .ZN(n1726) );
  INV_X1 U4248 ( .A(n14535), .ZN(n14664) );
  XNOR2_X1 U4249 ( .A(n13163), .B(n13162), .ZN(n14535) );
  AND2_X1 U4250 ( .A1(n20261), .A2(n19985), .ZN(n985) );
  OR2_X1 U4251 ( .A1(n20451), .A2(n14724), .ZN(n986) );
  XNOR2_X1 U4252 ( .A(n2046), .B(n10025), .ZN(n10746) );
  INV_X1 U4253 ( .A(n5941), .ZN(n1835) );
  AND2_X1 U4254 ( .A1(n6050), .A2(n6049), .ZN(n987) );
  INV_X1 U4255 ( .A(n5971), .ZN(n5700) );
  AND2_X1 U4256 ( .A1(n18590), .A2(n19656), .ZN(n988) );
  INV_X1 U4257 ( .A(n12658), .ZN(n15659) );
  OR2_X1 U4258 ( .A1(n5200), .A2(n5199), .ZN(n989) );
  OR2_X1 U4259 ( .A1(n11051), .A2(n11131), .ZN(n990) );
  OR2_X1 U4260 ( .A1(n11109), .A2(n11428), .ZN(n991) );
  AND2_X1 U4261 ( .A1(n19912), .A2(n5428), .ZN(n992) );
  AND3_X1 U4263 ( .A1(n18324), .A2(n18156), .A3(n2368), .ZN(n993) );
  INV_X1 U4264 ( .A(n12110), .ZN(n12441) );
  OR2_X2 U4265 ( .A1(n4759), .A2(n4760), .ZN(n6109) );
  AND2_X1 U4266 ( .A1(n18522), .A2(n18512), .ZN(n994) );
  OR2_X1 U4267 ( .A1(n8241), .A2(n8100), .ZN(n995) );
  AND2_X1 U4268 ( .A1(n14447), .A2(n14448), .ZN(n996) );
  AND2_X1 U4269 ( .A1(n16128), .A2(n16129), .ZN(n997) );
  INV_X1 U4271 ( .A(n15815), .ZN(n3534) );
  AND2_X1 U4273 ( .A1(n15742), .A2(n15521), .ZN(n1000) );
  AND2_X1 U4274 ( .A1(n1859), .A2(n12500), .ZN(n1001) );
  INV_X1 U4275 ( .A(n3366), .ZN(n2677) );
  INV_X1 U4276 ( .A(n14667), .ZN(n3366) );
  OR2_X1 U4277 ( .A1(n3055), .A2(n8194), .ZN(n1002) );
  INV_X1 U4278 ( .A(n8657), .ZN(n3518) );
  AND2_X1 U4279 ( .A1(n12499), .A2(n201), .ZN(n1003) );
  INV_X1 U4280 ( .A(n15607), .ZN(n15606) );
  INV_X1 U4281 ( .A(n9666), .ZN(n12103) );
  XOR2_X1 U4282 ( .A(n13843), .B(n17544), .Z(n1004) );
  OR2_X1 U4283 ( .A1(n11639), .A2(n12214), .ZN(n1005) );
  OR2_X1 U4284 ( .A1(n7633), .A2(n20511), .ZN(n1006) );
  INV_X1 U4286 ( .A(n9167), .ZN(n9082) );
  AND2_X1 U4287 ( .A1(n2928), .A2(n4057), .ZN(n1007) );
  OR2_X1 U4288 ( .A1(n11977), .A2(n250), .ZN(n1008) );
  OR2_X1 U4289 ( .A1(n12262), .A2(n3731), .ZN(n1009) );
  AND2_X1 U4290 ( .A1(n19922), .A2(n8203), .ZN(n1010) );
  AND2_X1 U4291 ( .A1(n284), .A2(n5953), .ZN(n1011) );
  OR2_X1 U4292 ( .A1(n9298), .A2(n891), .ZN(n1012) );
  NAND2_X1 U4293 ( .A1(n17097), .A2(n18111), .ZN(n1013) );
  OR2_X1 U4294 ( .A1(n13507), .A2(n14498), .ZN(n1014) );
  NOR2_X2 U4295 ( .A1(n11196), .A2(n11195), .ZN(n12480) );
  INV_X1 U4296 ( .A(n12480), .ZN(n2550) );
  AND2_X1 U4297 ( .A1(n9021), .A2(n9023), .ZN(n1015) );
  NAND2_X1 U4298 ( .A1(n19033), .A2(n19992), .ZN(n1016) );
  INV_X1 U4299 ( .A(n13939), .ZN(n14422) );
  INV_X1 U4300 ( .A(n15822), .ZN(n15507) );
  AND2_X1 U4301 ( .A1(n19524), .A2(n4528), .ZN(n1017) );
  INV_X1 U4302 ( .A(n7568), .ZN(n8263) );
  OR2_X1 U4303 ( .A1(n15674), .A2(n15673), .ZN(n1018) );
  AND2_X1 U4304 ( .A1(n14935), .A2(n15187), .ZN(n1019) );
  INV_X1 U4305 ( .A(n9048), .ZN(n3394) );
  INV_X1 U4306 ( .A(n9329), .ZN(n2174) );
  OR2_X1 U4307 ( .A1(n12647), .A2(n12684), .ZN(n1020) );
  BUF_X1 U4308 ( .A(n15220), .Z(n17479) );
  INV_X1 U4309 ( .A(n15187), .ZN(n15504) );
  OR2_X1 U4310 ( .A1(n14392), .A2(n14717), .ZN(n1021) );
  OR2_X1 U4311 ( .A1(n18072), .A2(n19753), .ZN(n1022) );
  INV_X1 U4312 ( .A(n9159), .ZN(n1230) );
  OR2_X1 U4313 ( .A1(n8958), .A2(n8959), .ZN(n1023) );
  OR2_X1 U4314 ( .A1(n14266), .A2(n14265), .ZN(n1024) );
  OR2_X1 U4315 ( .A1(n6220), .A2(n5758), .ZN(n1025) );
  INV_X1 U4316 ( .A(n4840), .ZN(n4223) );
  INV_X1 U4317 ( .A(n19208), .ZN(n2943) );
  INV_X1 U4318 ( .A(n8420), .ZN(n9214) );
  AND2_X1 U4319 ( .A1(n5300), .A2(n5428), .ZN(n1026) );
  INV_X1 U4321 ( .A(n8708), .ZN(n1041) );
  NAND2_X1 U4322 ( .A1(n9082), .A2(n9166), .ZN(n1027) );
  INV_X1 U4323 ( .A(n12549), .ZN(n3615) );
  NAND3_X1 U4324 ( .A1(n4841), .A2(n3978), .A3(n20105), .ZN(n1028) );
  INV_X1 U4325 ( .A(n19410), .ZN(n3749) );
  INV_X1 U4327 ( .A(n573), .ZN(n1259) );
  INV_X1 U4328 ( .A(n2275), .ZN(n2709) );
  INV_X1 U4329 ( .A(n1911), .ZN(n1780) );
  INV_X1 U4330 ( .A(n18146), .ZN(n1228) );
  INV_X1 U4331 ( .A(n2401), .ZN(n1781) );
  INV_X1 U4332 ( .A(n18819), .ZN(n1783) );
  XNOR2_X1 U4333 ( .A(n10163), .B(n2329), .ZN(n1031) );
  NAND2_X1 U4334 ( .A1(n14547), .A2(n20266), .ZN(n1033) );
  NAND2_X1 U4336 ( .A1(n14656), .A2(n14021), .ZN(n1034) );
  NOR2_X1 U4337 ( .A1(n18319), .A2(n1035), .ZN(n3776) );
  OAI21_X1 U4339 ( .B1(n18317), .B2(n1035), .A(n18157), .ZN(n18059) );
  OAI211_X1 U4341 ( .C1(n19174), .C2(n1035), .A(n19168), .B(n19169), .ZN(
        n19173) );
  AND2_X1 U4343 ( .A1(n1041), .A2(n1037), .ZN(n3058) );
  OR2_X1 U4344 ( .A1(n1041), .A2(n1037), .ZN(n8711) );
  OAI21_X1 U4345 ( .B1(n9233), .B2(n1037), .A(n1036), .ZN(n6215) );
  NAND2_X1 U4346 ( .A1(n8411), .A2(n1037), .ZN(n1036) );
  OAI21_X1 U4347 ( .B1(n11127), .B2(n1039), .A(n1038), .ZN(n10817) );
  NAND2_X1 U4348 ( .A1(n11127), .A2(n1040), .ZN(n1038) );
  NAND2_X1 U4349 ( .A1(n20099), .A2(n1040), .ZN(n2729) );
  NAND2_X1 U4350 ( .A1(n1040), .A2(n19725), .ZN(n11359) );
  NAND3_X1 U4351 ( .A1(n9238), .A2(n8411), .A3(n2653), .ZN(n8631) );
  AOI21_X1 U4352 ( .B1(n9180), .B2(n9238), .A(n2653), .ZN(n9185) );
  NOR2_X1 U4353 ( .A1(n248), .A2(n1042), .ZN(n1044) );
  NOR2_X1 U4354 ( .A1(n11061), .A2(n12261), .ZN(n1042) );
  NAND2_X1 U4355 ( .A1(n1045), .A2(n1044), .ZN(n1043) );
  NAND2_X1 U4357 ( .A1(n248), .A2(n12262), .ZN(n12565) );
  NAND2_X1 U4358 ( .A1(n1048), .A2(n1046), .ZN(n5304) );
  NAND2_X1 U4359 ( .A1(n1047), .A2(n4457), .ZN(n1046) );
  NAND2_X1 U4361 ( .A1(n4720), .A2(n4081), .ZN(n1048) );
  NAND2_X1 U4362 ( .A1(n1049), .A2(n1163), .ZN(n4720) );
  NAND2_X1 U4363 ( .A1(n19868), .A2(n5075), .ZN(n1049) );
  NAND2_X1 U4364 ( .A1(n1472), .A2(n4667), .ZN(n5255) );
  NAND3_X1 U4365 ( .A1(n1472), .A2(n4667), .A3(n19688), .ZN(n1050) );
  NAND2_X1 U4366 ( .A1(n5257), .A2(n4668), .ZN(n1051) );
  OR2_X1 U4367 ( .A1(n12334), .A2(n11992), .ZN(n11970) );
  INV_X1 U4368 ( .A(n11240), .ZN(n11346) );
  INV_X1 U4371 ( .A(n11829), .ZN(n1578) );
  OR2_X1 U4372 ( .A1(n7855), .A2(n6830), .ZN(n7857) );
  INV_X1 U4373 ( .A(n3959), .ZN(n5580) );
  OAI21_X1 U4374 ( .B1(n12416), .B2(n11312), .A(n2758), .ZN(n13031) );
  AND2_X1 U4375 ( .A1(n4901), .A2(n4856), .ZN(n3769) );
  INV_X1 U4376 ( .A(n5663), .ZN(n6098) );
  OR2_X1 U4377 ( .A1(n5663), .A2(n5953), .ZN(n6099) );
  NOR2_X1 U4378 ( .A1(n10513), .A2(n11034), .ZN(n10836) );
  OR2_X1 U4379 ( .A1(n10783), .A2(n11034), .ZN(n2485) );
  INV_X1 U4380 ( .A(n11034), .ZN(n11435) );
  INV_X1 U4381 ( .A(n8611), .ZN(n2781) );
  OR2_X1 U4382 ( .A1(n4197), .A2(n4755), .ZN(n2034) );
  INV_X1 U4383 ( .A(n15756), .ZN(n2103) );
  OR2_X1 U4384 ( .A1(n3986), .A2(n20459), .ZN(n1719) );
  AND2_X1 U4385 ( .A1(n16810), .A2(n19655), .ZN(n17927) );
  OR2_X1 U4386 ( .A1(n19737), .A2(n19672), .ZN(n17149) );
  AND2_X1 U4388 ( .A1(n11193), .A2(n11186), .ZN(n11083) );
  XNOR2_X1 U4389 ( .A(n2211), .B(n6772), .ZN(n7686) );
  NOR2_X1 U4390 ( .A1(n10745), .A2(n20233), .ZN(n1788) );
  INV_X1 U4391 ( .A(n8253), .ZN(n6704) );
  OR2_X1 U4392 ( .A1(n8253), .A2(n8251), .ZN(n8250) );
  AND2_X1 U4393 ( .A1(n1807), .A2(n4369), .ZN(n2936) );
  INV_X1 U4394 ( .A(n1807), .ZN(n1685) );
  INV_X1 U4395 ( .A(n17686), .ZN(n1605) );
  INV_X1 U4396 ( .A(n14813), .ZN(n14812) );
  OR2_X1 U4397 ( .A1(n15582), .A2(n3315), .ZN(n15811) );
  NOR2_X1 U4398 ( .A1(n905), .A2(n8742), .ZN(n2066) );
  OR2_X1 U4399 ( .A1(n8482), .A2(n8743), .ZN(n9370) );
  NAND2_X1 U4400 ( .A1(n5568), .A2(n2377), .ZN(n1052) );
  NAND2_X1 U4401 ( .A1(n5568), .A2(n2377), .ZN(n1053) );
  NAND2_X1 U4402 ( .A1(n5568), .A2(n2377), .ZN(n7287) );
  AND2_X1 U4403 ( .A1(n8162), .A2(n7852), .ZN(n8260) );
  AND2_X1 U4405 ( .A1(n11158), .A2(n11160), .ZN(n9555) );
  AND3_X1 U4406 ( .A1(n14870), .A2(n14869), .A3(n14868), .ZN(n1054) );
  OR2_X1 U4409 ( .A1(n18350), .A2(n18287), .ZN(n18354) );
  OR2_X1 U4410 ( .A1(n15457), .A2(n15050), .ZN(n15352) );
  MUX2_X1 U4411 ( .A(n15210), .B(n15209), .S(n3822), .Z(n15215) );
  NOR2_X1 U4412 ( .A1(n15559), .A2(n3822), .ZN(n15511) );
  OR2_X1 U4413 ( .A1(n3822), .A2(n15558), .ZN(n14964) );
  OR2_X1 U4414 ( .A1(n14236), .A2(n14148), .ZN(n14150) );
  INV_X1 U4415 ( .A(n11253), .ZN(n10803) );
  NAND2_X1 U4416 ( .A1(n3405), .A2(n10716), .ZN(n3404) );
  OR2_X1 U4417 ( .A1(n12003), .A2(n12001), .ZN(n3240) );
  OR2_X1 U4418 ( .A1(n3537), .A2(n12001), .ZN(n2184) );
  OR2_X1 U4419 ( .A1(n14150), .A2(n14239), .ZN(n14008) );
  OR2_X1 U4420 ( .A1(n14240), .A2(n14239), .ZN(n14241) );
  NOR2_X1 U4421 ( .A1(n9241), .A2(n9240), .ZN(n1777) );
  AND2_X1 U4422 ( .A1(n9189), .A2(n9240), .ZN(n2444) );
  AND2_X1 U4423 ( .A1(n9240), .A2(n8713), .ZN(n6656) );
  OR2_X1 U4424 ( .A1(n8569), .A2(n8568), .ZN(n3227) );
  OAI21_X1 U4425 ( .B1(n20490), .B2(n7466), .A(n3680), .ZN(n3679) );
  INV_X1 U4426 ( .A(n7797), .ZN(n8017) );
  OR2_X1 U4427 ( .A1(n5277), .A2(n5709), .ZN(n3467) );
  AOI21_X1 U4428 ( .B1(n5817), .B2(n5990), .A(n5815), .ZN(n3470) );
  AND2_X1 U4429 ( .A1(n12230), .A2(n12122), .ZN(n12235) );
  INV_X1 U4430 ( .A(n12230), .ZN(n12227) );
  AND2_X1 U4431 ( .A1(n15510), .A2(n14159), .ZN(n15210) );
  XNOR2_X1 U4432 ( .A(n9892), .B(n9893), .ZN(n3471) );
  INV_X1 U4433 ( .A(n3471), .ZN(n11474) );
  NOR2_X1 U4434 ( .A1(n11219), .A2(n3471), .ZN(n11217) );
  XNOR2_X1 U4435 ( .A(n19746), .B(n10425), .ZN(n10340) );
  INV_X1 U4436 ( .A(n18697), .ZN(n1055) );
  XNOR2_X1 U4437 ( .A(n13624), .B(n641), .ZN(n10793) );
  AND3_X1 U4438 ( .A1(n8207), .A2(n8206), .A3(n2885), .ZN(n1056) );
  BUF_X1 U4439 ( .A(n10154), .Z(n1057) );
  OR2_X1 U4440 ( .A1(n8208), .A2(n2886), .ZN(n2885) );
  OAI211_X1 U4441 ( .C1(n9118), .C2(n9218), .A(n9117), .B(n9116), .ZN(n10154)
         );
  NOR2_X1 U4442 ( .A1(n12609), .A2(n12601), .ZN(n12607) );
  AOI21_X1 U4444 ( .B1(n3898), .B2(n4005), .A(n2490), .ZN(n3901) );
  OAI21_X1 U4445 ( .B1(n1363), .B2(n1072), .A(n1071), .ZN(n1070) );
  AND2_X1 U4446 ( .A1(n11232), .A2(n10677), .ZN(n1600) );
  XNOR2_X1 U4447 ( .A(n10596), .B(n7663), .ZN(n2202) );
  NAND2_X1 U4448 ( .A1(n7427), .A2(n1791), .ZN(n1058) );
  NAND2_X1 U4449 ( .A1(n7426), .A2(n8232), .ZN(n1059) );
  NAND2_X1 U4450 ( .A1(n1058), .A2(n1059), .ZN(n7429) );
  AND2_X1 U4451 ( .A1(n20168), .A2(n19814), .ZN(n1060) );
  INV_X1 U4454 ( .A(n5022), .ZN(n4269) );
  INV_X1 U4455 ( .A(n14833), .ZN(n2779) );
  OR2_X1 U4457 ( .A1(n12100), .A2(n11381), .ZN(n3325) );
  XNOR2_X1 U4458 ( .A(n6455), .B(n6454), .ZN(n8076) );
  INV_X1 U4459 ( .A(n14648), .ZN(n3246) );
  AND2_X1 U4460 ( .A1(n20181), .A2(n14249), .ZN(n3685) );
  NOR2_X1 U4461 ( .A1(n1960), .A2(n9106), .ZN(n9104) );
  OR2_X1 U4462 ( .A1(n4899), .A2(n4963), .ZN(n3232) );
  OR2_X1 U4463 ( .A1(n18559), .A2(n18556), .ZN(n2960) );
  AND2_X1 U4464 ( .A1(n9147), .A2(n8790), .ZN(n8683) );
  OAI211_X1 U4465 ( .C1(n5704), .C2(n19562), .A(n5999), .B(n2051), .ZN(n5436)
         );
  NOR2_X1 U4466 ( .A1(n19756), .A2(n12240), .ZN(n12241) );
  NOR2_X1 U4467 ( .A1(n20445), .A2(n18592), .ZN(n18573) );
  AND2_X1 U4468 ( .A1(n12524), .A2(n11464), .ZN(n11768) );
  OAI21_X1 U4470 ( .B1(n14597), .B2(n14598), .A(n2926), .ZN(n3758) );
  INV_X1 U4471 ( .A(n14396), .ZN(n1527) );
  AND2_X1 U4472 ( .A1(n14154), .A2(n14396), .ZN(n13994) );
  INV_X1 U4473 ( .A(n11176), .ZN(n11173) );
  OR2_X1 U4474 ( .A1(n10657), .A2(n11176), .ZN(n2231) );
  OR2_X1 U4475 ( .A1(n11466), .A2(n11568), .ZN(n10885) );
  XNOR2_X1 U4476 ( .A(n9414), .B(n9854), .ZN(n10321) );
  NOR2_X1 U4478 ( .A1(n15459), .A2(n15350), .ZN(n14860) );
  AND2_X1 U4479 ( .A1(n190), .A2(n11321), .ZN(n1123) );
  OR2_X1 U4480 ( .A1(n11253), .A2(n19886), .ZN(n10310) );
  XNOR2_X1 U4481 ( .A(n17377), .B(n3209), .ZN(n17263) );
  XNOR2_X1 U4482 ( .A(n17377), .B(n3102), .ZN(n16296) );
  OR2_X1 U4484 ( .A1(n2984), .A2(n9304), .ZN(n3788) );
  XNOR2_X1 U4485 ( .A(n9799), .B(n9462), .ZN(n10481) );
  AND2_X1 U4486 ( .A1(n14662), .A2(n14663), .ZN(n2937) );
  INV_X1 U4487 ( .A(n14663), .ZN(n1552) );
  NAND2_X1 U4488 ( .A1(n20263), .A2(n14483), .ZN(n1062) );
  XOR2_X1 U4489 ( .A(n6252), .B(n6251), .Z(n1063) );
  XNOR2_X1 U4490 ( .A(n3744), .B(n13709), .ZN(n3743) );
  XNOR2_X1 U4491 ( .A(n13708), .B(n13704), .ZN(n3742) );
  XNOR2_X1 U4492 ( .A(n12861), .B(n13020), .ZN(n13708) );
  OR2_X1 U4493 ( .A1(n11553), .A2(n9017), .ZN(n10916) );
  INV_X1 U4494 ( .A(n20360), .ZN(n1452) );
  OR2_X1 U4495 ( .A1(n7519), .A2(n20359), .ZN(n3089) );
  AND2_X1 U4496 ( .A1(n9296), .A2(n9295), .ZN(n8520) );
  INV_X1 U4497 ( .A(n9296), .ZN(n3418) );
  NOR2_X1 U4499 ( .A1(n17223), .A2(n3573), .ZN(n16170) );
  AND2_X1 U4500 ( .A1(n18233), .A2(n20179), .ZN(n18120) );
  NOR2_X1 U4501 ( .A1(n17545), .A2(n18233), .ZN(n17973) );
  AND2_X1 U4502 ( .A1(n18233), .A2(n18226), .ZN(n2836) );
  INV_X1 U4503 ( .A(n19496), .ZN(n2697) );
  AND2_X1 U4504 ( .A1(n11292), .A2(n20235), .ZN(n3587) );
  INV_X1 U4505 ( .A(n11292), .ZN(n10978) );
  OR2_X1 U4506 ( .A1(n8325), .A2(n19856), .ZN(n7584) );
  INV_X1 U4507 ( .A(n3440), .ZN(n3497) );
  NOR2_X1 U4508 ( .A1(n244), .A2(n13147), .ZN(n13149) );
  OR2_X1 U4509 ( .A1(n7627), .A2(n20198), .ZN(n6212) );
  AND2_X1 U4510 ( .A1(n20198), .A2(n8192), .ZN(n7878) );
  INV_X1 U4511 ( .A(n12095), .ZN(n1091) );
  INV_X1 U4512 ( .A(n18311), .ZN(n19324) );
  INV_X1 U4513 ( .A(n14269), .ZN(n14574) );
  INV_X1 U4514 ( .A(n15167), .ZN(n15378) );
  AND2_X1 U4515 ( .A1(n13930), .A2(n12879), .ZN(n14334) );
  BUF_X1 U4516 ( .A(n13930), .Z(n14338) );
  XNOR2_X1 U4517 ( .A(n13341), .B(n13342), .ZN(n14692) );
  OR2_X1 U4519 ( .A1(n15162), .A2(n15501), .ZN(n2293) );
  OR2_X1 U4520 ( .A1(n14434), .A2(n14487), .ZN(n14433) );
  XNOR2_X1 U4521 ( .A(n13517), .B(n2296), .ZN(n2834) );
  OR2_X1 U4522 ( .A1(n5405), .A2(n5408), .ZN(n5146) );
  OAI211_X1 U4525 ( .C1(n12502), .C2(n12004), .A(n12500), .B(n12499), .ZN(
        n12006) );
  OR2_X1 U4527 ( .A1(n8981), .A2(n9267), .ZN(n3797) );
  INV_X1 U4529 ( .A(n17489), .ZN(n3347) );
  OR2_X1 U4530 ( .A1(n14529), .A2(n15018), .ZN(n15281) );
  OR2_X1 U4531 ( .A1(n5562), .A2(n6036), .ZN(n5534) );
  INV_X1 U4532 ( .A(n12284), .ZN(n13085) );
  AND2_X1 U4534 ( .A1(n10829), .A2(n11133), .ZN(n1165) );
  OR2_X1 U4535 ( .A1(n8958), .A2(n8960), .ZN(n1477) );
  AND2_X1 U4536 ( .A1(n4816), .A2(n5073), .ZN(n2022) );
  INV_X1 U4537 ( .A(n5073), .ZN(n2287) );
  OR2_X1 U4539 ( .A1(n15226), .A2(n15454), .ZN(n1987) );
  OAI22_X1 U4540 ( .A1(n19196), .A2(n19182), .B1(n19209), .B2(n19208), .ZN(
        n19212) );
  INV_X1 U4541 ( .A(n14450), .ZN(n1363) );
  AND2_X1 U4542 ( .A1(n19986), .A2(n19859), .ZN(n2316) );
  AOI21_X1 U4543 ( .B1(n13928), .B2(n3025), .A(n14448), .ZN(n14756) );
  AOI21_X1 U4544 ( .B1(n12407), .B2(n12408), .A(n12754), .ZN(n3012) );
  MUX2_X1 U4545 ( .A(n11595), .B(n12755), .S(n12754), .Z(n11596) );
  AND2_X1 U4546 ( .A1(n12754), .A2(n12407), .ZN(n1234) );
  NAND2_X1 U4547 ( .A1(n1064), .A2(n5200), .ZN(n3097) );
  OAI21_X1 U4548 ( .B1(n6089), .B2(n5176), .A(n4874), .ZN(n1064) );
  NAND2_X1 U4549 ( .A1(n1064), .A2(n5495), .ZN(n4875) );
  AOI21_X1 U4550 ( .B1(n269), .B2(n1065), .A(n9082), .ZN(n9083) );
  NAND2_X1 U4551 ( .A1(n3227), .A2(n1065), .ZN(n8403) );
  NAND2_X1 U4552 ( .A1(n8569), .A2(n9168), .ZN(n1065) );
  NOR2_X1 U4553 ( .A1(n273), .A2(n1560), .ZN(n7995) );
  AND2_X1 U4554 ( .A1(n19001), .A2(n19013), .ZN(n19023) );
  NAND3_X1 U4555 ( .A1(n1068), .A2(n18929), .A3(n2120), .ZN(n1066) );
  NAND2_X1 U4556 ( .A1(n18928), .A2(n17749), .ZN(n1067) );
  NAND2_X1 U4557 ( .A1(n20009), .A2(n20146), .ZN(n8278) );
  NAND2_X1 U4558 ( .A1(n251), .A2(n12437), .ZN(n11943) );
  NAND2_X1 U4559 ( .A1(n20365), .A2(n18592), .ZN(n17627) );
  NAND2_X1 U4560 ( .A1(n17096), .A2(n18633), .ZN(n1069) );
  NAND2_X1 U4561 ( .A1(n14455), .A2(n14453), .ZN(n1072) );
  INV_X1 U4562 ( .A(n1070), .ZN(n1359) );
  NAND3_X1 U4563 ( .A1(n13927), .A2(n14453), .A3(n14448), .ZN(n1071) );
  XNOR2_X1 U4564 ( .A(n20208), .B(n6514), .ZN(n1073) );
  XNOR2_X1 U4565 ( .A(n6730), .B(n6515), .ZN(n1074) );
  NAND2_X1 U4567 ( .A1(n1078), .A2(n15336), .ZN(n1077) );
  NAND2_X1 U4568 ( .A1(n15339), .A2(n15469), .ZN(n15466) );
  INV_X1 U4570 ( .A(n15466), .ZN(n1078) );
  NAND3_X1 U4571 ( .A1(n14897), .A2(n19888), .A3(n15466), .ZN(n1079) );
  NAND2_X1 U4572 ( .A1(n1080), .A2(n18619), .ZN(n18628) );
  NOR2_X1 U4573 ( .A1(n1080), .A2(n18619), .ZN(n18180) );
  XNOR2_X1 U4574 ( .A(n1081), .B(n7143), .ZN(n6374) );
  XNOR2_X1 U4575 ( .A(n1081), .B(n6839), .ZN(n6891) );
  XNOR2_X1 U4576 ( .A(n6307), .B(n1081), .ZN(n6309) );
  NAND2_X1 U4577 ( .A1(n1083), .A2(n989), .ZN(n1082) );
  INV_X1 U4578 ( .A(n5177), .ZN(n1083) );
  NAND2_X1 U4579 ( .A1(n1086), .A2(n1084), .ZN(n9151) );
  NAND2_X1 U4580 ( .A1(n1085), .A2(n7921), .ZN(n1084) );
  MUX2_X1 U4581 ( .A(n7984), .B(n7981), .S(n6312), .Z(n1085) );
  NAND3_X1 U4582 ( .A1(n7920), .A2(n7768), .A3(n1087), .ZN(n1086) );
  NAND2_X1 U4583 ( .A1(n7919), .A2(n1726), .ZN(n1087) );
  NAND2_X1 U4584 ( .A1(n19812), .A2(n7978), .ZN(n7920) );
  INV_X1 U4585 ( .A(n1089), .ZN(n14304) );
  NAND2_X1 U4586 ( .A1(n14506), .A2(n1089), .ZN(n14502) );
  OAI21_X1 U4588 ( .B1(n14498), .B2(n14506), .A(n1089), .ZN(n13974) );
  NAND2_X1 U4589 ( .A1(n15020), .A2(n1090), .ZN(n14960) );
  INV_X1 U4590 ( .A(n1656), .ZN(n1090) );
  NAND2_X1 U4591 ( .A1(n1091), .A2(n12686), .ZN(n12428) );
  NOR2_X1 U4592 ( .A1(n3649), .A2(n1094), .ZN(n11944) );
  OAI21_X1 U4593 ( .B1(n2805), .B2(n1094), .A(n12428), .ZN(n12434) );
  OAI21_X1 U4594 ( .B1(n12687), .B2(n1094), .A(n1092), .ZN(n1550) );
  OAI211_X1 U4595 ( .C1(n12651), .C2(n1094), .A(n12650), .B(n1093), .ZN(n13543) );
  OAI21_X1 U4596 ( .B1(n12646), .B2(n12685), .A(n1094), .ZN(n1093) );
  INV_X1 U4597 ( .A(n12095), .ZN(n1094) );
  NAND2_X1 U4598 ( .A1(n5823), .A2(n6017), .ZN(n1096) );
  OAI21_X1 U4599 ( .B1(n1098), .B2(n12442), .A(n1097), .ZN(n11067) );
  NAND2_X1 U4600 ( .A1(n12442), .A2(n12443), .ZN(n1097) );
  NAND2_X1 U4601 ( .A1(n1099), .A2(n11942), .ZN(n1098) );
  INV_X1 U4602 ( .A(n1101), .ZN(n1100) );
  OAI22_X1 U4603 ( .A1(n15614), .A2(n15546), .B1(n15619), .B2(n15547), .ZN(
        n1101) );
  NAND2_X1 U4604 ( .A1(n15071), .A2(n15615), .ZN(n15614) );
  INV_X1 U4605 ( .A(n15615), .ZN(n15619) );
  NAND2_X1 U4606 ( .A1(n9071), .A2(n9346), .ZN(n1102) );
  NAND2_X1 U4607 ( .A1(n9072), .A2(n9339), .ZN(n1103) );
  OAI21_X2 U4608 ( .B1(n9243), .B2(n268), .A(n2636), .ZN(n9854) );
  NAND2_X1 U4609 ( .A1(n1486), .A2(n1104), .ZN(n2717) );
  NAND3_X1 U4610 ( .A1(n14125), .A2(n14126), .A3(n1104), .ZN(n14129) );
  OR2_X1 U4611 ( .A1(n19731), .A2(n14394), .ZN(n2201) );
  AOI21_X1 U4612 ( .B1(n1661), .B2(n214), .A(n1660), .ZN(n1659) );
  OAI21_X1 U4613 ( .B1(n15919), .B2(n15420), .A(n3709), .ZN(n14259) );
  NAND2_X1 U4614 ( .A1(n1105), .A2(n8303), .ZN(n1242) );
  NAND2_X1 U4615 ( .A1(n1247), .A2(n7876), .ZN(n1105) );
  NAND2_X1 U4616 ( .A1(n1108), .A2(n1107), .ZN(n1106) );
  INV_X1 U4617 ( .A(n3389), .ZN(n1107) );
  NAND2_X1 U4618 ( .A1(n3391), .A2(n3390), .ZN(n1108) );
  NAND2_X1 U4620 ( .A1(n1111), .A2(n1110), .ZN(n1109) );
  AOI21_X1 U4621 ( .B1(n17868), .B2(n17676), .A(n17078), .ZN(n1110) );
  NAND2_X1 U4622 ( .A1(n17074), .A2(n1112), .ZN(n1111) );
  NAND2_X1 U4623 ( .A1(n1114), .A2(n1113), .ZN(n16631) );
  NAND2_X1 U4624 ( .A1(n16627), .A2(n16465), .ZN(n1113) );
  NAND2_X1 U4625 ( .A1(n16628), .A2(n1115), .ZN(n1114) );
  NAND3_X1 U4626 ( .A1(n9498), .A2(n11670), .A3(n11845), .ZN(n1116) );
  NAND2_X1 U4627 ( .A1(n9543), .A2(n12185), .ZN(n1117) );
  XNOR2_X1 U4628 ( .A(n12286), .B(n12287), .ZN(n3440) );
  OAI21_X1 U4629 ( .B1(n17911), .B2(n17912), .A(n18501), .ZN(n1118) );
  AOI21_X2 U4630 ( .B1(n15924), .B2(n15923), .A(n1119), .ZN(n16224) );
  AND2_X1 U4631 ( .A1(n7548), .A2(n7547), .ZN(n2778) );
  INV_X1 U4632 ( .A(n14571), .ZN(n14267) );
  NAND2_X1 U4633 ( .A1(n12348), .A2(n1120), .ZN(n13778) );
  NAND2_X1 U4634 ( .A1(n1001), .A2(n12497), .ZN(n1120) );
  NOR2_X1 U4637 ( .A1(n1123), .A2(n11327), .ZN(n1122) );
  NAND2_X1 U4639 ( .A1(n11488), .A2(n12530), .ZN(n11520) );
  NAND2_X1 U4640 ( .A1(n11209), .A2(n11443), .ZN(n10469) );
  NAND2_X1 U4641 ( .A1(n4401), .A2(n4400), .ZN(n6153) );
  NAND2_X1 U4642 ( .A1(n14076), .A2(n14780), .ZN(n14217) );
  OR2_X1 U4645 ( .A1(n17812), .A2(n19846), .ZN(n18949) );
  NAND2_X1 U4647 ( .A1(n8571), .A2(n9062), .ZN(n8572) );
  INV_X1 U4648 ( .A(n5845), .ZN(n5847) );
  INV_X1 U4649 ( .A(n3507), .ZN(n3711) );
  AND2_X1 U4650 ( .A1(n1336), .A2(n920), .ZN(n1872) );
  OAI211_X1 U4651 ( .C1(n7227), .C2(n8313), .A(n7226), .B(n7225), .ZN(n8925)
         );
  INV_X1 U4652 ( .A(n9313), .ZN(n9053) );
  AOI21_X1 U4653 ( .B1(n3796), .B2(n20568), .A(n2525), .ZN(n2524) );
  INV_X1 U4654 ( .A(n8813), .ZN(n8810) );
  AND3_X1 U4655 ( .A1(n11094), .A2(n11443), .A3(n11445), .ZN(n2656) );
  INV_X1 U4656 ( .A(n15422), .ZN(n3710) );
  INV_X1 U4657 ( .A(n8602), .ZN(n8956) );
  INV_X1 U4659 ( .A(n15521), .ZN(n15593) );
  INV_X1 U4660 ( .A(n13041), .ZN(n12697) );
  INV_X1 U4661 ( .A(n17494), .ZN(n17488) );
  XNOR2_X1 U4662 ( .A(n6719), .B(n6761), .ZN(n7079) );
  XNOR2_X1 U4663 ( .A(n16980), .B(n17109), .ZN(n16892) );
  NOR2_X1 U4664 ( .A1(n10919), .A2(n10755), .ZN(n10923) );
  OR2_X1 U4666 ( .A1(n9272), .A2(n9275), .ZN(n9282) );
  XNOR2_X1 U4667 ( .A(n3162), .B(n20064), .ZN(n15087) );
  INV_X1 U4668 ( .A(n11769), .ZN(n11792) );
  NAND2_X1 U4669 ( .A1(n2271), .A2(n2270), .ZN(n11769) );
  NAND2_X1 U4670 ( .A1(n7694), .A2(n7911), .ZN(n1679) );
  INV_X1 U4671 ( .A(n1770), .ZN(n5624) );
  NAND2_X1 U4674 ( .A1(n3429), .A2(n1126), .ZN(n3428) );
  NAND2_X1 U4675 ( .A1(n3431), .A2(n3427), .ZN(n1126) );
  XNOR2_X2 U4678 ( .A(n12789), .B(n12790), .ZN(n14335) );
  NAND2_X1 U4679 ( .A1(n1127), .A2(n2485), .ZN(n2484) );
  NAND2_X1 U4680 ( .A1(n11116), .A2(n11440), .ZN(n1127) );
  NOR2_X1 U4681 ( .A1(n3617), .A2(n12549), .ZN(n3613) );
  NAND2_X1 U4682 ( .A1(n1761), .A2(n1128), .ZN(n1759) );
  NAND2_X1 U4684 ( .A1(n5860), .A2(n6140), .ZN(n5620) );
  OAI21_X2 U4685 ( .B1(n4456), .B2(n153), .A(n4455), .ZN(n6140) );
  NAND2_X1 U4686 ( .A1(n15237), .A2(n15350), .ZN(n15353) );
  OAI21_X2 U4687 ( .B1(n13881), .B2(n13555), .A(n13554), .ZN(n15350) );
  NAND3_X2 U4688 ( .A1(n1129), .A2(n2730), .A3(n14147), .ZN(n15558) );
  NAND2_X1 U4691 ( .A1(n12226), .A2(n12228), .ZN(n11692) );
  NAND2_X1 U4692 ( .A1(n10927), .A2(n10928), .ZN(n10931) );
  NOR2_X1 U4693 ( .A1(n11549), .A2(n11546), .ZN(n10928) );
  NOR2_X1 U4694 ( .A1(n11371), .A2(n11372), .ZN(n13099) );
  XNOR2_X1 U4695 ( .A(n17005), .B(n16873), .ZN(n2994) );
  NOR2_X1 U4697 ( .A1(n11834), .A2(n12359), .ZN(n11835) );
  NAND2_X1 U4699 ( .A1(n9831), .A2(n11343), .ZN(n1133) );
  NAND2_X1 U4700 ( .A1(n12631), .A2(n3401), .ZN(n12632) );
  AND2_X1 U4702 ( .A1(n5496), .A2(n5741), .ZN(n2525) );
  AND2_X1 U4703 ( .A1(n8017), .A2(n7965), .ZN(n7811) );
  XNOR2_X1 U4704 ( .A(n7293), .B(n7292), .ZN(n7786) );
  AND2_X1 U4705 ( .A1(n19434), .A2(n19433), .ZN(n2450) );
  INV_X1 U4706 ( .A(n4021), .ZN(n4131) );
  INV_X1 U4707 ( .A(n12523), .ZN(n12288) );
  INV_X1 U4708 ( .A(n8890), .ZN(n9005) );
  NAND2_X1 U4712 ( .A1(n9331), .A2(n9330), .ZN(n9076) );
  NAND2_X1 U4713 ( .A1(n2924), .A2(n14394), .ZN(n2923) );
  NAND2_X2 U4714 ( .A1(n3412), .A2(n1136), .ZN(n16128) );
  OR2_X1 U4715 ( .A1(n14111), .A2(n20498), .ZN(n1136) );
  NAND2_X1 U4716 ( .A1(n2022), .A2(n5072), .ZN(n1137) );
  NAND2_X1 U4718 ( .A1(n874), .A2(n12616), .ZN(n12243) );
  AOI22_X1 U4720 ( .A1(n13865), .A2(n3516), .B1(n701), .B2(n14442), .ZN(n3174)
         );
  NAND2_X1 U4721 ( .A1(n11734), .A2(n1139), .ZN(n11737) );
  NAND2_X1 U4723 ( .A1(n7492), .A2(n7491), .ZN(n10028) );
  NOR2_X1 U4724 ( .A1(n17998), .A2(n1141), .ZN(n18000) );
  OAI21_X1 U4725 ( .B1(n2960), .B2(n18568), .A(n2957), .ZN(n1141) );
  NAND2_X1 U4726 ( .A1(n6587), .A2(n9189), .ZN(n9188) );
  NAND3_X1 U4727 ( .A1(n1238), .A2(n1237), .A3(n1143), .ZN(n1142) );
  NAND2_X1 U4728 ( .A1(n7845), .A2(n8114), .ZN(n1144) );
  NAND2_X1 U4729 ( .A1(n13671), .A2(n14716), .ZN(n14245) );
  NAND2_X1 U4730 ( .A1(n19456), .A2(n1145), .ZN(n18014) );
  NAND2_X1 U4731 ( .A1(n16402), .A2(n16401), .ZN(n1146) );
  NAND2_X1 U4732 ( .A1(n16403), .A2(n16404), .ZN(n1147) );
  XNOR2_X1 U4735 ( .A(n10370), .B(n2900), .ZN(n2046) );
  NAND2_X1 U4738 ( .A1(n4848), .A2(n3996), .ZN(n4849) );
  INV_X1 U4739 ( .A(n9616), .ZN(n3515) );
  NAND2_X1 U4740 ( .A1(n1858), .A2(n1861), .ZN(n1149) );
  NAND2_X1 U4743 ( .A1(n4899), .A2(n4962), .ZN(n3974) );
  OR2_X1 U4744 ( .A1(n9106), .A2(n9105), .ZN(n8780) );
  OAI211_X1 U4746 ( .C1(n19517), .C2(n8998), .A(n8657), .B(n3554), .ZN(n3553)
         );
  OAI22_X1 U4747 ( .A1(n15138), .A2(n15386), .B1(n15696), .B2(n15702), .ZN(
        n15039) );
  NAND2_X1 U4751 ( .A1(n5471), .A2(n6036), .ZN(n5472) );
  NAND2_X1 U4752 ( .A1(n5562), .A2(n5569), .ZN(n5471) );
  XNOR2_X1 U4753 ( .A(n13588), .B(n12770), .ZN(n13490) );
  OR2_X1 U4754 ( .A1(n17219), .A2(n19386), .ZN(n3391) );
  XNOR2_X1 U4755 ( .A(n16225), .B(n16134), .ZN(n17119) );
  XNOR2_X1 U4756 ( .A(n1153), .B(n13750), .ZN(n13751) );
  XNOR2_X1 U4757 ( .A(n13748), .B(n13749), .ZN(n1153) );
  NAND2_X1 U4758 ( .A1(n1155), .A2(n15049), .ZN(n1154) );
  NAND2_X1 U4759 ( .A1(n9190), .A2(n2443), .ZN(n9700) );
  OAI21_X1 U4761 ( .B1(n4131), .B2(n4293), .A(n1156), .ZN(n4135) );
  NAND2_X1 U4762 ( .A1(n4131), .A2(n4298), .ZN(n1156) );
  NOR2_X1 U4763 ( .A1(n11359), .A2(n20099), .ZN(n3667) );
  NAND2_X1 U4764 ( .A1(n19979), .A2(n5920), .ZN(n6011) );
  NAND2_X1 U4766 ( .A1(n1239), .A2(n4840), .ZN(n4839) );
  NAND2_X1 U4767 ( .A1(n11509), .A2(n20106), .ZN(n10007) );
  INV_X1 U4769 ( .A(n1159), .ZN(n1158) );
  NAND2_X1 U4771 ( .A1(n7859), .A2(n8232), .ZN(n1160) );
  OAI21_X1 U4772 ( .B1(n12376), .B2(n19504), .A(n12375), .ZN(n2332) );
  NAND3_X1 U4773 ( .A1(n5493), .A2(n5900), .A3(n6089), .ZN(n2098) );
  OAI21_X1 U4774 ( .B1(n1162), .B2(n1161), .A(n20417), .ZN(n17586) );
  NOR2_X1 U4775 ( .A1(n19661), .A2(n19655), .ZN(n1161) );
  INV_X1 U4776 ( .A(n18532), .ZN(n1162) );
  NAND3_X1 U4778 ( .A1(n8362), .A2(n8361), .A3(n8360), .ZN(n2934) );
  NAND3_X1 U4779 ( .A1(n14379), .A2(n2767), .A3(n20204), .ZN(n2766) );
  NAND2_X1 U4780 ( .A1(n14230), .A2(n14229), .ZN(n14379) );
  AOI22_X2 U4781 ( .A1(n15776), .A2(n15775), .B1(n15773), .B2(n15774), .ZN(
        n16939) );
  INV_X1 U4783 ( .A(n12208), .ZN(n12210) );
  AOI22_X1 U4784 ( .A1(n10799), .A2(n11348), .B1(n10800), .B2(n11346), .ZN(
        n1592) );
  OR2_X1 U4785 ( .A1(n14228), .A2(n14229), .ZN(n2304) );
  INV_X1 U4788 ( .A(n2627), .ZN(n1164) );
  NAND2_X1 U4789 ( .A1(n1680), .A2(n1165), .ZN(n11134) );
  NAND2_X1 U4790 ( .A1(n1167), .A2(n1166), .ZN(n16728) );
  NAND2_X1 U4791 ( .A1(n17677), .A2(n17074), .ZN(n1167) );
  INV_X1 U4793 ( .A(n14451), .ZN(n14180) );
  NOR2_X1 U4794 ( .A1(n10639), .A2(n10932), .ZN(n10737) );
  INV_X1 U4795 ( .A(n17214), .ZN(n1173) );
  NAND2_X1 U4796 ( .A1(n16466), .A2(n1395), .ZN(n16662) );
  NOR2_X1 U4797 ( .A1(n18496), .A2(n1174), .ZN(n18499) );
  XNOR2_X1 U4798 ( .A(n17443), .B(n16293), .ZN(n14895) );
  OAI22_X2 U4799 ( .A1(n14888), .A2(n14889), .B1(n15311), .B2(n14887), .ZN(
        n17443) );
  AOI21_X1 U4802 ( .B1(n9776), .B2(n10862), .A(n11302), .ZN(n1175) );
  NOR2_X1 U4803 ( .A1(n996), .A2(n1362), .ZN(n14459) );
  NAND2_X1 U4804 ( .A1(n5085), .A2(n1596), .ZN(n1360) );
  NAND2_X1 U4805 ( .A1(n19980), .A2(n5917), .ZN(n5588) );
  NOR2_X1 U4806 ( .A1(n1176), .A2(n15336), .ZN(n12874) );
  AND2_X1 U4807 ( .A1(n12841), .A2(n12840), .ZN(n1176) );
  NAND2_X1 U4808 ( .A1(n7992), .A2(n8010), .ZN(n7993) );
  NAND2_X1 U4811 ( .A1(n1179), .A2(n1178), .ZN(n14528) );
  NAND3_X1 U4812 ( .A1(n14648), .A2(n14525), .A3(n14522), .ZN(n1178) );
  NAND2_X1 U4813 ( .A1(n14523), .A2(n19831), .ZN(n1179) );
  NAND2_X1 U4815 ( .A1(n15714), .A2(n15871), .ZN(n1181) );
  NAND2_X1 U4817 ( .A1(n14192), .A2(n14620), .ZN(n1265) );
  OR2_X1 U4818 ( .A1(n15813), .A2(n15581), .ZN(n15816) );
  NAND3_X1 U4820 ( .A1(n5316), .A2(n5572), .A3(n5583), .ZN(n1182) );
  NAND2_X1 U4821 ( .A1(n5605), .A2(n5714), .ZN(n5243) );
  AOI21_X1 U4822 ( .B1(n15782), .B2(n15783), .A(n15686), .ZN(n1183) );
  NOR2_X1 U4823 ( .A1(n13912), .A2(n1184), .ZN(n13917) );
  AND2_X1 U4824 ( .A1(n15171), .A2(n15327), .ZN(n1184) );
  INV_X1 U4826 ( .A(n12059), .ZN(n2053) );
  XNOR2_X1 U4827 ( .A(n961), .B(n1185), .ZN(n1524) );
  INV_X1 U4828 ( .A(n8509), .ZN(n1185) );
  XNOR2_X1 U4832 ( .A(n1187), .B(n15225), .ZN(n15250) );
  XNOR2_X1 U4833 ( .A(n16887), .B(n16926), .ZN(n1187) );
  NAND3_X1 U4835 ( .A1(n1188), .A2(n15416), .A3(n15007), .ZN(n14372) );
  NAND2_X1 U4836 ( .A1(n15078), .A2(n15907), .ZN(n1188) );
  NOR2_X2 U4837 ( .A1(n3720), .A2(n11621), .ZN(n13776) );
  OAI21_X1 U4838 ( .B1(n8438), .B2(n9149), .A(n1736), .ZN(n1738) );
  OAI21_X1 U4839 ( .B1(n11160), .B2(n11159), .A(n11161), .ZN(n1903) );
  NAND2_X1 U4840 ( .A1(n15443), .A2(n15442), .ZN(n15312) );
  NAND3_X1 U4841 ( .A1(n10801), .A2(n11060), .A3(n11057), .ZN(n1189) );
  OR3_X1 U4842 ( .A1(n19776), .A2(n5086), .A3(n20202), .ZN(n4031) );
  NAND3_X1 U4843 ( .A1(n17155), .A2(n19675), .A3(n17489), .ZN(n2693) );
  AOI21_X1 U4844 ( .B1(n12205), .B2(n12589), .A(n1190), .ZN(n12977) );
  AND2_X2 U4845 ( .A1(n13862), .A2(n13863), .ZN(n17288) );
  NOR2_X1 U4846 ( .A1(n19509), .A2(n18600), .ZN(n1195) );
  OAI21_X1 U4847 ( .B1(n19509), .B2(n1192), .A(n1193), .ZN(n18219) );
  NAND2_X1 U4848 ( .A1(n3693), .A2(n18215), .ZN(n1192) );
  NAND2_X1 U4849 ( .A1(n1195), .A2(n18625), .ZN(n17576) );
  INV_X1 U4851 ( .A(n18215), .ZN(n1194) );
  NAND2_X1 U4852 ( .A1(n1196), .A2(n9006), .ZN(n8767) );
  NAND2_X1 U4853 ( .A1(n8890), .A2(n8895), .ZN(n1196) );
  MUX2_X1 U4854 ( .A(n6182), .B(n6181), .S(n2865), .Z(n6188) );
  MUX2_X2 U4855 ( .A(n6382), .B(n6383), .S(n6184), .Z(n7355) );
  NAND2_X1 U4856 ( .A1(n1198), .A2(n8372), .ZN(n3490) );
  NAND2_X1 U4857 ( .A1(n6733), .A2(n1199), .ZN(n1198) );
  OR2_X1 U4858 ( .A1(n6734), .A2(n8370), .ZN(n1199) );
  NAND3_X1 U4859 ( .A1(n20003), .A2(n15529), .A3(n18423), .ZN(n16490) );
  INV_X1 U4862 ( .A(n1201), .ZN(n9352) );
  INV_X1 U4863 ( .A(n9359), .ZN(n9356) );
  NAND2_X1 U4865 ( .A1(n9355), .A2(n1201), .ZN(n1200) );
  OAI21_X1 U4866 ( .B1(n1204), .B2(n9359), .A(n1203), .ZN(n1202) );
  NAND2_X1 U4867 ( .A1(n9358), .A2(n9359), .ZN(n1203) );
  NAND2_X1 U4868 ( .A1(n20447), .A2(n19269), .ZN(n2533) );
  INV_X1 U4869 ( .A(n1206), .ZN(n3558) );
  NAND2_X1 U4870 ( .A1(n11513), .A2(n11510), .ZN(n1206) );
  NAND2_X1 U4871 ( .A1(n11575), .A2(n1206), .ZN(n11512) );
  NAND2_X1 U4872 ( .A1(n20424), .A2(n14542), .ZN(n1208) );
  NAND2_X1 U4873 ( .A1(n13982), .A2(n14542), .ZN(n1209) );
  NAND2_X1 U4874 ( .A1(n1918), .A2(n1210), .ZN(n1917) );
  AOI21_X1 U4875 ( .B1(n11397), .B2(n11297), .A(n11399), .ZN(n1210) );
  NAND2_X1 U4876 ( .A1(n269), .A2(n8569), .ZN(n1211) );
  AND2_X1 U4877 ( .A1(n1212), .A2(n11990), .ZN(n12340) );
  INV_X1 U4878 ( .A(n12334), .ZN(n1212) );
  NOR2_X1 U4880 ( .A1(n12337), .A2(n1213), .ZN(n10315) );
  NAND2_X1 U4881 ( .A1(n5309), .A2(n1214), .ZN(n2466) );
  NOR2_X1 U4882 ( .A1(n5144), .A2(n1214), .ZN(n4052) );
  INV_X1 U4884 ( .A(n1215), .ZN(n14587) );
  NAND2_X1 U4885 ( .A1(n14811), .A2(n14593), .ZN(n1215) );
  NAND2_X1 U4886 ( .A1(n1215), .A2(n14812), .ZN(n11791) );
  NAND2_X1 U4887 ( .A1(n15271), .A2(n15274), .ZN(n1218) );
  NAND3_X1 U4888 ( .A1(n15604), .A2(n1221), .A3(n1216), .ZN(n1219) );
  NAND2_X1 U4889 ( .A1(n15271), .A2(n15601), .ZN(n1216) );
  NAND2_X1 U4891 ( .A1(n14986), .A2(n15274), .ZN(n1220) );
  NAND2_X1 U4892 ( .A1(n1217), .A2(n1220), .ZN(n14987) );
  NAND2_X1 U4893 ( .A1(n1218), .A2(n1219), .ZN(n1217) );
  NAND2_X1 U4894 ( .A1(n15270), .A2(n15600), .ZN(n1221) );
  NAND2_X1 U4895 ( .A1(n15275), .A2(n15276), .ZN(n15604) );
  NAND2_X1 U4896 ( .A1(n15035), .A2(n15034), .ZN(n1223) );
  NAND2_X1 U4897 ( .A1(n11843), .A2(n20201), .ZN(n1224) );
  NOR2_X1 U4899 ( .A1(n14620), .A2(n954), .ZN(n15315) );
  INV_X1 U4900 ( .A(n14619), .ZN(n15314) );
  NAND2_X1 U4901 ( .A1(n13858), .A2(n1226), .ZN(n15676) );
  XNOR2_X1 U4902 ( .A(n10563), .B(n1227), .ZN(n9526) );
  NAND2_X1 U4903 ( .A1(n12083), .A2(n1229), .ZN(n12085) );
  NAND2_X1 U4904 ( .A1(n12415), .A2(n12417), .ZN(n1229) );
  NAND2_X1 U4905 ( .A1(n10637), .A2(n20279), .ZN(n12415) );
  NAND2_X1 U4906 ( .A1(n1230), .A2(n9158), .ZN(n2782) );
  NAND2_X1 U4907 ( .A1(n8247), .A2(n8253), .ZN(n7562) );
  XNOR2_X2 U4908 ( .A(n6481), .B(n6482), .ZN(n8253) );
  NAND2_X1 U4909 ( .A1(n291), .A2(n4410), .ZN(n1232) );
  NAND2_X1 U4910 ( .A1(n8334), .A2(n3645), .ZN(n2301) );
  INV_X1 U4911 ( .A(n9123), .ZN(n1233) );
  NAND2_X1 U4912 ( .A1(n245), .A2(n1234), .ZN(n3702) );
  NAND2_X1 U4913 ( .A1(n12756), .A2(n12759), .ZN(n1235) );
  NAND2_X1 U4915 ( .A1(n8113), .A2(n8253), .ZN(n1237) );
  NAND2_X1 U4916 ( .A1(n6704), .A2(n3312), .ZN(n1238) );
  INV_X1 U4917 ( .A(n4656), .ZN(n1239) );
  NAND2_X1 U4918 ( .A1(n4841), .A2(n1239), .ZN(n4221) );
  NAND2_X1 U4919 ( .A1(n19859), .A2(n985), .ZN(n14831) );
  XNOR2_X1 U4920 ( .A(n12750), .B(n12749), .ZN(n2684) );
  NAND3_X1 U4921 ( .A1(n1241), .A2(n1688), .A3(n246), .ZN(n1240) );
  NAND2_X1 U4922 ( .A1(n10716), .A2(n12629), .ZN(n1241) );
  NAND2_X1 U4923 ( .A1(n8991), .A2(n8990), .ZN(n8650) );
  NAND2_X1 U4924 ( .A1(n1245), .A2(n20001), .ZN(n1243) );
  NAND2_X1 U4925 ( .A1(n8044), .A2(n8304), .ZN(n1245) );
  INV_X1 U4926 ( .A(n8304), .ZN(n8045) );
  NAND2_X1 U4927 ( .A1(n8304), .A2(n8305), .ZN(n1247) );
  NAND2_X1 U4929 ( .A1(n1250), .A2(n1252), .ZN(n1249) );
  NAND2_X1 U4930 ( .A1(n12060), .A2(n11979), .ZN(n1250) );
  INV_X1 U4931 ( .A(n4152), .ZN(n4354) );
  NAND3_X1 U4932 ( .A1(n4547), .A2(n4546), .A3(n4603), .ZN(n1253) );
  NAND2_X1 U4933 ( .A1(n2781), .A2(n9165), .ZN(n1254) );
  NOR2_X1 U4934 ( .A1(n9157), .A2(n1256), .ZN(n1255) );
  NAND2_X1 U4935 ( .A1(n9159), .A2(n9158), .ZN(n1256) );
  NAND2_X1 U4936 ( .A1(n11652), .A2(n11651), .ZN(n1258) );
  XNOR2_X1 U4937 ( .A(n13790), .B(n1259), .ZN(n12786) );
  XNOR2_X1 U4938 ( .A(n1260), .B(n13677), .ZN(n12014) );
  XNOR2_X1 U4939 ( .A(n13734), .B(n1260), .ZN(n13486) );
  NAND2_X1 U4940 ( .A1(n14251), .A2(n1261), .ZN(n14254) );
  OAI211_X2 U4943 ( .C1(n1264), .C2(n3329), .A(n2681), .B(n1263), .ZN(n15702)
         );
  NAND3_X1 U4944 ( .A1(n1264), .A2(n20181), .A3(n19918), .ZN(n1263) );
  NOR2_X1 U4947 ( .A1(n7653), .A2(n8960), .ZN(n1267) );
  NAND2_X1 U4950 ( .A1(n2071), .A2(n4845), .ZN(n1270) );
  OAI21_X1 U4951 ( .B1(n4845), .B2(n4421), .A(n1270), .ZN(n4422) );
  OR2_X1 U4952 ( .A1(n1270), .A2(n4844), .ZN(n5903) );
  NAND2_X1 U4953 ( .A1(n1271), .A2(n3775), .ZN(n2190) );
  NAND2_X1 U4954 ( .A1(n1271), .A2(n1502), .ZN(n1500) );
  NAND2_X1 U4955 ( .A1(n1803), .A2(n1272), .ZN(n4620) );
  OAI21_X1 U4956 ( .B1(n4006), .B2(n4003), .A(n1272), .ZN(n4007) );
  NAND3_X1 U4957 ( .A1(n4308), .A2(n4307), .A3(n1272), .ZN(n4309) );
  NAND2_X1 U4958 ( .A1(n4302), .A2(n4306), .ZN(n1272) );
  AND2_X2 U4959 ( .A1(n12465), .A2(n991), .ZN(n12138) );
  NAND2_X1 U4960 ( .A1(n1273), .A2(n8046), .ZN(n8050) );
  NAND3_X1 U4961 ( .A1(n1273), .A2(n8046), .A3(n2597), .ZN(n2635) );
  NAND2_X1 U4962 ( .A1(n20001), .A2(n8303), .ZN(n1273) );
  NOR2_X1 U4963 ( .A1(n6105), .A2(n6109), .ZN(n1275) );
  NOR2_X1 U4964 ( .A1(n5957), .A2(n6105), .ZN(n6111) );
  NAND2_X1 U4965 ( .A1(n5172), .A2(n1275), .ZN(n1274) );
  NAND2_X1 U4966 ( .A1(n1276), .A2(n6155), .ZN(n1347) );
  NAND2_X1 U4967 ( .A1(n6153), .A2(n1277), .ZN(n1276) );
  INV_X1 U4968 ( .A(n5349), .ZN(n1277) );
  OAI21_X2 U4969 ( .B1(n2585), .B2(n4380), .A(n2584), .ZN(n5349) );
  NAND3_X1 U4970 ( .A1(n12104), .A2(n11383), .A3(n20468), .ZN(n1278) );
  NAND2_X1 U4971 ( .A1(n10864), .A2(n11271), .ZN(n1279) );
  NAND2_X1 U4972 ( .A1(n1281), .A2(n10796), .ZN(n11810) );
  INV_X1 U4973 ( .A(n9832), .ZN(n1281) );
  INV_X1 U4974 ( .A(n10797), .ZN(n1282) );
  NAND2_X1 U4975 ( .A1(n15841), .A2(n1286), .ZN(n15264) );
  MUX2_X1 U4976 ( .A(n15625), .B(n15100), .S(n1288), .Z(n14417) );
  NAND2_X1 U4977 ( .A1(n2471), .A2(n1286), .ZN(n15631) );
  NAND2_X1 U4978 ( .A1(n1289), .A2(n1288), .ZN(n1287) );
  NAND2_X1 U4979 ( .A1(n15841), .A2(n1290), .ZN(n1289) );
  NAND2_X1 U4980 ( .A1(n15839), .A2(n15840), .ZN(n1290) );
  NAND2_X1 U4981 ( .A1(n15839), .A2(n15625), .ZN(n15841) );
  NAND2_X1 U4982 ( .A1(n15837), .A2(n15836), .ZN(n1291) );
  NAND2_X1 U4984 ( .A1(n3642), .A2(n14264), .ZN(n1292) );
  MUX2_X1 U4986 ( .A(n15538), .B(n15400), .S(n15898), .Z(n1293) );
  NAND2_X1 U4987 ( .A1(n14263), .A2(n14262), .ZN(n1294) );
  NAND3_X1 U4988 ( .A1(n1295), .A2(n14811), .A3(n14807), .ZN(n14140) );
  NAND2_X1 U4989 ( .A1(n1296), .A2(n18383), .ZN(n18387) );
  OAI21_X1 U4990 ( .B1(n1296), .B2(n18369), .A(n18392), .ZN(n18373) );
  NAND2_X2 U4992 ( .A1(n1297), .A2(n1301), .ZN(n13335) );
  NAND2_X1 U4993 ( .A1(n1298), .A2(n11167), .ZN(n1297) );
  NAND2_X1 U4994 ( .A1(n12282), .A2(n12042), .ZN(n1300) );
  NAND2_X1 U4995 ( .A1(n1302), .A2(n12041), .ZN(n1301) );
  OR2_X2 U4996 ( .A1(n3017), .A2(n3016), .ZN(n12041) );
  NAND2_X1 U4997 ( .A1(n12278), .A2(n12282), .ZN(n1302) );
  MUX2_X1 U4999 ( .A(n17391), .B(n17392), .S(n3066), .Z(n17393) );
  AOI22_X1 U5000 ( .A1(n12514), .A2(n12513), .B1(n11995), .B2(n13275), .ZN(
        n1305) );
  NAND2_X1 U5001 ( .A1(n10365), .A2(n11110), .ZN(n1306) );
  NAND2_X1 U5002 ( .A1(n7912), .A2(n7910), .ZN(n1308) );
  NAND2_X1 U5003 ( .A1(n18772), .A2(n19803), .ZN(n18713) );
  NAND3_X1 U5004 ( .A1(n18277), .A2(n18276), .A3(n1309), .ZN(n1310) );
  NAND3_X1 U5005 ( .A1(n18772), .A2(n19803), .A3(n18781), .ZN(n1309) );
  XNOR2_X1 U5006 ( .A(n1310), .B(n18279), .ZN(Ciphertext[82]) );
  NAND2_X1 U5007 ( .A1(n10980), .A2(n11290), .ZN(n1311) );
  AOI21_X1 U5008 ( .B1(n11292), .B2(n19506), .A(n3588), .ZN(n1312) );
  NAND3_X1 U5009 ( .A1(n10813), .A2(n19949), .A3(n1039), .ZN(n1314) );
  XNOR2_X1 U5010 ( .A(n10084), .B(n10083), .ZN(n10785) );
  OAI21_X1 U5011 ( .B1(n1039), .B2(n1317), .A(n1316), .ZN(n1315) );
  AOI21_X1 U5012 ( .B1(n19725), .B2(n1039), .A(n10813), .ZN(n1316) );
  OR2_X1 U5013 ( .A1(n11038), .A2(n19949), .ZN(n1318) );
  NAND2_X1 U5014 ( .A1(n10112), .A2(n11360), .ZN(n11038) );
  NAND2_X1 U5015 ( .A1(n1441), .A2(n1319), .ZN(n5311) );
  AND2_X1 U5016 ( .A1(n1320), .A2(n2468), .ZN(n1319) );
  NAND3_X2 U5017 ( .A1(n1501), .A2(n1503), .A3(n1321), .ZN(n9462) );
  NAND2_X1 U5018 ( .A1(n8979), .A2(n9265), .ZN(n9264) );
  NAND2_X1 U5020 ( .A1(n1325), .A2(n9214), .ZN(n1322) );
  NAND2_X1 U5021 ( .A1(n2726), .A2(n1326), .ZN(n1325) );
  NAND3_X1 U5022 ( .A1(n1332), .A2(n20496), .A3(n11384), .ZN(n1327) );
  NAND2_X1 U5023 ( .A1(n1331), .A2(n1330), .ZN(n1329) );
  NAND2_X1 U5024 ( .A1(n12101), .A2(n20468), .ZN(n11384) );
  INV_X1 U5025 ( .A(n11384), .ZN(n1331) );
  NAND2_X1 U5026 ( .A1(n3601), .A2(n10684), .ZN(n1332) );
  NAND2_X1 U5028 ( .A1(n7879), .A2(n8053), .ZN(n1335) );
  NAND2_X1 U5030 ( .A1(n5797), .A2(n5796), .ZN(n4182) );
  OAI21_X1 U5031 ( .B1(n12298), .B2(n12299), .A(n12274), .ZN(n1336) );
  NAND3_X1 U5032 ( .A1(n14576), .A2(n14574), .A3(n14575), .ZN(n14577) );
  NAND2_X1 U5033 ( .A1(n8070), .A2(n7420), .ZN(n8208) );
  NAND2_X1 U5034 ( .A1(n9317), .A2(n9065), .ZN(n8466) );
  NAND2_X1 U5037 ( .A1(n11572), .A2(n11573), .ZN(n1338) );
  OAI22_X1 U5039 ( .A1(n3458), .A2(n11125), .B1(n19949), .B2(n10813), .ZN(
        n3459) );
  OAI21_X1 U5041 ( .B1(n7671), .B2(n20252), .A(n8377), .ZN(n8145) );
  OR2_X1 U5042 ( .A1(n14213), .A2(n3497), .ZN(n3274) );
  NAND3_X1 U5043 ( .A1(n16442), .A2(n16167), .A3(n17505), .ZN(n2633) );
  NAND2_X1 U5044 ( .A1(n2732), .A2(n1339), .ZN(n2733) );
  AOI22_X1 U5045 ( .A1(n12470), .A2(n12466), .B1(n12467), .B2(n12468), .ZN(
        n1339) );
  NAND2_X1 U5046 ( .A1(n5682), .A2(n5410), .ZN(n5686) );
  NAND2_X1 U5048 ( .A1(n4621), .A2(n20143), .ZN(n4624) );
  NAND2_X1 U5049 ( .A1(n18214), .A2(n18213), .ZN(n17560) );
  NAND2_X1 U5050 ( .A1(n2951), .A2(n2950), .ZN(n18214) );
  NAND2_X1 U5051 ( .A1(n3306), .A2(n1723), .ZN(n1722) );
  NOR2_X1 U5052 ( .A1(n9255), .A2(n8974), .ZN(n8970) );
  INV_X1 U5053 ( .A(n11476), .ZN(n3482) );
  NOR2_X1 U5054 ( .A1(n15294), .A2(n14461), .ZN(n15107) );
  INV_X1 U5055 ( .A(n8941), .ZN(n8730) );
  OR2_X1 U5056 ( .A1(n9320), .A2(n9836), .ZN(n1855) );
  AND2_X1 U5057 ( .A1(n6379), .A2(n5728), .ZN(n5383) );
  OAI21_X1 U5058 ( .B1(n5383), .B2(n19476), .A(n5846), .ZN(n1568) );
  INV_X1 U5059 ( .A(n13891), .ZN(n14799) );
  INV_X1 U5060 ( .A(n1654), .ZN(n11155) );
  XNOR2_X1 U5061 ( .A(n6794), .B(n3590), .ZN(n6684) );
  INV_X1 U5062 ( .A(n7932), .ZN(n2031) );
  AOI21_X1 U5063 ( .B1(n17080), .B2(n3114), .A(n17825), .ZN(n3115) );
  AOI22_X1 U5064 ( .A1(n5433), .A2(n5432), .B1(n5996), .B2(n3627), .ZN(n5437)
         );
  XNOR2_X1 U5065 ( .A(n2582), .B(n13433), .ZN(n1756) );
  NAND3_X1 U5066 ( .A1(n5242), .A2(n3086), .A3(n5241), .ZN(n5245) );
  OAI211_X2 U5067 ( .C1(n5180), .C2(n4632), .A(n5179), .B(n5178), .ZN(n6985)
         );
  XNOR2_X1 U5068 ( .A(n13064), .B(n19337), .ZN(n13067) );
  OAI22_X1 U5069 ( .A1(n8763), .A2(n8693), .B1(n2243), .B2(n9177), .ZN(n8694)
         );
  OAI21_X2 U5070 ( .B1(n8585), .B2(n9304), .A(n1340), .ZN(n10612) );
  NAND2_X1 U5071 ( .A1(n2073), .A2(n2074), .ZN(n1340) );
  NAND2_X1 U5073 ( .A1(n19519), .A2(n9291), .ZN(n9051) );
  AND2_X2 U5074 ( .A1(n7896), .A2(n7895), .ZN(n8649) );
  OAI21_X1 U5075 ( .B1(n3711), .B2(n11216), .A(n1341), .ZN(n11477) );
  NAND2_X1 U5076 ( .A1(n3711), .A2(n11076), .ZN(n1341) );
  NAND3_X1 U5077 ( .A1(n14937), .A2(n1344), .A3(n1343), .ZN(n16045) );
  NAND2_X1 U5078 ( .A1(n1019), .A2(n13933), .ZN(n1343) );
  NAND2_X1 U5079 ( .A1(n14936), .A2(n15506), .ZN(n1344) );
  NAND2_X1 U5080 ( .A1(n1347), .A2(n1345), .ZN(n5247) );
  NAND2_X1 U5081 ( .A1(n5246), .A2(n20405), .ZN(n1345) );
  INV_X1 U5083 ( .A(n9188), .ZN(n1778) );
  NAND3_X1 U5084 ( .A1(n4222), .A2(n1028), .A3(n1348), .ZN(n6022) );
  NAND2_X1 U5085 ( .A1(n4840), .A2(n3977), .ZN(n1348) );
  NAND2_X1 U5086 ( .A1(n15257), .A2(n15256), .ZN(n1349) );
  OR2_X1 U5087 ( .A1(n11565), .A2(n11569), .ZN(n2948) );
  NAND2_X1 U5089 ( .A1(n13893), .A2(n1351), .ZN(n1350) );
  NAND2_X1 U5090 ( .A1(n14800), .A2(n14796), .ZN(n13893) );
  INV_X1 U5091 ( .A(n12141), .ZN(n11931) );
  NAND2_X1 U5093 ( .A1(n12288), .A2(n11792), .ZN(n1512) );
  NAND2_X1 U5094 ( .A1(n4170), .A2(n4169), .ZN(n4018) );
  NAND2_X1 U5096 ( .A1(n2482), .A2(n1883), .ZN(n1353) );
  INV_X1 U5097 ( .A(n2456), .ZN(n1354) );
  NAND2_X1 U5098 ( .A1(n19922), .A2(n7615), .ZN(n2456) );
  INV_X1 U5101 ( .A(n4696), .ZN(n2872) );
  NAND2_X1 U5102 ( .A1(n4439), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5103 ( .A1(n10815), .A2(n10814), .ZN(n1356) );
  NAND2_X1 U5104 ( .A1(n10816), .A2(n19949), .ZN(n1357) );
  OR2_X1 U5105 ( .A1(n7801), .A2(n8016), .ZN(n3211) );
  NAND2_X1 U5106 ( .A1(n8079), .A2(n8219), .ZN(n8077) );
  XNOR2_X2 U5107 ( .A(n6460), .B(n6459), .ZN(n8219) );
  NAND2_X1 U5109 ( .A1(n4872), .A2(n4873), .ZN(n5899) );
  NAND2_X1 U5111 ( .A1(n1359), .A2(n1358), .ZN(n15339) );
  OR2_X1 U5112 ( .A1(n12873), .A2(n14448), .ZN(n1358) );
  XNOR2_X2 U5113 ( .A(n5191), .B(n5190), .ZN(n8304) );
  OAI211_X1 U5114 ( .C1(n12352), .C2(n12354), .A(n3330), .B(n12355), .ZN(
        n12356) );
  XNOR2_X2 U5115 ( .A(n3944), .B(Key[182]), .ZN(n4355) );
  INV_X1 U5116 ( .A(Plaintext[29]), .ZN(n2036) );
  NAND3_X1 U5118 ( .A1(n8052), .A2(n8192), .A3(n8196), .ZN(n1361) );
  NAND2_X1 U5120 ( .A1(n2499), .A2(n8786), .ZN(n9147) );
  OAI21_X1 U5122 ( .B1(n11346), .B2(n11238), .A(n1365), .ZN(n10149) );
  NAND2_X1 U5123 ( .A1(n11346), .A2(n11239), .ZN(n1365) );
  NOR2_X1 U5124 ( .A1(n3733), .A2(n12562), .ZN(n11726) );
  OR2_X1 U5125 ( .A1(n11990), .A2(n12334), .ZN(n11667) );
  NAND2_X1 U5126 ( .A1(n1367), .A2(n3589), .ZN(n5665) );
  OAI21_X1 U5127 ( .B1(n283), .B2(n5663), .A(n5664), .ZN(n1367) );
  NAND2_X1 U5128 ( .A1(n14660), .A2(n14659), .ZN(n1368) );
  XNOR2_X1 U5129 ( .A(n6632), .B(n6686), .ZN(n1369) );
  XOR2_X1 U5130 ( .A(n13033), .B(n13032), .Z(n2240) );
  OAI21_X1 U5131 ( .B1(n4913), .B2(n4911), .A(n4477), .ZN(n3871) );
  AOI21_X1 U5132 ( .B1(n14506), .B2(n14498), .A(n14499), .ZN(n1762) );
  NAND2_X1 U5133 ( .A1(n1372), .A2(n1370), .ZN(n11896) );
  NAND2_X1 U5134 ( .A1(n11962), .A2(n1371), .ZN(n1370) );
  NAND2_X1 U5136 ( .A1(n1373), .A2(n180), .ZN(n1372) );
  NAND2_X1 U5137 ( .A1(n12629), .A2(n11618), .ZN(n1373) );
  XNOR2_X1 U5138 ( .A(n1374), .B(n18849), .ZN(Ciphertext[96]) );
  NAND2_X1 U5140 ( .A1(n12283), .A2(n20215), .ZN(n11580) );
  NAND2_X1 U5142 ( .A1(n11107), .A2(n19830), .ZN(n1376) );
  INV_X1 U5144 ( .A(n11431), .ZN(n1378) );
  NOR2_X1 U5145 ( .A1(n8957), .A2(n1379), .ZN(n9670) );
  OAI22_X1 U5146 ( .A1(n9370), .A2(n8602), .B1(n8951), .B2(n8950), .ZN(n1379)
         );
  NAND2_X1 U5148 ( .A1(n11708), .A2(n12479), .ZN(n1380) );
  XNOR2_X1 U5149 ( .A(n13409), .B(n13767), .ZN(n11029) );
  NOR2_X2 U5150 ( .A1(n11024), .A2(n11023), .ZN(n13409) );
  NAND2_X1 U5151 ( .A1(n1382), .A2(n1381), .ZN(n5341) );
  NAND2_X1 U5152 ( .A1(n6123), .A2(n5868), .ZN(n1381) );
  NAND2_X1 U5155 ( .A1(n1385), .A2(n1384), .ZN(n19228) );
  NAND2_X1 U5156 ( .A1(n19754), .A2(n19227), .ZN(n1384) );
  NAND2_X1 U5157 ( .A1(n20124), .A2(n19235), .ZN(n1385) );
  OAI21_X2 U5158 ( .B1(n4680), .B2(n169), .A(n4679), .ZN(n6166) );
  OAI21_X1 U5159 ( .B1(n11438), .B2(n11439), .A(n11437), .ZN(n11441) );
  NAND2_X1 U5160 ( .A1(n8674), .A2(n8672), .ZN(n7465) );
  NAND2_X1 U5161 ( .A1(n8960), .A2(n8959), .ZN(n8502) );
  NAND2_X1 U5162 ( .A1(n15101), .A2(n15838), .ZN(n15102) );
  NAND2_X1 U5163 ( .A1(n4764), .A2(n19788), .ZN(n5027) );
  NAND2_X1 U5164 ( .A1(n13506), .A2(n1014), .ZN(n13508) );
  NAND2_X1 U5165 ( .A1(n12451), .A2(n12452), .ZN(n12454) );
  OR2_X1 U5166 ( .A1(n19474), .A2(n8193), .ZN(n7881) );
  NAND2_X1 U5168 ( .A1(n11143), .A2(n10957), .ZN(n10702) );
  OR2_X1 U5169 ( .A1(n11256), .A2(n11321), .ZN(n10776) );
  NAND2_X2 U5171 ( .A1(n7884), .A2(n7883), .ZN(n9274) );
  OR2_X1 U5172 ( .A1(n4440), .A2(n4439), .ZN(n4795) );
  AOI22_X1 U5174 ( .A1(n3468), .A2(n5985), .B1(n5989), .B2(n5711), .ZN(n4113)
         );
  AOI21_X1 U5175 ( .B1(n1388), .B2(n20472), .A(n2225), .ZN(n9303) );
  NOR2_X1 U5176 ( .A1(n270), .A2(n9300), .ZN(n1388) );
  NAND3_X1 U5178 ( .A1(n3917), .A2(n3131), .A3(n4753), .ZN(n1389) );
  NAND2_X1 U5179 ( .A1(n3918), .A2(n1391), .ZN(n1390) );
  NAND2_X1 U5180 ( .A1(n2419), .A2(n9201), .ZN(n2418) );
  NAND2_X1 U5181 ( .A1(n20009), .A2(n9204), .ZN(n2419) );
  NAND3_X1 U5182 ( .A1(n5620), .A2(n6148), .A3(n6138), .ZN(n5343) );
  NAND2_X1 U5183 ( .A1(n2593), .A2(n2594), .ZN(n2592) );
  NAND2_X1 U5186 ( .A1(n1394), .A2(n6042), .ZN(n1393) );
  OAI21_X1 U5187 ( .B1(n6041), .B2(n5144), .A(n2149), .ZN(n1394) );
  NAND2_X1 U5188 ( .A1(n1213), .A2(n12334), .ZN(n1396) );
  NAND2_X1 U5189 ( .A1(n12335), .A2(n11990), .ZN(n1397) );
  OAI21_X1 U5190 ( .B1(n8424), .B2(n8423), .A(n8781), .ZN(n1398) );
  OAI211_X2 U5191 ( .C1(n8634), .C2(n8633), .A(n8632), .B(n8631), .ZN(n10359)
         );
  OAI21_X1 U5192 ( .B1(n11989), .B2(n14623), .A(n1399), .ZN(n14849) );
  NAND2_X1 U5193 ( .A1(n14195), .A2(n11988), .ZN(n1399) );
  NAND2_X1 U5194 ( .A1(n10995), .A2(n10946), .ZN(n9560) );
  AOI21_X1 U5195 ( .B1(n20165), .B2(n7770), .A(n2976), .ZN(n7772) );
  INV_X1 U5196 ( .A(n15503), .ZN(n1758) );
  XNOR2_X1 U5197 ( .A(n13464), .B(n2881), .ZN(n2264) );
  NAND2_X1 U5198 ( .A1(n1403), .A2(n11867), .ZN(n2365) );
  XNOR2_X1 U5199 ( .A(n7289), .B(n18170), .ZN(n6932) );
  NAND2_X1 U5201 ( .A1(n8602), .A2(n8482), .ZN(n9372) );
  NAND2_X1 U5202 ( .A1(n1405), .A2(n8093), .ZN(n1404) );
  NAND2_X1 U5203 ( .A1(n1407), .A2(n1406), .ZN(n10470) );
  NAND2_X1 U5204 ( .A1(n10468), .A2(n11201), .ZN(n1406) );
  NAND2_X1 U5205 ( .A1(n10469), .A2(n11093), .ZN(n1407) );
  NAND2_X1 U5206 ( .A1(n9931), .A2(n11523), .ZN(n9932) );
  NAND2_X1 U5207 ( .A1(n19270), .A2(n19271), .ZN(n19272) );
  NAND2_X1 U5209 ( .A1(n9328), .A2(n9330), .ZN(n1408) );
  XNOR2_X1 U5211 ( .A(n10610), .B(n10609), .ZN(n10730) );
  OR2_X1 U5212 ( .A1(n2527), .A2(n16306), .ZN(n17648) );
  NOR2_X1 U5213 ( .A1(n20000), .A2(n9105), .ZN(n8423) );
  MUX2_X1 U5214 ( .A(n14525), .B(n951), .S(n14648), .Z(n14310) );
  INV_X1 U5216 ( .A(n5046), .ZN(n4796) );
  INV_X1 U5217 ( .A(n1508), .ZN(n12130) );
  INV_X1 U5218 ( .A(n2005), .ZN(n1491) );
  NOR2_X1 U5219 ( .A1(n10911), .A2(n12606), .ZN(n3764) );
  AOI22_X1 U5220 ( .A1(n14944), .A2(n2645), .B1(n15107), .B2(n2644), .ZN(n2643) );
  NAND2_X1 U5221 ( .A1(n7618), .A2(n7420), .ZN(n1411) );
  NAND3_X1 U5223 ( .A1(n3404), .A2(n1414), .A3(n1413), .ZN(n12284) );
  NAND2_X1 U5224 ( .A1(n20184), .A2(n3402), .ZN(n1413) );
  NAND2_X1 U5225 ( .A1(n14509), .A2(n14644), .ZN(n14508) );
  NAND2_X1 U5226 ( .A1(n1415), .A2(n14354), .ZN(n15909) );
  NAND2_X1 U5227 ( .A1(n1572), .A2(n1571), .ZN(n1415) );
  NOR2_X1 U5229 ( .A1(n8315), .A2(n7475), .ZN(n7594) );
  AOI21_X1 U5230 ( .B1(n4543), .B2(n4544), .A(n4542), .ZN(n5538) );
  NAND3_X1 U5232 ( .A1(n8033), .A2(n20012), .A3(n8034), .ZN(n1416) );
  NAND3_X2 U5233 ( .A1(n2121), .A2(n11720), .A3(n967), .ZN(n13491) );
  OR2_X1 U5234 ( .A1(n11073), .A2(n10898), .ZN(n1418) );
  NAND2_X1 U5236 ( .A1(n2143), .A2(n11804), .ZN(n1419) );
  OR2_X1 U5237 ( .A1(n8200), .A2(n5762), .ZN(n7872) );
  INV_X1 U5238 ( .A(n5102), .ZN(n1421) );
  NAND2_X1 U5239 ( .A1(n10923), .A2(n11523), .ZN(n12222) );
  INV_X1 U5240 ( .A(n13017), .ZN(n13576) );
  INV_X1 U5241 ( .A(n1640), .ZN(n15395) );
  NAND2_X1 U5243 ( .A1(n1423), .A2(n4413), .ZN(n4414) );
  NAND2_X1 U5244 ( .A1(n4412), .A2(n4411), .ZN(n1423) );
  NAND2_X1 U5245 ( .A1(n8324), .A2(n19856), .ZN(n1424) );
  INV_X1 U5246 ( .A(n7786), .ZN(n1425) );
  OR2_X1 U5247 ( .A1(n12383), .A2(n12468), .ZN(n3783) );
  OR2_X1 U5248 ( .A1(n2628), .A2(n13891), .ZN(n14797) );
  NAND2_X1 U5249 ( .A1(n8619), .A2(n2243), .ZN(n2242) );
  AND2_X1 U5250 ( .A1(n2523), .A2(n12759), .ZN(n12411) );
  NAND2_X1 U5251 ( .A1(n1426), .A2(n6104), .ZN(n5956) );
  OAI22_X1 U5252 ( .A1(n5957), .A2(n6107), .B1(n6113), .B2(n6105), .ZN(n1426)
         );
  OR2_X1 U5253 ( .A1(n8650), .A2(n8649), .ZN(n9281) );
  AOI22_X1 U5254 ( .A1(n8252), .A2(n8251), .B1(n8253), .B2(n8254), .ZN(n8255)
         );
  XNOR2_X1 U5256 ( .A(n1427), .B(n12896), .ZN(n12898) );
  XNOR2_X1 U5257 ( .A(n12897), .B(n13126), .ZN(n1427) );
  AND3_X1 U5259 ( .A1(n14988), .A2(n14990), .A3(n14989), .ZN(n14991) );
  OAI21_X1 U5260 ( .B1(n12631), .B2(n12630), .A(n11619), .ZN(n11960) );
  INV_X1 U5261 ( .A(n15059), .ZN(n15061) );
  XNOR2_X1 U5262 ( .A(n2285), .B(n8508), .ZN(n10755) );
  OAI21_X1 U5263 ( .B1(n19657), .B2(n3522), .A(n19819), .ZN(n3253) );
  INV_X1 U5265 ( .A(n4233), .ZN(n4860) );
  XNOR2_X1 U5266 ( .A(n10151), .B(n10002), .ZN(n9261) );
  INV_X1 U5267 ( .A(n1746), .ZN(n6186) );
  INV_X1 U5268 ( .A(n1776), .ZN(n2407) );
  INV_X1 U5269 ( .A(n15683), .ZN(n15782) );
  INV_X1 U5270 ( .A(n12162), .ZN(n12535) );
  NAND3_X1 U5271 ( .A1(n19520), .A2(n7592), .A3(n8313), .ZN(n7597) );
  INV_X1 U5272 ( .A(n15266), .ZN(n15847) );
  INV_X1 U5273 ( .A(n8937), .ZN(n8940) );
  OAI21_X1 U5274 ( .B1(n19505), .B2(n19719), .A(n11490), .ZN(n2134) );
  XNOR2_X1 U5275 ( .A(n7303), .B(n3067), .ZN(n7310) );
  INV_X1 U5276 ( .A(n1603), .ZN(n1428) );
  NAND2_X1 U5277 ( .A1(n1430), .A2(n1429), .ZN(n8724) );
  NAND3_X1 U5278 ( .A1(n9358), .A2(n9359), .A3(n9528), .ZN(n1429) );
  NAND2_X1 U5279 ( .A1(n8723), .A2(n9356), .ZN(n1430) );
  XNOR2_X1 U5280 ( .A(n6867), .B(n6977), .ZN(n7353) );
  NOR2_X2 U5281 ( .A1(n8065), .A2(n1431), .ZN(n9065) );
  NAND2_X1 U5282 ( .A1(n1433), .A2(n1432), .ZN(n1431) );
  NAND2_X1 U5283 ( .A1(n8063), .A2(n8190), .ZN(n1432) );
  AOI21_X1 U5286 ( .B1(n4584), .B2(n4582), .A(n4271), .ZN(n2334) );
  NAND2_X1 U5287 ( .A1(n4269), .A2(n4095), .ZN(n4584) );
  OAI21_X1 U5289 ( .B1(n11145), .B2(n10642), .A(n1749), .ZN(n1670) );
  NAND2_X1 U5290 ( .A1(n5698), .A2(n5973), .ZN(n1435) );
  XNOR2_X1 U5291 ( .A(n17267), .B(n16508), .ZN(n1436) );
  NAND2_X1 U5294 ( .A1(n7724), .A2(n8159), .ZN(n8258) );
  NAND2_X1 U5296 ( .A1(n12522), .A2(n182), .ZN(n1439) );
  NAND2_X1 U5297 ( .A1(n17665), .A2(n17662), .ZN(n17086) );
  NAND3_X1 U5298 ( .A1(n4360), .A2(n4359), .A3(n2370), .ZN(n5483) );
  NOR2_X1 U5299 ( .A1(n4363), .A2(n5719), .ZN(n5240) );
  NOR2_X1 U5301 ( .A1(n1442), .A2(n4033), .ZN(n1441) );
  NAND2_X1 U5303 ( .A1(n15438), .A2(n15775), .ZN(n1444) );
  NAND2_X1 U5305 ( .A1(n4896), .A2(n4897), .ZN(n1445) );
  OAI22_X2 U5306 ( .A1(n6047), .A2(n5313), .B1(n5312), .B2(n5781), .ZN(n6728)
         );
  NAND2_X1 U5307 ( .A1(n10889), .A2(n10926), .ZN(n1446) );
  NAND2_X1 U5308 ( .A1(n10844), .A2(n193), .ZN(n1447) );
  NAND2_X1 U5309 ( .A1(n1448), .A2(n709), .ZN(n1485) );
  NOR2_X1 U5310 ( .A1(n1449), .A2(n9103), .ZN(n1448) );
  NAND2_X1 U5311 ( .A1(n9100), .A2(n9099), .ZN(n1449) );
  NOR2_X1 U5312 ( .A1(n20007), .A2(n3430), .ZN(n3429) );
  INV_X1 U5314 ( .A(n8917), .ZN(n8734) );
  INV_X1 U5315 ( .A(n4337), .ZN(n3753) );
  OR2_X1 U5316 ( .A1(n3753), .A2(n1017), .ZN(n3607) );
  NOR2_X1 U5317 ( .A1(n14790), .A2(n14103), .ZN(n2411) );
  NAND2_X1 U5319 ( .A1(n17944), .A2(n19105), .ZN(n1450) );
  NOR2_X2 U5321 ( .A1(n14107), .A2(n14108), .ZN(n16429) );
  NOR2_X1 U5322 ( .A1(n11534), .A2(n19915), .ZN(n11536) );
  NAND2_X1 U5325 ( .A1(n9204), .A2(n9201), .ZN(n8433) );
  NAND2_X1 U5327 ( .A1(n14237), .A2(n14406), .ZN(n14242) );
  NAND2_X1 U5328 ( .A1(n12531), .A2(n924), .ZN(n12530) );
  NAND2_X1 U5330 ( .A1(n2048), .A2(n5997), .ZN(n1455) );
  NAND2_X1 U5331 ( .A1(n1457), .A2(n1456), .ZN(n13568) );
  NAND2_X1 U5332 ( .A1(n14860), .A2(n15237), .ZN(n1456) );
  NAND2_X1 U5333 ( .A1(n13561), .A2(n1458), .ZN(n1457) );
  NAND2_X1 U5334 ( .A1(n12154), .A2(n12152), .ZN(n11711) );
  NAND2_X1 U5335 ( .A1(n11169), .A2(n11170), .ZN(n1459) );
  NAND2_X1 U5336 ( .A1(n8840), .A2(n1461), .ZN(n10422) );
  NAND3_X1 U5337 ( .A1(n1631), .A2(n1630), .A3(n8676), .ZN(n1461) );
  OAI21_X1 U5338 ( .B1(n10667), .B2(n11399), .A(n2044), .ZN(n2043) );
  NAND3_X1 U5339 ( .A1(n14430), .A2(n3154), .A3(n14494), .ZN(n2138) );
  NAND2_X1 U5340 ( .A1(n1462), .A2(n8205), .ZN(n7874) );
  NAND2_X1 U5341 ( .A1(n2378), .A2(n2379), .ZN(n1462) );
  NAND2_X1 U5342 ( .A1(n17891), .A2(n17890), .ZN(n17662) );
  XNOR2_X2 U5343 ( .A(n16109), .B(n16108), .ZN(n17890) );
  INV_X1 U5344 ( .A(n12211), .ZN(n2712) );
  NAND2_X1 U5345 ( .A1(n1464), .A2(n1463), .ZN(n9583) );
  NAND2_X1 U5346 ( .A1(n9287), .A2(n9576), .ZN(n1463) );
  NAND2_X1 U5347 ( .A1(n9288), .A2(n9289), .ZN(n1464) );
  INV_X1 U5349 ( .A(n1506), .ZN(n3182) );
  NAND2_X1 U5350 ( .A1(n8356), .A2(n1506), .ZN(n1480) );
  NAND2_X1 U5351 ( .A1(n3181), .A2(n7500), .ZN(n1506) );
  NAND2_X1 U5353 ( .A1(n9104), .A2(n8781), .ZN(n9109) );
  NAND2_X1 U5354 ( .A1(n1465), .A2(n4691), .ZN(n4688) );
  NAND2_X1 U5355 ( .A1(n1468), .A2(n1466), .ZN(n2396) );
  NAND2_X1 U5357 ( .A1(n1820), .A2(n14738), .ZN(n1469) );
  NAND2_X1 U5358 ( .A1(n1470), .A2(n8478), .ZN(n10497) );
  XNOR2_X2 U5363 ( .A(Key[35]), .B(Plaintext[35]), .ZN(n4954) );
  OR2_X1 U5366 ( .A1(n12579), .A2(n12576), .ZN(n11924) );
  XNOR2_X1 U5367 ( .A(n7325), .B(n2571), .ZN(n6881) );
  INV_X1 U5368 ( .A(n4524), .ZN(n4516) );
  INV_X1 U5369 ( .A(n8195), .ZN(n8054) );
  INV_X1 U5370 ( .A(n2749), .ZN(n2504) );
  NAND2_X1 U5371 ( .A1(n4426), .A2(n4827), .ZN(n1472) );
  OAI21_X1 U5372 ( .B1(n1039), .B2(n1317), .A(n1473), .ZN(n11362) );
  NOR2_X1 U5373 ( .A1(n11127), .A2(n19949), .ZN(n1473) );
  INV_X1 U5374 ( .A(n1475), .ZN(n1474) );
  OAI21_X1 U5375 ( .B1(n5748), .B2(n2482), .A(n5205), .ZN(n1475) );
  NAND2_X1 U5376 ( .A1(n15295), .A2(n15297), .ZN(n14770) );
  OAI22_X1 U5378 ( .A1(n1806), .A2(n5730), .B1(n5847), .B2(n1805), .ZN(n1476)
         );
  NAND2_X1 U5379 ( .A1(n2461), .A2(n5098), .ZN(n4712) );
  NAND2_X1 U5380 ( .A1(n8722), .A2(n9359), .ZN(n8721) );
  NAND2_X2 U5381 ( .A1(n3490), .A2(n7672), .ZN(n9359) );
  XNOR2_X1 U5382 ( .A(n6728), .B(n456), .ZN(n6729) );
  NAND2_X1 U5383 ( .A1(n207), .A2(n8958), .ZN(n1478) );
  INV_X1 U5384 ( .A(n12137), .ZN(n12385) );
  NAND3_X1 U5385 ( .A1(n12468), .A2(n12386), .A3(n12137), .ZN(n1946) );
  XNOR2_X1 U5386 ( .A(n6960), .B(n980), .ZN(n6227) );
  XNOR2_X1 U5387 ( .A(n7348), .B(n6226), .ZN(n6960) );
  XNOR2_X1 U5388 ( .A(n9773), .B(n9774), .ZN(n1479) );
  INV_X1 U5389 ( .A(n6109), .ZN(n5657) );
  NAND2_X1 U5390 ( .A1(n1899), .A2(n1901), .ZN(n14847) );
  NAND2_X1 U5391 ( .A1(n11094), .A2(n11443), .ZN(n11448) );
  NAND2_X1 U5393 ( .A1(n14275), .A2(n20498), .ZN(n13957) );
  NAND2_X1 U5394 ( .A1(n8093), .A2(n8212), .ZN(n7432) );
  NAND2_X1 U5395 ( .A1(n4186), .A2(n4185), .ZN(n3622) );
  NAND2_X1 U5396 ( .A1(n4156), .A2(n3623), .ZN(n4186) );
  NAND2_X1 U5397 ( .A1(n1480), .A2(n1565), .ZN(n2930) );
  OR2_X1 U5398 ( .A1(n9251), .A2(n8974), .ZN(n1481) );
  NOR2_X1 U5399 ( .A1(n3403), .A2(n180), .ZN(n3402) );
  OAI21_X1 U5400 ( .B1(n11578), .B2(n11739), .A(n11577), .ZN(n2367) );
  NAND3_X2 U5402 ( .A1(n1854), .A2(n11274), .A3(n974), .ZN(n12807) );
  OAI211_X1 U5403 ( .C1(n9004), .C2(n8890), .A(n19490), .B(n1484), .ZN(n8626)
         );
  NAND2_X1 U5404 ( .A1(n12545), .A2(n12542), .ZN(n12306) );
  INV_X1 U5405 ( .A(n13989), .ZN(n15302) );
  NAND2_X1 U5406 ( .A1(n15714), .A2(n15874), .ZN(n13989) );
  OAI21_X1 U5407 ( .B1(n19515), .B2(n20000), .A(n1485), .ZN(n9110) );
  OAI21_X1 U5409 ( .B1(n14688), .B2(n14690), .A(n14385), .ZN(n1486) );
  AOI21_X1 U5410 ( .B1(n9028), .B2(n8829), .A(n9029), .ZN(n1487) );
  NAND3_X1 U5411 ( .A1(n885), .A2(n9274), .A3(n9275), .ZN(n9280) );
  XNOR2_X2 U5412 ( .A(Key[21]), .B(Plaintext[21]), .ZN(n4297) );
  XOR2_X1 U5413 ( .A(n13550), .B(n13080), .Z(n1809) );
  OAI211_X2 U5414 ( .C1(n9069), .C2(n545), .A(n2502), .B(n2503), .ZN(n10220)
         );
  NAND2_X1 U5415 ( .A1(n18427), .A2(n15529), .ZN(n1701) );
  AND3_X2 U5416 ( .A1(n2643), .A2(n2646), .A3(n3308), .ZN(n17269) );
  OAI21_X1 U5417 ( .B1(n17483), .B2(n19823), .A(n1488), .ZN(n15177) );
  NAND2_X1 U5418 ( .A1(n1718), .A2(n17243), .ZN(n1488) );
  NOR2_X1 U5419 ( .A1(n15239), .A2(n3348), .ZN(n1489) );
  INV_X1 U5420 ( .A(n9563), .ZN(n9340) );
  NAND3_X1 U5421 ( .A1(n1493), .A2(n1492), .A3(n1491), .ZN(n1490) );
  NAND2_X1 U5422 ( .A1(n15443), .A2(n15228), .ZN(n1492) );
  NAND2_X1 U5423 ( .A1(n15446), .A2(n1494), .ZN(n1493) );
  NAND2_X1 U5424 ( .A1(n1495), .A2(n9023), .ZN(n2025) );
  OAI22_X1 U5425 ( .A1(n8515), .A2(n9021), .B1(n8841), .B2(n8672), .ZN(n1495)
         );
  AND3_X2 U5426 ( .A1(n17567), .A2(n1496), .A3(n17561), .ZN(n18600) );
  NAND2_X1 U5427 ( .A1(n17563), .A2(n17562), .ZN(n1496) );
  NAND2_X1 U5428 ( .A1(n9411), .A2(n19817), .ZN(n1497) );
  NAND3_X2 U5430 ( .A1(n1500), .A2(n3771), .A3(n1499), .ZN(n8979) );
  NAND2_X1 U5431 ( .A1(n8771), .A2(n8979), .ZN(n1501) );
  INV_X1 U5432 ( .A(n3775), .ZN(n1502) );
  NAND2_X1 U5433 ( .A1(n1504), .A2(n19880), .ZN(n1503) );
  NAND2_X1 U5434 ( .A1(n1505), .A2(n9266), .ZN(n1504) );
  NAND2_X1 U5435 ( .A1(n7866), .A2(n9262), .ZN(n1505) );
  NAND2_X1 U5436 ( .A1(n7742), .A2(n1506), .ZN(n7698) );
  NAND2_X1 U5440 ( .A1(n1507), .A2(n8126), .ZN(n6439) );
  NOR2_X1 U5441 ( .A1(n1507), .A2(n8470), .ZN(n9087) );
  NOR2_X1 U5442 ( .A1(n8565), .A2(n1507), .ZN(n1575) );
  NAND3_X1 U5443 ( .A1(n9091), .A2(n1507), .A3(n8884), .ZN(n8887) );
  NAND2_X1 U5444 ( .A1(n9090), .A2(n1507), .ZN(n1577) );
  MUX2_X1 U5445 ( .A(n1507), .B(n8565), .S(n9091), .Z(n8130) );
  NAND3_X1 U5446 ( .A1(n8471), .A2(n1507), .A3(n8470), .ZN(n8472) );
  OR2_X1 U5448 ( .A1(n11586), .A2(n1508), .ZN(n1547) );
  AND2_X1 U5449 ( .A1(n12127), .A2(n1508), .ZN(n1643) );
  NAND2_X1 U5450 ( .A1(n10967), .A2(n1508), .ZN(n10974) );
  OAI21_X1 U5451 ( .B1(n11763), .B2(n12126), .A(n1508), .ZN(n11587) );
  AOI21_X1 U5452 ( .B1(n10972), .B2(n1508), .A(n1735), .ZN(n10973) );
  NAND3_X1 U5453 ( .A1(n1512), .A2(n1511), .A3(n1510), .ZN(n1509) );
  NAND2_X1 U5454 ( .A1(n12520), .A2(n12523), .ZN(n1510) );
  NAND2_X1 U5455 ( .A1(n11793), .A2(n12523), .ZN(n1514) );
  OAI21_X1 U5456 ( .B1(n9220), .B2(n1516), .A(n1515), .ZN(n2452) );
  INV_X1 U5457 ( .A(n9218), .ZN(n1515) );
  NOR2_X1 U5458 ( .A1(n8797), .A2(n9113), .ZN(n1516) );
  NOR2_X1 U5459 ( .A1(n9112), .A2(n9114), .ZN(n9220) );
  NAND2_X1 U5460 ( .A1(n1517), .A2(n15364), .ZN(n15367) );
  NAND2_X1 U5461 ( .A1(n1520), .A2(n15577), .ZN(n1517) );
  NAND2_X1 U5462 ( .A1(n14643), .A2(n20473), .ZN(n1518) );
  NAND2_X1 U5463 ( .A1(n14646), .A2(n14645), .ZN(n1519) );
  NAND2_X1 U5464 ( .A1(n251), .A2(n12443), .ZN(n1521) );
  OAI211_X1 U5465 ( .C1(n12109), .C2(n1522), .A(n1521), .B(n12441), .ZN(n12112) );
  INV_X1 U5466 ( .A(n12442), .ZN(n1522) );
  OR2_X2 U5467 ( .A1(n10682), .A2(n10681), .ZN(n12442) );
  NAND2_X1 U5468 ( .A1(n12441), .A2(n12442), .ZN(n12444) );
  NAND2_X1 U5469 ( .A1(n12438), .A2(n1522), .ZN(n12113) );
  AOI22_X1 U5470 ( .A1(n12438), .A2(n12437), .B1(n1522), .B2(n12436), .ZN(
        n12447) );
  NAND2_X1 U5471 ( .A1(n15711), .A2(n15871), .ZN(n1525) );
  NOR2_X1 U5475 ( .A1(n14154), .A2(n20171), .ZN(n13996) );
  AND2_X1 U5476 ( .A1(n1527), .A2(n14394), .ZN(n14397) );
  NOR2_X1 U5477 ( .A1(n5630), .A2(n5631), .ZN(n1949) );
  OAI21_X2 U5478 ( .B1(n4330), .B2(n4331), .A(n4329), .ZN(n5631) );
  XNOR2_X1 U5479 ( .A(n17296), .B(n17302), .ZN(n1529) );
  XNOR2_X2 U5480 ( .A(n1530), .B(Plaintext[191]), .ZN(n4615) );
  INV_X1 U5481 ( .A(Key[191]), .ZN(n1530) );
  NAND2_X1 U5482 ( .A1(n1531), .A2(n18688), .ZN(n17988) );
  NAND2_X1 U5483 ( .A1(n17972), .A2(n1532), .ZN(n1531) );
  INV_X1 U5484 ( .A(n18667), .ZN(n18686) );
  NAND2_X1 U5485 ( .A1(n5393), .A2(n5322), .ZN(n5397) );
  NAND2_X1 U5486 ( .A1(n1536), .A2(n4614), .ZN(n1533) );
  NAND2_X1 U5487 ( .A1(n1538), .A2(n7746), .ZN(n2497) );
  NAND2_X1 U5488 ( .A1(n1540), .A2(n1539), .ZN(n1538) );
  NAND2_X1 U5489 ( .A1(n7749), .A2(n7750), .ZN(n1539) );
  INV_X1 U5490 ( .A(n7691), .ZN(n1541) );
  NAND2_X1 U5491 ( .A1(n9150), .A2(n9149), .ZN(n1543) );
  OAI21_X1 U5492 ( .B1(n8338), .B2(n2499), .A(n9145), .ZN(n1544) );
  INV_X1 U5493 ( .A(n7507), .ZN(n3445) );
  NAND3_X1 U5495 ( .A1(n1549), .A2(n7912), .A3(n1548), .ZN(n7913) );
  NAND2_X1 U5496 ( .A1(n7910), .A2(n3445), .ZN(n1549) );
  NOR2_X1 U5500 ( .A1(n1552), .A2(n14666), .ZN(n14669) );
  OAI21_X1 U5501 ( .B1(n2676), .B2(n1552), .A(n1551), .ZN(n2675) );
  NAND2_X1 U5502 ( .A1(n1552), .A2(n14662), .ZN(n1551) );
  AOI21_X1 U5503 ( .B1(n14536), .B2(n13164), .A(n1552), .ZN(n14537) );
  NAND2_X1 U5504 ( .A1(n15563), .A2(n3822), .ZN(n1553) );
  NAND2_X1 U5505 ( .A1(n15211), .A2(n15562), .ZN(n1554) );
  NAND2_X1 U5506 ( .A1(n921), .A2(n15510), .ZN(n15211) );
  NAND2_X1 U5507 ( .A1(n1555), .A2(n15866), .ZN(n15859) );
  OAI21_X1 U5508 ( .B1(n1555), .B2(n15866), .A(n2655), .ZN(n15172) );
  INV_X1 U5509 ( .A(n15857), .ZN(n1555) );
  OR2_X1 U5510 ( .A1(n16787), .A2(n16025), .ZN(n1556) );
  NAND2_X1 U5511 ( .A1(n1558), .A2(n16786), .ZN(n1557) );
  NAND2_X1 U5512 ( .A1(n1559), .A2(n16784), .ZN(n1558) );
  NAND2_X1 U5513 ( .A1(n1560), .A2(n8014), .ZN(n7827) );
  NOR2_X1 U5514 ( .A1(n1560), .A2(n20154), .ZN(n7086) );
  NAND2_X1 U5515 ( .A1(n7077), .A2(n1560), .ZN(n7107) );
  NAND2_X1 U5516 ( .A1(n5367), .A2(n1562), .ZN(n1561) );
  NOR2_X1 U5517 ( .A1(n5323), .A2(n5368), .ZN(n1562) );
  NAND3_X1 U5518 ( .A1(n4019), .A2(n5401), .A3(n1564), .ZN(n1563) );
  NAND2_X1 U5519 ( .A1(n5367), .A2(n5393), .ZN(n1564) );
  NAND3_X1 U5520 ( .A1(n15061), .A2(n15306), .A3(n1640), .ZN(n14187) );
  NAND2_X1 U5521 ( .A1(n8358), .A2(n1565), .ZN(n7696) );
  NAND2_X1 U5522 ( .A1(n8357), .A2(n1565), .ZN(n2931) );
  INV_X1 U5523 ( .A(n7741), .ZN(n1565) );
  INV_X1 U5524 ( .A(n4479), .ZN(n3967) );
  NAND2_X1 U5525 ( .A1(n4919), .A2(n1793), .ZN(n4239) );
  NAND2_X1 U5527 ( .A1(n1567), .A2(n9023), .ZN(n9024) );
  NAND2_X1 U5528 ( .A1(n8841), .A2(n1567), .ZN(n8839) );
  NAND2_X1 U5529 ( .A1(n1632), .A2(n1566), .ZN(n8587) );
  OR2_X1 U5530 ( .A1(n8836), .A2(n1567), .ZN(n1566) );
  NAND2_X1 U5531 ( .A1(n4721), .A2(n1569), .ZN(n5728) );
  NAND2_X2 U5532 ( .A1(n4704), .A2(n4703), .ZN(n6379) );
  INV_X1 U5533 ( .A(n14327), .ZN(n14350) );
  INV_X1 U5534 ( .A(n14819), .ZN(n1571) );
  NOR2_X1 U5535 ( .A1(n14353), .A2(n3444), .ZN(n1572) );
  NAND2_X1 U5536 ( .A1(n1574), .A2(n9090), .ZN(n8886) );
  INV_X1 U5539 ( .A(n9453), .ZN(n1576) );
  NAND2_X1 U5540 ( .A1(n8562), .A2(n1577), .ZN(n9454) );
  NAND2_X1 U5541 ( .A1(n11953), .A2(n11598), .ZN(n11599) );
  OAI21_X1 U5542 ( .B1(n10953), .B2(n11009), .A(n1579), .ZN(n9552) );
  NAND2_X1 U5543 ( .A1(n11009), .A2(n11149), .ZN(n1579) );
  INV_X1 U5544 ( .A(n10953), .ZN(n1580) );
  INV_X1 U5545 ( .A(Plaintext[76]), .ZN(n1581) );
  MUX2_X1 U5547 ( .A(n5024), .B(n19788), .S(n5022), .Z(n5028) );
  MUX2_X1 U5548 ( .A(n8824), .B(n8825), .S(n9313), .Z(n8826) );
  AND2_X1 U5552 ( .A1(n4217), .A2(n4219), .ZN(n1586) );
  NOR2_X1 U5553 ( .A1(n5826), .A2(n3569), .ZN(n1585) );
  NAND2_X1 U5554 ( .A1(n5823), .A2(n1585), .ZN(n3568) );
  NAND3_X1 U5555 ( .A1(n7866), .A2(n1587), .A3(n9264), .ZN(n8454) );
  MUX2_X1 U5556 ( .A(n9262), .B(n7866), .S(n9266), .Z(n8983) );
  NAND2_X1 U5557 ( .A1(n10876), .A2(n1588), .ZN(n10877) );
  NOR2_X1 U5558 ( .A1(n1591), .A2(n1589), .ZN(n1588) );
  NAND2_X1 U5559 ( .A1(n11633), .A2(n19755), .ZN(n1589) );
  NAND2_X1 U5560 ( .A1(n14248), .A2(n20377), .ZN(n2790) );
  INV_X1 U5561 ( .A(n4574), .ZN(n4371) );
  NAND2_X1 U5562 ( .A1(n12208), .A2(n11808), .ZN(n10821) );
  INV_X1 U5563 ( .A(n14656), .ZN(n1593) );
  NAND3_X1 U5564 ( .A1(n5096), .A2(n5098), .A3(n4788), .ZN(n1595) );
  NAND2_X1 U5565 ( .A1(n5097), .A2(n5096), .ZN(n1594) );
  NAND2_X1 U5566 ( .A1(n20202), .A2(n5088), .ZN(n1596) );
  XNOR2_X2 U5567 ( .A(Key[110]), .B(Plaintext[110]), .ZN(n5088) );
  NAND2_X1 U5568 ( .A1(n1598), .A2(n2460), .ZN(n1597) );
  NAND2_X1 U5569 ( .A1(n2461), .A2(n5094), .ZN(n1598) );
  INV_X1 U5570 ( .A(n10677), .ZN(n1601) );
  INV_X1 U5572 ( .A(n9221), .ZN(n1603) );
  NAND2_X1 U5573 ( .A1(n1603), .A2(n1604), .ZN(n8226) );
  INV_X1 U5574 ( .A(n9217), .ZN(n1604) );
  NAND3_X1 U5575 ( .A1(n5172), .A2(n5657), .A3(n6105), .ZN(n2558) );
  NAND2_X1 U5576 ( .A1(n11093), .A2(n11445), .ZN(n1606) );
  OAI21_X1 U5577 ( .B1(n11093), .B2(n10845), .A(n1606), .ZN(n10727) );
  AOI21_X1 U5578 ( .B1(n1606), .B2(n11444), .A(n19920), .ZN(n11450) );
  NAND2_X1 U5579 ( .A1(n8271), .A2(n1607), .ZN(n7720) );
  NAND2_X1 U5580 ( .A1(n1608), .A2(n8141), .ZN(n2156) );
  NAND3_X1 U5583 ( .A1(n11509), .A2(n10935), .A3(n259), .ZN(n10908) );
  MUX2_X1 U5584 ( .A(n10937), .B(n259), .S(n19864), .Z(n10938) );
  INV_X1 U5586 ( .A(n14935), .ZN(n1614) );
  NAND2_X1 U5588 ( .A1(n15188), .A2(n1611), .ZN(n1610) );
  AND2_X1 U5589 ( .A1(n15503), .A2(n15822), .ZN(n1611) );
  NAND2_X1 U5591 ( .A1(n15504), .A2(n15505), .ZN(n1615) );
  NAND2_X1 U5593 ( .A1(n1620), .A2(n5660), .ZN(n1619) );
  NAND2_X1 U5594 ( .A1(n6111), .A2(n6109), .ZN(n1621) );
  NAND2_X1 U5595 ( .A1(n5658), .A2(n5657), .ZN(n1622) );
  NAND2_X1 U5596 ( .A1(n5659), .A2(n6105), .ZN(n1623) );
  OAI21_X1 U5597 ( .B1(n14303), .B2(n14481), .A(n14434), .ZN(n1628) );
  NAND2_X1 U5598 ( .A1(n14311), .A2(n237), .ZN(n1624) );
  NAND2_X1 U5599 ( .A1(n14310), .A2(n14522), .ZN(n1625) );
  OAI22_X1 U5600 ( .A1(n15553), .A2(n1626), .B1(n14978), .B2(n15413), .ZN(
        n14907) );
  NAND2_X1 U5601 ( .A1(n15413), .A2(n15551), .ZN(n1626) );
  NAND2_X1 U5602 ( .A1(n1628), .A2(n1627), .ZN(n15409) );
  NAND2_X1 U5603 ( .A1(n1629), .A2(n14487), .ZN(n1627) );
  NAND2_X1 U5604 ( .A1(n14302), .A2(n14482), .ZN(n1629) );
  INV_X1 U5605 ( .A(n15551), .ZN(n14905) );
  NAND2_X1 U5606 ( .A1(n1632), .A2(n19857), .ZN(n1630) );
  INV_X1 U5607 ( .A(n8672), .ZN(n1632) );
  NAND2_X1 U5608 ( .A1(n8515), .A2(n1632), .ZN(n2024) );
  MUX2_X1 U5609 ( .A(n1632), .B(n9024), .S(n19857), .Z(n9025) );
  NAND2_X1 U5610 ( .A1(n249), .A2(n12352), .ZN(n1633) );
  NOR2_X2 U5611 ( .A1(n1635), .A2(n1634), .ZN(n13070) );
  NOR2_X1 U5612 ( .A1(n11032), .A2(n1637), .ZN(n1636) );
  INV_X1 U5613 ( .A(n19769), .ZN(n1637) );
  INV_X1 U5614 ( .A(n1638), .ZN(n13414) );
  NAND2_X1 U5615 ( .A1(n2902), .A2(n2905), .ZN(n1638) );
  NAND2_X1 U5616 ( .A1(n1638), .A2(n15221), .ZN(n15770) );
  NAND2_X1 U5617 ( .A1(n1639), .A2(n15666), .ZN(n15668) );
  AND2_X1 U5618 ( .A1(n234), .A2(n1638), .ZN(n15664) );
  NAND2_X1 U5619 ( .A1(n15772), .A2(n1638), .ZN(n15774) );
  AOI22_X2 U5620 ( .A1(n3254), .A2(n14369), .B1(n3253), .B2(n3299), .ZN(n1640)
         );
  NAND2_X1 U5621 ( .A1(n1640), .A2(n15309), .ZN(n14177) );
  OR2_X1 U5622 ( .A1(n15310), .A2(n1640), .ZN(n14188) );
  NAND3_X1 U5623 ( .A1(n3649), .A2(n12685), .A3(n12647), .ZN(n1641) );
  INV_X1 U5624 ( .A(n14731), .ZN(n14726) );
  XNOR2_X2 U5625 ( .A(n13402), .B(n13401), .ZN(n14731) );
  NAND2_X1 U5626 ( .A1(n255), .A2(n1643), .ZN(n12132) );
  NAND2_X1 U5627 ( .A1(n15498), .A2(n15497), .ZN(n1644) );
  NOR2_X1 U5628 ( .A1(n19512), .A2(n15195), .ZN(n15498) );
  NAND3_X1 U5629 ( .A1(n1647), .A2(n1649), .A3(n19512), .ZN(n1645) );
  NAND4_X1 U5630 ( .A1(n15508), .A2(n15821), .A3(n15820), .A4(n1646), .ZN(
        n16374) );
  NAND3_X1 U5631 ( .A1(n15822), .A2(n13933), .A3(n1758), .ZN(n1646) );
  NAND2_X1 U5632 ( .A1(n15192), .A2(n15501), .ZN(n1647) );
  NAND2_X1 U5633 ( .A1(n15499), .A2(n15500), .ZN(n1649) );
  NAND2_X1 U5634 ( .A1(n3819), .A2(n15501), .ZN(n1650) );
  NAND3_X2 U5635 ( .A1(n6402), .A2(n3808), .A3(n6401), .ZN(n9453) );
  NAND2_X1 U5636 ( .A1(n1652), .A2(n1576), .ZN(n1651) );
  NAND2_X1 U5638 ( .A1(n10650), .A2(n20516), .ZN(n8400) );
  MUX2_X1 U5639 ( .A(n11161), .B(n10649), .S(n20516), .Z(n10652) );
  MUX2_X1 U5640 ( .A(n10945), .B(n11159), .S(n11155), .Z(n9557) );
  NOR2_X1 U5641 ( .A1(n19872), .A2(n20516), .ZN(n9556) );
  OAI211_X2 U5642 ( .C1(n15133), .C2(n19848), .A(n2105), .B(n1655), .ZN(n16893) );
  NAND2_X1 U5643 ( .A1(n1656), .A2(n15132), .ZN(n1655) );
  NAND2_X1 U5644 ( .A1(n9010), .A2(n19490), .ZN(n1658) );
  NAND2_X1 U5645 ( .A1(n9006), .A2(n8895), .ZN(n9010) );
  XNOR2_X1 U5647 ( .A(n1659), .B(n2423), .ZN(Ciphertext[30]) );
  NAND2_X1 U5648 ( .A1(n18518), .A2(n19773), .ZN(n18505) );
  NAND2_X1 U5649 ( .A1(n1662), .A2(n18505), .ZN(n1661) );
  NAND2_X1 U5650 ( .A1(n18504), .A2(n20492), .ZN(n1662) );
  NAND2_X1 U5651 ( .A1(n11091), .A2(n11090), .ZN(n1663) );
  NAND2_X1 U5652 ( .A1(n11086), .A2(n11110), .ZN(n1664) );
  NAND2_X1 U5653 ( .A1(n1665), .A2(n289), .ZN(n4871) );
  NAND2_X1 U5654 ( .A1(n4381), .A2(n4866), .ZN(n1665) );
  INV_X1 U5655 ( .A(n4864), .ZN(n4865) );
  XNOR2_X2 U5657 ( .A(n1666), .B(n1667), .ZN(n14148) );
  XNOR2_X1 U5658 ( .A(n13754), .B(n13753), .ZN(n1666) );
  XNOR2_X1 U5659 ( .A(n13758), .B(n13759), .ZN(n1667) );
  NAND2_X1 U5660 ( .A1(n19154), .A2(n19708), .ZN(n1668) );
  NAND2_X1 U5663 ( .A1(n10970), .A2(n11553), .ZN(n3488) );
  OR2_X1 U5664 ( .A1(n18498), .A2(n18497), .ZN(n1675) );
  NAND3_X1 U5665 ( .A1(n16257), .A2(n16256), .A3(n1674), .ZN(n16259) );
  OAI211_X1 U5666 ( .C1(n1676), .C2(n17640), .A(n18500), .B(n1675), .ZN(n1674)
         );
  INV_X1 U5667 ( .A(n18498), .ZN(n1676) );
  NAND2_X1 U5668 ( .A1(n7691), .A2(n7746), .ZN(n1677) );
  NAND2_X1 U5669 ( .A1(n3447), .A2(n7750), .ZN(n1678) );
  AOI21_X1 U5670 ( .B1(n11418), .B2(n10829), .A(n1680), .ZN(n3046) );
  INV_X1 U5671 ( .A(n11131), .ZN(n1680) );
  NAND2_X1 U5672 ( .A1(n1681), .A2(n990), .ZN(n11423) );
  NAND2_X1 U5673 ( .A1(n11418), .A2(n11051), .ZN(n1681) );
  INV_X1 U5674 ( .A(n15754), .ZN(n1683) );
  NAND2_X1 U5676 ( .A1(n15589), .A2(n14039), .ZN(n1682) );
  NAND2_X1 U5677 ( .A1(n1683), .A2(n15758), .ZN(n15589) );
  NAND2_X1 U5679 ( .A1(n1686), .A2(n14288), .ZN(n14024) );
  INV_X1 U5680 ( .A(n14659), .ZN(n1686) );
  NAND2_X1 U5681 ( .A1(n199), .A2(n20266), .ZN(n14659) );
  INV_X1 U5682 ( .A(n14547), .ZN(n14023) );
  NAND2_X1 U5683 ( .A1(n2467), .A2(n6046), .ZN(n1687) );
  NAND2_X1 U5684 ( .A1(n12634), .A2(n180), .ZN(n1688) );
  NAND2_X1 U5685 ( .A1(n12633), .A2(n12634), .ZN(n1689) );
  NOR2_X2 U5686 ( .A1(n8796), .A2(n8793), .ZN(n9218) );
  OAI21_X1 U5687 ( .B1(n8176), .B2(n19901), .A(n1691), .ZN(n1690) );
  NAND2_X1 U5688 ( .A1(n1692), .A2(n19901), .ZN(n1691) );
  INV_X1 U5689 ( .A(n8178), .ZN(n1692) );
  NAND2_X1 U5690 ( .A1(n282), .A2(n8157), .ZN(n8256) );
  XNOR2_X1 U5691 ( .A(n1694), .B(n6840), .ZN(n1693) );
  XNOR2_X1 U5692 ( .A(n6842), .B(n6843), .ZN(n1694) );
  NAND2_X1 U5693 ( .A1(n1695), .A2(n5743), .ZN(n5203) );
  AOI21_X1 U5694 ( .B1(n1695), .B2(n5749), .A(n5743), .ZN(n5180) );
  NOR2_X1 U5695 ( .A1(n15645), .A2(n15256), .ZN(n15258) );
  NAND2_X1 U5696 ( .A1(n1699), .A2(n20266), .ZN(n1696) );
  NAND2_X1 U5697 ( .A1(n1698), .A2(n14653), .ZN(n1697) );
  NAND2_X1 U5698 ( .A1(n14653), .A2(n14656), .ZN(n3281) );
  NAND2_X1 U5700 ( .A1(n18425), .A2(n19997), .ZN(n2545) );
  NOR2_X1 U5701 ( .A1(n18427), .A2(n19997), .ZN(n18415) );
  NAND2_X1 U5702 ( .A1(n18427), .A2(n19997), .ZN(n18404) );
  OAI21_X1 U5703 ( .B1(n18412), .B2(n19997), .A(n18425), .ZN(n16491) );
  NAND2_X1 U5704 ( .A1(n18406), .A2(n1701), .ZN(n18408) );
  AND2_X1 U5705 ( .A1(n9532), .A2(n1703), .ZN(n1704) );
  NAND3_X1 U5706 ( .A1(n8592), .A2(n9531), .A3(n9358), .ZN(n1703) );
  NAND2_X1 U5707 ( .A1(n9533), .A2(n1704), .ZN(n9534) );
  NAND2_X1 U5708 ( .A1(n1706), .A2(n5529), .ZN(n1705) );
  NAND2_X1 U5709 ( .A1(n5562), .A2(n1707), .ZN(n1706) );
  NAND2_X1 U5710 ( .A1(n5563), .A2(n5569), .ZN(n1707) );
  NAND2_X1 U5711 ( .A1(n6036), .A2(n5532), .ZN(n6035) );
  NAND2_X1 U5712 ( .A1(n5562), .A2(n5563), .ZN(n6037) );
  NAND2_X1 U5713 ( .A1(n10958), .A2(n11145), .ZN(n1710) );
  NAND2_X1 U5714 ( .A1(n10959), .A2(n1721), .ZN(n1711) );
  AOI21_X1 U5715 ( .B1(n3486), .B2(n17236), .A(n19374), .ZN(n1712) );
  NAND2_X1 U5716 ( .A1(n1716), .A2(n1715), .ZN(n1714) );
  NAND2_X1 U5717 ( .A1(n18077), .A2(n20111), .ZN(n1715) );
  NAND2_X1 U5718 ( .A1(n2794), .A2(n1717), .ZN(n1716) );
  INV_X1 U5719 ( .A(n18394), .ZN(n1717) );
  OAI22_X1 U5720 ( .A1(n17241), .A2(n19823), .B1(n812), .B2(n20354), .ZN(
        n17242) );
  NOR2_X1 U5721 ( .A1(n17243), .A2(n1718), .ZN(n16463) );
  NAND2_X1 U5722 ( .A1(n20354), .A2(n19823), .ZN(n16461) );
  NAND2_X1 U5723 ( .A1(n19823), .A2(n17245), .ZN(n18541) );
  AND3_X1 U5724 ( .A1(n17480), .A2(n17479), .A3(n1718), .ZN(n17481) );
  MUX2_X1 U5725 ( .A(n20354), .B(n17480), .S(n1718), .Z(n16809) );
  INV_X1 U5726 ( .A(n5879), .ZN(n5980) );
  NAND2_X1 U5727 ( .A1(n5320), .A2(n6068), .ZN(n5879) );
  INV_X1 U5728 ( .A(n11145), .ZN(n1721) );
  NAND2_X1 U5729 ( .A1(n14442), .A2(n14168), .ZN(n1724) );
  NAND3_X1 U5730 ( .A1(n1726), .A2(n7978), .A3(n7981), .ZN(n6318) );
  NAND2_X1 U5731 ( .A1(n1730), .A2(n18078), .ZN(n1729) );
  NAND3_X1 U5732 ( .A1(n1732), .A2(n18376), .A3(n1733), .ZN(n1730) );
  NAND2_X1 U5733 ( .A1(n19763), .A2(n20361), .ZN(n1732) );
  NAND2_X1 U5734 ( .A1(n11586), .A2(n12128), .ZN(n11759) );
  NAND2_X1 U5735 ( .A1(n11642), .A2(n1734), .ZN(n11644) );
  AND2_X1 U5736 ( .A1(n11586), .A2(n12126), .ZN(n1734) );
  NAND3_X1 U5737 ( .A1(n11642), .A2(n11586), .A3(n882), .ZN(n11643) );
  NAND3_X1 U5738 ( .A1(n2499), .A2(n8786), .A3(n9145), .ZN(n1736) );
  NAND2_X1 U5739 ( .A1(n1740), .A2(n3281), .ZN(n1739) );
  NAND2_X1 U5740 ( .A1(n1742), .A2(n14023), .ZN(n1741) );
  NAND2_X1 U5741 ( .A1(n3281), .A2(n3280), .ZN(n1742) );
  NAND2_X1 U5742 ( .A1(n13221), .A2(n1744), .ZN(n1743) );
  NAND2_X1 U5743 ( .A1(n5844), .A2(n1746), .ZN(n5850) );
  NAND3_X1 U5744 ( .A1(n11142), .A2(n20366), .A3(n10960), .ZN(n1747) );
  NAND2_X1 U5746 ( .A1(n1749), .A2(n11145), .ZN(n1748) );
  XNOR2_X2 U5747 ( .A(n9505), .B(n9504), .ZN(n11145) );
  INV_X1 U5749 ( .A(n8823), .ZN(n1751) );
  NAND3_X1 U5750 ( .A1(n9307), .A2(n9313), .A3(n1754), .ZN(n1753) );
  NAND2_X1 U5752 ( .A1(n12500), .A2(n12499), .ZN(n12347) );
  AND2_X1 U5753 ( .A1(n1763), .A2(n1762), .ZN(n14308) );
  NAND2_X1 U5754 ( .A1(n14307), .A2(n13868), .ZN(n1763) );
  NAND2_X1 U5755 ( .A1(n1764), .A2(n5115), .ZN(n4838) );
  OAI21_X1 U5756 ( .B1(n169), .B2(n2042), .A(n4417), .ZN(n1764) );
  NAND2_X1 U5757 ( .A1(n8380), .A2(n8132), .ZN(n8389) );
  NAND2_X1 U5758 ( .A1(n8829), .A2(n9029), .ZN(n1765) );
  NAND2_X1 U5760 ( .A1(n5826), .A2(n3569), .ZN(n1832) );
  NAND2_X1 U5762 ( .A1(n4235), .A2(n4234), .ZN(n1769) );
  NAND2_X1 U5763 ( .A1(n4236), .A2(n4905), .ZN(n1768) );
  OAI21_X1 U5764 ( .B1(n5621), .B2(n6129), .A(n1770), .ZN(n5262) );
  NAND2_X1 U5766 ( .A1(n1774), .A2(n1773), .ZN(n1772) );
  INV_X1 U5767 ( .A(n19302), .ZN(n1773) );
  MUX2_X1 U5768 ( .A(n19292), .B(n19284), .S(n19299), .Z(n1774) );
  NAND2_X1 U5769 ( .A1(n19912), .A2(n1776), .ZN(n4181) );
  NAND2_X1 U5770 ( .A1(n1776), .A2(n5796), .ZN(n5793) );
  OAI22_X1 U5771 ( .A1(n5301), .A2(n5791), .B1(n5428), .B2(n1776), .ZN(n4184)
         );
  NAND2_X1 U5773 ( .A1(n1778), .A2(n19663), .ZN(n8714) );
  OAI21_X1 U5775 ( .B1(n11769), .B2(n1779), .A(n12288), .ZN(n11465) );
  INV_X1 U5776 ( .A(n182), .ZN(n1779) );
  XNOR2_X1 U5777 ( .A(n15739), .B(n1780), .ZN(n16094) );
  AND3_X2 U5778 ( .A1(n15278), .A2(n15279), .A3(n15280), .ZN(n15739) );
  XNOR2_X1 U5779 ( .A(n15739), .B(n1781), .ZN(n16689) );
  XNOR2_X1 U5780 ( .A(n15739), .B(n1782), .ZN(n15291) );
  XNOR2_X1 U5781 ( .A(n15739), .B(n1783), .ZN(n16907) );
  XNOR2_X1 U5782 ( .A(n15739), .B(n2417), .ZN(n17412) );
  NAND2_X1 U5783 ( .A1(n19521), .A2(n1785), .ZN(n1784) );
  XNOR2_X1 U5784 ( .A(n1786), .B(n13570), .ZN(n13402) );
  INV_X1 U5785 ( .A(n13428), .ZN(n1786) );
  XNOR2_X1 U5786 ( .A(n1787), .B(n13428), .ZN(n11901) );
  INV_X1 U5787 ( .A(n11862), .ZN(n1787) );
  NAND2_X1 U5788 ( .A1(n11480), .A2(n1788), .ZN(n2897) );
  NAND3_X1 U5791 ( .A1(n20206), .A2(n15121), .A3(n14514), .ZN(n1790) );
  INV_X1 U5792 ( .A(n8232), .ZN(n1791) );
  NAND2_X1 U5794 ( .A1(n4966), .A2(n3593), .ZN(n1792) );
  NAND2_X1 U5795 ( .A1(n1793), .A2(n4482), .ZN(n4966) );
  INV_X1 U5796 ( .A(n4479), .ZN(n1793) );
  NOR2_X1 U5797 ( .A1(n14450), .A2(n14449), .ZN(n1795) );
  XNOR2_X2 U5799 ( .A(n12867), .B(n12866), .ZN(n14450) );
  AOI22_X2 U5800 ( .A1(n1794), .A2(n14179), .B1(n14450), .B2(n13560), .ZN(
        n15237) );
  AND2_X1 U5801 ( .A1(n19510), .A2(n18682), .ZN(n18669) );
  AND2_X1 U5802 ( .A1(n18688), .A2(n18682), .ZN(n1796) );
  NAND2_X1 U5803 ( .A1(n19510), .A2(n1796), .ZN(n1800) );
  XNOR2_X1 U5804 ( .A(n1797), .B(n17024), .ZN(Ciphertext[68]) );
  NAND3_X1 U5805 ( .A1(n1800), .A2(n1799), .A3(n1798), .ZN(n1797) );
  NAND2_X1 U5806 ( .A1(n18668), .A2(n19510), .ZN(n1798) );
  OAI21_X1 U5807 ( .B1(n5697), .B2(n19804), .A(n1801), .ZN(n5698) );
  NAND2_X1 U5808 ( .A1(n5699), .A2(n5968), .ZN(n1801) );
  NAND3_X1 U5809 ( .A1(n20272), .A2(n15121), .A3(n1802), .ZN(n15123) );
  AOI22_X1 U5810 ( .A1(n20206), .A2(n1802), .B1(n15121), .B2(n14520), .ZN(
        n14185) );
  MUX2_X1 U5811 ( .A(n14516), .B(n20206), .S(n15120), .Z(n14521) );
  MUX2_X1 U5812 ( .A(n14514), .B(n13562), .S(n15120), .Z(n13565) );
  INV_X1 U5814 ( .A(n6184), .ZN(n2865) );
  OR2_X1 U5815 ( .A1(n5846), .A2(n6184), .ZN(n1805) );
  NAND2_X1 U5816 ( .A1(n288), .A2(n6184), .ZN(n1806) );
  NAND2_X1 U5817 ( .A1(n13856), .A2(n954), .ZN(n14195) );
  NAND2_X1 U5820 ( .A1(n1807), .A2(n5717), .ZN(n3605) );
  NAND2_X1 U5821 ( .A1(n14355), .A2(n1808), .ZN(n13938) );
  NAND2_X1 U5822 ( .A1(n14419), .A2(n1808), .ZN(n3180) );
  NAND2_X1 U5823 ( .A1(n8811), .A2(n8813), .ZN(n9121) );
  NAND2_X1 U5824 ( .A1(n11114), .A2(n11458), .ZN(n11453) );
  INV_X1 U5825 ( .A(n11458), .ZN(n1812) );
  INV_X1 U5826 ( .A(n11110), .ZN(n11451) );
  MUX2_X1 U5827 ( .A(n11454), .B(n11088), .S(n11110), .Z(n1814) );
  NAND2_X1 U5828 ( .A1(n15885), .A2(n15335), .ZN(n1815) );
  NAND2_X1 U5829 ( .A1(n1817), .A2(n16016), .ZN(n1816) );
  AOI22_X1 U5830 ( .A1(n13968), .A2(n3473), .B1(n15334), .B2(n16009), .ZN(
        n1818) );
  INV_X1 U5831 ( .A(n14736), .ZN(n1819) );
  NAND2_X1 U5833 ( .A1(n14270), .A2(n1821), .ZN(n1820) );
  OR2_X1 U5834 ( .A1(n14569), .A2(n14736), .ZN(n1821) );
  NAND2_X1 U5835 ( .A1(n18327), .A2(n19168), .ZN(n18320) );
  NAND2_X1 U5836 ( .A1(n9326), .A2(n9331), .ZN(n1822) );
  OR2_X1 U5838 ( .A1(n954), .A2(n15313), .ZN(n11988) );
  XNOR2_X1 U5839 ( .A(n3787), .B(n9315), .ZN(n1823) );
  MUX2_X1 U5840 ( .A(n7976), .B(n7975), .S(n7974), .Z(n1825) );
  OAI21_X1 U5841 ( .B1(n12351), .B2(n19768), .A(n12350), .ZN(n12357) );
  NAND2_X1 U5842 ( .A1(n12755), .A2(n245), .ZN(n1827) );
  INV_X1 U5843 ( .A(n4034), .ZN(n2468) );
  NAND3_X1 U5845 ( .A1(n3164), .A2(n20363), .A3(n12537), .ZN(n11806) );
  NAND2_X1 U5846 ( .A1(n11547), .A2(n11548), .ZN(n10068) );
  NAND3_X1 U5847 ( .A1(n19530), .A2(n20424), .A3(n14020), .ZN(n15757) );
  NAND2_X1 U5848 ( .A1(n5824), .A2(n1832), .ZN(n5831) );
  OR2_X1 U5849 ( .A1(n6129), .A2(n5623), .ZN(n5694) );
  NAND2_X1 U5851 ( .A1(n317), .A2(n8937), .ZN(n8944) );
  NAND2_X1 U5852 ( .A1(n1834), .A2(n1833), .ZN(n7583) );
  NAND2_X1 U5853 ( .A1(n8297), .A2(n5941), .ZN(n1833) );
  NAND2_X1 U5855 ( .A1(n11395), .A2(n11297), .ZN(n10860) );
  NAND2_X1 U5856 ( .A1(n1837), .A2(n1836), .ZN(n5254) );
  NAND2_X1 U5857 ( .A1(n5401), .A2(n5323), .ZN(n1836) );
  NAND2_X1 U5858 ( .A1(n5393), .A2(n1838), .ZN(n1837) );
  NAND3_X1 U5859 ( .A1(n7716), .A2(n7687), .A3(n8131), .ZN(n1839) );
  OR2_X1 U5860 ( .A1(n4866), .A2(n4651), .ZN(n4870) );
  AND2_X1 U5861 ( .A1(n8291), .A2(n8292), .ZN(n3406) );
  NOR2_X1 U5862 ( .A1(n8381), .A2(n163), .ZN(n7714) );
  OR2_X1 U5864 ( .A1(n12207), .A2(n247), .ZN(n12188) );
  INV_X1 U5866 ( .A(n9580), .ZN(n9578) );
  NAND2_X1 U5867 ( .A1(n19519), .A2(n1841), .ZN(n9580) );
  XNOR2_X1 U5870 ( .A(n7040), .B(n1842), .ZN(n4939) );
  XNOR2_X1 U5871 ( .A(n4780), .B(n4781), .ZN(n1842) );
  XNOR2_X1 U5872 ( .A(n1843), .B(n18503), .ZN(Ciphertext[29]) );
  NAND2_X1 U5875 ( .A1(n7606), .A2(n8184), .ZN(n7892) );
  NAND2_X1 U5876 ( .A1(n2614), .A2(n2615), .ZN(n5982) );
  NAND2_X1 U5877 ( .A1(n19752), .A2(n15531), .ZN(n15082) );
  INV_X1 U5878 ( .A(n3241), .ZN(n12358) );
  NAND2_X1 U5879 ( .A1(n14516), .A2(n14321), .ZN(n13562) );
  NAND2_X1 U5880 ( .A1(n17518), .A2(n17517), .ZN(n17581) );
  XNOR2_X1 U5881 ( .A(n1845), .B(n18587), .ZN(Ciphertext[51]) );
  NAND3_X1 U5882 ( .A1(n3411), .A2(n18586), .A3(n18582), .ZN(n1845) );
  OAI21_X1 U5883 ( .B1(n5995), .B2(n5999), .A(n1846), .ZN(n5275) );
  NAND2_X1 U5884 ( .A1(n5995), .A2(n5998), .ZN(n1846) );
  NAND2_X1 U5885 ( .A1(n1371), .A2(n11722), .ZN(n3676) );
  NAND3_X1 U5886 ( .A1(n11284), .A2(n19779), .A3(n11282), .ZN(n1847) );
  NAND2_X1 U5887 ( .A1(n10999), .A2(n10947), .ZN(n1848) );
  XOR2_X1 U5888 ( .A(n10441), .B(n10299), .Z(n2900) );
  XNOR2_X1 U5889 ( .A(n13239), .B(n3237), .ZN(n13240) );
  NAND2_X1 U5891 ( .A1(n14578), .A2(n14740), .ZN(n1849) );
  NAND2_X2 U5893 ( .A1(n9078), .A2(n9079), .ZN(n10382) );
  NAND2_X1 U5894 ( .A1(n8180), .A2(n8179), .ZN(n1851) );
  NAND3_X1 U5896 ( .A1(n2931), .A2(n2932), .A3(n8359), .ZN(n2933) );
  XNOR2_X2 U5897 ( .A(Key[19]), .B(Plaintext[19]), .ZN(n4979) );
  NAND2_X1 U5898 ( .A1(n1853), .A2(n1852), .ZN(n10857) );
  NAND2_X1 U5899 ( .A1(n11329), .A2(n11330), .ZN(n1852) );
  OAI21_X1 U5903 ( .B1(n14401), .B2(n19908), .A(n14400), .ZN(n3047) );
  NAND3_X1 U5904 ( .A1(n12758), .A2(n3702), .A3(n1856), .ZN(n13002) );
  AOI22_X1 U5905 ( .A1(n12755), .A2(n12754), .B1(n12756), .B2(n12759), .ZN(
        n1856) );
  XOR2_X1 U5906 ( .A(n7305), .B(n6484), .Z(n1863) );
  NAND3_X2 U5907 ( .A1(n2798), .A2(n2802), .A3(n2801), .ZN(n17098) );
  NAND3_X1 U5908 ( .A1(n12813), .A2(n19626), .A3(n11803), .ZN(n3169) );
  NOR2_X1 U5909 ( .A1(n9137), .A2(n263), .ZN(n9138) );
  NOR2_X1 U5910 ( .A1(n15545), .A2(n15406), .ZN(n2799) );
  NAND2_X1 U5911 ( .A1(n4950), .A2(n4912), .ZN(n4909) );
  NAND2_X1 U5913 ( .A1(n1860), .A2(n1859), .ZN(n1858) );
  NAND2_X1 U5914 ( .A1(n201), .A2(n12502), .ZN(n1860) );
  NAND2_X1 U5915 ( .A1(n19775), .A2(n1862), .ZN(n18004) );
  INV_X1 U5916 ( .A(n15394), .ZN(n2968) );
  NAND2_X1 U5917 ( .A1(n7420), .A2(n2886), .ZN(n7873) );
  NAND3_X1 U5918 ( .A1(n20157), .A2(n1819), .A3(n14574), .ZN(n13263) );
  NAND2_X2 U5919 ( .A1(n2403), .A2(n1864), .ZN(n7296) );
  NAND2_X1 U5920 ( .A1(n5417), .A2(n5226), .ZN(n1864) );
  INV_X1 U5922 ( .A(n1866), .ZN(n1865) );
  NAND2_X1 U5923 ( .A1(n5842), .A2(n6166), .ZN(n1868) );
  NAND2_X1 U5925 ( .A1(n957), .A2(n5700), .ZN(n1870) );
  OAI21_X1 U5926 ( .B1(n5450), .B2(n5449), .A(n5971), .ZN(n1871) );
  NAND2_X1 U5927 ( .A1(n12010), .A2(n12364), .ZN(n12011) );
  NAND3_X2 U5930 ( .A1(n8393), .A2(n8394), .A3(n966), .ZN(n10236) );
  NAND2_X1 U5931 ( .A1(n12340), .A2(n11974), .ZN(n11824) );
  OAI211_X2 U5932 ( .C1(n14201), .C2(n1262), .A(n2790), .B(n1873), .ZN(n15071)
         );
  NAND2_X1 U5933 ( .A1(n14604), .A2(n20513), .ZN(n1873) );
  INV_X1 U5934 ( .A(n4347), .ZN(n4540) );
  INV_X1 U5935 ( .A(n10685), .ZN(n12101) );
  XNOR2_X2 U5936 ( .A(n3916), .B(Key[150]), .ZN(n4754) );
  INV_X1 U5938 ( .A(n12686), .ZN(n12647) );
  XNOR2_X1 U5939 ( .A(n1874), .B(n18405), .ZN(Ciphertext[12]) );
  NAND3_X1 U5940 ( .A1(n18403), .A2(n18402), .A3(n1875), .ZN(n1874) );
  XNOR2_X1 U5941 ( .A(n10411), .B(n10412), .ZN(n11129) );
  AOI21_X1 U5943 ( .B1(n19971), .B2(n12072), .A(n12601), .ZN(n2911) );
  INV_X1 U5944 ( .A(n12800), .ZN(n14342) );
  OAI22_X1 U5945 ( .A1(n14306), .A2(n14305), .B1(n19742), .B2(n1876), .ZN(
        n14309) );
  INV_X1 U5946 ( .A(n14729), .ZN(n14728) );
  INV_X1 U5947 ( .A(n5868), .ZN(n5386) );
  INV_X1 U5948 ( .A(n5116), .ZN(n1916) );
  OAI21_X1 U5950 ( .B1(n7968), .B2(n7927), .A(n7969), .ZN(n3386) );
  NAND2_X1 U5952 ( .A1(n12067), .A2(n1879), .ZN(n1878) );
  NAND2_X1 U5954 ( .A1(n1880), .A2(n8804), .ZN(n3501) );
  NAND2_X1 U5955 ( .A1(n2631), .A2(n9209), .ZN(n1880) );
  INV_X1 U5956 ( .A(n1903), .ZN(n1902) );
  NOR2_X2 U5957 ( .A1(n4001), .A2(n1881), .ZN(n7264) );
  AOI21_X1 U5958 ( .B1(n2616), .B2(n4000), .A(n3999), .ZN(n1881) );
  NAND2_X1 U5959 ( .A1(n2974), .A2(n15431), .ZN(n15084) );
  NAND2_X1 U5960 ( .A1(n3980), .A2(n2071), .ZN(n1882) );
  NAND2_X1 U5962 ( .A1(n4887), .A2(n4945), .ZN(n4116) );
  OR2_X1 U5964 ( .A1(n11884), .A2(n11120), .ZN(n11461) );
  NAND2_X1 U5966 ( .A1(n11495), .A2(n888), .ZN(n10729) );
  NAND3_X1 U5967 ( .A1(n5473), .A2(n5472), .A3(n6034), .ZN(n1886) );
  NAND2_X1 U5968 ( .A1(n1888), .A2(n1887), .ZN(n11085) );
  NAND2_X1 U5969 ( .A1(n11081), .A2(n11499), .ZN(n1887) );
  NAND2_X1 U5970 ( .A1(n11505), .A2(n11188), .ZN(n1888) );
  NAND2_X1 U5971 ( .A1(n6217), .A2(n1890), .ZN(n6970) );
  NAND2_X1 U5972 ( .A1(n6203), .A2(n1891), .ZN(n6217) );
  NAND2_X1 U5973 ( .A1(n10890), .A2(n11549), .ZN(n1893) );
  NAND2_X1 U5975 ( .A1(n6033), .A2(n2940), .ZN(n1895) );
  OAI211_X1 U5978 ( .C1(n3389), .C2(n20463), .A(n1896), .B(n17219), .ZN(n18344) );
  NAND2_X1 U5979 ( .A1(n19383), .A2(n1897), .ZN(n1896) );
  OR2_X1 U5980 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  NAND3_X1 U5981 ( .A1(n2174), .A2(n9333), .A3(n9330), .ZN(n9336) );
  NAND2_X1 U5982 ( .A1(n1939), .A2(n3313), .ZN(n1898) );
  NAND2_X1 U5985 ( .A1(n14846), .A2(n3573), .ZN(n1901) );
  XNOR2_X1 U5986 ( .A(n7348), .B(n7163), .ZN(n6744) );
  OR2_X1 U5987 ( .A1(n4355), .A2(n4313), .ZN(n1908) );
  NAND2_X1 U5988 ( .A1(n17888), .A2(n19947), .ZN(n1905) );
  NAND2_X1 U5989 ( .A1(n17889), .A2(n1907), .ZN(n1906) );
  NAND2_X1 U5991 ( .A1(n11199), .A2(n3051), .ZN(n3048) );
  NAND2_X1 U5992 ( .A1(n10730), .A2(n11493), .ZN(n11199) );
  NAND3_X1 U5994 ( .A1(n4361), .A2(n4358), .A3(n4547), .ZN(n4359) );
  NAND2_X1 U5995 ( .A1(n1910), .A2(n1909), .ZN(n7636) );
  NAND2_X1 U5996 ( .A1(n7634), .A2(n8212), .ZN(n1909) );
  NAND2_X1 U5998 ( .A1(n9119), .A2(n8328), .ZN(n1912) );
  AND3_X1 U5999 ( .A1(n12629), .A2(n11722), .A3(n11618), .ZN(n11621) );
  NAND2_X1 U6000 ( .A1(n4066), .A2(n1914), .ZN(n4067) );
  NAND2_X1 U6002 ( .A1(n11296), .A2(n2724), .ZN(n1918) );
  NAND2_X2 U6003 ( .A1(n3591), .A2(n3043), .ZN(n6206) );
  NAND2_X1 U6004 ( .A1(n1919), .A2(n2115), .ZN(n5264) );
  NAND3_X1 U6005 ( .A1(n5804), .A2(n6194), .A3(n5805), .ZN(n2868) );
  NAND2_X1 U6006 ( .A1(n8375), .A2(n8376), .ZN(n8369) );
  NAND3_X1 U6007 ( .A1(n9327), .A2(n262), .A3(n20008), .ZN(n9337) );
  NAND2_X1 U6008 ( .A1(n3265), .A2(n3872), .ZN(n1920) );
  NAND3_X2 U6009 ( .A1(n1922), .A2(n4443), .A3(n4444), .ZN(n6138) );
  NOR2_X1 U6011 ( .A1(n17899), .A2(n1923), .ZN(n17900) );
  NOR2_X1 U6012 ( .A1(n17897), .A2(n1924), .ZN(n1923) );
  NAND2_X1 U6013 ( .A1(n15148), .A2(n15874), .ZN(n1925) );
  NAND3_X1 U6014 ( .A1(n1926), .A2(n1005), .A3(n2742), .ZN(n11640) );
  NAND2_X1 U6015 ( .A1(n2743), .A2(n3692), .ZN(n1926) );
  NOR2_X1 U6018 ( .A1(n983), .A2(n2874), .ZN(n2873) );
  OAI21_X1 U6019 ( .B1(n8078), .B2(n3654), .A(n3653), .ZN(n8082) );
  OAI21_X1 U6020 ( .B1(n3041), .B2(n15412), .A(n14980), .ZN(n1968) );
  NAND2_X1 U6021 ( .A1(n11147), .A2(n11148), .ZN(n10708) );
  XNOR2_X1 U6022 ( .A(n13102), .B(n13101), .ZN(n3373) );
  XNOR2_X2 U6023 ( .A(n3856), .B(Key[95]), .ZN(n5098) );
  NOR2_X1 U6024 ( .A1(n8510), .A2(n9021), .ZN(n8674) );
  INV_X1 U6025 ( .A(n5612), .ZN(n6159) );
  INV_X1 U6026 ( .A(n2523), .ZN(n12409) );
  INV_X1 U6028 ( .A(n6300), .ZN(n7241) );
  INV_X1 U6029 ( .A(n3995), .ZN(n4687) );
  OAI21_X1 U6030 ( .B1(n10935), .B2(n19864), .A(n1928), .ZN(n10744) );
  NAND2_X1 U6031 ( .A1(n10935), .A2(n11573), .ZN(n1928) );
  NAND2_X1 U6036 ( .A1(n1015), .A2(n8841), .ZN(n1929) );
  OAI211_X2 U6037 ( .C1(n12381), .C2(n11732), .A(n1931), .B(n1930), .ZN(n13642) );
  NAND2_X1 U6038 ( .A1(n11731), .A2(n12381), .ZN(n1930) );
  NAND2_X1 U6039 ( .A1(n12371), .A2(n20497), .ZN(n1931) );
  MUX2_X1 U6040 ( .A(n9114), .B(n9221), .S(n9113), .Z(n9115) );
  OAI21_X1 U6041 ( .B1(n4646), .B2(n4647), .A(n4645), .ZN(n4649) );
  NAND2_X1 U6042 ( .A1(n4646), .A2(n4319), .ZN(n4645) );
  NAND2_X1 U6043 ( .A1(n12007), .A2(n12008), .ZN(n12012) );
  NAND2_X1 U6044 ( .A1(n1934), .A2(n1933), .ZN(n1932) );
  INV_X1 U6045 ( .A(n9046), .ZN(n1933) );
  INV_X1 U6046 ( .A(n9045), .ZN(n1934) );
  NAND2_X1 U6048 ( .A1(n1935), .A2(n13877), .ZN(n14496) );
  OAI21_X1 U6049 ( .B1(n14492), .B2(n14491), .A(n1936), .ZN(n1935) );
  NAND3_X1 U6050 ( .A1(n10661), .A2(n11244), .A3(n10662), .ZN(n2859) );
  NAND2_X1 U6051 ( .A1(n10856), .A2(n20095), .ZN(n10662) );
  XNOR2_X2 U6052 ( .A(Key[141]), .B(Plaintext[141]), .ZN(n4734) );
  AND2_X1 U6053 ( .A1(n4633), .A2(n4185), .ZN(n3728) );
  OAI211_X1 U6054 ( .C1(n14081), .C2(n20500), .A(n1937), .B(n3497), .ZN(n3496)
         );
  NAND2_X1 U6055 ( .A1(n1938), .A2(n14801), .ZN(n1937) );
  INV_X1 U6056 ( .A(n2628), .ZN(n1938) );
  NAND2_X1 U6058 ( .A1(n3385), .A2(n9046), .ZN(n9037) );
  INV_X1 U6059 ( .A(n4708), .ZN(n4771) );
  NOR2_X1 U6060 ( .A1(n19958), .A2(n3315), .ZN(n1939) );
  XNOR2_X1 U6061 ( .A(n1940), .B(n7213), .ZN(n7215) );
  XNOR2_X1 U6062 ( .A(n7210), .B(n7360), .ZN(n1940) );
  NAND2_X1 U6063 ( .A1(n19507), .A2(n4969), .ZN(n4480) );
  OR2_X1 U6064 ( .A1(n4908), .A2(n4907), .ZN(n1942) );
  NAND2_X1 U6065 ( .A1(n11111), .A2(n11114), .ZN(n1943) );
  NAND2_X1 U6066 ( .A1(n11112), .A2(n11454), .ZN(n1944) );
  NAND2_X1 U6067 ( .A1(n12387), .A2(n12470), .ZN(n1945) );
  NAND2_X1 U6068 ( .A1(n1948), .A2(n1947), .ZN(n6808) );
  NAND2_X1 U6069 ( .A1(n5215), .A2(n1949), .ZN(n1948) );
  NAND2_X1 U6070 ( .A1(n10710), .A2(n20160), .ZN(n10714) );
  AOI21_X1 U6071 ( .B1(n1950), .B2(n8217), .A(n8216), .ZN(n8224) );
  NAND2_X1 U6072 ( .A1(n8219), .A2(n8215), .ZN(n1950) );
  NAND3_X2 U6074 ( .A1(n1954), .A2(n11691), .A3(n1951), .ZN(n13193) );
  NAND2_X1 U6077 ( .A1(n12123), .A2(n12230), .ZN(n1954) );
  OAI211_X2 U6078 ( .C1(n19809), .C2(n8217), .A(n6475), .B(n6474), .ZN(n9240)
         );
  NOR2_X1 U6079 ( .A1(n15468), .A2(n15469), .ZN(n1955) );
  NAND2_X1 U6080 ( .A1(n4171), .A2(n20143), .ZN(n4288) );
  NAND3_X1 U6081 ( .A1(n151), .A2(n19037), .A3(n1016), .ZN(n19039) );
  OAI21_X1 U6082 ( .B1(n13275), .B2(n12325), .A(n1956), .ZN(n11678) );
  NAND2_X1 U6083 ( .A1(n13275), .A2(n12513), .ZN(n1956) );
  OAI21_X2 U6084 ( .B1(n6112), .B2(n6113), .A(n1957), .ZN(n7221) );
  NAND2_X1 U6085 ( .A1(n6110), .A2(n6109), .ZN(n1958) );
  INV_X1 U6086 ( .A(n7711), .ZN(n6952) );
  NAND2_X1 U6087 ( .A1(n6091), .A2(n6088), .ZN(n1959) );
  NAND2_X1 U6088 ( .A1(n2692), .A2(n2693), .ZN(n2691) );
  AND2_X1 U6089 ( .A1(n12417), .A2(n20352), .ZN(n12427) );
  INV_X1 U6092 ( .A(n16171), .ZN(n3573) );
  NAND2_X1 U6093 ( .A1(n1963), .A2(n1961), .ZN(n9242) );
  NAND2_X1 U6094 ( .A1(n6610), .A2(n8090), .ZN(n1963) );
  AND2_X1 U6097 ( .A1(n19472), .A2(n17946), .ZN(n17774) );
  OR2_X1 U6098 ( .A1(n7930), .A2(n7933), .ZN(n7941) );
  INV_X1 U6099 ( .A(n11211), .ZN(n11486) );
  AND3_X2 U6100 ( .A1(n1965), .A2(n8816), .A3(n1964), .ZN(n10404) );
  NAND2_X1 U6101 ( .A1(n8819), .A2(n8818), .ZN(n1965) );
  OAI21_X1 U6102 ( .B1(n12535), .B2(n3477), .A(n12531), .ZN(n3476) );
  XNOR2_X1 U6103 ( .A(n13136), .B(n20170), .ZN(n12517) );
  INV_X1 U6105 ( .A(n15127), .ZN(n15017) );
  INV_X1 U6106 ( .A(n6031), .ZN(n5928) );
  OAI211_X1 U6107 ( .C1(n14195), .C2(n2731), .A(n14194), .B(n14193), .ZN(
        n15615) );
  NOR2_X1 U6108 ( .A1(n15846), .A2(n15267), .ZN(n2529) );
  XNOR2_X1 U6110 ( .A(n3619), .B(n6719), .ZN(n7286) );
  XNOR2_X1 U6111 ( .A(n2520), .B(n2519), .ZN(n14012) );
  OR2_X1 U6112 ( .A1(n15277), .A2(n15601), .ZN(n15278) );
  XNOR2_X1 U6113 ( .A(n1966), .B(n18428), .ZN(Ciphertext[17]) );
  OAI22_X1 U6114 ( .A1(n2546), .A2(n18427), .B1(n18426), .B2(n18425), .ZN(
        n1966) );
  AOI21_X1 U6115 ( .B1(n8072), .B2(n2456), .A(n585), .ZN(n1967) );
  NAND2_X1 U6118 ( .A1(n12591), .A2(n12200), .ZN(n11978) );
  NAND2_X1 U6119 ( .A1(n1968), .A2(n3042), .ZN(n16944) );
  NAND3_X1 U6120 ( .A1(n20313), .A2(n8537), .A3(n9073), .ZN(n8464) );
  NAND2_X1 U6121 ( .A1(n11429), .A2(n1970), .ZN(n10827) );
  NAND2_X1 U6124 ( .A1(n11151), .A2(n11152), .ZN(n1971) );
  INV_X1 U6125 ( .A(n4510), .ZN(n4513) );
  INV_X1 U6126 ( .A(n11880), .ZN(n3441) );
  XNOR2_X1 U6127 ( .A(n13345), .B(n13346), .ZN(n1973) );
  NAND2_X1 U6128 ( .A1(n15860), .A2(n1974), .ZN(n15867) );
  NAND2_X1 U6129 ( .A1(n8263), .A2(n8153), .ZN(n8104) );
  OAI21_X1 U6131 ( .B1(n11976), .B2(n11977), .A(n2160), .ZN(n1975) );
  NAND2_X1 U6132 ( .A1(n6010), .A2(n19979), .ZN(n5502) );
  NAND2_X1 U6133 ( .A1(n5804), .A2(n5805), .ZN(n5808) );
  NAND2_X1 U6134 ( .A1(n3345), .A2(n17879), .ZN(n3344) );
  NAND2_X2 U6135 ( .A1(n2497), .A2(n7913), .ZN(n2499) );
  NAND2_X1 U6136 ( .A1(n4540), .A2(n4541), .ZN(n4543) );
  NAND2_X1 U6137 ( .A1(n3259), .A2(n5101), .ZN(n5103) );
  NAND3_X1 U6138 ( .A1(n7929), .A2(n9149), .A3(n7928), .ZN(n7943) );
  OAI21_X1 U6140 ( .B1(n5122), .B2(n5917), .A(n5916), .ZN(n1978) );
  INV_X1 U6141 ( .A(n11377), .ZN(n11329) );
  OAI211_X1 U6142 ( .C1(n8529), .C2(n9038), .A(n1979), .B(n7657), .ZN(n7658)
         );
  AOI22_X2 U6143 ( .A1(n11393), .A2(n11392), .B1(n19750), .B2(n11391), .ZN(
        n12545) );
  NOR2_X1 U6144 ( .A1(n3764), .A2(n3762), .ZN(n3761) );
  NOR2_X1 U6145 ( .A1(n3030), .A2(n18869), .ZN(n18051) );
  OR2_X1 U6148 ( .A1(n4171), .A2(n4622), .ZN(n4627) );
  NAND2_X1 U6149 ( .A1(n2291), .A2(n3316), .ZN(n1983) );
  OAI21_X1 U6150 ( .B1(n9451), .B2(n8884), .A(n8563), .ZN(n9455) );
  INV_X1 U6151 ( .A(n7931), .ZN(n2030) );
  INV_X1 U6152 ( .A(n10849), .ZN(n13114) );
  INV_X1 U6153 ( .A(n4355), .ZN(n4547) );
  AND2_X1 U6154 ( .A1(n5571), .A2(n5581), .ZN(n3533) );
  XNOR2_X2 U6155 ( .A(n3881), .B(Key[2]), .ZN(n4171) );
  NAND2_X1 U6156 ( .A1(n11674), .A2(n11670), .ZN(n11843) );
  NAND2_X1 U6157 ( .A1(n15745), .A2(n15521), .ZN(n14982) );
  NAND3_X1 U6158 ( .A1(n14486), .A2(n14302), .A3(n14480), .ZN(n13554) );
  NAND2_X1 U6159 ( .A1(n20263), .A2(n14482), .ZN(n14486) );
  NAND2_X1 U6160 ( .A1(n5804), .A2(n1986), .ZN(n5380) );
  AND2_X1 U6163 ( .A1(n11500), .A2(n11193), .ZN(n1988) );
  AND2_X1 U6164 ( .A1(n14673), .A2(n20424), .ZN(n13982) );
  INV_X1 U6165 ( .A(n7443), .ZN(n8280) );
  OR2_X2 U6166 ( .A1(n9195), .A2(n9194), .ZN(n10107) );
  NAND2_X1 U6168 ( .A1(n1989), .A2(n3660), .ZN(n3659) );
  INV_X1 U6170 ( .A(n2183), .ZN(n12564) );
  NAND2_X1 U6171 ( .A1(n1991), .A2(n1990), .ZN(n2183) );
  NAND2_X1 U6172 ( .A1(n12263), .A2(n12262), .ZN(n1990) );
  NAND2_X1 U6173 ( .A1(n12261), .A2(n12264), .ZN(n1991) );
  NAND2_X1 U6174 ( .A1(n14721), .A2(n1992), .ZN(n15566) );
  OR2_X1 U6175 ( .A1(n14723), .A2(n19843), .ZN(n1992) );
  OR2_X1 U6177 ( .A1(n4541), .A2(n4347), .ZN(n4254) );
  NAND2_X1 U6178 ( .A1(n1995), .A2(n1993), .ZN(n7677) );
  NAND2_X1 U6179 ( .A1(n7676), .A2(n1994), .ZN(n1993) );
  NAND2_X1 U6180 ( .A1(n8362), .A2(n7675), .ZN(n1995) );
  NAND2_X1 U6182 ( .A1(n15700), .A2(n20145), .ZN(n1997) );
  OAI21_X1 U6183 ( .B1(n14344), .B2(n14789), .A(n1999), .ZN(n14104) );
  NAND2_X1 U6184 ( .A1(n2411), .A2(n2412), .ZN(n1999) );
  OAI21_X1 U6185 ( .B1(n2001), .B2(n2000), .A(n18996), .ZN(n18998) );
  NAND2_X1 U6186 ( .A1(n18991), .A2(n18993), .ZN(n2000) );
  NAND2_X1 U6187 ( .A1(n18994), .A2(n18992), .ZN(n2001) );
  NAND2_X1 U6188 ( .A1(n14723), .A2(n14717), .ZN(n14719) );
  XNOR2_X2 U6189 ( .A(n6949), .B(n7270), .ZN(n8341) );
  NAND2_X1 U6190 ( .A1(n1062), .A2(n3818), .ZN(n2002) );
  NOR2_X1 U6191 ( .A1(n2813), .A2(n14461), .ZN(n2812) );
  NAND3_X1 U6192 ( .A1(n4593), .A2(n4594), .A3(n6194), .ZN(n4595) );
  OAI21_X1 U6194 ( .B1(n14939), .B2(n14940), .A(n20449), .ZN(n2006) );
  OAI21_X1 U6196 ( .B1(n15160), .B2(n15159), .A(n15195), .ZN(n2007) );
  NAND2_X1 U6198 ( .A1(n20180), .A2(n20441), .ZN(n8217) );
  NAND2_X1 U6199 ( .A1(n11417), .A2(n11129), .ZN(n11419) );
  NAND2_X1 U6200 ( .A1(n16580), .A2(n2008), .ZN(n19338) );
  OR2_X1 U6201 ( .A1(n16657), .A2(n19372), .ZN(n2008) );
  NAND2_X1 U6203 ( .A1(n2009), .A2(n11410), .ZN(n3612) );
  NAND2_X1 U6204 ( .A1(n11408), .A2(n19736), .ZN(n2009) );
  OAI21_X2 U6205 ( .B1(n3879), .B2(n2010), .A(n3878), .ZN(n5796) );
  NAND2_X1 U6206 ( .A1(n4980), .A2(n4978), .ZN(n2010) );
  NAND3_X1 U6210 ( .A1(n3626), .A2(n2013), .A3(n2011), .ZN(n13041) );
  NAND2_X1 U6211 ( .A1(n12120), .A2(n2012), .ZN(n2011) );
  INV_X1 U6212 ( .A(n12124), .ZN(n2012) );
  NAND2_X1 U6213 ( .A1(n12123), .A2(n12227), .ZN(n2013) );
  NAND2_X1 U6215 ( .A1(n19663), .A2(n2476), .ZN(n2015) );
  OAI21_X1 U6216 ( .B1(n1859), .B2(n12500), .A(n2016), .ZN(n2864) );
  NAND2_X1 U6217 ( .A1(n9189), .A2(n6656), .ZN(n2425) );
  NAND2_X1 U6218 ( .A1(n3846), .A2(n4676), .ZN(n5114) );
  OAI21_X1 U6219 ( .B1(n8466), .B2(n8545), .A(n2330), .ZN(n8468) );
  OAI22_X1 U6220 ( .A1(n2017), .A2(n8602), .B1(n8949), .B2(n8951), .ZN(n7652)
         );
  NAND2_X1 U6221 ( .A1(n8949), .A2(n905), .ZN(n2017) );
  XNOR2_X1 U6222 ( .A(n13253), .B(n13750), .ZN(n2189) );
  NAND3_X1 U6223 ( .A1(n12148), .A2(n3260), .A3(n19952), .ZN(n2104) );
  INV_X1 U6226 ( .A(n18424), .ZN(n2019) );
  XNOR2_X1 U6227 ( .A(n2020), .B(n10297), .ZN(n10302) );
  XNOR2_X1 U6228 ( .A(n10295), .B(n10612), .ZN(n2020) );
  MUX2_X1 U6229 ( .A(n8194), .B(n7456), .S(n8051), .Z(n2021) );
  NAND2_X1 U6231 ( .A1(n5115), .A2(n4676), .ZN(n3848) );
  OAI21_X1 U6233 ( .B1(n8215), .B2(n8219), .A(n2026), .ZN(n3793) );
  NAND2_X1 U6234 ( .A1(n8220), .A2(n8219), .ZN(n2026) );
  NAND2_X1 U6236 ( .A1(n2028), .A2(n2027), .ZN(n4266) );
  OAI21_X1 U6237 ( .B1(n4754), .B2(n4563), .A(n4567), .ZN(n2027) );
  NAND2_X1 U6238 ( .A1(n4265), .A2(n3131), .ZN(n2028) );
  NAND2_X1 U6239 ( .A1(n12004), .A2(n12005), .ZN(n2901) );
  INV_X1 U6240 ( .A(n5483), .ZN(n4363) );
  AOI21_X1 U6243 ( .B1(n11358), .B2(n11127), .A(n1039), .ZN(n2029) );
  NAND2_X1 U6244 ( .A1(n4687), .A2(n178), .ZN(n4392) );
  NAND3_X2 U6245 ( .A1(n2034), .A2(n4758), .A3(n3129), .ZN(n5669) );
  NOR2_X1 U6246 ( .A1(n3112), .A2(n11177), .ZN(n3111) );
  INV_X1 U6247 ( .A(n15644), .ZN(n2223) );
  INV_X1 U6249 ( .A(n18033), .ZN(n18268) );
  XNOR2_X1 U6251 ( .A(n10324), .B(n10323), .ZN(n11088) );
  INV_X1 U6252 ( .A(n15341), .ZN(n15337) );
  XNOR2_X2 U6253 ( .A(Key[33]), .B(Plaintext[33]), .ZN(n4912) );
  NAND2_X1 U6254 ( .A1(n5324), .A2(n5373), .ZN(n5325) );
  NAND2_X1 U6255 ( .A1(n1838), .A2(n5401), .ZN(n5373) );
  OAI21_X1 U6256 ( .B1(n2548), .B2(n7585), .A(n2037), .ZN(n3611) );
  NAND2_X1 U6257 ( .A1(n7312), .A2(n2548), .ZN(n2037) );
  NAND2_X1 U6258 ( .A1(n2040), .A2(n2038), .ZN(n14754) );
  NAND3_X1 U6259 ( .A1(n14054), .A2(n13938), .A3(n2039), .ZN(n2038) );
  NAND2_X1 U6260 ( .A1(n13941), .A2(n13940), .ZN(n2040) );
  OAI21_X1 U6261 ( .B1(n4675), .B2(n2042), .A(n2041), .ZN(n3842) );
  NAND2_X1 U6262 ( .A1(n4675), .A2(n4835), .ZN(n2041) );
  AOI21_X1 U6263 ( .B1(n11399), .B2(n11395), .A(n11397), .ZN(n2044) );
  NAND2_X1 U6266 ( .A1(n7645), .A2(n8221), .ZN(n7648) );
  XNOR2_X1 U6267 ( .A(n16885), .B(n16331), .ZN(n16332) );
  NOR2_X1 U6268 ( .A1(n9371), .A2(n2066), .ZN(n2065) );
  NAND2_X1 U6269 ( .A1(n3500), .A2(n11480), .ZN(n11487) );
  NAND3_X2 U6270 ( .A1(n14158), .A2(n2047), .A3(n3815), .ZN(n14159) );
  NAND2_X1 U6271 ( .A1(n14248), .A2(n20513), .ZN(n2047) );
  NAND3_X2 U6272 ( .A1(n7596), .A2(n7597), .A3(n7595), .ZN(n8937) );
  OAI21_X1 U6273 ( .B1(n5996), .B2(n6000), .A(n5995), .ZN(n2048) );
  NAND2_X1 U6274 ( .A1(n216), .A2(n3030), .ZN(n2049) );
  NAND2_X1 U6275 ( .A1(n5704), .A2(n5434), .ZN(n2051) );
  NAND2_X1 U6276 ( .A1(n2053), .A2(n1591), .ZN(n2052) );
  NAND2_X1 U6277 ( .A1(n12056), .A2(n12619), .ZN(n2054) );
  NAND2_X1 U6278 ( .A1(n11880), .A2(n11460), .ZN(n11879) );
  XNOR2_X2 U6279 ( .A(n10218), .B(n10217), .ZN(n11880) );
  NOR2_X1 U6280 ( .A1(n12201), .A2(n12594), .ZN(n2056) );
  NAND2_X1 U6281 ( .A1(n2059), .A2(n2057), .ZN(n19006) );
  NAND2_X1 U6282 ( .A1(n19724), .A2(n2058), .ZN(n2057) );
  NAND2_X1 U6283 ( .A1(n18999), .A2(n19013), .ZN(n2059) );
  NAND2_X1 U6284 ( .A1(n14490), .A2(n20453), .ZN(n13877) );
  NAND2_X1 U6285 ( .A1(n11206), .A2(n11094), .ZN(n2060) );
  NAND2_X1 U6286 ( .A1(n10846), .A2(n11203), .ZN(n2061) );
  NAND2_X1 U6288 ( .A1(n18940), .A2(n18936), .ZN(n18933) );
  NAND3_X1 U6290 ( .A1(n11327), .A2(n11255), .A3(n19886), .ZN(n10309) );
  OAI211_X2 U6292 ( .C1(n12875), .C2(n20502), .A(n2069), .B(n2068), .ZN(n17411) );
  NAND2_X1 U6293 ( .A1(n12874), .A2(n19888), .ZN(n2068) );
  NAND2_X1 U6294 ( .A1(n3979), .A2(n3978), .ZN(n2070) );
  NAND2_X1 U6295 ( .A1(n4420), .A2(n4220), .ZN(n3979) );
  INV_X1 U6296 ( .A(n3978), .ZN(n2071) );
  INV_X1 U6297 ( .A(n12544), .ZN(n12305) );
  NAND2_X1 U6298 ( .A1(n4866), .A2(n4865), .ZN(n2072) );
  AOI22_X1 U6300 ( .A1(n11405), .A2(n11404), .B1(n11406), .B2(n19506), .ZN(
        n2810) );
  NAND2_X1 U6301 ( .A1(n8583), .A2(n9298), .ZN(n2073) );
  NAND2_X1 U6302 ( .A1(n8584), .A2(n8846), .ZN(n2074) );
  XNOR2_X2 U6303 ( .A(n16056), .B(n16055), .ZN(n17876) );
  OAI21_X1 U6304 ( .B1(n988), .B2(n2075), .A(n18597), .ZN(n17626) );
  NOR2_X1 U6305 ( .A1(n17624), .A2(n19656), .ZN(n2075) );
  INV_X1 U6306 ( .A(n3588), .ZN(n11403) );
  NAND3_X1 U6307 ( .A1(n4146), .A2(n4645), .A3(n4325), .ZN(n2076) );
  NAND2_X1 U6308 ( .A1(n4016), .A2(n4642), .ZN(n2077) );
  OR2_X1 U6310 ( .A1(n3634), .A2(n3551), .ZN(n3550) );
  INV_X1 U6311 ( .A(n8074), .ZN(n3703) );
  INV_X1 U6312 ( .A(n4638), .ZN(n2919) );
  INV_X1 U6313 ( .A(Plaintext[143]), .ZN(n3153) );
  INV_X1 U6314 ( .A(n18774), .ZN(n18749) );
  XOR2_X1 U6315 ( .A(n10552), .B(n1969), .Z(n3424) );
  AOI22_X1 U6316 ( .A1(n4276), .A2(n5018), .B1(n5014), .B2(n4111), .ZN(n5276)
         );
  XNOR2_X1 U6317 ( .A(n9605), .B(n10549), .ZN(n2570) );
  XNOR2_X1 U6318 ( .A(n4247), .B(n4246), .ZN(n8060) );
  XNOR2_X1 U6319 ( .A(n13533), .B(n2078), .ZN(n13140) );
  XNOR2_X1 U6320 ( .A(n13137), .B(n13616), .ZN(n2078) );
  NAND2_X1 U6322 ( .A1(n19590), .A2(n9564), .ZN(n8703) );
  OR2_X2 U6323 ( .A1(n14459), .A2(n14458), .ZN(n15295) );
  NAND2_X1 U6324 ( .A1(n2441), .A2(n8384), .ZN(n8135) );
  NAND2_X1 U6325 ( .A1(n7684), .A2(n8380), .ZN(n8384) );
  NAND2_X1 U6326 ( .A1(n2081), .A2(n2080), .ZN(n5561) );
  NAND2_X1 U6327 ( .A1(n5557), .A2(n6048), .ZN(n2080) );
  NAND2_X1 U6329 ( .A1(n5010), .A2(n4204), .ZN(n4206) );
  NOR2_X1 U6330 ( .A1(n14768), .A2(n15107), .ZN(n14771) );
  AOI22_X1 U6331 ( .A1(n17581), .A2(n20433), .B1(n17582), .B2(n19773), .ZN(
        n17583) );
  AOI21_X1 U6332 ( .B1(n20618), .B2(n12147), .A(n3666), .ZN(n12314) );
  OAI211_X1 U6333 ( .C1(n14678), .C2(n20120), .A(n14279), .B(n14677), .ZN(
        n14683) );
  NAND3_X1 U6334 ( .A1(n19752), .A2(n15421), .A3(n15420), .ZN(n15083) );
  NAND2_X1 U6335 ( .A1(n12369), .A2(n12374), .ZN(n11856) );
  NAND2_X1 U6336 ( .A1(n893), .A2(n300), .ZN(n2084) );
  NAND2_X1 U6337 ( .A1(n17737), .A2(n18501), .ZN(n17739) );
  NAND3_X1 U6339 ( .A1(n14210), .A2(n2086), .A3(n2085), .ZN(n15070) );
  NAND2_X1 U6340 ( .A1(n14207), .A2(n14206), .ZN(n2085) );
  NAND2_X1 U6341 ( .A1(n14209), .A2(n14208), .ZN(n2086) );
  OAI22_X1 U6344 ( .A1(n15500), .A2(n15502), .B1(n15192), .B2(n15496), .ZN(
        n14042) );
  AND3_X2 U6345 ( .A1(n2088), .A2(n3173), .A3(n3172), .ZN(n15500) );
  NAND2_X1 U6347 ( .A1(n7890), .A2(n8190), .ZN(n2089) );
  OR2_X1 U6349 ( .A1(n4094), .A2(n4268), .ZN(n4582) );
  NAND2_X1 U6350 ( .A1(n2093), .A2(n2091), .ZN(n4436) );
  NAND2_X1 U6351 ( .A1(n2092), .A2(n6124), .ZN(n2091) );
  OR2_X1 U6352 ( .A1(n19921), .A2(n14690), .ZN(n2094) );
  XNOR2_X1 U6355 ( .A(n13850), .B(n13851), .ZN(n2095) );
  NAND3_X1 U6357 ( .A1(n1041), .A2(n9234), .A3(n2097), .ZN(n3059) );
  NAND2_X1 U6358 ( .A1(n2254), .A2(n2255), .ZN(n12644) );
  XNOR2_X1 U6359 ( .A(n13078), .B(n19904), .ZN(n2200) );
  XNOR2_X1 U6360 ( .A(n13154), .B(n13027), .ZN(n13078) );
  NAND2_X1 U6361 ( .A1(n16319), .A2(n2945), .ZN(n2127) );
  NAND2_X1 U6362 ( .A1(n12483), .A2(n12472), .ZN(n2552) );
  XNOR2_X2 U6363 ( .A(n15988), .B(n15987), .ZN(n17676) );
  AOI21_X1 U6364 ( .B1(n15755), .B2(n2247), .A(n2101), .ZN(n2374) );
  NAND2_X1 U6366 ( .A1(n15760), .A2(n15754), .ZN(n2102) );
  OAI21_X1 U6367 ( .B1(n11363), .B2(n19952), .A(n2104), .ZN(n11372) );
  NAND2_X1 U6368 ( .A1(n15131), .A2(n15285), .ZN(n2105) );
  NAND2_X1 U6369 ( .A1(n8195), .A2(n8055), .ZN(n8194) );
  XNOR2_X1 U6372 ( .A(n13052), .B(n13051), .ZN(n14497) );
  OR2_X1 U6373 ( .A1(n9081), .A2(n9166), .ZN(n2941) );
  INV_X1 U6374 ( .A(n4706), .ZN(n3203) );
  INV_X1 U6375 ( .A(Plaintext[124]), .ZN(n3204) );
  NOR2_X1 U6376 ( .A1(n11051), .A2(n10829), .ZN(n2162) );
  NOR2_X1 U6377 ( .A1(n15303), .A2(n15302), .ZN(n2581) );
  XNOR2_X1 U6378 ( .A(n10351), .B(n9908), .ZN(n10395) );
  XNOR2_X1 U6379 ( .A(n16555), .B(n16236), .ZN(n16871) );
  XNOR2_X1 U6380 ( .A(n6410), .B(n7288), .ZN(n6864) );
  NAND3_X1 U6381 ( .A1(n5770), .A2(n5766), .A3(n5546), .ZN(n5738) );
  NAND2_X1 U6383 ( .A1(n2267), .A2(n15338), .ZN(n2109) );
  AOI22_X1 U6386 ( .A1(n20117), .A2(n18850), .B1(n19989), .B2(n18869), .ZN(
        n18871) );
  XNOR2_X1 U6387 ( .A(n10247), .B(n10248), .ZN(n10251) );
  NAND2_X1 U6388 ( .A1(n15039), .A2(n15141), .ZN(n2111) );
  NAND2_X1 U6389 ( .A1(n2113), .A2(n2112), .ZN(n14858) );
  NAND2_X1 U6390 ( .A1(n14857), .A2(n15766), .ZN(n2112) );
  NAND2_X1 U6391 ( .A1(n11155), .A2(n11159), .ZN(n2970) );
  NAND2_X1 U6394 ( .A1(n19710), .A2(n9262), .ZN(n2116) );
  INV_X1 U6395 ( .A(n9262), .ZN(n2118) );
  INV_X1 U6398 ( .A(n18025), .ZN(n2120) );
  NAND2_X1 U6399 ( .A1(n6143), .A2(n6140), .ZN(n4462) );
  NAND2_X1 U6400 ( .A1(n11718), .A2(n12282), .ZN(n2121) );
  NAND2_X1 U6401 ( .A1(n8071), .A2(n5762), .ZN(n8202) );
  NAND2_X1 U6402 ( .A1(n15664), .A2(n15773), .ZN(n15670) );
  XNOR2_X1 U6404 ( .A(n17127), .B(n2280), .ZN(n15951) );
  OAI21_X1 U6406 ( .B1(n12392), .B2(n3082), .A(n12391), .ZN(n12831) );
  NAND2_X1 U6407 ( .A1(n4927), .A2(n4932), .ZN(n4930) );
  OAI21_X1 U6408 ( .B1(n13977), .B2(n14284), .A(n2125), .ZN(n13978) );
  NAND3_X1 U6409 ( .A1(n5605), .A2(n5604), .A3(n5714), .ZN(n5607) );
  OAI21_X1 U6410 ( .B1(n8288), .B2(n7807), .A(n2126), .ZN(n7400) );
  NAND2_X1 U6411 ( .A1(n7807), .A2(n8289), .ZN(n2126) );
  OR3_X1 U6412 ( .A1(n8998), .A2(n8997), .A3(n7752), .ZN(n7774) );
  XNOR2_X2 U6413 ( .A(n3875), .B(Key[18]), .ZN(n4296) );
  AND2_X1 U6414 ( .A1(n8760), .A2(n265), .ZN(n8766) );
  OAI22_X1 U6416 ( .A1(n17662), .A2(n20185), .B1(n3214), .B2(n17890), .ZN(
        n3213) );
  OAI21_X1 U6417 ( .B1(n9299), .B2(n3418), .A(n2786), .ZN(n3201) );
  NAND2_X1 U6418 ( .A1(n3652), .A2(n4418), .ZN(n3651) );
  XNOR2_X1 U6419 ( .A(n2127), .B(n2263), .ZN(Ciphertext[152]) );
  OAI21_X1 U6420 ( .B1(n9172), .B2(n8617), .A(n8619), .ZN(n7806) );
  NAND3_X1 U6422 ( .A1(n15411), .A2(n15551), .A3(n2129), .ZN(n16050) );
  NAND2_X1 U6423 ( .A1(n20147), .A2(n15056), .ZN(n15411) );
  NAND2_X1 U6424 ( .A1(n256), .A2(n12179), .ZN(n9498) );
  NOR3_X1 U6426 ( .A1(n12267), .A2(n3734), .A3(n12562), .ZN(n11062) );
  NAND2_X1 U6428 ( .A1(n2133), .A2(n2132), .ZN(n10316) );
  NAND2_X1 U6429 ( .A1(n12337), .A2(n12336), .ZN(n2132) );
  NAND2_X1 U6430 ( .A1(n11974), .A2(n12334), .ZN(n2133) );
  NOR2_X1 U6431 ( .A1(n2135), .A2(n2134), .ZN(n11498) );
  NAND2_X1 U6432 ( .A1(n2137), .A2(n2136), .ZN(n6711) );
  NAND2_X1 U6433 ( .A1(n5707), .A2(n6002), .ZN(n2137) );
  NAND2_X1 U6434 ( .A1(n3319), .A2(n5880), .ZN(n5153) );
  NAND2_X1 U6435 ( .A1(n19329), .A2(n19324), .ZN(n19310) );
  NAND2_X1 U6436 ( .A1(n12632), .A2(n246), .ZN(n2139) );
  NAND2_X1 U6437 ( .A1(n11618), .A2(n1371), .ZN(n2140) );
  AND3_X2 U6438 ( .A1(n8043), .A2(n2142), .A3(n2141), .ZN(n8542) );
  NAND2_X1 U6439 ( .A1(n8296), .A2(n8300), .ZN(n2141) );
  NAND2_X1 U6440 ( .A1(n8042), .A2(n1835), .ZN(n2142) );
  OR2_X1 U6442 ( .A1(n5781), .A2(n6046), .ZN(n2144) );
  AOI22_X1 U6444 ( .A1(n12072), .A2(n12609), .B1(n12606), .B2(n12073), .ZN(
        n12076) );
  XNOR2_X1 U6445 ( .A(n929), .B(n10369), .ZN(n2145) );
  MUX2_X1 U6446 ( .A(n5880), .B(n5881), .S(n3319), .Z(n5882) );
  OAI21_X2 U6447 ( .B1(n12026), .B2(n12377), .A(n12025), .ZN(n13369) );
  NAND2_X1 U6449 ( .A1(n891), .A2(n9300), .ZN(n8584) );
  NAND2_X1 U6451 ( .A1(n14609), .A2(n14608), .ZN(n3226) );
  NAND2_X1 U6452 ( .A1(n15862), .A2(n15864), .ZN(n15860) );
  NAND2_X1 U6453 ( .A1(n12477), .A2(n12142), .ZN(n2148) );
  AND2_X1 U6454 ( .A1(n14203), .A2(n14012), .ZN(n14143) );
  INV_X1 U6456 ( .A(n12542), .ZN(n2600) );
  OR2_X1 U6457 ( .A1(n20357), .A2(n4867), .ZN(n4227) );
  NAND2_X1 U6459 ( .A1(n11569), .A2(n11564), .ZN(n2949) );
  OAI21_X1 U6460 ( .B1(n14159), .B2(n15509), .A(n2908), .ZN(n15514) );
  OAI22_X1 U6461 ( .A1(n8665), .A2(n9204), .B1(n20009), .B2(n9130), .ZN(n9779)
         );
  NAND2_X1 U6464 ( .A1(n6041), .A2(n5888), .ZN(n2149) );
  NAND2_X1 U6465 ( .A1(n14649), .A2(n19831), .ZN(n2153) );
  NAND2_X1 U6466 ( .A1(n2154), .A2(n8904), .ZN(n8592) );
  NAND2_X1 U6467 ( .A1(n2756), .A2(n19941), .ZN(n2154) );
  NAND2_X1 U6468 ( .A1(n5865), .A2(n2157), .ZN(n6786) );
  NAND2_X1 U6469 ( .A1(n2158), .A2(n5864), .ZN(n2157) );
  OAI22_X1 U6470 ( .A1(n20464), .A2(n4440), .B1(n5040), .B2(n4439), .ZN(n4441)
         );
  NOR2_X1 U6471 ( .A1(n9883), .A2(n11234), .ZN(n11367) );
  NAND2_X1 U6473 ( .A1(n12685), .A2(n12684), .ZN(n12687) );
  AOI21_X1 U6474 ( .B1(n5510), .B2(n5070), .A(n5071), .ZN(n4665) );
  NAND2_X1 U6475 ( .A1(n5069), .A2(n4410), .ZN(n5510) );
  NAND2_X1 U6476 ( .A1(n12307), .A2(n12543), .ZN(n2159) );
  OAI21_X1 U6477 ( .B1(n11418), .B2(n11417), .A(n2161), .ZN(n10725) );
  OAI21_X2 U6479 ( .B1(n6203), .B2(n5230), .A(n5229), .ZN(n7249) );
  NAND2_X1 U6482 ( .A1(n2236), .A2(n2237), .ZN(n18157) );
  XNOR2_X1 U6483 ( .A(n2163), .B(n16131), .ZN(n16133) );
  XNOR2_X1 U6484 ( .A(n16130), .B(n16988), .ZN(n2163) );
  NAND2_X1 U6485 ( .A1(n8032), .A2(n8284), .ZN(n2166) );
  OAI21_X1 U6486 ( .B1(n6139), .B2(n5866), .A(n5265), .ZN(n5267) );
  OR2_X1 U6488 ( .A1(n6951), .A2(n8365), .ZN(n7676) );
  OR2_X1 U6489 ( .A1(n11477), .A2(n3482), .ZN(n3480) );
  INV_X1 U6490 ( .A(n11311), .ZN(n2759) );
  NAND2_X1 U6492 ( .A1(n2698), .A2(n2167), .ZN(n2723) );
  NAND2_X1 U6493 ( .A1(n2171), .A2(n2168), .ZN(n9570) );
  NAND2_X1 U6494 ( .A1(n9564), .A2(n9563), .ZN(n2169) );
  OR2_X1 U6495 ( .A1(n20105), .A2(n3978), .ZN(n4658) );
  AND2_X1 U6496 ( .A1(n20235), .A2(n11292), .ZN(n10979) );
  INV_X1 U6497 ( .A(n3741), .ZN(n3103) );
  XNOR2_X1 U6498 ( .A(n17380), .B(n2172), .ZN(n17381) );
  XNOR2_X1 U6499 ( .A(n17377), .B(n17378), .ZN(n2172) );
  XNOR2_X1 U6501 ( .A(n10604), .B(n2349), .ZN(n10606) );
  AND2_X1 U6502 ( .A1(n8653), .A2(n9265), .ZN(n7867) );
  INV_X1 U6504 ( .A(n5815), .ZN(n3468) );
  XNOR2_X1 U6505 ( .A(n941), .B(n7296), .ZN(n7064) );
  OR2_X1 U6506 ( .A1(n17773), .A2(n18333), .ZN(n2177) );
  OAI21_X1 U6507 ( .B1(n5419), .B2(n5226), .A(n5418), .ZN(n2404) );
  XNOR2_X1 U6508 ( .A(n16566), .B(n17276), .ZN(n16091) );
  NAND2_X1 U6511 ( .A1(n2179), .A2(n2178), .ZN(n18798) );
  NAND2_X1 U6512 ( .A1(n18796), .A2(n18795), .ZN(n2178) );
  INV_X1 U6514 ( .A(n18814), .ZN(n18811) );
  NAND2_X1 U6515 ( .A1(n2182), .A2(n2180), .ZN(n17058) );
  NAND2_X1 U6516 ( .A1(n18916), .A2(n2181), .ZN(n2180) );
  NOR2_X1 U6517 ( .A1(n18921), .A2(n18899), .ZN(n2181) );
  NAND2_X1 U6518 ( .A1(n18874), .A2(n19874), .ZN(n2182) );
  INV_X1 U6522 ( .A(n17303), .ZN(n3205) );
  OR2_X1 U6523 ( .A1(n11954), .A2(n11951), .ZN(n11956) );
  NOR2_X1 U6524 ( .A1(n3839), .A2(n5782), .ZN(n3249) );
  NOR2_X1 U6525 ( .A1(n3671), .A2(n11145), .ZN(n3670) );
  AND2_X1 U6526 ( .A1(n14465), .A2(n14462), .ZN(n14176) );
  INV_X1 U6527 ( .A(n9164), .ZN(n8609) );
  XNOR2_X1 U6528 ( .A(n2312), .B(n13624), .ZN(n13533) );
  OAI21_X1 U6529 ( .B1(n9158), .B2(n8696), .A(n8610), .ZN(n8614) );
  XNOR2_X1 U6530 ( .A(n5884), .B(n7118), .ZN(n6659) );
  NAND2_X1 U6531 ( .A1(n12565), .A2(n2183), .ZN(n12566) );
  NAND3_X2 U6532 ( .A1(n3536), .A2(n2185), .A3(n2184), .ZN(n13715) );
  NAND2_X1 U6533 ( .A1(n2737), .A2(n12002), .ZN(n2185) );
  OAI211_X2 U6534 ( .C1(n14696), .C2(n14695), .A(n14694), .B(n2186), .ZN(
        n15567) );
  NAND3_X1 U6535 ( .A1(n2187), .A2(n11639), .A3(n12209), .ZN(n2714) );
  NAND2_X1 U6536 ( .A1(n12067), .A2(n12206), .ZN(n2187) );
  NAND2_X1 U6537 ( .A1(n9276), .A2(n8991), .ZN(n7897) );
  NAND2_X1 U6538 ( .A1(n11939), .A2(n12110), .ZN(n12099) );
  NAND2_X1 U6540 ( .A1(n8083), .A2(n8232), .ZN(n2188) );
  NAND2_X1 U6542 ( .A1(n6584), .A2(n6585), .ZN(n2191) );
  NOR2_X1 U6543 ( .A1(n4185), .A2(n4633), .ZN(n4159) );
  AOI22_X1 U6544 ( .A1(n15372), .A2(n15567), .B1(n15564), .B2(n20183), .ZN(
        n15373) );
  OAI211_X1 U6545 ( .C1(n11329), .C2(n2858), .A(n2861), .B(n2857), .ZN(n2856)
         );
  NAND2_X1 U6546 ( .A1(n3393), .A2(n3457), .ZN(n3392) );
  INV_X1 U6548 ( .A(n19113), .ZN(n2195) );
  INV_X1 U6550 ( .A(n17533), .ZN(n2197) );
  NAND2_X1 U6551 ( .A1(n4771), .A2(n5035), .ZN(n5038) );
  INV_X1 U6552 ( .A(n19386), .ZN(n17220) );
  INV_X1 U6553 ( .A(n8167), .ZN(n3121) );
  NAND3_X1 U6554 ( .A1(n19789), .A2(n5926), .A3(n6026), .ZN(n2342) );
  INV_X1 U6556 ( .A(n7750), .ZN(n3446) );
  XNOR2_X1 U6557 ( .A(n2199), .B(n10588), .ZN(n9428) );
  XNOR2_X1 U6558 ( .A(n3184), .B(n10430), .ZN(n2199) );
  NAND2_X1 U6559 ( .A1(n3632), .A2(n11599), .ZN(n3631) );
  NAND2_X1 U6561 ( .A1(n1527), .A2(n2201), .ZN(n14234) );
  OAI211_X2 U6563 ( .C1(n5669), .C2(n4880), .A(n5677), .B(n4879), .ZN(n7337)
         );
  AND2_X1 U6565 ( .A1(n14556), .A2(n14553), .ZN(n14551) );
  NAND2_X1 U6567 ( .A1(n4588), .A2(n4585), .ZN(n5054) );
  OAI21_X1 U6569 ( .B1(n11421), .B2(n11420), .A(n11422), .ZN(n2440) );
  NAND2_X1 U6570 ( .A1(n2205), .A2(n2204), .ZN(n17056) );
  NAND2_X1 U6571 ( .A1(n19684), .A2(n18961), .ZN(n2204) );
  NAND2_X1 U6572 ( .A1(n17055), .A2(n220), .ZN(n2205) );
  NAND2_X1 U6573 ( .A1(n16674), .A2(n19352), .ZN(n2206) );
  OAI21_X1 U6574 ( .B1(n4368), .B2(n5240), .A(n5720), .ZN(n2207) );
  NOR2_X2 U6575 ( .A1(n11068), .A2(n11067), .ZN(n13319) );
  OR2_X2 U6577 ( .A1(n10812), .A2(n10811), .ZN(n12211) );
  NAND2_X1 U6579 ( .A1(n2209), .A2(n11570), .ZN(n10752) );
  NAND2_X1 U6580 ( .A1(n10751), .A2(n2210), .ZN(n2209) );
  INV_X1 U6581 ( .A(n11568), .ZN(n2210) );
  XNOR2_X1 U6582 ( .A(n6771), .B(n6770), .ZN(n2211) );
  NAND2_X1 U6583 ( .A1(n2213), .A2(n2212), .ZN(n15359) );
  NAND2_X1 U6584 ( .A1(n15357), .A2(n15815), .ZN(n2212) );
  NAND2_X1 U6585 ( .A1(n15358), .A2(n3534), .ZN(n2213) );
  NAND2_X1 U6589 ( .A1(n5032), .A2(n4706), .ZN(n4709) );
  NAND2_X1 U6591 ( .A1(n8282), .A2(n8286), .ZN(n2217) );
  XNOR2_X1 U6593 ( .A(n13031), .B(n12986), .ZN(n13733) );
  INV_X1 U6594 ( .A(n18046), .ZN(n2586) );
  INV_X1 U6595 ( .A(n5087), .ZN(n4801) );
  OR2_X1 U6596 ( .A1(n4979), .A2(n4296), .ZN(n4020) );
  INV_X1 U6597 ( .A(n3305), .ZN(n12610) );
  INV_X1 U6598 ( .A(n15295), .ZN(n3307) );
  INV_X1 U6599 ( .A(n10926), .ZN(n11545) );
  XNOR2_X1 U6600 ( .A(n13707), .B(n13002), .ZN(n3460) );
  OAI21_X1 U6601 ( .B1(n5972), .B2(n5971), .A(n5970), .ZN(n5975) );
  NAND2_X1 U6602 ( .A1(n5967), .A2(n5697), .ZN(n5970) );
  XNOR2_X1 U6604 ( .A(n2224), .B(n16518), .ZN(n16520) );
  XNOR2_X1 U6605 ( .A(n16602), .B(n16517), .ZN(n2224) );
  NAND2_X1 U6606 ( .A1(n8193), .A2(n8197), .ZN(n7627) );
  NAND2_X1 U6608 ( .A1(n18165), .A2(n19292), .ZN(n2226) );
  XNOR2_X1 U6609 ( .A(n9946), .B(n10071), .ZN(n10621) );
  XNOR2_X1 U6611 ( .A(n13513), .B(n2228), .ZN(n13515) );
  XNOR2_X1 U6612 ( .A(n13514), .B(n13512), .ZN(n2228) );
  OAI21_X1 U6613 ( .B1(n10854), .B2(n11230), .A(n2229), .ZN(n11233) );
  NAND2_X1 U6614 ( .A1(n11230), .A2(n11365), .ZN(n2229) );
  XNOR2_X1 U6615 ( .A(n2230), .B(n13852), .ZN(n12249) );
  XNOR2_X1 U6616 ( .A(n13757), .B(n12219), .ZN(n2230) );
  INV_X1 U6617 ( .A(n873), .ZN(n2929) );
  XNOR2_X2 U6618 ( .A(n12783), .B(n12782), .ZN(n13931) );
  INV_X1 U6619 ( .A(n11176), .ZN(n2232) );
  NAND2_X1 U6620 ( .A1(n10997), .A2(n11289), .ZN(n2235) );
  INV_X1 U6621 ( .A(Plaintext[53]), .ZN(n3543) );
  OAI21_X1 U6624 ( .B1(n16152), .B2(n20423), .A(n16151), .ZN(n2237) );
  NAND2_X1 U6625 ( .A1(n4545), .A2(n2239), .ZN(n4551) );
  NAND3_X1 U6627 ( .A1(n3710), .A2(n15921), .A3(n15421), .ZN(n14899) );
  NOR2_X1 U6628 ( .A1(n12212), .A2(n12211), .ZN(n2743) );
  NAND2_X1 U6630 ( .A1(n10854), .A2(n11230), .ZN(n9884) );
  NAND2_X1 U6631 ( .A1(n8618), .A2(n8987), .ZN(n2241) );
  INV_X1 U6632 ( .A(n8987), .ZN(n2243) );
  NAND3_X2 U6633 ( .A1(n14628), .A2(n14621), .A3(n14622), .ZN(n15600) );
  MUX2_X1 U6635 ( .A(n8525), .B(n8526), .S(n9038), .Z(n8531) );
  NAND2_X1 U6636 ( .A1(n15761), .A2(n2247), .ZN(n2246) );
  INV_X1 U6637 ( .A(n15760), .ZN(n2247) );
  NAND2_X2 U6638 ( .A1(n3165), .A2(n4794), .ZN(n5663) );
  NAND2_X1 U6639 ( .A1(n12443), .A2(n12440), .ZN(n12435) );
  NAND3_X1 U6640 ( .A1(n20261), .A2(n2697), .A3(n14828), .ZN(n2696) );
  NOR2_X1 U6641 ( .A1(n7311), .A2(n7312), .ZN(n7998) );
  NAND2_X1 U6642 ( .A1(n210), .A2(n2596), .ZN(n2576) );
  XNOR2_X1 U6643 ( .A(n2250), .B(n13470), .ZN(n13473) );
  XNOR2_X1 U6644 ( .A(n13469), .B(n13818), .ZN(n2250) );
  NAND2_X1 U6646 ( .A1(n7905), .A2(n280), .ZN(n2252) );
  AOI21_X1 U6647 ( .B1(n2253), .B2(n4509), .A(n4371), .ZN(n4374) );
  NAND2_X1 U6648 ( .A1(n4372), .A2(n4577), .ZN(n2253) );
  INV_X1 U6649 ( .A(n15188), .ZN(n13933) );
  XOR2_X1 U6650 ( .A(n13778), .B(n13059), .Z(n2620) );
  NAND2_X1 U6651 ( .A1(n12637), .A2(n19861), .ZN(n2254) );
  NAND2_X1 U6652 ( .A1(n12638), .A2(n2256), .ZN(n2255) );
  MUX2_X2 U6653 ( .A(n10807), .B(n10806), .S(n11257), .Z(n12209) );
  XNOR2_X2 U6654 ( .A(n12764), .B(n12763), .ZN(n14827) );
  NAND2_X1 U6655 ( .A1(n2688), .A2(n2703), .ZN(n2702) );
  INV_X1 U6656 ( .A(n15052), .ZN(n15458) );
  INV_X1 U6657 ( .A(n8993), .ZN(n9278) );
  NAND2_X1 U6658 ( .A1(n13961), .A2(n14924), .ZN(n13970) );
  NAND2_X1 U6659 ( .A1(n6905), .A2(n7909), .ZN(n2258) );
  NAND2_X1 U6661 ( .A1(n19268), .A2(n19267), .ZN(n2261) );
  NAND2_X1 U6662 ( .A1(n19266), .A2(n20444), .ZN(n2262) );
  INV_X1 U6663 ( .A(n18354), .ZN(n18289) );
  NOR2_X2 U6664 ( .A1(n6898), .A2(n6897), .ZN(n10252) );
  INV_X1 U6665 ( .A(n6107), .ZN(n3010) );
  OAI21_X1 U6666 ( .B1(n11931), .B2(n12480), .A(n2265), .ZN(n11708) );
  NAND2_X1 U6667 ( .A1(n12478), .A2(n12142), .ZN(n2265) );
  NAND4_X2 U6668 ( .A1(n2266), .A2(n3132), .A3(n5062), .A4(n5061), .ZN(n5930)
         );
  OAI21_X1 U6669 ( .B1(n13166), .B2(n14664), .A(n3367), .ZN(n14671) );
  NAND2_X1 U6671 ( .A1(n15337), .A2(n15336), .ZN(n2267) );
  NAND3_X1 U6672 ( .A1(n14130), .A2(n14129), .A3(n14128), .ZN(n15607) );
  INV_X1 U6674 ( .A(n2269), .ZN(n2268) );
  OAI22_X1 U6675 ( .A1(n17832), .A2(n17831), .B1(n17833), .B2(n18959), .ZN(
        n2269) );
  NAND2_X1 U6676 ( .A1(n11441), .A2(n11440), .ZN(n2270) );
  NAND2_X1 U6677 ( .A1(n11442), .A2(n2272), .ZN(n2271) );
  XNOR2_X2 U6678 ( .A(n3930), .B(Key[164]), .ZN(n4347) );
  NOR2_X1 U6679 ( .A1(n15664), .A2(n2273), .ZN(n13460) );
  INV_X1 U6680 ( .A(n15772), .ZN(n2273) );
  NOR2_X2 U6681 ( .A1(n15398), .A2(n15399), .ZN(n16761) );
  AOI21_X1 U6682 ( .B1(n2761), .B2(n2760), .A(n2759), .ZN(n2758) );
  NOR2_X1 U6683 ( .A1(n209), .A2(n6068), .ZN(n3767) );
  XNOR2_X1 U6684 ( .A(n10507), .B(n2506), .ZN(n10509) );
  NAND2_X1 U6685 ( .A1(n4485), .A2(n3996), .ZN(n4681) );
  XNOR2_X2 U6687 ( .A(n13728), .B(n13729), .ZN(n14381) );
  NOR2_X1 U6688 ( .A1(n20611), .A2(n20361), .ZN(n18381) );
  XNOR2_X1 U6689 ( .A(n13191), .B(n12825), .ZN(n2783) );
  AOI21_X1 U6690 ( .B1(n2276), .B2(n14502), .A(n13040), .ZN(n13056) );
  NAND2_X1 U6691 ( .A1(n9307), .A2(n9310), .ZN(n8824) );
  NAND2_X1 U6692 ( .A1(n2277), .A2(n20434), .ZN(n17615) );
  INV_X1 U6693 ( .A(n19298), .ZN(n2277) );
  AOI21_X2 U6694 ( .B1(n17605), .B2(n17604), .A(n17603), .ZN(n19298) );
  NAND2_X1 U6695 ( .A1(n5749), .A2(n5747), .ZN(n2482) );
  AOI21_X1 U6696 ( .B1(n11369), .B2(n10680), .A(n11364), .ZN(n10681) );
  NOR2_X2 U6698 ( .A1(n7652), .A2(n7651), .ZN(n10566) );
  NAND2_X1 U6700 ( .A1(n5546), .A2(n5736), .ZN(n4545) );
  NAND2_X1 U6702 ( .A1(n15453), .A2(n15683), .ZN(n2279) );
  NAND3_X1 U6705 ( .A1(n4151), .A2(n4312), .A3(n4361), .ZN(n4155) );
  NAND2_X1 U6708 ( .A1(n13308), .A2(n2282), .ZN(n2281) );
  OAI211_X2 U6709 ( .C1(n7470), .C2(n8031), .A(n2283), .B(n8030), .ZN(n9060)
         );
  NAND2_X1 U6710 ( .A1(n8028), .A2(n8029), .ZN(n2283) );
  XNOR2_X1 U6711 ( .A(n8509), .B(n9445), .ZN(n2285) );
  NAND2_X1 U6712 ( .A1(n16730), .A2(n3755), .ZN(n3283) );
  AOI21_X1 U6713 ( .B1(n6070), .B2(n6072), .A(n2286), .ZN(n6074) );
  BUF_X1 U6714 ( .A(n3843), .Z(n4676) );
  OAI211_X1 U6715 ( .C1(n5072), .C2(n5071), .A(n4816), .B(n2287), .ZN(n4818)
         );
  AND3_X2 U6716 ( .A1(n3650), .A2(n3651), .A3(n4419), .ZN(n5868) );
  XNOR2_X2 U6717 ( .A(n16124), .B(n16125), .ZN(n17840) );
  INV_X1 U6718 ( .A(n15188), .ZN(n2288) );
  INV_X1 U6719 ( .A(n2561), .ZN(n3385) );
  XNOR2_X1 U6720 ( .A(n3620), .B(n7381), .ZN(n7388) );
  MUX2_X1 U6721 ( .A(n12532), .B(n12534), .S(n12162), .Z(n11807) );
  INV_X1 U6722 ( .A(n15660), .ZN(n15653) );
  NAND2_X1 U6723 ( .A1(n17774), .A2(n17777), .ZN(n2289) );
  NAND2_X1 U6724 ( .A1(n17449), .A2(n18129), .ZN(n2290) );
  NAND2_X1 U6725 ( .A1(n2292), .A2(n6075), .ZN(n2291) );
  NAND2_X1 U6726 ( .A1(n3318), .A2(n209), .ZN(n2292) );
  NOR2_X2 U6727 ( .A1(n8487), .A2(n8486), .ZN(n10402) );
  NAND2_X1 U6728 ( .A1(n3995), .A2(n4684), .ZN(n4226) );
  NAND2_X1 U6729 ( .A1(n15078), .A2(n15077), .ZN(n14371) );
  NAND2_X1 U6731 ( .A1(n2919), .A2(n20487), .ZN(n3634) );
  INV_X1 U6733 ( .A(n15465), .ZN(n12768) );
  OAI211_X2 U6734 ( .C1(n12726), .C2(n12727), .A(n13924), .B(n3190), .ZN(
        n15465) );
  OAI21_X1 U6736 ( .B1(n16461), .B2(n17479), .A(n960), .ZN(n2297) );
  OAI21_X1 U6738 ( .B1(n5717), .B2(n5716), .A(n5718), .ZN(n3664) );
  OR2_X1 U6739 ( .A1(n3995), .A2(n3996), .ZN(n4851) );
  XNOR2_X2 U6742 ( .A(Key[75]), .B(Plaintext[75]), .ZN(n4824) );
  XNOR2_X1 U6743 ( .A(n6982), .B(n7050), .ZN(n6328) );
  NAND3_X1 U6744 ( .A1(n619), .A2(n4612), .A3(n3716), .ZN(n3714) );
  OAI21_X2 U6747 ( .B1(n9063), .B2(n9036), .A(n9035), .ZN(n9991) );
  NAND3_X2 U6748 ( .A1(n11308), .A2(n11309), .A3(n11307), .ZN(n12809) );
  OAI21_X1 U6749 ( .B1(n17601), .B2(n17890), .A(n2302), .ZN(n17889) );
  NAND2_X1 U6750 ( .A1(n20019), .A2(n17890), .ZN(n2302) );
  AOI21_X1 U6751 ( .B1(n7853), .B2(n7854), .A(n7852), .ZN(n2303) );
  NAND2_X1 U6752 ( .A1(n9029), .A2(n9062), .ZN(n8677) );
  INV_X1 U6753 ( .A(n2800), .ZN(n15073) );
  INV_X1 U6755 ( .A(n4615), .ZN(n3717) );
  OAI211_X2 U6756 ( .C1(n15797), .C2(n15796), .A(n2309), .B(n2308), .ZN(n17426) );
  NAND2_X1 U6757 ( .A1(n15793), .A2(n15796), .ZN(n2308) );
  NAND2_X1 U6758 ( .A1(n16810), .A2(n18546), .ZN(n18532) );
  NAND2_X1 U6759 ( .A1(n13274), .A2(n12324), .ZN(n12329) );
  NAND2_X1 U6760 ( .A1(n12322), .A2(n12323), .ZN(n13274) );
  NAND2_X1 U6761 ( .A1(n13859), .A2(n15443), .ZN(n2311) );
  OAI21_X1 U6763 ( .B1(n14601), .B2(n19918), .A(n1262), .ZN(n2314) );
  NAND2_X1 U6764 ( .A1(n9491), .A2(n12180), .ZN(n11845) );
  OAI21_X1 U6767 ( .B1(n2316), .B2(n14833), .A(n14828), .ZN(n12767) );
  NAND4_X2 U6768 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), .ZN(n7365)
         );
  INV_X1 U6769 ( .A(n2955), .ZN(n7610) );
  OR2_X1 U6770 ( .A1(n14420), .A2(n14355), .ZN(n14356) );
  AND2_X1 U6771 ( .A1(n12315), .A2(n2612), .ZN(n2338) );
  INV_X1 U6773 ( .A(n14461), .ZN(n15111) );
  NAND2_X1 U6774 ( .A1(n16780), .A2(n870), .ZN(n16779) );
  XNOR2_X1 U6775 ( .A(n2318), .B(n16788), .ZN(Ciphertext[135]) );
  NAND3_X1 U6776 ( .A1(n3139), .A2(n3142), .A3(n3143), .ZN(n2318) );
  OAI21_X2 U6777 ( .B1(n11037), .B2(n10523), .A(n10522), .ZN(n12514) );
  NAND3_X1 U6778 ( .A1(n12243), .A2(n12619), .A3(n894), .ZN(n12244) );
  NAND2_X1 U6779 ( .A1(n14236), .A2(n14239), .ZN(n14401) );
  NAND2_X1 U6780 ( .A1(n3048), .A2(n3052), .ZN(n2319) );
  NAND3_X1 U6781 ( .A1(n4160), .A2(n4517), .A3(n4523), .ZN(n4161) );
  NAND2_X1 U6782 ( .A1(n12313), .A2(n12153), .ZN(n2320) );
  NAND2_X1 U6783 ( .A1(n3235), .A2(n18104), .ZN(n18110) );
  AND3_X2 U6784 ( .A1(n14152), .A2(n14151), .A3(n14150), .ZN(n3822) );
  NAND3_X2 U6785 ( .A1(n2322), .A2(n2321), .A3(n5290), .ZN(n7006) );
  NAND3_X1 U6786 ( .A1(n5289), .A2(n5291), .A3(n5443), .ZN(n2322) );
  OR2_X2 U6787 ( .A1(n4408), .A2(n4407), .ZN(n5873) );
  INV_X1 U6788 ( .A(n7405), .ZN(n7402) );
  NAND2_X1 U6790 ( .A1(n7479), .A2(n7953), .ZN(n2324) );
  INV_X1 U6791 ( .A(n7951), .ZN(n2325) );
  INV_X1 U6792 ( .A(n7952), .ZN(n2326) );
  MUX2_X1 U6793 ( .A(n15282), .B(n15128), .S(n15127), .Z(n15129) );
  NOR2_X2 U6794 ( .A1(n14528), .A2(n14527), .ZN(n15127) );
  XNOR2_X1 U6795 ( .A(n7123), .B(n7119), .ZN(n3572) );
  INV_X1 U6796 ( .A(n2661), .ZN(n2659) );
  OAI211_X2 U6798 ( .C1(n19789), .C2(n6030), .A(n6029), .B(n6028), .ZN(n7042)
         );
  OAI211_X2 U6799 ( .C1(n12539), .C2(n12538), .A(n2328), .B(n2327), .ZN(n3159)
         );
  NAND2_X1 U6800 ( .A1(n12536), .A2(n12535), .ZN(n2327) );
  NOR2_X1 U6802 ( .A1(n14494), .A2(n3155), .ZN(n14495) );
  NAND3_X1 U6804 ( .A1(n9837), .A2(n20476), .A3(n8542), .ZN(n2330) );
  INV_X1 U6808 ( .A(n12377), .ZN(n2333) );
  XOR2_X1 U6809 ( .A(n13581), .B(n13582), .Z(n3062) );
  INV_X1 U6810 ( .A(n11604), .ZN(n11605) );
  NOR2_X1 U6811 ( .A1(n3669), .A2(n11339), .ZN(n11266) );
  AOI22_X1 U6812 ( .A1(n8068), .A2(n7622), .B1(n8067), .B2(n8179), .ZN(n3526)
         );
  AOI22_X2 U6813 ( .A1(n12876), .A2(n14050), .B1(n13932), .B2(n13931), .ZN(
        n15188) );
  OR2_X2 U6814 ( .A1(n2334), .A2(n4038), .ZN(n5888) );
  NAND3_X1 U6815 ( .A1(n3729), .A2(n3730), .A3(n18033), .ZN(n3691) );
  NAND2_X1 U6817 ( .A1(n8617), .A2(n19827), .ZN(n8618) );
  INV_X1 U6818 ( .A(n12484), .ZN(n12477) );
  NAND3_X1 U6819 ( .A1(n14275), .A2(n14562), .A3(n14705), .ZN(n2541) );
  NAND2_X1 U6820 ( .A1(n15635), .A2(n15636), .ZN(n15637) );
  NAND2_X1 U6821 ( .A1(n18593), .A2(n20365), .ZN(n17919) );
  NAND2_X1 U6824 ( .A1(n8873), .A2(n9107), .ZN(n8874) );
  AOI22_X2 U6825 ( .A1(n17162), .A2(n17163), .B1(n17160), .B2(n17161), .ZN(
        n18589) );
  INV_X1 U6826 ( .A(n13312), .ZN(n13161) );
  OAI211_X1 U6828 ( .C1(n8312), .C2(n8313), .A(n2339), .B(n20144), .ZN(n8320)
         );
  NAND2_X1 U6829 ( .A1(n8312), .A2(n19520), .ZN(n2339) );
  NAND2_X1 U6831 ( .A1(n13141), .A2(n13147), .ZN(n12572) );
  NAND2_X1 U6832 ( .A1(n20157), .A2(n14268), .ZN(n14576) );
  NAND3_X2 U6833 ( .A1(n2717), .A2(n2716), .A3(n14386), .ZN(n15625) );
  OR2_X1 U6834 ( .A1(n12934), .A2(n14327), .ZN(n2535) );
  OAI211_X2 U6835 ( .C1(n5597), .C2(n6026), .A(n2343), .B(n2342), .ZN(n6819)
         );
  NAND2_X1 U6836 ( .A1(n5928), .A2(n5596), .ZN(n2343) );
  NAND2_X1 U6837 ( .A1(n11008), .A2(n12576), .ZN(n2346) );
  OAI21_X2 U6838 ( .B1(n4347), .B2(n4203), .A(n4202), .ZN(n5670) );
  NAND3_X1 U6839 ( .A1(n2348), .A2(n18579), .A3(n18578), .ZN(n18580) );
  OAI21_X1 U6840 ( .B1(n18575), .B2(n18576), .A(n19665), .ZN(n2348) );
  NOR2_X1 U6842 ( .A1(n12082), .A2(n12427), .ZN(n12086) );
  XNOR2_X1 U6843 ( .A(n13266), .B(n19854), .ZN(n13579) );
  AND2_X1 U6845 ( .A1(n2350), .A2(n12110), .ZN(n11622) );
  INV_X1 U6846 ( .A(n12443), .ZN(n2350) );
  MUX2_X1 U6847 ( .A(n8671), .B(n8586), .S(n19857), .Z(n2351) );
  XNOR2_X1 U6848 ( .A(n2352), .B(n16755), .ZN(n16757) );
  XNOR2_X1 U6849 ( .A(n17335), .B(n17989), .ZN(n2352) );
  NAND3_X1 U6850 ( .A1(n5735), .A2(n5763), .A3(n5736), .ZN(n5737) );
  OAI211_X1 U6852 ( .C1(n11193), .C2(n10903), .A(n2355), .B(n2354), .ZN(n10625) );
  NAND2_X1 U6853 ( .A1(n10577), .A2(n11193), .ZN(n2354) );
  NAND2_X1 U6854 ( .A1(n10576), .A2(n11186), .ZN(n2355) );
  OR2_X1 U6856 ( .A1(n7908), .A2(n6904), .ZN(n7003) );
  INV_X1 U6857 ( .A(n13180), .ZN(n15778) );
  XNOR2_X1 U6858 ( .A(n10574), .B(n10568), .ZN(n2496) );
  NAND2_X1 U6859 ( .A1(n15336), .A2(n15341), .ZN(n15467) );
  AND3_X2 U6861 ( .A1(n2358), .A2(n14333), .A3(n2357), .ZN(n16300) );
  NAND2_X1 U6862 ( .A1(n14332), .A2(n20502), .ZN(n2357) );
  OAI21_X1 U6864 ( .B1(n18120), .B2(n19876), .A(n2359), .ZN(n18125) );
  NAND2_X1 U6865 ( .A1(n19876), .A2(n18121), .ZN(n2359) );
  NAND2_X1 U6866 ( .A1(n19069), .A2(n19685), .ZN(n19055) );
  MUX2_X1 U6867 ( .A(n10731), .B(n10732), .S(n11493), .Z(n2360) );
  NAND2_X1 U6868 ( .A1(n3117), .A2(n17828), .ZN(n3116) );
  OR2_X1 U6869 ( .A1(n4602), .A2(n4355), .ZN(n4605) );
  NAND2_X1 U6870 ( .A1(n11204), .A2(n11209), .ZN(n11097) );
  NAND2_X1 U6871 ( .A1(n3297), .A2(n3298), .ZN(n9381) );
  XNOR2_X1 U6872 ( .A(n2362), .B(n2361), .ZN(Ciphertext[120]) );
  NAND3_X1 U6873 ( .A1(n20467), .A2(n15167), .A3(n3621), .ZN(n2363) );
  NAND2_X1 U6874 ( .A1(n15382), .A2(n20103), .ZN(n2364) );
  NAND2_X1 U6875 ( .A1(n17488), .A2(n16800), .ZN(n2692) );
  NAND2_X1 U6876 ( .A1(n2365), .A2(n10862), .ZN(n10868) );
  INV_X1 U6877 ( .A(n14518), .ZN(n13564) );
  NAND2_X1 U6878 ( .A1(n20272), .A2(n15121), .ZN(n14518) );
  NAND2_X1 U6880 ( .A1(n2367), .A2(n2366), .ZN(n13063) );
  NAND3_X1 U6881 ( .A1(n4909), .A2(n4910), .A3(n4954), .ZN(n4918) );
  OAI211_X1 U6883 ( .C1(n4136), .C2(n3231), .A(n3230), .B(n4377), .ZN(n3229)
         );
  AOI21_X1 U6885 ( .B1(n8239), .B2(n7862), .A(n8111), .ZN(n3772) );
  NAND3_X1 U6886 ( .A1(n7779), .A2(n8007), .A3(n8313), .ZN(n7778) );
  OR2_X1 U6887 ( .A1(n4361), .A2(n4362), .ZN(n2370) );
  NAND2_X1 U6888 ( .A1(n9176), .A2(n8761), .ZN(n8760) );
  OAI21_X1 U6891 ( .B1(n11960), .B2(n1371), .A(n3721), .ZN(n3720) );
  NOR2_X1 U6892 ( .A1(n16636), .A2(n2372), .ZN(n16637) );
  NAND2_X1 U6893 ( .A1(n16635), .A2(n19348), .ZN(n2372) );
  NAND2_X1 U6894 ( .A1(n14849), .A2(n15655), .ZN(n15243) );
  NOR2_X1 U6896 ( .A1(n15562), .A2(n15510), .ZN(n2373) );
  MUX2_X1 U6897 ( .A(n18763), .B(n18773), .S(n18774), .Z(n18767) );
  AOI22_X2 U6899 ( .A1(n13975), .A2(n14306), .B1(n13871), .B2(n13870), .ZN(
        n15192) );
  NOR2_X2 U6900 ( .A1(n2374), .A2(n2814), .ZN(n17410) );
  NOR2_X1 U6901 ( .A1(n3689), .A2(n3690), .ZN(n15765) );
  OAI22_X1 U6902 ( .A1(n12095), .A2(n2805), .B1(n12429), .B2(n12645), .ZN(
        n2804) );
  INV_X1 U6903 ( .A(n4910), .ZN(n3079) );
  NAND2_X1 U6906 ( .A1(n8203), .A2(n8070), .ZN(n2378) );
  AND2_X1 U6907 ( .A1(n15454), .A2(n15777), .ZN(n13095) );
  AND2_X1 U6908 ( .A1(n231), .A2(n15379), .ZN(n15030) );
  NAND2_X1 U6909 ( .A1(n14418), .A2(n13937), .ZN(n14054) );
  NAND2_X1 U6910 ( .A1(n14377), .A2(n15846), .ZN(n2380) );
  INV_X1 U6911 ( .A(n6113), .ZN(n6108) );
  INV_X1 U6912 ( .A(n14449), .ZN(n14455) );
  NOR2_X1 U6913 ( .A1(n11646), .A2(n12121), .ZN(n12123) );
  NOR2_X1 U6915 ( .A1(n12919), .A2(n701), .ZN(n12926) );
  INV_X1 U6916 ( .A(n7632), .ZN(n8094) );
  INV_X1 U6919 ( .A(n5674), .ZN(n5673) );
  OR3_X1 U6920 ( .A1(n8741), .A2(n8743), .A3(n8742), .ZN(n7649) );
  NAND3_X1 U6921 ( .A1(n12226), .A2(n12224), .A3(n12220), .ZN(n10934) );
  NAND2_X1 U6922 ( .A1(n7623), .A2(n8067), .ZN(n2387) );
  NAND4_X2 U6923 ( .A1(n12218), .A2(n12216), .A3(n12215), .A4(n12217), .ZN(
        n13295) );
  NAND2_X1 U6926 ( .A1(n4116), .A2(n2389), .ZN(n4885) );
  AOI21_X1 U6927 ( .B1(n12646), .B2(n2805), .A(n3647), .ZN(n3646) );
  NAND2_X1 U6928 ( .A1(n4508), .A2(n4509), .ZN(n4515) );
  NAND2_X1 U6929 ( .A1(n14423), .A2(n14422), .ZN(n2390) );
  NAND2_X1 U6930 ( .A1(n14421), .A2(n2039), .ZN(n2391) );
  OAI21_X1 U6931 ( .B1(n1055), .B2(n1022), .A(n2393), .ZN(n17632) );
  NAND2_X1 U6932 ( .A1(n17631), .A2(n1055), .ZN(n2393) );
  NAND2_X1 U6933 ( .A1(n5767), .A2(n5766), .ZN(n5225) );
  OAI21_X2 U6934 ( .B1(n12564), .B2(n12267), .A(n12266), .ZN(n13616) );
  INV_X1 U6937 ( .A(n17878), .ZN(n3345) );
  NAND2_X1 U6939 ( .A1(n8734), .A2(n8736), .ZN(n8921) );
  OAI21_X1 U6940 ( .B1(n7934), .B2(n20195), .A(n7936), .ZN(n7520) );
  XNOR2_X1 U6941 ( .A(n17400), .B(n3091), .ZN(n3090) );
  XNOR2_X2 U6942 ( .A(n6934), .B(n2397), .ZN(n8166) );
  XNOR2_X1 U6943 ( .A(n6932), .B(n6933), .ZN(n2397) );
  NAND2_X1 U6946 ( .A1(n4358), .A2(n4546), .ZN(n4311) );
  AOI21_X1 U6947 ( .B1(n8729), .B2(n2400), .A(n8947), .ZN(n8594) );
  INV_X1 U6950 ( .A(n11399), .ZN(n2725) );
  NAND2_X1 U6951 ( .A1(n20097), .A2(n18813), .ZN(n17991) );
  NAND2_X1 U6952 ( .A1(n14673), .A2(n3373), .ZN(n2402) );
  INV_X1 U6953 ( .A(n2404), .ZN(n2403) );
  NAND2_X1 U6954 ( .A1(n5024), .A2(n4271), .ZN(n4581) );
  AOI21_X2 U6955 ( .B1(n7410), .B2(n7409), .A(n2405), .ZN(n8749) );
  OAI211_X2 U6956 ( .C1(n4584), .C2(n5026), .A(n4583), .B(n4582), .ZN(n6189)
         );
  OAI21_X1 U6957 ( .B1(n5796), .B2(n2407), .A(n2406), .ZN(n5431) );
  NAND2_X1 U6958 ( .A1(n5790), .A2(n5796), .ZN(n2406) );
  OAI21_X1 U6959 ( .B1(n20377), .B2(n19918), .A(n2408), .ZN(n3329) );
  NAND2_X1 U6960 ( .A1(n1262), .A2(n19918), .ZN(n2408) );
  NAND2_X1 U6961 ( .A1(n17592), .A2(n20150), .ZN(n17593) );
  INV_X1 U6962 ( .A(n20141), .ZN(n2412) );
  NAND2_X1 U6963 ( .A1(n19361), .A2(n19366), .ZN(n2414) );
  NAND2_X1 U6964 ( .A1(n2415), .A2(n5686), .ZN(n5183) );
  NAND2_X1 U6965 ( .A1(n6084), .A2(n5683), .ZN(n2415) );
  AND3_X1 U6966 ( .A1(n5485), .A2(n5486), .A3(n5487), .ZN(n3746) );
  INV_X1 U6967 ( .A(n10897), .ZN(n11210) );
  INV_X1 U6968 ( .A(n5888), .ZN(n5309) );
  OR2_X1 U6969 ( .A1(n14823), .A2(n12931), .ZN(n3442) );
  INV_X1 U6970 ( .A(n14556), .ZN(n14677) );
  INV_X1 U6971 ( .A(n5720), .ZN(n3086) );
  OAI21_X1 U6972 ( .B1(n2419), .B2(n20146), .A(n2418), .ZN(n9133) );
  OAI21_X1 U6973 ( .B1(n11482), .B2(n11211), .A(n10059), .ZN(n11073) );
  OAI21_X1 U6974 ( .B1(n17496), .B2(n17495), .A(n2421), .ZN(n3217) );
  NAND2_X1 U6975 ( .A1(n2422), .A2(n17495), .ZN(n2421) );
  INV_X1 U6976 ( .A(n14722), .ZN(n13671) );
  XNOR2_X1 U6977 ( .A(n2542), .B(n16695), .ZN(n16835) );
  INV_X1 U6978 ( .A(n6744), .ZN(n6552) );
  INV_X1 U6979 ( .A(n9564), .ZN(n9342) );
  XNOR2_X1 U6980 ( .A(n13697), .B(n12448), .ZN(n12458) );
  INV_X1 U6981 ( .A(n8905), .ZN(n3493) );
  NAND2_X1 U6982 ( .A1(n8720), .A2(n9354), .ZN(n8905) );
  OAI211_X2 U6983 ( .C1(n6656), .C2(n6655), .A(n3288), .B(n2425), .ZN(n10445)
         );
  INV_X1 U6984 ( .A(n15744), .ZN(n15749) );
  NAND2_X1 U6985 ( .A1(n15593), .A2(n19502), .ZN(n15744) );
  NAND2_X1 U6987 ( .A1(n2429), .A2(n2427), .ZN(n2426) );
  NAND2_X1 U6988 ( .A1(n12207), .A2(n2428), .ZN(n2427) );
  INV_X1 U6989 ( .A(n12209), .ZN(n2428) );
  NAND2_X1 U6990 ( .A1(n12189), .A2(n12209), .ZN(n2429) );
  XNOR2_X1 U6991 ( .A(n2430), .B(n19853), .ZN(n8936) );
  XNOR2_X1 U6992 ( .A(n10039), .B(n17637), .ZN(n2430) );
  INV_X1 U6993 ( .A(n9241), .ZN(n8628) );
  INV_X1 U6994 ( .A(n12350), .ZN(n2737) );
  NAND2_X1 U6995 ( .A1(n12467), .A2(n12138), .ZN(n2431) );
  NAND2_X1 U6996 ( .A1(n12139), .A2(n12466), .ZN(n2432) );
  NOR2_X1 U6997 ( .A1(n14327), .A2(n14087), .ZN(n14819) );
  XNOR2_X1 U6998 ( .A(n2433), .B(n7162), .ZN(n7167) );
  XNOR2_X1 U6999 ( .A(n7161), .B(n7202), .ZN(n2433) );
  AND2_X2 U7000 ( .A1(n16663), .A2(n16664), .ZN(n19453) );
  OAI21_X1 U7001 ( .B1(n2435), .B2(n2434), .A(n5945), .ZN(n5461) );
  INV_X1 U7003 ( .A(n15449), .ZN(n2438) );
  NAND2_X1 U7004 ( .A1(n2606), .A2(n10858), .ZN(n2602) );
  NAND2_X1 U7005 ( .A1(n15111), .A2(n15294), .ZN(n15108) );
  NAND2_X1 U7006 ( .A1(n8135), .A2(n8382), .ZN(n7498) );
  AOI21_X1 U7008 ( .B1(n3503), .B2(n9215), .A(n9210), .ZN(n3502) );
  NAND2_X1 U7009 ( .A1(n18172), .A2(n19766), .ZN(n18812) );
  NAND2_X1 U7010 ( .A1(n9242), .A2(n2444), .ZN(n2443) );
  OAI22_X1 U7012 ( .A1(n2450), .A2(n2449), .B1(n19435), .B2(n19448), .ZN(
        n19438) );
  NOR2_X1 U7013 ( .A1(n3828), .A2(n19434), .ZN(n2449) );
  NOR2_X1 U7014 ( .A1(n3769), .A2(n4499), .ZN(n2585) );
  INV_X1 U7015 ( .A(n10833), .ZN(n10837) );
  NAND3_X1 U7016 ( .A1(n2936), .A2(n5346), .A3(n3745), .ZN(n4376) );
  INV_X1 U7017 ( .A(n11527), .ZN(n2470) );
  NAND2_X1 U7018 ( .A1(n3053), .A2(n8054), .ZN(n6211) );
  NAND2_X1 U7019 ( .A1(n16210), .A2(n16790), .ZN(n16211) );
  NAND2_X1 U7020 ( .A1(n7606), .A2(n8185), .ZN(n8182) );
  NAND2_X1 U7021 ( .A1(n3180), .A2(n14358), .ZN(n2451) );
  OAI21_X1 U7023 ( .B1(n15811), .B2(n15815), .A(n3374), .ZN(n15819) );
  NOR2_X1 U7024 ( .A1(n8055), .A2(n8192), .ZN(n3054) );
  AOI22_X1 U7025 ( .A1(n10825), .A2(n11489), .B1(n10824), .B2(n11069), .ZN(
        n12061) );
  OR3_X1 U7027 ( .A1(n8993), .A2(n9274), .A3(n20265), .ZN(n9279) );
  NAND2_X1 U7029 ( .A1(n9115), .A2(n9218), .ZN(n9116) );
  OAI21_X1 U7032 ( .B1(n14439), .B2(n14441), .A(n238), .ZN(n13557) );
  NAND2_X1 U7033 ( .A1(n8201), .A2(n8070), .ZN(n8072) );
  NAND2_X1 U7034 ( .A1(n2458), .A2(n11173), .ZN(n3359) );
  OAI21_X1 U7035 ( .B1(n3789), .B2(n11174), .A(n3362), .ZN(n2458) );
  NAND2_X1 U7036 ( .A1(n3358), .A2(n2457), .ZN(n12224) );
  OR2_X1 U7037 ( .A1(n11176), .A2(n2458), .ZN(n2457) );
  OAI21_X1 U7040 ( .B1(n6013), .B2(n6007), .A(n6011), .ZN(n5208) );
  INV_X1 U7041 ( .A(n5098), .ZN(n2460) );
  INV_X1 U7042 ( .A(n5092), .ZN(n2461) );
  AND2_X1 U7043 ( .A1(n5092), .A2(n5093), .ZN(n2462) );
  NAND3_X1 U7044 ( .A1(n2464), .A2(n11080), .A3(n2463), .ZN(n12258) );
  NAND3_X1 U7045 ( .A1(n11077), .A2(n11474), .A3(n11079), .ZN(n2463) );
  NAND2_X1 U7046 ( .A1(n3507), .A2(n11076), .ZN(n11079) );
  NAND3_X1 U7047 ( .A1(n2466), .A2(n5311), .A3(n5144), .ZN(n2465) );
  INV_X1 U7048 ( .A(n5781), .ZN(n2467) );
  NAND2_X1 U7049 ( .A1(n11530), .A2(n11528), .ZN(n2469) );
  NAND2_X1 U7050 ( .A1(n15626), .A2(n2472), .ZN(n2471) );
  NAND2_X1 U7051 ( .A1(n15840), .A2(n15625), .ZN(n15626) );
  NAND2_X1 U7052 ( .A1(n2475), .A2(n2473), .ZN(n2797) );
  NAND2_X1 U7053 ( .A1(n2474), .A2(n18130), .ZN(n2473) );
  NAND2_X1 U7054 ( .A1(n18131), .A2(n17946), .ZN(n2474) );
  INV_X1 U7055 ( .A(n19974), .ZN(n2475) );
  NAND4_X2 U7056 ( .A1(n7662), .A2(n2479), .A3(n7660), .A4(n2478), .ZN(n10163)
         );
  NAND2_X1 U7057 ( .A1(n8747), .A2(n8932), .ZN(n8924) );
  NAND2_X1 U7059 ( .A1(n4491), .A2(n4899), .ZN(n2480) );
  AND2_X1 U7060 ( .A1(n4883), .A2(n2482), .ZN(n2481) );
  NAND2_X1 U7061 ( .A1(n2483), .A2(n2487), .ZN(n11892) );
  NAND2_X1 U7062 ( .A1(n2484), .A2(n2486), .ZN(n2483) );
  INV_X1 U7063 ( .A(n11119), .ZN(n2486) );
  NAND2_X1 U7064 ( .A1(n11036), .A2(n11119), .ZN(n2487) );
  INV_X1 U7066 ( .A(Plaintext[17]), .ZN(n2488) );
  NAND2_X1 U7067 ( .A1(n4986), .A2(n2489), .ZN(n4991) );
  INV_X1 U7068 ( .A(n4302), .ZN(n2490) );
  NAND2_X1 U7069 ( .A1(n12513), .A2(n10625), .ZN(n13270) );
  NAND2_X1 U7071 ( .A1(n13275), .A2(n20073), .ZN(n2491) );
  NAND2_X1 U7072 ( .A1(n2493), .A2(n5455), .ZN(n2559) );
  NAND4_X2 U7073 ( .A1(n5173), .A2(n2493), .A3(n5175), .A4(n5174), .ZN(n6634)
         );
  NAND2_X1 U7074 ( .A1(n6108), .A2(n5656), .ZN(n2493) );
  XNOR2_X1 U7075 ( .A(n10569), .B(n10573), .ZN(n2495) );
  NAND2_X1 U7076 ( .A1(n2499), .A2(n8790), .ZN(n7928) );
  NAND2_X1 U7077 ( .A1(n9148), .A2(n2499), .ZN(n8785) );
  NOR2_X1 U7078 ( .A1(n9148), .A2(n2499), .ZN(n9150) );
  NAND2_X1 U7079 ( .A1(n20019), .A2(n17886), .ZN(n17665) );
  AND2_X1 U7080 ( .A1(n20019), .A2(n19947), .ZN(n17599) );
  NAND2_X1 U7081 ( .A1(n3247), .A2(n2500), .ZN(n14888) );
  NAND2_X1 U7082 ( .A1(n2501), .A2(n9145), .ZN(n7929) );
  NAND3_X1 U7083 ( .A1(n9145), .A2(n8786), .A3(n2501), .ZN(n8787) );
  XNOR2_X1 U7084 ( .A(n9960), .B(n2505), .ZN(n9324) );
  INV_X1 U7085 ( .A(n10026), .ZN(n2505) );
  OR2_X1 U7086 ( .A1(n17094), .A2(n2507), .ZN(n2513) );
  NAND2_X1 U7087 ( .A1(n2517), .A2(n17095), .ZN(n2507) );
  NAND2_X1 U7088 ( .A1(n17092), .A2(n212), .ZN(n2517) );
  OAI21_X1 U7089 ( .B1(n2508), .B2(n17094), .A(n2511), .ZN(n2510) );
  INV_X1 U7090 ( .A(n2517), .ZN(n2508) );
  OAI211_X1 U7091 ( .C1(n2513), .C2(n2512), .A(n2510), .B(n2509), .ZN(
        Ciphertext[190]) );
  INV_X1 U7092 ( .A(n17095), .ZN(n2511) );
  INV_X1 U7093 ( .A(n2514), .ZN(n2512) );
  NAND2_X1 U7094 ( .A1(n2516), .A2(n2515), .ZN(n2514) );
  XNOR2_X1 U7095 ( .A(n12559), .B(n2518), .ZN(n2519) );
  XNOR2_X1 U7096 ( .A(n12826), .B(n12027), .ZN(n13213) );
  XNOR2_X1 U7097 ( .A(n12826), .B(n2521), .ZN(n2520) );
  NAND2_X1 U7099 ( .A1(n2523), .A2(n12389), .ZN(n12391) );
  OAI211_X1 U7100 ( .C1(n245), .C2(n2523), .A(n12389), .B(n11313), .ZN(n11314)
         );
  NAND2_X1 U7101 ( .A1(n12757), .A2(n2523), .ZN(n12758) );
  NAND2_X1 U7102 ( .A1(n19404), .A2(n17650), .ZN(n2527) );
  INV_X1 U7104 ( .A(n15636), .ZN(n2530) );
  XNOR2_X1 U7105 ( .A(n2531), .B(n17686), .ZN(Ciphertext[164]) );
  OAI211_X1 U7106 ( .C1(n20444), .C2(n19261), .A(n2534), .B(n2532), .ZN(n2531)
         );
  OAI211_X1 U7107 ( .C1(n2816), .C2(n19269), .A(n2533), .B(n19267), .ZN(n2532)
         );
  NAND2_X1 U7108 ( .A1(n17685), .A2(n19276), .ZN(n2534) );
  XNOR2_X1 U7110 ( .A(n13259), .B(n13602), .ZN(n12834) );
  NAND2_X1 U7112 ( .A1(n12393), .A2(n12479), .ZN(n2538) );
  INV_X1 U7113 ( .A(n7935), .ZN(n2540) );
  NAND2_X1 U7114 ( .A1(n2540), .A2(n20359), .ZN(n7930) );
  XNOR2_X1 U7117 ( .A(n2542), .B(n16980), .ZN(n16756) );
  XNOR2_X1 U7118 ( .A(n16507), .B(n20121), .ZN(n16142) );
  XNOR2_X1 U7119 ( .A(n20121), .B(n16081), .ZN(n16083) );
  NAND3_X1 U7120 ( .A1(n19802), .A2(n7879), .A3(n3055), .ZN(n2543) );
  OAI21_X1 U7121 ( .B1(n2546), .B2(n18409), .A(n18408), .ZN(n18411) );
  NAND2_X1 U7122 ( .A1(n8325), .A2(n2548), .ZN(n7442) );
  AOI21_X1 U7123 ( .B1(n7590), .B2(n2548), .A(n8322), .ZN(n3221) );
  OAI211_X2 U7125 ( .C1(n2553), .C2(n12394), .A(n2549), .B(n2554), .ZN(n13528)
         );
  NAND3_X1 U7126 ( .A1(n2552), .A2(n2551), .A3(n2550), .ZN(n2549) );
  NAND2_X1 U7127 ( .A1(n11931), .A2(n12478), .ZN(n2551) );
  NAND2_X1 U7128 ( .A1(n12141), .A2(n12480), .ZN(n12394) );
  NAND2_X1 U7129 ( .A1(n11932), .A2(n11931), .ZN(n2554) );
  OR2_X1 U7130 ( .A1(n5458), .A2(n6097), .ZN(n2555) );
  NAND2_X1 U7131 ( .A1(n1011), .A2(n6097), .ZN(n2556) );
  XNOR2_X1 U7132 ( .A(n7070), .B(n2557), .ZN(n6225) );
  NAND3_X1 U7133 ( .A1(n2559), .A2(n2560), .A3(n2558), .ZN(n2557) );
  NAND3_X1 U7134 ( .A1(n6108), .A2(n5656), .A3(n6109), .ZN(n2560) );
  OAI21_X2 U7136 ( .B1(n13875), .B2(n13874), .A(n13873), .ZN(n15496) );
  XNOR2_X2 U7137 ( .A(n10364), .B(n10363), .ZN(n11110) );
  XNOR2_X2 U7139 ( .A(n10355), .B(n10354), .ZN(n11452) );
  NAND2_X1 U7142 ( .A1(n3386), .A2(n7820), .ZN(n3384) );
  MUX2_X1 U7143 ( .A(n3387), .B(n3386), .S(n7820), .Z(n2561) );
  NOR2_X1 U7144 ( .A1(n981), .A2(n2562), .ZN(n11831) );
  NOR2_X1 U7145 ( .A1(n13973), .A2(n2563), .ZN(n2564) );
  NAND2_X1 U7146 ( .A1(n2566), .A2(n20443), .ZN(n2565) );
  NAND2_X1 U7147 ( .A1(n2568), .A2(n2567), .ZN(n2566) );
  NAND2_X1 U7148 ( .A1(n951), .A2(n14525), .ZN(n2567) );
  NAND2_X1 U7149 ( .A1(n19634), .A2(n14648), .ZN(n2568) );
  XNOR2_X1 U7150 ( .A(n20216), .B(n7035), .ZN(n7229) );
  XNOR2_X1 U7151 ( .A(n20216), .B(n6735), .ZN(n6423) );
  XNOR2_X1 U7152 ( .A(n20216), .B(n7360), .ZN(n7362) );
  INV_X1 U7154 ( .A(n5611), .ZN(n6151) );
  NAND2_X1 U7155 ( .A1(n2576), .A2(n2595), .ZN(n2572) );
  NAND2_X1 U7157 ( .A1(n2579), .A2(n20533), .ZN(n2577) );
  NAND2_X1 U7158 ( .A1(n2580), .A2(n15905), .ZN(n2579) );
  NAND2_X1 U7159 ( .A1(n15907), .A2(n15909), .ZN(n2580) );
  INV_X1 U7162 ( .A(n13838), .ZN(n2582) );
  NAND3_X1 U7163 ( .A1(n2583), .A2(n6153), .A3(n6150), .ZN(n5614) );
  NAND2_X1 U7164 ( .A1(n5611), .A2(n5349), .ZN(n2583) );
  NAND2_X1 U7165 ( .A1(n4379), .A2(n4857), .ZN(n2584) );
  OR2_X1 U7166 ( .A1(n19933), .A2(n17812), .ZN(n17690) );
  NAND2_X1 U7167 ( .A1(n2587), .A2(n18046), .ZN(n17317) );
  NAND2_X1 U7168 ( .A1(n19933), .A2(n17812), .ZN(n2587) );
  INV_X1 U7173 ( .A(n17812), .ZN(n2590) );
  NAND2_X1 U7174 ( .A1(n2592), .A2(n14787), .ZN(n2591) );
  NAND2_X1 U7175 ( .A1(n14343), .A2(n14790), .ZN(n2593) );
  NAND2_X1 U7176 ( .A1(n14103), .A2(n14791), .ZN(n2594) );
  NAND2_X1 U7177 ( .A1(n4377), .A2(n4899), .ZN(n2595) );
  NAND2_X1 U7178 ( .A1(n20205), .A2(n4960), .ZN(n2596) );
  NAND2_X1 U7180 ( .A1(n20057), .A2(n19865), .ZN(n2597) );
  NAND2_X1 U7181 ( .A1(n2598), .A2(n12542), .ZN(n12547) );
  INV_X1 U7182 ( .A(n12545), .ZN(n2598) );
  NOR2_X1 U7183 ( .A1(n2601), .A2(n3978), .ZN(n3977) );
  INV_X1 U7184 ( .A(n4657), .ZN(n2601) );
  NAND2_X1 U7185 ( .A1(n2603), .A2(n2602), .ZN(n12619) );
  NAND2_X1 U7186 ( .A1(n2610), .A2(n10858), .ZN(n2603) );
  NAND2_X1 U7187 ( .A1(n2604), .A2(n894), .ZN(n2608) );
  NAND2_X1 U7189 ( .A1(n2607), .A2(n10858), .ZN(n12057) );
  NAND3_X1 U7190 ( .A1(n12059), .A2(n12053), .A3(n2608), .ZN(n11634) );
  AOI21_X1 U7191 ( .B1(n2612), .B2(n11773), .A(n3260), .ZN(n11774) );
  NAND2_X1 U7192 ( .A1(n12313), .A2(n12148), .ZN(n2612) );
  OAI21_X1 U7193 ( .B1(n6069), .B2(n5879), .A(n2613), .ZN(n5883) );
  NAND3_X1 U7194 ( .A1(n6069), .A2(n6075), .A3(n6067), .ZN(n2613) );
  NAND2_X1 U7195 ( .A1(n6069), .A2(n6067), .ZN(n2616) );
  NAND2_X1 U7196 ( .A1(n2616), .A2(n6070), .ZN(n2614) );
  NAND2_X1 U7197 ( .A1(n5979), .A2(n5320), .ZN(n2615) );
  NAND2_X1 U7198 ( .A1(n969), .A2(n2617), .ZN(n9643) );
  XNOR2_X1 U7199 ( .A(n10594), .B(n10105), .ZN(n10106) );
  XNOR2_X1 U7200 ( .A(n2619), .B(n12862), .ZN(n14452) );
  XNOR2_X1 U7201 ( .A(n13708), .B(n2620), .ZN(n2619) );
  XNOR2_X1 U7202 ( .A(n2621), .B(n6659), .ZN(n2622) );
  INV_X1 U7203 ( .A(n6588), .ZN(n2621) );
  XNOR2_X1 U7205 ( .A(n13771), .B(n13769), .ZN(n2624) );
  NAND2_X1 U7206 ( .A1(n8644), .A2(n8937), .ZN(n2955) );
  OAI211_X1 U7207 ( .C1(n15885), .C2(n2625), .A(n16017), .B(n14926), .ZN(
        n14927) );
  NAND2_X1 U7208 ( .A1(n16012), .A2(n19740), .ZN(n2625) );
  NAND2_X1 U7209 ( .A1(n2627), .A2(n8018), .ZN(n7804) );
  INV_X1 U7210 ( .A(n14584), .ZN(n2628) );
  NAND2_X1 U7211 ( .A1(n2629), .A2(n6166), .ZN(n5462) );
  MUX2_X1 U7212 ( .A(n1867), .B(n170), .S(n6172), .Z(n4692) );
  NAND2_X1 U7213 ( .A1(n5843), .A2(n2630), .ZN(n7274) );
  NOR2_X1 U7214 ( .A1(n9135), .A2(n2727), .ZN(n2631) );
  OR2_X1 U7215 ( .A1(n5073), .A2(n291), .ZN(n4662) );
  INV_X1 U7216 ( .A(n4816), .ZN(n2632) );
  NAND2_X1 U7217 ( .A1(n20168), .A2(n19814), .ZN(n16442) );
  NAND2_X1 U7218 ( .A1(n2634), .A2(n9218), .ZN(n8429) );
  INV_X1 U7219 ( .A(n9118), .ZN(n2634) );
  NAND2_X1 U7220 ( .A1(n9217), .A2(n9221), .ZN(n9118) );
  AOI22_X1 U7221 ( .A1(n267), .A2(n9189), .B1(n8713), .B2(n9241), .ZN(n9243)
         );
  NAND2_X1 U7223 ( .A1(n2637), .A2(n6587), .ZN(n2636) );
  NAND2_X1 U7224 ( .A1(n987), .A2(n5328), .ZN(n2638) );
  NAND2_X1 U7225 ( .A1(n2641), .A2(n5328), .ZN(n2640) );
  NOR2_X1 U7228 ( .A1(n15297), .A2(n15111), .ZN(n2645) );
  OR2_X1 U7229 ( .A1(n15108), .A2(n15109), .ZN(n2646) );
  INV_X1 U7230 ( .A(n12047), .ZN(n2647) );
  NAND2_X1 U7231 ( .A1(n2647), .A2(n12122), .ZN(n11647) );
  INV_X1 U7232 ( .A(n12047), .ZN(n12229) );
  NAND2_X1 U7234 ( .A1(n3156), .A2(n14746), .ZN(n3155) );
  OAI21_X1 U7235 ( .B1(n8183), .B2(n8059), .A(n2648), .ZN(n8065) );
  NAND2_X1 U7236 ( .A1(n4730), .A2(n2649), .ZN(n2648) );
  NAND2_X1 U7237 ( .A1(n19716), .A2(n8630), .ZN(n2652) );
  OR2_X1 U7238 ( .A1(n13911), .A2(n13907), .ZN(n2654) );
  NOR2_X1 U7239 ( .A1(n15857), .A2(n2655), .ZN(n15858) );
  AOI22_X1 U7240 ( .A1(n15722), .A2(n15864), .B1(n15721), .B2(n2655), .ZN(
        n13916) );
  NAND2_X1 U7241 ( .A1(n15859), .A2(n2655), .ZN(n15725) );
  INV_X1 U7243 ( .A(n10450), .ZN(n11094) );
  NAND3_X1 U7246 ( .A1(n2662), .A2(n2664), .A3(n2660), .ZN(n16810) );
  NAND2_X1 U7247 ( .A1(n2661), .A2(n19658), .ZN(n2660) );
  NAND3_X1 U7248 ( .A1(n17552), .A2(n18103), .A3(n2665), .ZN(n2664) );
  OR2_X1 U7249 ( .A1(n17959), .A2(n17954), .ZN(n2665) );
  INV_X1 U7250 ( .A(n16805), .ZN(n18105) );
  NAND2_X1 U7251 ( .A1(n6096), .A2(n6101), .ZN(n3589) );
  NAND2_X1 U7253 ( .A1(n3685), .A2(n2682), .ZN(n2666) );
  NAND2_X1 U7254 ( .A1(n19354), .A2(n20244), .ZN(n2668) );
  AOI21_X2 U7255 ( .B1(n15929), .B2(n2669), .A(n15928), .ZN(n18423) );
  NOR2_X1 U7256 ( .A1(n4797), .A2(n5047), .ZN(n2671) );
  NAND2_X1 U7257 ( .A1(n2675), .A2(n2677), .ZN(n2673) );
  NOR2_X1 U7259 ( .A1(n15870), .A2(n15876), .ZN(n15873) );
  MUX2_X1 U7260 ( .A(n14664), .B(n14316), .S(n14662), .Z(n2678) );
  XNOR2_X1 U7261 ( .A(n13842), .B(n1004), .ZN(n2679) );
  NAND2_X1 U7262 ( .A1(n2680), .A2(n11475), .ZN(n3135) );
  NAND2_X1 U7263 ( .A1(n984), .A2(n2682), .ZN(n2681) );
  NAND2_X1 U7267 ( .A1(n5662), .A2(n6101), .ZN(n5948) );
  INV_X1 U7268 ( .A(n8095), .ZN(n2687) );
  OAI21_X1 U7269 ( .B1(n8094), .B2(n8211), .A(n2686), .ZN(n2688) );
  NAND2_X1 U7270 ( .A1(n2687), .A2(n8212), .ZN(n2686) );
  XNOR2_X2 U7271 ( .A(n6609), .B(n6608), .ZN(n8212) );
  XNOR2_X1 U7272 ( .A(n10351), .B(n2689), .ZN(n9724) );
  NAND2_X1 U7273 ( .A1(n8759), .A2(n8650), .ZN(n2690) );
  NAND2_X1 U7277 ( .A1(n14348), .A2(n19496), .ZN(n2695) );
  NAND2_X1 U7278 ( .A1(n14349), .A2(n19985), .ZN(n2698) );
  NAND2_X1 U7279 ( .A1(n4089), .A2(n2701), .ZN(n2699) );
  NAND2_X1 U7281 ( .A1(n4697), .A2(n5040), .ZN(n4799) );
  AND2_X1 U7282 ( .A1(n4440), .A2(n4439), .ZN(n2701) );
  OAI21_X1 U7283 ( .B1(n11469), .B2(n11568), .A(n2705), .ZN(n2704) );
  AOI21_X1 U7284 ( .B1(n10883), .B2(n11568), .A(n11566), .ZN(n2705) );
  XNOR2_X2 U7285 ( .A(n9951), .B(n9950), .ZN(n11568) );
  NAND2_X1 U7286 ( .A1(n2707), .A2(n12352), .ZN(n3330) );
  INV_X1 U7287 ( .A(n12353), .ZN(n2707) );
  XNOR2_X1 U7290 ( .A(n12713), .B(n2709), .ZN(n12728) );
  MUX2_X1 U7291 ( .A(n7969), .B(n7970), .S(n7922), .Z(n7977) );
  NAND2_X1 U7292 ( .A1(n2714), .A2(n2711), .ZN(n10849) );
  NAND2_X1 U7293 ( .A1(n15838), .A2(n15625), .ZN(n2715) );
  INV_X1 U7294 ( .A(n5279), .ZN(n3398) );
  NAND2_X1 U7295 ( .A1(n5669), .A2(n5425), .ZN(n2719) );
  OAI22_X1 U7296 ( .A1(n14340), .A2(n13931), .B1(n14337), .B2(n14342), .ZN(
        n3331) );
  NAND2_X1 U7297 ( .A1(n2722), .A2(n20533), .ZN(n2721) );
  NAND2_X1 U7298 ( .A1(n2725), .A2(n11395), .ZN(n11401) );
  MUX2_X1 U7299 ( .A(n10859), .B(n10860), .S(n11399), .Z(n10861) );
  NAND3_X1 U7300 ( .A1(n9214), .A2(n9209), .A3(n263), .ZN(n8394) );
  NAND3_X1 U7301 ( .A1(n2731), .A2(n14620), .A3(n14192), .ZN(n2730) );
  INV_X1 U7302 ( .A(n14627), .ZN(n2731) );
  XNOR2_X1 U7303 ( .A(n13295), .B(n2733), .ZN(n13135) );
  OR2_X1 U7304 ( .A1(n12469), .A2(n12470), .ZN(n2732) );
  XNOR2_X1 U7305 ( .A(n13063), .B(n855), .ZN(n13400) );
  XNOR2_X1 U7306 ( .A(n855), .B(n13848), .ZN(n13851) );
  XNOR2_X1 U7307 ( .A(n13343), .B(n2733), .ZN(n12864) );
  INV_X1 U7308 ( .A(n10694), .ZN(n10995) );
  NAND2_X1 U7310 ( .A1(n19817), .A2(n19779), .ZN(n2734) );
  OAI21_X1 U7312 ( .B1(n19651), .B2(n7743), .A(n2751), .ZN(n7742) );
  AOI22_X2 U7314 ( .A1(n7744), .A2(n7743), .B1(n7742), .B2(n7741), .ZN(n7752)
         );
  NAND2_X1 U7315 ( .A1(n11535), .A2(n11538), .ZN(n2736) );
  OAI21_X1 U7316 ( .B1(n11170), .B2(n11535), .A(n2736), .ZN(n8902) );
  INV_X1 U7317 ( .A(Plaintext[79]), .ZN(n2738) );
  NAND2_X1 U7318 ( .A1(n3904), .A2(n4554), .ZN(n5015) );
  NAND2_X1 U7319 ( .A1(n3905), .A2(n2740), .ZN(n2739) );
  NAND2_X1 U7320 ( .A1(n5021), .A2(n5018), .ZN(n2740) );
  NAND2_X1 U7321 ( .A1(n3904), .A2(n4555), .ZN(n5021) );
  AOI21_X2 U7322 ( .B1(n15493), .B2(n15587), .A(n2741), .ZN(n17109) );
  MUX2_X1 U7323 ( .A(n15492), .B(n15761), .S(n15760), .Z(n2741) );
  NAND2_X1 U7324 ( .A1(n12209), .A2(n12211), .ZN(n2742) );
  XNOR2_X1 U7325 ( .A(n9852), .B(n10182), .ZN(n2745) );
  NAND2_X1 U7326 ( .A1(n8733), .A2(n8736), .ZN(n8920) );
  NAND2_X1 U7327 ( .A1(n8733), .A2(n8735), .ZN(n8332) );
  NAND2_X1 U7328 ( .A1(n14706), .A2(n20113), .ZN(n14564) );
  AOI21_X1 U7329 ( .B1(n14704), .B2(n20113), .A(n14563), .ZN(n14111) );
  NOR2_X1 U7330 ( .A1(n919), .A2(n20113), .ZN(n14709) );
  OAI21_X1 U7331 ( .B1(n9318), .B2(n2749), .A(n9320), .ZN(n9319) );
  NOR2_X1 U7332 ( .A1(n8860), .A2(n2749), .ZN(n8864) );
  NAND2_X1 U7333 ( .A1(n9322), .A2(n2749), .ZN(n9838) );
  NAND2_X1 U7334 ( .A1(n8354), .A2(n7739), .ZN(n2751) );
  NAND2_X1 U7335 ( .A1(n2754), .A2(n2753), .ZN(n17309) );
  OR2_X1 U7336 ( .A1(n18221), .A2(n18016), .ZN(n2753) );
  NAND2_X1 U7337 ( .A1(n17308), .A2(n18221), .ZN(n2754) );
  OAI21_X1 U7338 ( .B1(n224), .B2(n20421), .A(n18977), .ZN(n18980) );
  OAI21_X1 U7339 ( .B1(n18224), .B2(n18223), .A(n20421), .ZN(n18721) );
  NAND2_X1 U7340 ( .A1(n9353), .A2(n8904), .ZN(n9357) );
  INV_X1 U7341 ( .A(n8720), .ZN(n9353) );
  OAI21_X1 U7342 ( .B1(n12600), .B2(n12606), .A(n2757), .ZN(n11630) );
  NAND2_X1 U7343 ( .A1(n12609), .A2(n12600), .ZN(n2757) );
  NAND2_X1 U7344 ( .A1(n2762), .A2(n12241), .ZN(n12620) );
  INV_X1 U7345 ( .A(n12619), .ZN(n2762) );
  XNOR2_X1 U7346 ( .A(n2763), .B(n13735), .ZN(n13313) );
  INV_X1 U7347 ( .A(n13120), .ZN(n2763) );
  XNOR2_X1 U7348 ( .A(n13792), .B(n2764), .ZN(n13793) );
  NAND2_X1 U7349 ( .A1(n10818), .A2(n10677), .ZN(n11369) );
  NOR2_X1 U7350 ( .A1(n10676), .A2(n10677), .ZN(n9875) );
  INV_X1 U7351 ( .A(n14229), .ZN(n2769) );
  NAND2_X1 U7353 ( .A1(n2769), .A2(n14381), .ZN(n2767) );
  NAND2_X1 U7354 ( .A1(n14697), .A2(n14232), .ZN(n2768) );
  NAND2_X1 U7355 ( .A1(n19503), .A2(n14381), .ZN(n14697) );
  XNOR2_X1 U7357 ( .A(n10165), .B(n20176), .ZN(n2771) );
  XNOR2_X1 U7358 ( .A(n9586), .B(n9588), .ZN(n2772) );
  NAND2_X1 U7359 ( .A1(n13919), .A2(n14167), .ZN(n2774) );
  AOI21_X1 U7362 ( .B1(n8568), .B2(n9168), .A(n9082), .ZN(n2777) );
  NAND2_X1 U7364 ( .A1(n235), .A2(n14818), .ZN(n14823) );
  XNOR2_X1 U7365 ( .A(n12824), .B(n12823), .ZN(n2784) );
  NAND2_X1 U7368 ( .A1(n2787), .A2(n9297), .ZN(n2786) );
  NOR2_X1 U7369 ( .A1(n8846), .A2(n9018), .ZN(n2787) );
  NAND2_X1 U7370 ( .A1(n11208), .A2(n2788), .ZN(n12142) );
  NAND2_X1 U7371 ( .A1(n958), .A2(n11445), .ZN(n2788) );
  NAND2_X1 U7373 ( .A1(n15406), .A2(n15547), .ZN(n2791) );
  NAND2_X1 U7374 ( .A1(n15546), .A2(n15071), .ZN(n15616) );
  NAND2_X1 U7375 ( .A1(n15618), .A2(n15405), .ZN(n15547) );
  NAND2_X1 U7376 ( .A1(n8305), .A2(n2792), .ZN(n8306) );
  OAI211_X1 U7377 ( .C1(n8303), .C2(n8301), .A(n8044), .B(n2792), .ZN(n7599)
         );
  NAND2_X1 U7379 ( .A1(n5272), .A2(n2792), .ZN(n3718) );
  INV_X1 U7380 ( .A(n20361), .ZN(n2793) );
  OAI21_X1 U7381 ( .B1(n5856), .B2(n5855), .A(n2796), .ZN(n2795) );
  NAND2_X1 U7383 ( .A1(n2799), .A2(n2800), .ZN(n2798) );
  NAND2_X1 U7384 ( .A1(n15072), .A2(n15620), .ZN(n2801) );
  INV_X1 U7385 ( .A(n15546), .ZN(n2803) );
  NAND3_X1 U7386 ( .A1(n19668), .A2(n19682), .A3(n18552), .ZN(n17931) );
  NAND2_X1 U7388 ( .A1(n2809), .A2(n2807), .ZN(n2806) );
  NAND2_X1 U7389 ( .A1(n13888), .A2(n14593), .ZN(n2807) );
  INV_X1 U7390 ( .A(n14590), .ZN(n2808) );
  AND2_X1 U7391 ( .A1(n12544), .A2(n250), .ZN(n3462) );
  AOI21_X2 U7392 ( .B1(n15299), .B2(n15298), .A(n2812), .ZN(n16095) );
  MUX2_X1 U7393 ( .A(n15297), .B(n15296), .S(n15295), .Z(n2813) );
  INV_X1 U7394 ( .A(n15759), .ZN(n2815) );
  NAND3_X1 U7395 ( .A1(n17661), .A2(n17662), .A3(n17890), .ZN(n2817) );
  NAND3_X1 U7396 ( .A1(n17665), .A2(n17661), .A3(n17662), .ZN(n2818) );
  NAND2_X1 U7397 ( .A1(n14027), .A2(n2820), .ZN(n15488) );
  NAND2_X1 U7398 ( .A1(n14574), .A2(n2821), .ZN(n2820) );
  NAND2_X1 U7399 ( .A1(n14268), .A2(n14569), .ZN(n2821) );
  NAND2_X1 U7400 ( .A1(n16262), .A2(n16777), .ZN(n2822) );
  NAND2_X1 U7401 ( .A1(n16264), .A2(n17824), .ZN(n2823) );
  XNOR2_X1 U7403 ( .A(n7079), .B(n6718), .ZN(n2825) );
  OR2_X1 U7409 ( .A1(n18603), .A2(n18630), .ZN(n2830) );
  XNOR2_X1 U7411 ( .A(n13291), .B(n2834), .ZN(n2833) );
  NAND2_X1 U7412 ( .A1(n2837), .A2(n2835), .ZN(n17551) );
  XNOR2_X2 U7413 ( .A(n17115), .B(n17114), .ZN(n18233) );
  NAND2_X1 U7415 ( .A1(n17548), .A2(n19771), .ZN(n2837) );
  NAND2_X1 U7416 ( .A1(n9209), .A2(n2727), .ZN(n9212) );
  NAND3_X1 U7417 ( .A1(n9209), .A2(n9135), .A3(n2727), .ZN(n3454) );
  INV_X1 U7418 ( .A(n14800), .ZN(n14081) );
  AOI21_X1 U7419 ( .B1(n3497), .B2(n14796), .A(n14584), .ZN(n2838) );
  NAND2_X1 U7420 ( .A1(n20380), .A2(n14522), .ZN(n14652) );
  NAND3_X1 U7421 ( .A1(n20380), .A2(n14522), .A3(n19831), .ZN(n2839) );
  XNOR2_X2 U7422 ( .A(n13001), .B(n13000), .ZN(n14522) );
  NOR2_X1 U7423 ( .A1(n2840), .A2(n8162), .ZN(n8163) );
  NAND2_X1 U7426 ( .A1(n19872), .A2(n2843), .ZN(n2842) );
  NOR2_X1 U7427 ( .A1(n11160), .A2(n11161), .ZN(n2843) );
  NAND2_X1 U7428 ( .A1(n11161), .A2(n11155), .ZN(n2846) );
  NAND2_X1 U7429 ( .A1(n2848), .A2(n9366), .ZN(n2847) );
  NAND2_X1 U7431 ( .A1(n9364), .A2(n2849), .ZN(n2848) );
  NAND2_X1 U7432 ( .A1(n8960), .A2(n8961), .ZN(n2849) );
  NAND2_X1 U7433 ( .A1(n8961), .A2(n8500), .ZN(n9364) );
  NAND2_X1 U7434 ( .A1(n9361), .A2(n9362), .ZN(n8727) );
  NAND3_X1 U7435 ( .A1(n3421), .A2(n2853), .A3(n2851), .ZN(Ciphertext[28]) );
  NAND2_X1 U7436 ( .A1(n2852), .A2(n2854), .ZN(n2851) );
  NAND2_X1 U7437 ( .A1(n17639), .A2(n19729), .ZN(n17647) );
  NAND3_X1 U7438 ( .A1(n17639), .A2(n19729), .A3(n15134), .ZN(n2853) );
  NAND2_X1 U7439 ( .A1(n2855), .A2(n893), .ZN(n2854) );
  INV_X1 U7440 ( .A(n17914), .ZN(n2855) );
  NAND2_X1 U7441 ( .A1(n18592), .A2(n18585), .ZN(n18596) );
  INV_X1 U7442 ( .A(n11376), .ZN(n2858) );
  OR2_X1 U7443 ( .A1(n11330), .A2(n11376), .ZN(n2857) );
  INV_X1 U7444 ( .A(n20095), .ZN(n2860) );
  NAND2_X1 U7445 ( .A1(n2860), .A2(n11376), .ZN(n10661) );
  INV_X1 U7446 ( .A(n11328), .ZN(n11378) );
  NOR2_X1 U7447 ( .A1(n14811), .A2(n14810), .ZN(n14588) );
  OAI21_X1 U7449 ( .B1(n14589), .B2(n14590), .A(n14588), .ZN(n14591) );
  NAND2_X1 U7450 ( .A1(n2864), .A2(n12498), .ZN(n2863) );
  NAND2_X1 U7451 ( .A1(n5732), .A2(n5802), .ZN(n2867) );
  INV_X1 U7452 ( .A(n5045), .ZN(n5043) );
  OAI21_X1 U7453 ( .B1(n2872), .B2(n2871), .A(n4796), .ZN(n2870) );
  NOR2_X1 U7454 ( .A1(n4697), .A2(n5040), .ZN(n2871) );
  NOR2_X1 U7455 ( .A1(n3061), .A2(n5045), .ZN(n2874) );
  INV_X1 U7456 ( .A(n20247), .ZN(n8186) );
  MUX2_X1 U7457 ( .A(n20465), .B(n8190), .S(n8061), .Z(n2875) );
  XNOR2_X1 U7458 ( .A(n3902), .B(n7202), .ZN(n3963) );
  NAND2_X1 U7459 ( .A1(n2878), .A2(n2877), .ZN(n2876) );
  NAND2_X1 U7460 ( .A1(n992), .A2(n5429), .ZN(n2877) );
  NAND2_X1 U7461 ( .A1(n2879), .A2(n5793), .ZN(n2878) );
  INV_X1 U7463 ( .A(n13243), .ZN(n2881) );
  OAI21_X1 U7464 ( .B1(n19958), .B2(n15583), .A(n15811), .ZN(n15584) );
  INV_X1 U7465 ( .A(n8995), .ZN(n2883) );
  NAND2_X1 U7466 ( .A1(n19517), .A2(n8997), .ZN(n2884) );
  NAND2_X1 U7467 ( .A1(n11431), .A2(n11430), .ZN(n11042) );
  MUX2_X1 U7469 ( .A(n12269), .B(n12374), .S(n20497), .Z(n11732) );
  NAND2_X1 U7473 ( .A1(n14697), .A2(n2891), .ZN(n2890) );
  AOI22_X1 U7474 ( .A1(n17903), .A2(n17904), .B1(n19229), .B2(n2892), .ZN(
        n17905) );
  AOI22_X1 U7475 ( .A1(n17915), .A2(n19236), .B1(n17916), .B2(n2892), .ZN(
        n17917) );
  OAI22_X1 U7476 ( .A1(n19236), .A2(n20124), .B1(n18190), .B2(n19754), .ZN(
        n2892) );
  NOR2_X1 U7477 ( .A1(n19166), .A2(n2893), .ZN(n17797) );
  NAND2_X1 U7478 ( .A1(n2895), .A2(n2894), .ZN(n2893) );
  NAND2_X1 U7479 ( .A1(n2918), .A2(n17790), .ZN(n2894) );
  AOI21_X1 U7480 ( .B1(n19165), .B2(n17790), .A(n17791), .ZN(n2895) );
  INV_X1 U7481 ( .A(n17791), .ZN(n2896) );
  NAND2_X1 U7483 ( .A1(n10899), .A2(n19897), .ZN(n2899) );
  NAND2_X1 U7484 ( .A1(n11482), .A2(n10746), .ZN(n10898) );
  OAI21_X1 U7485 ( .B1(n12497), .B2(n12499), .A(n2901), .ZN(n12503) );
  INV_X1 U7486 ( .A(n2903), .ZN(n2902) );
  NAND2_X1 U7489 ( .A1(n13953), .A2(n14408), .ZN(n2905) );
  NAND2_X1 U7490 ( .A1(n18957), .A2(n2906), .ZN(n17068) );
  NAND2_X1 U7493 ( .A1(n15509), .A2(n3822), .ZN(n2908) );
  NAND3_X1 U7494 ( .A1(n921), .A2(n15559), .A3(n15509), .ZN(n14765) );
  NOR2_X1 U7495 ( .A1(n15560), .A2(n921), .ZN(n15561) );
  MUX2_X1 U7496 ( .A(n15559), .B(n921), .S(n15558), .Z(n15563) );
  XNOR2_X1 U7499 ( .A(n2913), .B(n2912), .ZN(Ciphertext[142]) );
  INV_X1 U7500 ( .A(n2410), .ZN(n2912) );
  NAND3_X1 U7501 ( .A1(n2917), .A2(n2916), .A3(n2914), .ZN(n2913) );
  OAI211_X1 U7502 ( .C1(n19692), .C2(n19708), .A(n2915), .B(n19948), .ZN(n2914) );
  NAND2_X1 U7503 ( .A1(n19692), .A2(n19154), .ZN(n2915) );
  NAND3_X1 U7504 ( .A1(n195), .A2(n19683), .A3(n19165), .ZN(n2916) );
  NAND2_X1 U7505 ( .A1(n18307), .A2(n2918), .ZN(n2917) );
  AOI21_X1 U7506 ( .B1(n3551), .B2(n2919), .A(n4528), .ZN(n3624) );
  NAND2_X1 U7507 ( .A1(n13557), .A2(n13558), .ZN(n2920) );
  NAND2_X1 U7508 ( .A1(n14442), .A2(n14440), .ZN(n2921) );
  AOI21_X2 U7509 ( .B1(n2927), .B2(n2926), .A(n2922), .ZN(n15559) );
  OAI22_X1 U7510 ( .A1(n2925), .A2(n1527), .B1(n2926), .B2(n2923), .ZN(n2922)
         );
  INV_X1 U7511 ( .A(n14393), .ZN(n2924) );
  NAND2_X1 U7512 ( .A1(n14594), .A2(n19731), .ZN(n2925) );
  NAND2_X1 U7513 ( .A1(n14156), .A2(n14155), .ZN(n2927) );
  NAND2_X1 U7514 ( .A1(n1527), .A2(n14594), .ZN(n14156) );
  INV_X1 U7515 ( .A(n9240), .ZN(n9186) );
  NAND2_X1 U7516 ( .A1(n9266), .A2(n9265), .ZN(n8981) );
  NAND2_X1 U7518 ( .A1(n5056), .A2(n4100), .ZN(n4590) );
  NAND2_X1 U7519 ( .A1(n2929), .A2(n5053), .ZN(n2928) );
  NAND2_X1 U7520 ( .A1(n8358), .A2(n8357), .ZN(n2932) );
  NAND2_X1 U7521 ( .A1(n2935), .A2(n8347), .ZN(n8273) );
  NAND2_X1 U7522 ( .A1(n8272), .A2(n8350), .ZN(n2935) );
  XNOR2_X1 U7523 ( .A(n9811), .B(n9995), .ZN(n2938) );
  MUX2_X1 U7524 ( .A(n11418), .B(n11051), .S(n11417), .Z(n11130) );
  MUX2_X1 U7525 ( .A(n11417), .B(n11051), .S(n205), .Z(n10832) );
  NAND3_X1 U7526 ( .A1(n8707), .A2(n1027), .A3(n2941), .ZN(n9908) );
  XNOR2_X1 U7527 ( .A(n6293), .B(n7232), .ZN(n7057) );
  XNOR2_X1 U7528 ( .A(n6494), .B(n6293), .ZN(n6625) );
  NAND2_X1 U7529 ( .A1(n2944), .A2(n2942), .ZN(n2945) );
  AOI21_X1 U7530 ( .B1(n19197), .B2(n2943), .A(n19189), .ZN(n2942) );
  NAND2_X1 U7531 ( .A1(n19190), .A2(n19202), .ZN(n2944) );
  OAI21_X1 U7532 ( .B1(n8298), .B2(n8040), .A(n1835), .ZN(n5965) );
  NOR2_X1 U7533 ( .A1(n7455), .A2(n1835), .ZN(n8514) );
  NAND2_X1 U7534 ( .A1(n12385), .A2(n2946), .ZN(n3530) );
  NOR2_X1 U7535 ( .A1(n12382), .A2(n11915), .ZN(n2946) );
  NAND2_X1 U7536 ( .A1(n898), .A2(n11568), .ZN(n11565) );
  NAND3_X1 U7537 ( .A1(n20349), .A2(n18111), .A3(n18112), .ZN(n2950) );
  INV_X1 U7539 ( .A(n16016), .ZN(n15885) );
  INV_X1 U7540 ( .A(n16016), .ZN(n3473) );
  XNOR2_X1 U7541 ( .A(n13082), .B(n2953), .ZN(n13083) );
  XNOR2_X1 U7542 ( .A(n12713), .B(n2954), .ZN(n2953) );
  OAI21_X1 U7543 ( .B1(n8004), .B2(n8315), .A(n281), .ZN(n7593) );
  NAND2_X1 U7544 ( .A1(n19690), .A2(n17927), .ZN(n17928) );
  OAI211_X2 U7545 ( .C1(n5303), .C2(n5302), .A(n5301), .B(n2956), .ZN(n7338)
         );
  NAND2_X1 U7546 ( .A1(n2958), .A2(n18568), .ZN(n2957) );
  NOR2_X1 U7547 ( .A1(n18555), .A2(n18565), .ZN(n2958) );
  AND2_X2 U7548 ( .A1(n2959), .A2(n16445), .ZN(n18565) );
  OAI211_X1 U7549 ( .C1(n1060), .C2(n16444), .A(n16797), .B(n16443), .ZN(n2959) );
  INV_X1 U7550 ( .A(n7728), .ZN(n8343) );
  INV_X1 U7551 ( .A(n8166), .ZN(n8340) );
  NAND2_X1 U7552 ( .A1(n2962), .A2(n8166), .ZN(n2961) );
  OAI21_X1 U7553 ( .B1(n7728), .B2(n2964), .A(n20274), .ZN(n2962) );
  INV_X1 U7555 ( .A(n8342), .ZN(n2964) );
  NAND2_X1 U7556 ( .A1(n2966), .A2(n2965), .ZN(n19405) );
  NAND2_X1 U7557 ( .A1(n16496), .A2(n2966), .ZN(n16501) );
  NAND2_X1 U7558 ( .A1(n17606), .A2(n19404), .ZN(n2966) );
  XNOR2_X1 U7560 ( .A(n17002), .B(n16555), .ZN(n17141) );
  AOI22_X1 U7563 ( .A1(n11158), .A2(n11157), .B1(n11156), .B2(n11155), .ZN(
        n12037) );
  INV_X1 U7564 ( .A(n5069), .ZN(n5072) );
  XNOR2_X2 U7565 ( .A(n3836), .B(Key[89]), .ZN(n5069) );
  INV_X1 U7566 ( .A(n5071), .ZN(n2971) );
  NAND2_X1 U7567 ( .A1(n3824), .A2(n2973), .ZN(n15414) );
  OAI21_X1 U7568 ( .B1(n15412), .B2(n2973), .A(n15411), .ZN(n15415) );
  OAI21_X1 U7569 ( .B1(n10855), .B2(n9883), .A(n11230), .ZN(n10873) );
  NAND2_X1 U7571 ( .A1(n14898), .A2(n2974), .ZN(n14900) );
  MUX2_X1 U7572 ( .A(n7958), .B(n7956), .S(n277), .Z(n7962) );
  NAND2_X1 U7573 ( .A1(n8906), .A2(n2976), .ZN(n7959) );
  NAND2_X1 U7574 ( .A1(n7915), .A2(n2975), .ZN(n7839) );
  AND2_X1 U7575 ( .A1(n7956), .A2(n2977), .ZN(n2975) );
  OAI21_X1 U7576 ( .B1(n7835), .B2(n7834), .A(n2977), .ZN(n7837) );
  XNOR2_X1 U7577 ( .A(n7178), .B(n2087), .ZN(n6375) );
  NAND2_X1 U7578 ( .A1(n14236), .A2(n19907), .ZN(n2979) );
  XNOR2_X1 U7579 ( .A(n2980), .B(n1228), .ZN(Ciphertext[64]) );
  AOI22_X1 U7581 ( .A1(n19935), .A2(n18143), .B1(n18144), .B2(n19934), .ZN(
        n2981) );
  NOR2_X1 U7583 ( .A1(n2984), .A2(n9296), .ZN(n3806) );
  INV_X1 U7584 ( .A(n9295), .ZN(n2984) );
  NAND2_X1 U7585 ( .A1(n2985), .A2(n8845), .ZN(n7438) );
  OAI21_X1 U7586 ( .B1(n20472), .B2(n3418), .A(n9018), .ZN(n8522) );
  NAND2_X1 U7587 ( .A1(n995), .A2(n2987), .ZN(n2986) );
  INV_X1 U7588 ( .A(n15379), .ZN(n15163) );
  INV_X1 U7589 ( .A(n9158), .ZN(n9160) );
  NAND2_X1 U7590 ( .A1(n9159), .A2(n8696), .ZN(n2989) );
  XNOR2_X1 U7591 ( .A(n16744), .B(n2993), .ZN(n2992) );
  OAI211_X1 U7593 ( .C1(n3002), .C2(n3000), .A(n2998), .B(n2995), .ZN(
        Ciphertext[176]) );
  NAND4_X1 U7594 ( .A1(n2997), .A2(n17543), .A3(n2996), .A4(n17544), .ZN(n2995) );
  INV_X1 U7595 ( .A(n3004), .ZN(n2997) );
  NAND3_X1 U7596 ( .A1(n2999), .A2(n3003), .A3(n298), .ZN(n2998) );
  INV_X1 U7597 ( .A(n17543), .ZN(n2999) );
  NOR2_X1 U7598 ( .A1(n3004), .A2(n3001), .ZN(n3000) );
  OR2_X1 U7599 ( .A1(n17542), .A2(n17544), .ZN(n3001) );
  XNOR2_X1 U7600 ( .A(n3003), .B(n17544), .ZN(n3002) );
  NAND2_X1 U7601 ( .A1(n19316), .A2(n19340), .ZN(n3003) );
  OAI21_X1 U7602 ( .B1(n19324), .B2(n19955), .A(n17541), .ZN(n3004) );
  NAND2_X1 U7603 ( .A1(n14809), .A2(n19781), .ZN(n3005) );
  NAND2_X1 U7604 ( .A1(n3007), .A2(n8241), .ZN(n8242) );
  INV_X1 U7605 ( .A(n7436), .ZN(n3007) );
  NAND2_X1 U7607 ( .A1(n16684), .A2(n17654), .ZN(n17538) );
  AND2_X1 U7608 ( .A1(n19388), .A2(n20004), .ZN(n16684) );
  AND2_X1 U7609 ( .A1(n3010), .A2(n6113), .ZN(n6110) );
  NAND2_X1 U7610 ( .A1(n4733), .A2(n4732), .ZN(n3009) );
  NAND2_X1 U7611 ( .A1(n3013), .A2(n3011), .ZN(n12414) );
  NAND2_X1 U7612 ( .A1(n12412), .A2(n3012), .ZN(n3011) );
  NAND2_X1 U7613 ( .A1(n12411), .A2(n12754), .ZN(n3013) );
  INV_X1 U7614 ( .A(n11174), .ZN(n3015) );
  AOI21_X1 U7615 ( .B1(n11178), .B2(n3789), .A(n3014), .ZN(n3016) );
  OAI21_X1 U7616 ( .B1(n11176), .B2(n11178), .A(n3015), .ZN(n3014) );
  MUX2_X1 U7617 ( .A(n3018), .B(n11179), .S(n9486), .Z(n3017) );
  NOR2_X1 U7618 ( .A1(n3015), .A2(n11177), .ZN(n3018) );
  NAND2_X1 U7619 ( .A1(n3019), .A2(n15504), .ZN(n15820) );
  OAI21_X1 U7620 ( .B1(n3019), .B2(n14069), .A(n15822), .ZN(n14072) );
  XNOR2_X1 U7621 ( .A(n3021), .B(n6992), .ZN(n3020) );
  XNOR2_X1 U7622 ( .A(n3022), .B(n6991), .ZN(n3021) );
  INV_X1 U7623 ( .A(n7333), .ZN(n3022) );
  AOI22_X2 U7625 ( .A1(n10660), .A2(n11952), .B1(n11828), .B2(n3024), .ZN(
        n13192) );
  NAND2_X1 U7626 ( .A1(n13927), .A2(n1364), .ZN(n3025) );
  INV_X1 U7627 ( .A(n18868), .ZN(n3028) );
  INV_X1 U7628 ( .A(n18868), .ZN(n3031) );
  MUX2_X1 U7630 ( .A(n15873), .B(n15872), .S(n19514), .Z(n15878) );
  XNOR2_X1 U7631 ( .A(n3035), .B(n1780), .ZN(Ciphertext[129]) );
  NAND3_X1 U7632 ( .A1(n20214), .A2(n19109), .A3(n19094), .ZN(n3036) );
  INV_X1 U7633 ( .A(n19089), .ZN(n3038) );
  NAND3_X1 U7634 ( .A1(n18358), .A2(n18341), .A3(n18344), .ZN(n18349) );
  NAND2_X1 U7635 ( .A1(n17236), .A2(n3461), .ZN(n3039) );
  NAND2_X1 U7636 ( .A1(n10103), .A2(n3040), .ZN(n3629) );
  INV_X1 U7637 ( .A(n19949), .ZN(n3040) );
  NAND2_X1 U7638 ( .A1(n14979), .A2(n14978), .ZN(n3041) );
  NAND2_X1 U7639 ( .A1(n6206), .A2(n19492), .ZN(n3044) );
  NAND2_X1 U7640 ( .A1(n4473), .A2(n4472), .ZN(n6205) );
  INV_X1 U7641 ( .A(n18442), .ZN(n3045) );
  NAND2_X1 U7642 ( .A1(n20139), .A2(n18467), .ZN(n18442) );
  NAND2_X1 U7645 ( .A1(n8925), .A2(n8748), .ZN(n3433) );
  AOI22_X2 U7646 ( .A1(n7405), .A2(n7948), .B1(n20367), .B2(n7404), .ZN(n8748)
         );
  OR2_X2 U7647 ( .A1(n14407), .A2(n3047), .ZN(n15628) );
  NAND2_X1 U7648 ( .A1(n937), .A2(n11278), .ZN(n9546) );
  NAND2_X1 U7649 ( .A1(n10729), .A2(n19913), .ZN(n3052) );
  NOR2_X1 U7650 ( .A1(n8193), .A2(n3054), .ZN(n3053) );
  INV_X1 U7651 ( .A(n8193), .ZN(n3055) );
  INV_X1 U7652 ( .A(n14714), .ZN(n3057) );
  NAND2_X1 U7653 ( .A1(n3057), .A2(n19843), .ZN(n3056) );
  OAI21_X1 U7654 ( .B1(n3058), .B2(n9238), .A(n9233), .ZN(n3060) );
  XNOR2_X1 U7655 ( .A(n10319), .B(n10029), .ZN(n10035) );
  NAND2_X1 U7656 ( .A1(n20464), .A2(n5046), .ZN(n3061) );
  XNOR2_X1 U7658 ( .A(n13762), .B(n13616), .ZN(n13303) );
  MUX2_X1 U7659 ( .A(n14395), .B(n14598), .S(n14396), .Z(n14398) );
  NAND3_X1 U7661 ( .A1(n18229), .A2(n18232), .A3(n3066), .ZN(n3064) );
  NAND3_X1 U7662 ( .A1(n19876), .A2(n18233), .A3(n3066), .ZN(n3065) );
  NAND3_X1 U7663 ( .A1(n1025), .A2(n3069), .A3(n3070), .ZN(n3068) );
  NAND2_X1 U7664 ( .A1(n5756), .A2(n287), .ZN(n3069) );
  NAND2_X1 U7665 ( .A1(n5757), .A2(n3071), .ZN(n3070) );
  NAND2_X1 U7667 ( .A1(n8000), .A2(n3074), .ZN(n3073) );
  NAND3_X1 U7669 ( .A1(n14439), .A2(n14442), .A3(n14441), .ZN(n12928) );
  NAND2_X1 U7670 ( .A1(n139), .A2(n14442), .ZN(n3173) );
  INV_X1 U7671 ( .A(n4953), .ZN(n3078) );
  INV_X1 U7672 ( .A(n4952), .ZN(n4475) );
  OAI21_X1 U7673 ( .B1(n4399), .B2(n3079), .A(n4916), .ZN(n4400) );
  INV_X1 U7674 ( .A(n18467), .ZN(n18461) );
  NAND2_X1 U7675 ( .A1(n18465), .A2(n18467), .ZN(n3512) );
  INV_X1 U7676 ( .A(n16469), .ZN(n3081) );
  MUX2_X1 U7677 ( .A(n14338), .B(n14335), .S(n12879), .Z(n12880) );
  MUX2_X1 U7679 ( .A(n7948), .B(n7949), .S(n7479), .Z(n7955) );
  NAND3_X1 U7680 ( .A1(n3583), .A2(n7950), .A3(n20367), .ZN(n3581) );
  INV_X1 U7681 ( .A(n16166), .ZN(n17505) );
  NAND3_X1 U7682 ( .A1(n5714), .A2(n3086), .A3(n5715), .ZN(n5724) );
  NAND2_X1 U7683 ( .A1(n14168), .A2(n14167), .ZN(n3088) );
  NAND2_X1 U7685 ( .A1(n7936), .A2(n7763), .ZN(n7519) );
  XNOR2_X1 U7687 ( .A(n3092), .B(n20126), .ZN(n3091) );
  INV_X1 U7688 ( .A(n16900), .ZN(n3092) );
  XNOR2_X1 U7689 ( .A(n16284), .B(n16285), .ZN(n3093) );
  OAI22_X1 U7691 ( .A1(n3095), .A2(n4361), .B1(n4608), .B2(n4601), .ZN(n3094)
         );
  NAND2_X1 U7692 ( .A1(n3097), .A2(n3096), .ZN(n6300) );
  INV_X1 U7693 ( .A(n6089), .ZN(n5199) );
  AOI21_X1 U7694 ( .B1(n6087), .B2(n20149), .A(n6089), .ZN(n3098) );
  INV_X1 U7696 ( .A(n12374), .ZN(n12376) );
  OAI21_X1 U7697 ( .B1(n11856), .B2(n12020), .A(n3099), .ZN(n11857) );
  NAND2_X1 U7698 ( .A1(n3100), .A2(n12369), .ZN(n3099) );
  NOR2_X1 U7699 ( .A1(n19504), .A2(n12374), .ZN(n3100) );
  INV_X1 U7700 ( .A(n10640), .ZN(n11534) );
  NAND3_X1 U7701 ( .A1(n11535), .A2(n11168), .A3(n11171), .ZN(n3104) );
  INV_X1 U7702 ( .A(n10638), .ZN(n11535) );
  NAND3_X1 U7703 ( .A1(n10640), .A2(n11538), .A3(n11539), .ZN(n3105) );
  NOR2_X1 U7704 ( .A1(n11535), .A2(n10640), .ZN(n11169) );
  NAND3_X1 U7705 ( .A1(n20146), .A2(n9129), .A3(n9201), .ZN(n3106) );
  NAND2_X1 U7706 ( .A1(n8276), .A2(n9782), .ZN(n3107) );
  OAI211_X2 U7707 ( .C1(n8244), .C2(n3775), .A(n8243), .B(n8242), .ZN(n9201)
         );
  NOR2_X2 U7709 ( .A1(n3113), .A2(n3111), .ZN(n12001) );
  MUX2_X1 U7710 ( .A(n9486), .B(n11176), .S(n11174), .Z(n3112) );
  MUX2_X1 U7711 ( .A(n9379), .B(n9378), .S(n2232), .Z(n3113) );
  XNOR2_X2 U7712 ( .A(n9225), .B(n9224), .ZN(n11176) );
  INV_X1 U7713 ( .A(n17172), .ZN(n17826) );
  NAND2_X1 U7714 ( .A1(n17824), .A2(n17823), .ZN(n3114) );
  INV_X1 U7715 ( .A(n17080), .ZN(n17822) );
  NAND2_X1 U7716 ( .A1(n17826), .A2(n17825), .ZN(n3117) );
  AOI22_X1 U7718 ( .A1(n8343), .A2(n2964), .B1(n8166), .B2(n8344), .ZN(n3118)
         );
  NAND2_X1 U7719 ( .A1(n3121), .A2(n20274), .ZN(n3119) );
  XNOR2_X1 U7721 ( .A(n6946), .B(n6945), .ZN(n6948) );
  NAND3_X2 U7722 ( .A1(n3124), .A2(n5281), .A3(n3123), .ZN(n6945) );
  NAND2_X1 U7723 ( .A1(n3125), .A2(n3128), .ZN(n3123) );
  NAND2_X1 U7724 ( .A1(n3125), .A2(n3126), .ZN(n3124) );
  OR2_X1 U7725 ( .A1(n5280), .A2(n3127), .ZN(n3126) );
  NAND2_X1 U7726 ( .A1(n5282), .A2(n3127), .ZN(n3125) );
  INV_X1 U7727 ( .A(n5424), .ZN(n3127) );
  NAND2_X1 U7728 ( .A1(n3130), .A2(n4754), .ZN(n3129) );
  NOR2_X1 U7729 ( .A1(n4565), .A2(n3131), .ZN(n3130) );
  INV_X1 U7730 ( .A(n4567), .ZN(n3131) );
  NAND2_X1 U7731 ( .A1(n5518), .A2(n5929), .ZN(n3371) );
  NAND2_X1 U7732 ( .A1(n5053), .A2(n20461), .ZN(n3132) );
  NAND2_X1 U7733 ( .A1(n204), .A2(n11076), .ZN(n3133) );
  NAND2_X1 U7734 ( .A1(n11476), .A2(n3471), .ZN(n3134) );
  NAND3_X1 U7735 ( .A1(n3138), .A2(n15702), .A3(n15696), .ZN(n3137) );
  NOR2_X1 U7736 ( .A1(n3141), .A2(n3140), .ZN(n3139) );
  NOR2_X1 U7737 ( .A1(n16779), .A2(n19144), .ZN(n3140) );
  NAND2_X1 U7739 ( .A1(n19147), .A2(n19145), .ZN(n3143) );
  NAND2_X1 U7742 ( .A1(n3148), .A2(n14905), .ZN(n3146) );
  NAND3_X1 U7743 ( .A1(n14903), .A2(n15056), .A3(n15413), .ZN(n3147) );
  INV_X1 U7744 ( .A(n14312), .ZN(n15549) );
  NOR2_X1 U7745 ( .A1(n15413), .A2(n15553), .ZN(n3148) );
  INV_X1 U7746 ( .A(n14236), .ZN(n14114) );
  NAND2_X1 U7747 ( .A1(n5659), .A2(n6113), .ZN(n5660) );
  NAND2_X1 U7748 ( .A1(n3150), .A2(n17835), .ZN(n17844) );
  NAND2_X1 U7749 ( .A1(n3150), .A2(n3755), .ZN(n3285) );
  NAND2_X1 U7750 ( .A1(n3558), .A2(n11572), .ZN(n3151) );
  NOR2_X1 U7751 ( .A1(n12299), .A2(n12273), .ZN(n12033) );
  OAI21_X1 U7752 ( .B1(n14747), .B2(n1936), .A(n3158), .ZN(n13934) );
  OAI211_X1 U7753 ( .C1(n14427), .C2(n1936), .A(n14747), .B(n3158), .ZN(n14428) );
  INV_X1 U7754 ( .A(n14747), .ZN(n3156) );
  NAND2_X1 U7755 ( .A1(n14752), .A2(n3157), .ZN(n15189) );
  OR2_X1 U7756 ( .A1(n14753), .A2(n3158), .ZN(n3157) );
  XNOR2_X1 U7757 ( .A(n3159), .B(n875), .ZN(n13474) );
  XNOR2_X1 U7758 ( .A(n3159), .B(n18691), .ZN(n13360) );
  XNOR2_X1 U7759 ( .A(n3159), .B(n538), .ZN(n13824) );
  XNOR2_X1 U7760 ( .A(n3159), .B(n19467), .ZN(n12540) );
  XNOR2_X1 U7761 ( .A(n13368), .B(n3159), .ZN(n13530) );
  NAND2_X1 U7762 ( .A1(n11117), .A2(n11435), .ZN(n3161) );
  XNOR2_X1 U7763 ( .A(n3162), .B(n16019), .ZN(n16020) );
  XNOR2_X1 U7764 ( .A(n17406), .B(n3162), .ZN(n16908) );
  XNOR2_X1 U7765 ( .A(n16770), .B(n3162), .ZN(n16829) );
  OAI211_X2 U7766 ( .C1(n15085), .C2(n15086), .A(n15084), .B(n15083), .ZN(
        n3162) );
  NAND2_X1 U7767 ( .A1(n12295), .A2(n3164), .ZN(n12163) );
  MUX2_X1 U7768 ( .A(n12534), .B(n12531), .S(n924), .Z(n11772) );
  INV_X1 U7769 ( .A(n3166), .ZN(n3165) );
  NAND2_X1 U7770 ( .A1(n5105), .A2(n5099), .ZN(n4792) );
  NAND2_X1 U7771 ( .A1(n5102), .A2(n5107), .ZN(n3598) );
  NAND2_X1 U7772 ( .A1(n12813), .A2(n11803), .ZN(n3171) );
  OAI211_X1 U7773 ( .C1(n12813), .C2(n19626), .A(n3169), .B(n3168), .ZN(n12119) );
  XNOR2_X1 U7775 ( .A(n3171), .B(n2151), .ZN(n13699) );
  XNOR2_X1 U7776 ( .A(n3171), .B(n18716), .ZN(n11817) );
  XNOR2_X1 U7777 ( .A(n13588), .B(n3171), .ZN(n12894) );
  OAI211_X2 U7778 ( .C1(n3177), .C2(n11005), .A(n3176), .B(n3175), .ZN(n11952)
         );
  MUX2_X1 U7779 ( .A(n937), .B(n19736), .S(n9547), .Z(n3177) );
  NAND2_X1 U7780 ( .A1(n14053), .A2(n14422), .ZN(n3178) );
  NAND2_X1 U7781 ( .A1(n2039), .A2(n14359), .ZN(n14358) );
  INV_X1 U7782 ( .A(n6345), .ZN(n3181) );
  INV_X1 U7783 ( .A(n6345), .ZN(n7743) );
  AOI22_X1 U7784 ( .A1(n3182), .A2(n7741), .B1(n6900), .B2(n8355), .ZN(n6901)
         );
  XNOR2_X1 U7785 ( .A(n10280), .B(n17095), .ZN(n3184) );
  NOR2_X1 U7786 ( .A1(n8697), .A2(n9161), .ZN(n3183) );
  NAND2_X1 U7787 ( .A1(n8698), .A2(n8697), .ZN(n3185) );
  NOR2_X1 U7788 ( .A1(n12103), .A2(n12101), .ZN(n3186) );
  NAND2_X1 U7789 ( .A1(n3449), .A2(n3189), .ZN(n3188) );
  OAI21_X1 U7791 ( .B1(n6148), .B2(n6138), .A(n3187), .ZN(n5266) );
  NAND2_X1 U7792 ( .A1(n6138), .A2(n5859), .ZN(n3187) );
  NAND2_X1 U7793 ( .A1(n5616), .A2(n3188), .ZN(n5617) );
  NAND2_X1 U7795 ( .A1(n14176), .A2(n12725), .ZN(n3190) );
  XNOR2_X2 U7797 ( .A(Key[101]), .B(Plaintext[101]), .ZN(n5080) );
  NAND2_X1 U7798 ( .A1(n4459), .A2(n5078), .ZN(n3450) );
  NAND3_X1 U7800 ( .A1(n4671), .A2(n4669), .A3(n4670), .ZN(n3192) );
  NAND2_X1 U7801 ( .A1(n4824), .A2(n4827), .ZN(n4670) );
  XNOR2_X2 U7802 ( .A(Key[73]), .B(Plaintext[73]), .ZN(n4827) );
  NAND2_X1 U7803 ( .A1(n3197), .A2(n3195), .ZN(n3194) );
  NAND2_X1 U7804 ( .A1(n3196), .A2(n6184), .ZN(n3195) );
  OAI21_X1 U7805 ( .B1(n6380), .B2(n19476), .A(n2865), .ZN(n3197) );
  NAND2_X1 U7806 ( .A1(n3198), .A2(n20270), .ZN(n8020) );
  NAND2_X1 U7807 ( .A1(n208), .A2(n3198), .ZN(n7812) );
  INV_X1 U7808 ( .A(n7801), .ZN(n3198) );
  NAND2_X1 U7809 ( .A1(n8927), .A2(n8928), .ZN(n3199) );
  NAND2_X1 U7810 ( .A1(n8926), .A2(n8925), .ZN(n3200) );
  NAND2_X1 U7811 ( .A1(n5035), .A2(n3203), .ZN(n5036) );
  NAND2_X1 U7812 ( .A1(n4771), .A2(n3203), .ZN(n4772) );
  NAND2_X1 U7813 ( .A1(n4770), .A2(n3203), .ZN(n4774) );
  XNOR2_X1 U7814 ( .A(n17266), .B(n17265), .ZN(n18038) );
  NAND2_X1 U7815 ( .A1(n3205), .A2(n18038), .ZN(n18237) );
  INV_X1 U7816 ( .A(n17303), .ZN(n17753) );
  OAI211_X1 U7819 ( .C1(n630), .C2(n3198), .A(n3212), .B(n3211), .ZN(n3210) );
  INV_X1 U7820 ( .A(n7466), .ZN(n3212) );
  OAI22_X1 U7821 ( .A1(n16260), .A2(n19947), .B1(n17663), .B2(n3216), .ZN(
        n3215) );
  NOR2_X1 U7824 ( .A1(n8323), .A2(n3809), .ZN(n3220) );
  OAI211_X1 U7827 ( .C1(n19496), .C2(n14828), .A(n3224), .B(n3223), .ZN(n3222)
         );
  NAND2_X1 U7828 ( .A1(n14828), .A2(n14827), .ZN(n3224) );
  NAND2_X1 U7829 ( .A1(n3225), .A2(n14203), .ZN(n14609) );
  INV_X1 U7830 ( .A(n14012), .ZN(n3225) );
  NAND2_X1 U7831 ( .A1(n3226), .A2(n14611), .ZN(n14616) );
  OAI21_X2 U7832 ( .B1(n3228), .B2(n5564), .A(n4993), .ZN(n7371) );
  MUX2_X1 U7833 ( .A(n5532), .B(n6033), .S(n5531), .Z(n3228) );
  NAND2_X1 U7834 ( .A1(n4136), .A2(n4960), .ZN(n3230) );
  AND4_X2 U7837 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n13795)
         );
  OR2_X1 U7838 ( .A1(n12175), .A2(n19768), .ZN(n3238) );
  INV_X1 U7839 ( .A(n8014), .ZN(n7826) );
  AOI21_X1 U7842 ( .B1(n7829), .B2(n7991), .A(n8014), .ZN(n3243) );
  NAND2_X1 U7844 ( .A1(n13008), .A2(n3246), .ZN(n3245) );
  NAND2_X1 U7846 ( .A1(n18762), .A2(n18774), .ZN(n18255) );
  NAND2_X1 U7847 ( .A1(n18250), .A2(n18249), .ZN(n3248) );
  NAND2_X1 U7848 ( .A1(n3249), .A2(n906), .ZN(n3867) );
  NAND2_X1 U7849 ( .A1(n8139), .A2(n8352), .ZN(n3251) );
  INV_X1 U7850 ( .A(n13921), .ZN(n3252) );
  INV_X1 U7853 ( .A(n11792), .ZN(n3256) );
  NAND2_X1 U7854 ( .A1(n3258), .A2(n3257), .ZN(n5846) );
  NAND2_X1 U7855 ( .A1(n4695), .A2(n3259), .ZN(n3257) );
  NAND2_X1 U7856 ( .A1(n4694), .A2(n5107), .ZN(n3258) );
  NOR2_X1 U7857 ( .A1(n12155), .A2(n3260), .ZN(n11908) );
  NAND2_X1 U7858 ( .A1(n12315), .A2(n3260), .ZN(n11712) );
  OAI21_X1 U7860 ( .B1(n8295), .B2(n7789), .A(n7454), .ZN(n3261) );
  NOR2_X1 U7861 ( .A1(n8676), .A2(n8513), .ZN(n8516) );
  XNOR2_X1 U7862 ( .A(n10125), .B(n10356), .ZN(n10130) );
  NAND3_X1 U7863 ( .A1(n3262), .A2(n5697), .A3(n5522), .ZN(n5523) );
  NAND2_X1 U7864 ( .A1(n3264), .A2(n3263), .ZN(n3262) );
  NAND2_X1 U7865 ( .A1(n4950), .A2(n4142), .ZN(n3263) );
  NAND2_X1 U7866 ( .A1(n4143), .A2(n3265), .ZN(n3264) );
  NAND2_X1 U7867 ( .A1(n14165), .A2(n14427), .ZN(n3266) );
  NAND2_X1 U7868 ( .A1(n14166), .A2(n14424), .ZN(n3268) );
  INV_X1 U7869 ( .A(n12607), .ZN(n3269) );
  XNOR2_X1 U7870 ( .A(n12713), .B(n18660), .ZN(n13392) );
  NAND3_X1 U7871 ( .A1(n3271), .A2(n280), .A3(n274), .ZN(n3270) );
  XNOR2_X2 U7872 ( .A(n6282), .B(n6281), .ZN(n7754) );
  XNOR2_X1 U7873 ( .A(n17377), .B(n3273), .ZN(n16918) );
  NAND2_X1 U7874 ( .A1(n14200), .A2(n14590), .ZN(n3275) );
  NAND2_X1 U7875 ( .A1(n11656), .A2(n19768), .ZN(n3277) );
  NAND2_X1 U7876 ( .A1(n14807), .A2(n14813), .ZN(n14196) );
  NAND2_X1 U7877 ( .A1(n12354), .A2(n19768), .ZN(n3537) );
  NAND3_X1 U7878 ( .A1(n3282), .A2(n16734), .A3(n3287), .ZN(n3284) );
  INV_X1 U7879 ( .A(n16730), .ZN(n3282) );
  NAND2_X1 U7881 ( .A1(n3286), .A2(n3284), .ZN(n19151) );
  NAND2_X1 U7882 ( .A1(n16734), .A2(n20423), .ZN(n3286) );
  XNOR2_X1 U7883 ( .A(n19760), .B(n10445), .ZN(n6657) );
  NAND2_X1 U7884 ( .A1(n3290), .A2(n5035), .ZN(n3289) );
  NAND2_X1 U7885 ( .A1(n3431), .A2(n16128), .ZN(n3291) );
  NAND2_X1 U7886 ( .A1(n15611), .A2(n3291), .ZN(n16932) );
  OAI21_X1 U7887 ( .B1(n9275), .B2(n9278), .A(n9272), .ZN(n8759) );
  INV_X1 U7888 ( .A(n19144), .ZN(n18337) );
  AND2_X1 U7891 ( .A1(n12429), .A2(n12686), .ZN(n12094) );
  NAND2_X1 U7892 ( .A1(n10718), .A2(n11474), .ZN(n3296) );
  XNOR2_X1 U7893 ( .A(n9902), .B(n10579), .ZN(n8740) );
  NAND2_X1 U7894 ( .A1(n8731), .A2(n8730), .ZN(n3297) );
  NAND2_X1 U7895 ( .A1(n8732), .A2(n8941), .ZN(n3298) );
  NAND2_X1 U7896 ( .A1(n3301), .A2(n3300), .ZN(n12039) );
  NAND2_X1 U7897 ( .A1(n11169), .A2(n19915), .ZN(n3300) );
  OAI21_X1 U7898 ( .B1(n3303), .B2(n11171), .A(n3302), .ZN(n3301) );
  NAND2_X1 U7899 ( .A1(n3304), .A2(n11171), .ZN(n3302) );
  NOR2_X1 U7900 ( .A1(n11170), .A2(n11168), .ZN(n3303) );
  NAND2_X1 U7901 ( .A1(n11534), .A2(n11170), .ZN(n3304) );
  NAND2_X1 U7902 ( .A1(n3305), .A2(n12237), .ZN(n12073) );
  MUX2_X1 U7904 ( .A(n12604), .B(n12605), .S(n12610), .Z(n12613) );
  XNOR2_X2 U7905 ( .A(n12909), .B(n12908), .ZN(n14442) );
  NAND2_X1 U7906 ( .A1(n14440), .A2(n14441), .ZN(n3306) );
  NAND3_X1 U7907 ( .A1(n15294), .A2(n15295), .A3(n15109), .ZN(n3308) );
  OAI211_X2 U7908 ( .C1(n5029), .C2(n5028), .A(n3310), .B(n3309), .ZN(n5927)
         );
  NAND3_X1 U7909 ( .A1(n5029), .A2(n5026), .A3(n5025), .ZN(n3310) );
  NAND2_X1 U7910 ( .A1(n14962), .A2(n3315), .ZN(n3314) );
  INV_X1 U7911 ( .A(n15581), .ZN(n3315) );
  NAND2_X1 U7912 ( .A1(n5320), .A2(n3319), .ZN(n3318) );
  INV_X1 U7913 ( .A(n5320), .ZN(n6070) );
  NAND2_X1 U7914 ( .A1(n3317), .A2(n5978), .ZN(n3316) );
  NAND2_X1 U7915 ( .A1(n3319), .A2(n6072), .ZN(n3317) );
  AOI21_X1 U7916 ( .B1(n4421), .B2(n20105), .A(n3977), .ZN(n3320) );
  XNOR2_X1 U7917 ( .A(n6506), .B(n6505), .ZN(n3321) );
  NAND2_X1 U7919 ( .A1(n15617), .A2(n15071), .ZN(n14892) );
  INV_X1 U7920 ( .A(n5692), .ZN(n4275) );
  AOI21_X1 U7921 ( .B1(n4254), .B2(n4348), .A(n4349), .ZN(n3322) );
  AOI21_X1 U7922 ( .B1(n4256), .B2(n4255), .A(n4540), .ZN(n3323) );
  AOI21_X1 U7923 ( .B1(n9884), .B2(n11235), .A(n9883), .ZN(n3326) );
  MUX2_X1 U7924 ( .A(n12505), .B(n12508), .S(n12506), .Z(n3565) );
  NAND2_X1 U7925 ( .A1(n9659), .A2(n1330), .ZN(n3324) );
  NOR2_X1 U7926 ( .A1(n12359), .A2(n12509), .ZN(n12505) );
  NOR2_X2 U7927 ( .A1(n3327), .A2(n3326), .ZN(n12509) );
  NAND2_X1 U7928 ( .A1(n9875), .A2(n10818), .ZN(n3328) );
  OAI21_X1 U7929 ( .B1(n14341), .B2(n14339), .A(n3333), .ZN(n3332) );
  NAND2_X1 U7930 ( .A1(n14334), .A2(n19485), .ZN(n3333) );
  NOR2_X1 U7932 ( .A1(n3335), .A2(n7762), .ZN(n3334) );
  NOR2_X1 U7933 ( .A1(n7934), .A2(n7760), .ZN(n3335) );
  MUX2_X1 U7935 ( .A(n7765), .B(n3337), .S(n7932), .Z(n3336) );
  NAND2_X1 U7936 ( .A1(n7934), .A2(n2540), .ZN(n3337) );
  INV_X1 U7937 ( .A(n7763), .ZN(n7934) );
  NAND3_X1 U7938 ( .A1(n3339), .A2(n19240), .A3(n3338), .ZN(n19245) );
  NAND2_X1 U7939 ( .A1(n3340), .A2(n19236), .ZN(n3339) );
  NAND2_X1 U7940 ( .A1(n3341), .A2(n19234), .ZN(n3340) );
  OR2_X1 U7941 ( .A1(n19237), .A2(n19235), .ZN(n3341) );
  NAND2_X1 U7942 ( .A1(n19227), .A2(n19237), .ZN(n19234) );
  OAI22_X2 U7943 ( .A1(n5694), .A2(n5695), .B1(n5693), .B2(n4275), .ZN(n7097)
         );
  NAND3_X1 U7947 ( .A1(n16801), .A2(n17489), .A3(n19675), .ZN(n3346) );
  OAI21_X1 U7949 ( .B1(n1458), .B2(n15052), .A(n15350), .ZN(n3348) );
  OR2_X1 U7951 ( .A1(n4538), .A2(n4539), .ZN(n3349) );
  NAND2_X1 U7952 ( .A1(n3933), .A2(n3932), .ZN(n3350) );
  XNOR2_X1 U7954 ( .A(n13440), .B(n3352), .ZN(n11852) );
  INV_X1 U7955 ( .A(n12993), .ZN(n3352) );
  XNOR2_X1 U7956 ( .A(n3353), .B(n12993), .ZN(n12858) );
  INV_X1 U7957 ( .A(n13078), .ZN(n3353) );
  OAI21_X1 U7958 ( .B1(n3356), .B2(n9255), .A(n9252), .ZN(n3355) );
  NAND2_X1 U7960 ( .A1(n11176), .A2(n10912), .ZN(n3358) );
  INV_X1 U7963 ( .A(n11177), .ZN(n3362) );
  XNOR2_X1 U7964 ( .A(n13569), .B(n13134), .ZN(n3363) );
  AND2_X1 U7965 ( .A1(n18489), .A2(n18498), .ZN(n17911) );
  NAND2_X1 U7966 ( .A1(n16166), .A2(n17501), .ZN(n16797) );
  NAND2_X1 U7967 ( .A1(n13166), .A2(n3366), .ZN(n13179) );
  NAND2_X1 U7968 ( .A1(n14665), .A2(n14664), .ZN(n3367) );
  NAND2_X1 U7969 ( .A1(n3369), .A2(n3445), .ZN(n3368) );
  OAI21_X1 U7970 ( .B1(n7748), .B2(n7750), .A(n3370), .ZN(n3369) );
  NAND2_X1 U7971 ( .A1(n7749), .A2(n7748), .ZN(n3370) );
  NAND2_X1 U7972 ( .A1(n3948), .A2(n4539), .ZN(n4200) );
  OAI21_X1 U7973 ( .B1(n4350), .B2(n4199), .A(n3948), .ZN(n3949) );
  MUX2_X1 U7974 ( .A(n4541), .B(n3948), .S(n4350), .Z(n4203) );
  NAND3_X1 U7975 ( .A1(n4536), .A2(n3948), .A3(n4350), .ZN(n4351) );
  INV_X1 U7976 ( .A(n3373), .ZN(n14262) );
  NOR2_X1 U7977 ( .A1(n13981), .A2(n3373), .ZN(n14539) );
  NOR2_X1 U7980 ( .A1(n7979), .A2(n7921), .ZN(n3375) );
  NAND2_X1 U7981 ( .A1(n7984), .A2(n7981), .ZN(n7979) );
  INV_X1 U7983 ( .A(n7921), .ZN(n7768) );
  NAND2_X1 U7984 ( .A1(n7768), .A2(n7978), .ZN(n3376) );
  AND2_X2 U7987 ( .A1(n3380), .A2(n3378), .ZN(n10350) );
  NAND2_X1 U7988 ( .A1(n9050), .A2(n3379), .ZN(n3378) );
  NAND3_X1 U7989 ( .A1(n3395), .A2(n9579), .A3(n3394), .ZN(n3379) );
  NAND2_X1 U7990 ( .A1(n9052), .A2(n9051), .ZN(n3380) );
  OAI22_X1 U7991 ( .A1(n19519), .A2(n9579), .B1(n8577), .B2(n19715), .ZN(n9052) );
  NAND2_X1 U7992 ( .A1(n11013), .A2(n3382), .ZN(n3381) );
  OAI22_X1 U7993 ( .A1(n4187), .A2(n4520), .B1(n4343), .B2(n4524), .ZN(n3943)
         );
  XNOR2_X2 U7994 ( .A(Key[173]), .B(Plaintext[173]), .ZN(n4524) );
  NAND2_X1 U7996 ( .A1(n3387), .A2(n7974), .ZN(n3383) );
  MUX2_X1 U7997 ( .A(n278), .B(n7922), .S(n7967), .Z(n3387) );
  NAND2_X1 U7998 ( .A1(n17222), .A2(n3389), .ZN(n3388) );
  NAND2_X1 U7999 ( .A1(n17219), .A2(n1897), .ZN(n3390) );
  INV_X1 U8000 ( .A(n15767), .ZN(n15656) );
  OR2_X2 U8001 ( .A1(n14856), .A2(n11594), .ZN(n15767) );
  NOR2_X1 U8003 ( .A1(n15657), .A2(n15767), .ZN(n3393) );
  AND2_X1 U8005 ( .A1(n13905), .A2(n14782), .ZN(n11320) );
  AND2_X1 U8006 ( .A1(n3397), .A2(n5279), .ZN(n5672) );
  INV_X1 U8007 ( .A(n5668), .ZN(n3397) );
  NAND3_X1 U8008 ( .A1(n3398), .A2(n5670), .A3(n5668), .ZN(n5281) );
  MUX2_X1 U8009 ( .A(n3398), .B(n5669), .S(n5670), .Z(n5426) );
  OAI21_X1 U8010 ( .B1(n5673), .B2(n3398), .A(n5670), .ZN(n5187) );
  NAND2_X1 U8011 ( .A1(n4209), .A2(n4208), .ZN(n3399) );
  NAND2_X1 U8012 ( .A1(n12630), .A2(n3401), .ZN(n3400) );
  INV_X1 U8014 ( .A(n12630), .ZN(n3403) );
  AOI21_X2 U8015 ( .B1(n8294), .B2(n8293), .A(n3406), .ZN(n9106) );
  XNOR2_X1 U8016 ( .A(n16707), .B(n17143), .ZN(n16822) );
  INV_X1 U8018 ( .A(n3408), .ZN(n3407) );
  OAI21_X1 U8019 ( .B1(n6028), .B2(n3410), .A(n3409), .ZN(n3408) );
  NAND2_X1 U8021 ( .A1(n3434), .A2(n19790), .ZN(n6028) );
  NAND2_X1 U8022 ( .A1(n16802), .A2(n17492), .ZN(n16803) );
  NAND2_X1 U8023 ( .A1(n16471), .A2(n17492), .ZN(n16472) );
  NAND2_X1 U8024 ( .A1(n7416), .A2(n3525), .ZN(n3524) );
  NAND2_X1 U8025 ( .A1(n3694), .A2(n14562), .ZN(n3412) );
  OAI21_X2 U8026 ( .B1(n14123), .B2(n14122), .A(n14121), .ZN(n15608) );
  NAND2_X1 U8027 ( .A1(n3427), .A2(n997), .ZN(n3413) );
  MUX2_X1 U8028 ( .A(n3431), .B(n16127), .S(n16128), .Z(n3415) );
  XNOR2_X1 U8029 ( .A(n10558), .B(n10430), .ZN(n10242) );
  NAND2_X1 U8031 ( .A1(n3418), .A2(n9020), .ZN(n3416) );
  NAND3_X1 U8032 ( .A1(n9019), .A2(n9296), .A3(n20159), .ZN(n3417) );
  XNOR2_X1 U8033 ( .A(n13649), .B(n3420), .ZN(n3419) );
  INV_X1 U8034 ( .A(n13650), .ZN(n3420) );
  NAND3_X1 U8035 ( .A1(n17646), .A2(n3422), .A3(n17647), .ZN(n3421) );
  NAND2_X1 U8036 ( .A1(n3423), .A2(n17737), .ZN(n3422) );
  NAND2_X1 U8037 ( .A1(n17645), .A2(n17644), .ZN(n3423) );
  XNOR2_X1 U8038 ( .A(n10125), .B(n3424), .ZN(n10412) );
  NAND2_X1 U8039 ( .A1(n3427), .A2(n3425), .ZN(n3426) );
  OAI21_X1 U8040 ( .B1(n8925), .B2(n8932), .A(n3433), .ZN(n8754) );
  NAND3_X1 U8044 ( .A1(n19735), .A2(n18672), .A3(n18666), .ZN(n3436) );
  NAND3_X1 U8045 ( .A1(n18686), .A2(n19735), .A3(n18671), .ZN(n3437) );
  NAND2_X1 U8047 ( .A1(n13891), .A2(n3440), .ZN(n13892) );
  NAND3_X1 U8048 ( .A1(n20500), .A2(n14800), .A3(n3440), .ZN(n14802) );
  OAI22_X1 U8049 ( .A1(n12321), .A2(n3439), .B1(n14797), .B2(n3440), .ZN(
        n14851) );
  INV_X1 U8050 ( .A(n14801), .ZN(n3439) );
  NAND2_X1 U8051 ( .A1(n11282), .A2(n19779), .ZN(n9413) );
  MUX2_X1 U8052 ( .A(n4746), .B(n4744), .S(n4204), .Z(n4751) );
  NAND2_X1 U8053 ( .A1(n4559), .A2(n4204), .ZN(n4250) );
  MUX2_X1 U8054 ( .A(n11881), .B(n11048), .S(n11880), .Z(n11049) );
  MUX2_X1 U8055 ( .A(n11460), .B(n11461), .S(n11880), .Z(n11462) );
  NAND2_X1 U8056 ( .A1(n14819), .A2(n3444), .ZN(n3443) );
  MUX2_X1 U8057 ( .A(n7749), .B(n7748), .S(n7508), .Z(n3447) );
  XNOR2_X1 U8058 ( .A(n3448), .B(n16067), .ZN(n16068) );
  XNOR2_X1 U8059 ( .A(n16860), .B(n3448), .ZN(n16765) );
  XNOR2_X1 U8060 ( .A(n16214), .B(n3448), .ZN(n15855) );
  OR2_X1 U8061 ( .A1(n15636), .A2(n15846), .ZN(n15848) );
  NAND2_X1 U8062 ( .A1(n3450), .A2(n5077), .ZN(n3449) );
  AOI21_X1 U8064 ( .B1(n20111), .B2(n20361), .A(n18384), .ZN(n3456) );
  INV_X1 U8066 ( .A(n15768), .ZN(n3457) );
  OAI21_X1 U8067 ( .B1(n4520), .B2(n4524), .A(n4519), .ZN(n4521) );
  NAND2_X1 U8070 ( .A1(n3461), .A2(n19374), .ZN(n17598) );
  OAI22_X1 U8071 ( .A1(n19647), .A2(n19372), .B1(n19380), .B2(n19666), .ZN(
        n3461) );
  OAI21_X1 U8072 ( .B1(n3463), .B2(n3462), .A(n11757), .ZN(n3464) );
  INV_X1 U8073 ( .A(n12306), .ZN(n3463) );
  INV_X1 U8074 ( .A(n9771), .ZN(n10298) );
  NAND2_X1 U8075 ( .A1(n8791), .A2(n9149), .ZN(n3465) );
  NAND2_X1 U8076 ( .A1(n8792), .A2(n8338), .ZN(n3466) );
  NAND2_X1 U8077 ( .A1(n3470), .A2(n5993), .ZN(n3469) );
  NAND2_X1 U8078 ( .A1(n5088), .A2(n5083), .ZN(n4090) );
  NAND3_X1 U8079 ( .A1(n4802), .A2(n5088), .A3(n19777), .ZN(n4700) );
  NAND3_X1 U8080 ( .A1(n4807), .A2(n5088), .A3(n4804), .ZN(n4805) );
  INV_X1 U8081 ( .A(n8192), .ZN(n8051) );
  NAND2_X1 U8083 ( .A1(n8053), .A2(n8192), .ZN(n3472) );
  XNOR2_X1 U8084 ( .A(n6116), .B(n6115), .ZN(n7457) );
  AND2_X1 U8085 ( .A1(n15333), .A2(n3473), .ZN(n15706) );
  NAND2_X1 U8086 ( .A1(n2475), .A2(n3475), .ZN(n18127) );
  NAND2_X1 U8087 ( .A1(n17945), .A2(n3475), .ZN(n17952) );
  AND2_X1 U8088 ( .A1(n12532), .A2(n12534), .ZN(n3477) );
  NAND2_X1 U8089 ( .A1(n11477), .A2(n3481), .ZN(n3478) );
  NAND2_X1 U8090 ( .A1(n11478), .A2(n3482), .ZN(n3479) );
  NAND2_X1 U8091 ( .A1(n3483), .A2(n6120), .ZN(n5390) );
  NAND3_X1 U8092 ( .A1(n6128), .A2(n5868), .A3(n3483), .ZN(n4433) );
  AND2_X1 U8093 ( .A1(n3484), .A2(n20252), .ZN(n8146) );
  NAND2_X1 U8094 ( .A1(n3484), .A2(n7671), .ZN(n8371) );
  NOR2_X1 U8095 ( .A1(n3484), .A2(n20252), .ZN(n6750) );
  NAND2_X1 U8097 ( .A1(n7677), .A2(n3491), .ZN(n8722) );
  NAND2_X1 U8099 ( .A1(n9359), .A2(n3493), .ZN(n3492) );
  MUX2_X1 U8100 ( .A(n9358), .B(n8904), .S(n9359), .Z(n3494) );
  NAND2_X1 U8101 ( .A1(n9352), .A2(n9358), .ZN(n3495) );
  INV_X1 U8102 ( .A(n6786), .ZN(n6511) );
  XNOR2_X2 U8103 ( .A(Key[68]), .B(Plaintext[68]), .ZN(n3978) );
  INV_X1 U8104 ( .A(n13617), .ZN(n3498) );
  OR2_X1 U8105 ( .A1(n11315), .A2(n12409), .ZN(n3499) );
  INV_X1 U8106 ( .A(n10746), .ZN(n3500) );
  XNOR2_X1 U8107 ( .A(n856), .B(n10296), .ZN(n10406) );
  NAND2_X1 U8109 ( .A1(n9211), .A2(n9135), .ZN(n3503) );
  NAND3_X1 U8112 ( .A1(n8923), .A2(n3506), .A3(n3505), .ZN(n3504) );
  NAND2_X1 U8113 ( .A1(n8733), .A2(n8734), .ZN(n3505) );
  NAND2_X1 U8114 ( .A1(n8916), .A2(n8497), .ZN(n3506) );
  AND2_X1 U8116 ( .A1(n204), .A2(n3711), .ZN(n9913) );
  NAND2_X1 U8117 ( .A1(n11476), .A2(n3507), .ZN(n9920) );
  NAND2_X1 U8118 ( .A1(n204), .A2(n3507), .ZN(n10717) );
  NOR2_X1 U8119 ( .A1(n204), .A2(n3507), .ZN(n10894) );
  OAI21_X1 U8120 ( .B1(n3711), .B2(n11474), .A(n3508), .ZN(n11478) );
  NAND2_X1 U8121 ( .A1(n11474), .A2(n11475), .ZN(n3508) );
  NAND2_X1 U8122 ( .A1(n3509), .A2(n18436), .ZN(n16486) );
  NAND2_X1 U8123 ( .A1(n3512), .A2(n3510), .ZN(n3509) );
  NAND2_X1 U8124 ( .A1(n18453), .A2(n20231), .ZN(n3510) );
  NAND3_X1 U8125 ( .A1(n14574), .A2(n14267), .A3(n14570), .ZN(n14272) );
  OAI21_X1 U8126 ( .B1(n12430), .B2(n12686), .A(n3514), .ZN(n11613) );
  MUX2_X1 U8127 ( .A(n11142), .B(n11144), .S(n9616), .Z(n10958) );
  MUX2_X1 U8128 ( .A(n3515), .B(n20366), .S(n10960), .Z(n3671) );
  INV_X1 U8129 ( .A(n12911), .ZN(n13865) );
  OAI21_X1 U8130 ( .B1(n4976), .B2(n4975), .A(n4977), .ZN(n3517) );
  NAND3_X1 U8131 ( .A1(n7751), .A2(n3520), .A3(n7752), .ZN(n8658) );
  INV_X1 U8132 ( .A(n7752), .ZN(n8999) );
  NAND2_X1 U8134 ( .A1(n11070), .A2(n3521), .ZN(n3638) );
  INV_X1 U8135 ( .A(n14465), .ZN(n3522) );
  NOR2_X1 U8136 ( .A1(n19531), .A2(n3522), .ZN(n14364) );
  NAND2_X1 U8137 ( .A1(n19657), .A2(n3522), .ZN(n12726) );
  OAI22_X1 U8138 ( .A1(n13924), .A2(n3522), .B1(n14363), .B2(n19538), .ZN(
        n13925) );
  OAI211_X2 U8139 ( .C1(n3526), .C2(n3525), .A(n3524), .B(n3523), .ZN(n9837)
         );
  INV_X1 U8140 ( .A(n8069), .ZN(n3525) );
  NAND3_X1 U8142 ( .A1(n5683), .A2(n5682), .A3(n3529), .ZN(n3527) );
  NAND2_X1 U8143 ( .A1(n5687), .A2(n5686), .ZN(n3528) );
  NAND2_X1 U8145 ( .A1(n11944), .A2(n11945), .ZN(n3531) );
  NAND2_X1 U8147 ( .A1(n3535), .A2(n17538), .ZN(n18311) );
  INV_X1 U8148 ( .A(n12001), .ZN(n11030) );
  NAND3_X1 U8149 ( .A1(n14078), .A2(n14217), .A3(n877), .ZN(n3539) );
  NAND2_X1 U8150 ( .A1(n8235), .A2(n8083), .ZN(n3540) );
  NAND2_X1 U8151 ( .A1(n8234), .A2(n19826), .ZN(n3541) );
  INV_X1 U8152 ( .A(n9204), .ZN(n3542) );
  NAND2_X1 U8153 ( .A1(n4233), .A2(n4907), .ZN(n4378) );
  OR2_X1 U8154 ( .A1(n18950), .A2(n18946), .ZN(n3548) );
  INV_X1 U8155 ( .A(n18043), .ZN(n18047) );
  NAND2_X1 U8156 ( .A1(n18047), .A2(n3546), .ZN(n3545) );
  NAND2_X1 U8157 ( .A1(n3728), .A2(n20369), .ZN(n3549) );
  XNOR2_X1 U8158 ( .A(n8339), .B(n9994), .ZN(n8396) );
  NOR2_X1 U8159 ( .A1(n8999), .A2(n8997), .ZN(n3557) );
  NAND2_X1 U8162 ( .A1(n8773), .A2(n3557), .ZN(n3556) );
  NAND3_X1 U8163 ( .A1(n4865), .A2(n4652), .A3(n20356), .ZN(n3561) );
  AOI21_X1 U8165 ( .B1(n4867), .B2(n4870), .A(n4865), .ZN(n3564) );
  OAI21_X1 U8166 ( .B1(n4651), .B2(n3560), .A(n3559), .ZN(n4655) );
  NAND2_X1 U8167 ( .A1(n4381), .A2(n20357), .ZN(n3559) );
  INV_X1 U8168 ( .A(n4867), .ZN(n3560) );
  OAI21_X1 U8169 ( .B1(n4651), .B2(n3562), .A(n3561), .ZN(n3563) );
  NAND2_X1 U8171 ( .A1(n12001), .A2(n12353), .ZN(n12350) );
  NAND2_X1 U8173 ( .A1(n164), .A2(n3978), .ZN(n4659) );
  NAND2_X1 U8174 ( .A1(n9660), .A2(n11383), .ZN(n3566) );
  NAND3_X1 U8175 ( .A1(n5447), .A2(n5825), .A3(n5826), .ZN(n3567) );
  OAI21_X2 U8176 ( .B1(n4231), .B2(n4230), .A(n4229), .ZN(n5823) );
  XNOR2_X1 U8179 ( .A(n13864), .B(n13184), .ZN(n3575) );
  XNOR2_X1 U8181 ( .A(n3578), .B(n18012), .ZN(Ciphertext[34]) );
  OAI211_X1 U8182 ( .C1(n18010), .C2(n19526), .A(n3580), .B(n3579), .ZN(n3578)
         );
  NAND2_X1 U8183 ( .A1(n994), .A2(n18518), .ZN(n3580) );
  INV_X1 U8185 ( .A(n7815), .ZN(n3583) );
  NAND2_X1 U8186 ( .A1(n3587), .A2(n19506), .ZN(n3584) );
  NAND2_X1 U8187 ( .A1(n3588), .A2(n11290), .ZN(n11293) );
  XNOR2_X1 U8188 ( .A(n6927), .B(n7143), .ZN(n3590) );
  INV_X1 U8189 ( .A(n4483), .ZN(n3592) );
  NAND2_X1 U8190 ( .A1(n4968), .A2(n4482), .ZN(n3593) );
  NAND2_X1 U8191 ( .A1(n8265), .A2(n8264), .ZN(n3594) );
  NAND3_X1 U8192 ( .A1(n3596), .A2(n8266), .A3(n3597), .ZN(n3595) );
  NAND2_X1 U8193 ( .A1(n7864), .A2(n3766), .ZN(n3596) );
  AOI21_X1 U8194 ( .B1(n3598), .B2(n4449), .A(n4077), .ZN(n4078) );
  INV_X1 U8195 ( .A(n14176), .ZN(n3599) );
  NAND2_X1 U8198 ( .A1(n20496), .A2(n3601), .ZN(n11274) );
  NAND2_X1 U8199 ( .A1(n5813), .A2(n19562), .ZN(n3603) );
  NAND2_X1 U8200 ( .A1(n5716), .A2(n3608), .ZN(n5722) );
  NAND3_X2 U8201 ( .A1(n7478), .A2(n3610), .A3(n3609), .ZN(n8815) );
  NAND2_X1 U8202 ( .A1(n7476), .A2(n20144), .ZN(n3610) );
  NAND2_X1 U8203 ( .A1(n3612), .A2(n11412), .ZN(n3616) );
  NAND2_X1 U8204 ( .A1(n3614), .A2(n3616), .ZN(n12553) );
  NAND2_X1 U8205 ( .A1(n11977), .A2(n12544), .ZN(n11796) );
  INV_X1 U8206 ( .A(n8990), .ZN(n9276) );
  OAI21_X1 U8207 ( .B1(n8649), .B2(n9276), .A(n9278), .ZN(n3618) );
  XNOR2_X1 U8208 ( .A(n10204), .B(n10114), .ZN(n9644) );
  INV_X1 U8209 ( .A(n7286), .ZN(n6095) );
  XNOR2_X1 U8210 ( .A(n7286), .B(n7285), .ZN(n7293) );
  INV_X1 U8211 ( .A(n7026), .ZN(n3619) );
  INV_X1 U8212 ( .A(n3620), .ZN(n7380) );
  XNOR2_X1 U8213 ( .A(n6918), .B(n6917), .ZN(n3620) );
  AOI21_X1 U8214 ( .B1(n15031), .B2(n15379), .A(n3621), .ZN(n15032) );
  MUX2_X1 U8215 ( .A(n19513), .B(n15167), .S(n15028), .Z(n12936) );
  NAND2_X1 U8216 ( .A1(n14873), .A2(n3621), .ZN(n14878) );
  OR2_X1 U8217 ( .A1(n4532), .A2(n4528), .ZN(n3623) );
  NAND2_X1 U8218 ( .A1(n12125), .A2(n12230), .ZN(n3626) );
  AND2_X1 U8219 ( .A1(n5435), .A2(n6000), .ZN(n3627) );
  NAND2_X1 U8220 ( .A1(n5996), .A2(n6000), .ZN(n5705) );
  XNOR2_X1 U8221 ( .A(n7122), .B(n7081), .ZN(n6621) );
  XNOR2_X1 U8222 ( .A(n6621), .B(n6620), .ZN(n6622) );
  NAND2_X1 U8224 ( .A1(n10921), .A2(n10919), .ZN(n10924) );
  NAND2_X1 U8226 ( .A1(n12222), .A2(n12221), .ZN(n10925) );
  XNOR2_X1 U8227 ( .A(n10348), .B(n10085), .ZN(n3628) );
  INV_X1 U8228 ( .A(n10348), .ZN(n10086) );
  NAND2_X1 U8229 ( .A1(n10104), .A2(n19949), .ZN(n3630) );
  NOR2_X1 U8230 ( .A1(n11658), .A2(n11955), .ZN(n3632) );
  XOR2_X1 U8231 ( .A(n13530), .B(n13579), .Z(n12682) );
  NAND4_X2 U8232 ( .A1(n12344), .A2(n12343), .A3(n12341), .A4(n12342), .ZN(
        n13266) );
  OAI21_X2 U8233 ( .B1(n4535), .B2(n4159), .A(n3634), .ZN(n5575) );
  NAND3_X1 U8234 ( .A1(n14357), .A2(n2039), .A3(n14422), .ZN(n3635) );
  AND2_X2 U8235 ( .A1(n12257), .A2(n3637), .ZN(n12250) );
  NAND2_X1 U8236 ( .A1(n11071), .A2(n11493), .ZN(n3639) );
  INV_X1 U8237 ( .A(n5841), .ZN(n3640) );
  NAND2_X1 U8238 ( .A1(n4490), .A2(n210), .ZN(n3641) );
  NAND2_X1 U8239 ( .A1(n14263), .A2(n3642), .ZN(n3643) );
  INV_X1 U8240 ( .A(n14262), .ZN(n3642) );
  NAND2_X1 U8241 ( .A1(n14019), .A2(n14262), .ZN(n3644) );
  NAND2_X1 U8242 ( .A1(n3643), .A2(n3644), .ZN(n15759) );
  NAND2_X1 U8243 ( .A1(n15756), .A2(n15754), .ZN(n15587) );
  NAND2_X1 U8244 ( .A1(n3645), .A2(n8917), .ZN(n7668) );
  NAND2_X1 U8245 ( .A1(n4835), .A2(n3846), .ZN(n4417) );
  OAI21_X1 U8246 ( .B1(n20256), .B2(n4676), .A(n4417), .ZN(n3652) );
  NAND2_X1 U8247 ( .A1(n2042), .A2(n19508), .ZN(n4418) );
  NAND2_X1 U8248 ( .A1(n8080), .A2(n20174), .ZN(n3653) );
  NAND2_X1 U8249 ( .A1(n8077), .A2(n3655), .ZN(n3654) );
  NAND2_X1 U8250 ( .A1(n4960), .A2(n292), .ZN(n3656) );
  NAND2_X1 U8251 ( .A1(n3656), .A2(n20205), .ZN(n4138) );
  OAI211_X1 U8252 ( .C1(n3657), .C2(n4899), .A(n4898), .B(n4892), .ZN(n4900)
         );
  AND2_X1 U8253 ( .A1(n3658), .A2(n4375), .ZN(n3745) );
  NOR2_X2 U8254 ( .A1(n8422), .A2(n8421), .ZN(n9111) );
  NAND2_X1 U8255 ( .A1(n3659), .A2(n3661), .ZN(n8422) );
  NAND2_X1 U8256 ( .A1(n8285), .A2(n8284), .ZN(n3661) );
  INV_X1 U8257 ( .A(n5984), .ZN(n3663) );
  NOR2_X1 U8258 ( .A1(n3665), .A2(n5558), .ZN(n5560) );
  NAND2_X1 U8259 ( .A1(n3665), .A2(n6051), .ZN(n5141) );
  NAND2_X1 U8260 ( .A1(n13164), .A2(n14535), .ZN(n13165) );
  NAND2_X1 U8261 ( .A1(n12311), .A2(n12312), .ZN(n3666) );
  OAI21_X1 U8263 ( .B1(n11340), .B2(n9830), .A(n3669), .ZN(n9831) );
  INV_X1 U8264 ( .A(n10673), .ZN(n3669) );
  INV_X1 U8266 ( .A(n13618), .ZN(n3675) );
  XNOR2_X1 U8267 ( .A(n13085), .B(n3675), .ZN(n13415) );
  NAND3_X1 U8268 ( .A1(n10990), .A2(n11869), .A3(n11302), .ZN(n10715) );
  NAND2_X1 U8269 ( .A1(n3681), .A2(n3678), .ZN(n3677) );
  NAND2_X1 U8270 ( .A1(n3679), .A2(n208), .ZN(n3678) );
  NAND2_X1 U8271 ( .A1(n20490), .A2(n20270), .ZN(n3680) );
  OAI21_X1 U8274 ( .B1(n3689), .B2(n3690), .A(n15769), .ZN(n3687) );
  AND2_X2 U8275 ( .A1(n3687), .A2(n3686), .ZN(n16742) );
  AOI21_X1 U8276 ( .B1(n15766), .B2(n15767), .A(n229), .ZN(n3688) );
  OAI22_X1 U8277 ( .A1(n14273), .A2(n14566), .B1(n14275), .B2(n14563), .ZN(
        n3694) );
  AND2_X2 U8278 ( .A1(n3698), .A2(n3695), .ZN(n15866) );
  NAND2_X1 U8279 ( .A1(n3699), .A2(n20518), .ZN(n3698) );
  NAND2_X1 U8280 ( .A1(n13903), .A2(n13902), .ZN(n3699) );
  NAND2_X1 U8283 ( .A1(n14703), .A2(n3705), .ZN(n3704) );
  OAI21_X1 U8284 ( .B1(n6090), .B2(n6089), .A(n890), .ZN(n6093) );
  NAND2_X1 U8285 ( .A1(n5905), .A2(n4862), .ZN(n6089) );
  NAND2_X1 U8286 ( .A1(n4859), .A2(n3706), .ZN(n5905) );
  NAND2_X1 U8287 ( .A1(n11707), .A2(n12480), .ZN(n3707) );
  XNOR2_X1 U8288 ( .A(n12849), .B(n13048), .ZN(n12998) );
  NAND2_X1 U8289 ( .A1(n15081), .A2(n15531), .ZN(n15916) );
  NAND2_X1 U8290 ( .A1(n15919), .A2(n15081), .ZN(n3709) );
  NAND2_X1 U8292 ( .A1(n11219), .A2(n204), .ZN(n3713) );
  NAND2_X1 U8293 ( .A1(n4612), .A2(n3716), .ZN(n3715) );
  NAND2_X1 U8294 ( .A1(n20509), .A2(n5742), .ZN(n5202) );
  NAND2_X1 U8295 ( .A1(n5271), .A2(n19865), .ZN(n3719) );
  NAND2_X1 U8296 ( .A1(n11620), .A2(n1371), .ZN(n3721) );
  INV_X1 U8297 ( .A(n5743), .ZN(n5746) );
  NAND2_X1 U8298 ( .A1(n15642), .A2(n15256), .ZN(n15835) );
  NAND2_X1 U8299 ( .A1(n15642), .A2(n3722), .ZN(n3723) );
  NAND2_X1 U8300 ( .A1(n3724), .A2(n3723), .ZN(n15099) );
  NAND2_X1 U8301 ( .A1(n15095), .A2(n3725), .ZN(n3724) );
  INV_X1 U8302 ( .A(n19931), .ZN(n3725) );
  OR2_X1 U8303 ( .A1(n14664), .A2(n14662), .ZN(n14536) );
  INV_X1 U8304 ( .A(n14662), .ZN(n3726) );
  NOR2_X1 U8305 ( .A1(n3726), .A2(n13164), .ZN(n14668) );
  AND3_X1 U8306 ( .A1(n3727), .A2(n14662), .A3(n14664), .ZN(n13178) );
  NAND2_X1 U8307 ( .A1(n14666), .A2(n14667), .ZN(n3727) );
  NAND2_X1 U8308 ( .A1(n20369), .A2(n4633), .ZN(n4637) );
  INV_X1 U8309 ( .A(n18842), .ZN(n18813) );
  NAND2_X1 U8310 ( .A1(n18275), .A2(n221), .ZN(n3729) );
  OR2_X1 U8311 ( .A1(n18275), .A2(n17769), .ZN(n3730) );
  NAND2_X1 U8312 ( .A1(n11888), .A2(n3732), .ZN(n3731) );
  INV_X1 U8313 ( .A(n12264), .ZN(n3733) );
  OAI21_X1 U8314 ( .B1(n12261), .B2(n3734), .A(n12016), .ZN(n11894) );
  NOR2_X1 U8315 ( .A1(n11727), .A2(n3734), .ZN(n11728) );
  XNOR2_X1 U8316 ( .A(n14914), .B(n3735), .ZN(n14915) );
  NAND2_X1 U8317 ( .A1(n3739), .A2(n3737), .ZN(n3736) );
  NAND2_X1 U8318 ( .A1(n3738), .A2(n14900), .ZN(n3737) );
  NOR2_X1 U8319 ( .A1(n3741), .A2(n14901), .ZN(n3738) );
  OAI21_X1 U8320 ( .B1(n3740), .B2(n3741), .A(n14901), .ZN(n3739) );
  INV_X1 U8321 ( .A(n14900), .ZN(n3740) );
  OAI21_X1 U8322 ( .B1(n15916), .B2(n15420), .A(n14899), .ZN(n3741) );
  INV_X1 U8323 ( .A(n14120), .ZN(n14230) );
  XNOR2_X1 U8324 ( .A(n13705), .B(n2257), .ZN(n3744) );
  NAND2_X1 U8325 ( .A1(n5484), .A2(n3746), .ZN(n7163) );
  NAND2_X1 U8327 ( .A1(n3748), .A2(n8301), .ZN(n7876) );
  NAND2_X1 U8328 ( .A1(n3747), .A2(n20057), .ZN(n5299) );
  AND2_X1 U8329 ( .A1(n19865), .A2(n8044), .ZN(n3747) );
  NAND3_X1 U8330 ( .A1(n8308), .A2(n8306), .A3(n8307), .ZN(n3750) );
  NAND2_X1 U8332 ( .A1(n4338), .A2(n3753), .ZN(n3752) );
  NAND2_X1 U8333 ( .A1(n11628), .A2(n11627), .ZN(n11969) );
  INV_X1 U8334 ( .A(n17836), .ZN(n3755) );
  INV_X1 U8335 ( .A(n16731), .ZN(n17838) );
  OAI21_X1 U8336 ( .B1(n16731), .B2(n3755), .A(n17840), .ZN(n16733) );
  NAND2_X1 U8338 ( .A1(n3951), .A2(n3759), .ZN(n5148) );
  NAND2_X1 U8340 ( .A1(n8264), .A2(n7864), .ZN(n3765) );
  NAND2_X1 U8341 ( .A1(n7569), .A2(n3766), .ZN(n7574) );
  MUX2_X1 U8342 ( .A(n6698), .B(n6699), .S(n8262), .Z(n6700) );
  AOI21_X2 U8343 ( .B1(n5585), .B2(n5586), .A(n5584), .ZN(n5884) );
  MUX2_X1 U8345 ( .A(n6071), .B(n6072), .S(n6068), .Z(n6073) );
  OAI21_X1 U8346 ( .B1(n3768), .B2(n9913), .A(n9921), .ZN(n9930) );
  MUX2_X1 U8347 ( .A(n4902), .B(n4497), .S(n4856), .Z(n3991) );
  AND2_X1 U8348 ( .A1(n4904), .A2(n4856), .ZN(n5901) );
  AND2_X1 U8349 ( .A1(n4497), .A2(n4498), .ZN(n3770) );
  NAND2_X1 U8350 ( .A1(n4856), .A2(n4907), .ZN(n4498) );
  NAND2_X1 U8351 ( .A1(n3774), .A2(n3772), .ZN(n3771) );
  NAND2_X1 U8352 ( .A1(n20493), .A2(n8099), .ZN(n3774) );
  OR2_X1 U8353 ( .A1(n3776), .A2(n19171), .ZN(n16115) );
  INV_X1 U8354 ( .A(n19171), .ZN(n18088) );
  INV_X1 U8355 ( .A(n16115), .ZN(n16154) );
  NAND2_X1 U8356 ( .A1(n1003), .A2(n12497), .ZN(n3777) );
  XNOR2_X1 U8357 ( .A(n3779), .B(n14164), .ZN(n16171) );
  XNOR2_X1 U8358 ( .A(n16185), .B(n16396), .ZN(n3779) );
  OR2_X1 U8359 ( .A1(n12382), .A2(n12386), .ZN(n3782) );
  NOR2_X1 U8360 ( .A1(n3782), .A2(n11915), .ZN(n3781) );
  NAND2_X1 U8363 ( .A1(n7935), .A2(n7932), .ZN(n3784) );
  NAND2_X1 U8364 ( .A1(n6244), .A2(n20359), .ZN(n3785) );
  NAND2_X1 U8365 ( .A1(n19936), .A2(n19362), .ZN(n17860) );
  MUX2_X1 U8367 ( .A(n17863), .B(n20212), .S(n17672), .Z(n17673) );
  XNOR2_X1 U8369 ( .A(n10514), .B(n10052), .ZN(n3787) );
  AND2_X1 U8370 ( .A1(n3789), .A2(n11177), .ZN(n9378) );
  INV_X1 U8371 ( .A(n10962), .ZN(n3789) );
  INV_X1 U8374 ( .A(n7645), .ZN(n3795) );
  INV_X1 U8375 ( .A(n4343), .ZN(n3925) );
  OR2_X1 U8378 ( .A1(n12600), .A2(n12601), .ZN(n11627) );
  BUF_X1 U8380 ( .A(n19098), .Z(n19094) );
  AND2_X1 U8381 ( .A1(n18834), .A2(n18829), .ZN(n18833) );
  OR2_X1 U8383 ( .A1(n18061), .A2(n19040), .ZN(n18081) );
  XNOR2_X1 U8384 ( .A(n16411), .B(n16410), .ZN(n18097) );
  OR2_X1 U8386 ( .A1(n15785), .A2(n15783), .ZN(n15691) );
  XNOR2_X1 U8387 ( .A(n10180), .B(n10030), .ZN(n10290) );
  OR2_X1 U8388 ( .A1(n12209), .A2(n12208), .ZN(n12187) );
  BUF_X1 U8389 ( .A(n19441), .Z(n19448) );
  INV_X1 U8390 ( .A(n18140), .ZN(n17384) );
  OR2_X1 U8392 ( .A1(n18568), .A2(n18199), .ZN(n18561) );
  OR2_X1 U8393 ( .A1(n18532), .A2(n18529), .ZN(n16816) );
  INV_X1 U8394 ( .A(n17705), .ZN(n17706) );
  XNOR2_X1 U8395 ( .A(n16082), .B(n2392), .ZN(n15798) );
  XNOR2_X1 U8396 ( .A(n6829), .B(n6828), .ZN(n6837) );
  AND2_X1 U8397 ( .A1(n5967), .A2(n5699), .ZN(n5449) );
  OAI21_X1 U8398 ( .B1(n854), .B2(n17186), .A(n17185), .ZN(n19092) );
  XNOR2_X1 U8399 ( .A(n16121), .B(n16120), .ZN(n17835) );
  AND2_X1 U8401 ( .A1(n14327), .A2(n14818), .ZN(n14086) );
  XNOR2_X1 U8403 ( .A(n13521), .B(n13520), .ZN(n13522) );
  OR2_X1 U8406 ( .A1(n15153), .A2(n192), .ZN(n15704) );
  AND2_X1 U8407 ( .A1(n15380), .A2(n15379), .ZN(n15382) );
  INV_X1 U8408 ( .A(n6010), .ZN(n5590) );
  NOR2_X2 U8409 ( .A1(n15186), .A2(n15185), .ZN(n16608) );
  AND2_X1 U8410 ( .A1(n14811), .A2(n14810), .ZN(n14814) );
  NAND2_X1 U8412 ( .A1(n12767), .A2(n12766), .ZN(n12842) );
  OR2_X1 U8413 ( .A1(n18495), .A2(n18498), .ZN(n17644) );
  OAI22_X1 U8414 ( .A1(n17617), .A2(n17616), .B1(n17615), .B2(n1773), .ZN(
        n17621) );
  OR2_X1 U8415 ( .A1(n19396), .A2(n17656), .ZN(n16683) );
  OR2_X1 U8416 ( .A1(n10663), .A2(n11321), .ZN(n10666) );
  XNOR2_X1 U8417 ( .A(n8567), .B(n8566), .ZN(n10761) );
  NOR2_X1 U8419 ( .A1(n18358), .A2(n18290), .ZN(n18288) );
  AND2_X1 U8420 ( .A1(n18489), .A2(n18500), .ZN(n17735) );
  AND2_X1 U8421 ( .A1(n18322), .A2(n18321), .ZN(n18326) );
  OR2_X1 U8423 ( .A1(n18700), .A2(n18699), .ZN(n18705) );
  NOR2_X1 U8424 ( .A1(n16493), .A2(n16492), .ZN(n16494) );
  AND3_X1 U8425 ( .A1(n17234), .A2(n17235), .A3(n17233), .ZN(n18382) );
  AND2_X1 U8426 ( .A1(n16544), .A2(n19955), .ZN(n19315) );
  XNOR2_X1 U8427 ( .A(n17044), .B(n17043), .ZN(n17187) );
  AND2_X1 U8428 ( .A1(n18362), .A2(n18365), .ZN(n17937) );
  NOR3_X1 U8431 ( .A1(n228), .A2(n19958), .A3(n15581), .ZN(n14834) );
  OR2_X1 U8433 ( .A1(n17896), .A2(n19707), .ZN(n16782) );
  XNOR2_X1 U8435 ( .A(n13235), .B(n13236), .ZN(n14269) );
  XNOR2_X1 U8436 ( .A(n10244), .B(n10243), .ZN(n11120) );
  OR2_X1 U8437 ( .A1(n4827), .A2(n5258), .ZN(n4671) );
  OR2_X1 U8438 ( .A1(n19227), .A2(n19754), .ZN(n19219) );
  OR2_X1 U8439 ( .A1(n11120), .A2(n11880), .ZN(n10810) );
  INV_X1 U8442 ( .A(n15295), .ZN(n14944) );
  AND2_X1 U8443 ( .A1(n11871), .A2(n11390), .ZN(n11303) );
  OAI211_X2 U8445 ( .C1(n10193), .C2(n11427), .A(n10192), .B(n10191), .ZN(
        n11990) );
  AOI21_X2 U8447 ( .B1(n9003), .B2(n7776), .A(n7775), .ZN(n9667) );
  NOR2_X1 U8448 ( .A1(n12648), .A2(n12686), .ZN(n12093) );
  AOI22_X1 U8451 ( .A1(n16497), .A2(n19403), .B1(n19402), .B2(n16307), .ZN(
        n19182) );
  AND2_X1 U8452 ( .A1(n19952), .A2(n12311), .ZN(n11905) );
  AND2_X1 U8453 ( .A1(n4632), .A2(n5743), .ZN(n3796) );
  AND3_X1 U8454 ( .A1(n12362), .A2(n12363), .A3(n12510), .ZN(n3798) );
  OR2_X1 U8455 ( .A1(n8934), .A2(n8933), .ZN(n3799) );
  AND2_X1 U8456 ( .A1(n9330), .A2(n9328), .ZN(n3800) );
  AND3_X1 U8457 ( .A1(n20215), .A2(n12281), .A3(n12042), .ZN(n3801) );
  AND2_X1 U8458 ( .A1(n5219), .A2(n5217), .ZN(n3802) );
  XNOR2_X1 U8459 ( .A(n3803), .B(n7351), .ZN(n7470) );
  XOR2_X1 U8460 ( .A(n7350), .B(n7349), .Z(n3803) );
  AND2_X1 U8461 ( .A1(n6059), .A2(n906), .ZN(n3804) );
  XOR2_X1 U8462 ( .A(n6737), .B(n6209), .Z(n3805) );
  OR2_X1 U8463 ( .A1(n7510), .A2(n7675), .ZN(n3808) );
  OR2_X1 U8464 ( .A1(n8325), .A2(n7585), .ZN(n3809) );
  XOR2_X1 U8465 ( .A(n9989), .B(n9988), .Z(n3810) );
  XOR2_X1 U8466 ( .A(n10616), .B(n10615), .Z(n3812) );
  OR2_X1 U8467 ( .A1(n12334), .A2(n12332), .ZN(n3813) );
  AND2_X1 U8468 ( .A1(n11495), .A2(n11493), .ZN(n3814) );
  OR2_X1 U8470 ( .A1(n15430), .A2(n15531), .ZN(n3817) );
  OR2_X1 U8471 ( .A1(n20263), .A2(n14482), .ZN(n3818) );
  AND2_X1 U8472 ( .A1(n15496), .A2(n15500), .ZN(n3819) );
  AND3_X1 U8473 ( .A1(n14637), .A2(n20473), .A3(n14512), .ZN(n3820) );
  AND2_X1 U8474 ( .A1(n19502), .A2(n15516), .ZN(n3821) );
  INV_X1 U8475 ( .A(n14316), .ZN(n13164) );
  XOR2_X1 U8476 ( .A(n13573), .B(n13574), .Z(n3823) );
  AND2_X1 U8477 ( .A1(n15413), .A2(n15553), .ZN(n3824) );
  XNOR2_X1 U8478 ( .A(n16074), .B(n16073), .ZN(n17878) );
  INV_X1 U8479 ( .A(n18519), .ZN(n18184) );
  OR2_X1 U8480 ( .A1(n16101), .A2(n17891), .ZN(n3825) );
  BUF_X1 U8481 ( .A(n16155), .Z(n18319) );
  OR2_X1 U8482 ( .A1(n17715), .A2(n17835), .ZN(n3826) );
  OR2_X1 U8483 ( .A1(n19381), .A2(n19439), .ZN(n3827) );
  AND2_X1 U8484 ( .A1(n19441), .A2(n19444), .ZN(n3828) );
  BUF_X1 U8485 ( .A(n19182), .Z(n19189) );
  NAND3_X1 U8486 ( .A1(n18666), .A2(n17964), .A3(n19735), .ZN(n3829) );
  OR2_X1 U8487 ( .A1(n5107), .A2(n5101), .ZN(n4450) );
  OR2_X1 U8489 ( .A1(n5095), .A2(n4405), .ZN(n3859) );
  INV_X1 U8490 ( .A(n4319), .ZN(n4127) );
  OR2_X1 U8491 ( .A1(n4518), .A2(n4343), .ZN(n4344) );
  INV_X1 U8492 ( .A(Plaintext[23]), .ZN(n3874) );
  OR2_X1 U8493 ( .A1(n4011), .A2(n4611), .ZN(n4612) );
  XNOR2_X1 U8494 ( .A(Key[159]), .B(Plaintext[159]), .ZN(n4575) );
  OR2_X1 U8496 ( .A1(n4669), .A2(n4214), .ZN(n4425) );
  OR2_X1 U8497 ( .A1(n4627), .A2(n4626), .ZN(n4628) );
  OAI21_X1 U8498 ( .B1(n4125), .B2(n4127), .A(n4126), .ZN(n4130) );
  NAND2_X1 U8500 ( .A1(n4838), .A2(n4837), .ZN(n5492) );
  INV_X1 U8501 ( .A(n5766), .ZN(n5545) );
  OR2_X1 U8502 ( .A1(n5088), .A2(n19776), .ZN(n4438) );
  OR2_X1 U8504 ( .A1(n4954), .A2(n4953), .ZN(n4477) );
  INV_X1 U8505 ( .A(n5559), .ZN(n3929) );
  OR2_X1 U8506 ( .A1(n5997), .A2(n5998), .ZN(n5813) );
  INV_X1 U8507 ( .A(n6129), .ZN(n5356) );
  OR2_X1 U8508 ( .A1(n5802), .A2(n5382), .ZN(n6190) );
  INV_X1 U8509 ( .A(n6379), .ZN(n5730) );
  AND2_X1 U8510 ( .A1(n6052), .A2(n6048), .ZN(n5558) );
  INV_X1 U8511 ( .A(n5393), .ZN(n5368) );
  INV_X1 U8513 ( .A(n5502), .ZN(n5122) );
  OR2_X1 U8516 ( .A1(n5317), .A2(n5581), .ZN(n5150) );
  INV_X1 U8517 ( .A(n5899), .ZN(n5908) );
  NOR2_X1 U8518 ( .A1(n284), .A2(n5953), .ZN(n5950) );
  OAI211_X1 U8519 ( .C1(n5593), .C2(n5594), .A(n5592), .B(n5591), .ZN(n7115)
         );
  OR2_X1 U8520 ( .A1(n5855), .A2(n5612), .ZN(n5353) );
  OR2_X1 U8521 ( .A1(n5363), .A2(n4598), .ZN(n5215) );
  OR2_X1 U8522 ( .A1(n7948), .A2(n7953), .ZN(n7168) );
  XNOR2_X1 U8523 ( .A(n6605), .B(n6604), .ZN(n7632) );
  OR2_X1 U8525 ( .A1(n20360), .A2(n7936), .ZN(n7761) );
  XNOR2_X1 U8526 ( .A(n6671), .B(n6670), .ZN(n7568) );
  BUF_X1 U8527 ( .A(n7632), .Z(n7633) );
  INV_X1 U8528 ( .A(n8029), .ZN(n7469) );
  INV_X1 U8529 ( .A(n8011), .ZN(n8012) );
  INV_X1 U8531 ( .A(n7407), .ZN(n7077) );
  XNOR2_X1 U8532 ( .A(n5238), .B(n5239), .ZN(n7877) );
  OR2_X1 U8533 ( .A1(n20180), .A2(n7644), .ZN(n6468) );
  INV_X1 U8535 ( .A(n8055), .ZN(n8052) );
  OR2_X1 U8536 ( .A1(n7003), .A2(n7903), .ZN(n6284) );
  XNOR2_X1 U8537 ( .A(n6493), .B(n6492), .ZN(n6702) );
  INV_X1 U8538 ( .A(n6837), .ZN(n7724) );
  INV_X1 U8539 ( .A(n8131), .ZN(n8138) );
  XNOR2_X1 U8540 ( .A(n6781), .B(n6780), .ZN(n7684) );
  OR2_X1 U8541 ( .A1(n7958), .A2(n7956), .ZN(n7917) );
  AND2_X1 U8542 ( .A1(n7749), .A2(n7508), .ZN(n6908) );
  OR2_X1 U8543 ( .A1(n7676), .A2(n7673), .ZN(n7513) );
  AOI22_X1 U8544 ( .A1(n20012), .A2(n7445), .B1(n8280), .B2(n8286), .ZN(n7796)
         );
  AOI22_X1 U8545 ( .A1(n8154), .A2(n8153), .B1(n8262), .B2(n8152), .ZN(n8156)
         );
  AND2_X1 U8546 ( .A1(n8185), .A2(n8184), .ZN(n8187) );
  INV_X1 U8547 ( .A(n9346), .ZN(n9567) );
  INV_X1 U8548 ( .A(n8482), .ZN(n9368) );
  NOR2_X1 U8549 ( .A1(n8423), .A2(n19515), .ZN(n8327) );
  INV_X1 U8550 ( .A(n9934), .ZN(n10037) );
  INV_X1 U8551 ( .A(n11339), .ZN(n11340) );
  XNOR2_X1 U8552 ( .A(n9878), .B(n9635), .ZN(n10462) );
  INV_X1 U8553 ( .A(n11489), .ZN(n11494) );
  INV_X1 U8554 ( .A(n9294), .ZN(n8680) );
  XNOR2_X1 U8555 ( .A(n9653), .B(n9652), .ZN(n10684) );
  AOI21_X1 U8556 ( .B1(n11564), .B2(n11567), .A(n11469), .ZN(n11470) );
  XNOR2_X1 U8557 ( .A(n10433), .B(n9387), .ZN(n9390) );
  NOR2_X1 U8558 ( .A1(n11253), .A2(n11255), .ZN(n11323) );
  XNOR2_X1 U8559 ( .A(n10075), .B(n10076), .ZN(n10112) );
  OR2_X1 U8560 ( .A1(n19750), .A2(n11866), .ZN(n11304) );
  OR2_X1 U8561 ( .A1(n11452), .A2(n11110), .ZN(n10734) );
  XNOR2_X1 U8563 ( .A(n9990), .B(n3810), .ZN(n10742) );
  BUF_X1 U8564 ( .A(n10783), .Z(n11116) );
  NOR2_X1 U8565 ( .A1(n19959), .A2(n11133), .ZN(n11421) );
  INV_X1 U8566 ( .A(n11445), .ZN(n11209) );
  NOR2_X1 U8567 ( .A1(n11513), .A2(n19864), .ZN(n11574) );
  AND2_X1 U8568 ( .A1(n10704), .A2(n11152), .ZN(n10707) );
  BUF_X1 U8569 ( .A(n9666), .Z(n11383) );
  OR2_X1 U8570 ( .A1(n12616), .A2(n12053), .ZN(n12055) );
  NOR2_X1 U8571 ( .A1(n12545), .A2(n12544), .ZN(n12555) );
  INV_X1 U8572 ( .A(n12809), .ZN(n12487) );
  OR2_X1 U8573 ( .A1(n12508), .A2(n12359), .ZN(n9886) );
  AND2_X1 U8574 ( .A1(n11686), .A2(n11863), .ZN(n11730) );
  INV_X1 U8575 ( .A(n11841), .ZN(n12181) );
  XNOR2_X1 U8576 ( .A(n13481), .B(n457), .ZN(n13432) );
  OAI21_X1 U8577 ( .B1(n11908), .B2(n11907), .A(n11906), .ZN(n13451) );
  AND2_X1 U8578 ( .A1(n12383), .A2(n12382), .ZN(n12388) );
  OR2_X1 U8579 ( .A1(n12595), .A2(n12201), .ZN(n12060) );
  OR2_X1 U8580 ( .A1(n12333), .A2(n12332), .ZN(n12344) );
  AND2_X1 U8581 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  INV_X1 U8582 ( .A(n13481), .ZN(n12984) );
  OAI21_X1 U8584 ( .B1(n11974), .B2(n11667), .A(n11666), .ZN(n11668) );
  XNOR2_X1 U8585 ( .A(n13432), .B(n13797), .ZN(n13434) );
  XNOR2_X1 U8586 ( .A(n12962), .B(n2347), .ZN(n12964) );
  XNOR2_X1 U8587 ( .A(n13714), .B(n13499), .ZN(n11789) );
  XNOR2_X1 U8588 ( .A(n13477), .B(n13279), .ZN(n13316) );
  OR2_X1 U8589 ( .A1(n14279), .A2(n14555), .ZN(n14280) );
  OR2_X1 U8591 ( .A1(n14132), .A2(n14729), .ZN(n14133) );
  XNOR2_X1 U8592 ( .A(n12970), .B(n13207), .ZN(n12972) );
  XNOR2_X1 U8594 ( .A(n13015), .B(n13014), .ZN(n13872) );
  BUF_X1 U8595 ( .A(n13980), .Z(n14542) );
  INV_X1 U8596 ( .A(n14543), .ZN(n14544) );
  OR2_X1 U8598 ( .A1(n14304), .A2(n14506), .ZN(n13506) );
  XNOR2_X1 U8599 ( .A(n13639), .B(n13638), .ZN(n14388) );
  INV_X1 U8600 ( .A(n14104), .ZN(n14105) );
  AND2_X1 U8601 ( .A1(n3307), .A2(n15296), .ZN(n14768) );
  OR2_X1 U8602 ( .A1(n15696), .A2(n15695), .ZN(n14938) );
  AND2_X1 U8603 ( .A1(n13907), .A2(n14611), .ZN(n14207) );
  AND2_X1 U8604 ( .A1(n19485), .A2(n12877), .ZN(n12878) );
  INV_X1 U8605 ( .A(n14699), .ZN(n14122) );
  AND2_X1 U8606 ( .A1(n14089), .A2(n14088), .ZN(n14090) );
  BUF_X1 U8607 ( .A(n12910), .Z(n14168) );
  XNOR2_X1 U8608 ( .A(n13472), .B(n13473), .ZN(n14425) );
  AND2_X1 U8609 ( .A1(n14508), .A2(n14507), .ZN(n14513) );
  INV_X1 U8610 ( .A(n15600), .ZN(n15271) );
  AND2_X1 U8611 ( .A1(n14434), .A2(n14487), .ZN(n13881) );
  NOR2_X1 U8612 ( .A1(n15606), .A2(n16128), .ZN(n15201) );
  INV_X1 U8613 ( .A(n13982), .ZN(n13133) );
  BUF_X1 U8614 ( .A(n14497), .Z(n14501) );
  OR2_X1 U8615 ( .A1(n15595), .A2(n15748), .ZN(n15519) );
  AND2_X1 U8616 ( .A1(n15636), .A2(n15843), .ZN(n15092) );
  OR2_X1 U8617 ( .A1(n15704), .A2(n13968), .ZN(n13969) );
  OR2_X1 U8618 ( .A1(n15909), .A2(n15907), .ZN(n15416) );
  INV_X1 U8619 ( .A(n14964), .ZN(n14969) );
  BUF_X1 U8620 ( .A(n15655), .Z(n15768) );
  INV_X1 U8621 ( .A(n15532), .ZN(n15086) );
  NAND4_X1 U8622 ( .A1(n15649), .A2(n15648), .A3(n15647), .A4(n15646), .ZN(
        n15994) );
  NOR2_X1 U8623 ( .A1(n14876), .A2(n14875), .ZN(n14877) );
  OR2_X1 U8624 ( .A1(n13861), .A2(n13860), .ZN(n13862) );
  OAI21_X1 U8625 ( .B1(n14959), .B2(n15284), .A(n14958), .ZN(n15020) );
  OAI21_X1 U8626 ( .B1(n15290), .B2(n15289), .A(n15288), .ZN(n16992) );
  OR2_X1 U8627 ( .A1(n2005), .A2(n15445), .ZN(n15324) );
  OR2_X1 U8628 ( .A1(n15540), .A2(n15898), .ZN(n15541) );
  XNOR2_X1 U8629 ( .A(n16419), .B(n16418), .ZN(n16422) );
  INV_X1 U8630 ( .A(n18946), .ZN(n17687) );
  XNOR2_X1 U8631 ( .A(n16593), .B(n16706), .ZN(n17357) );
  BUF_X1 U8632 ( .A(n19782), .Z(n16420) );
  XNOR2_X1 U8633 ( .A(n15798), .B(n17426), .ZN(n15810) );
  AND2_X1 U8634 ( .A1(n17492), .A2(n17491), .ZN(n17496) );
  AND2_X1 U8635 ( .A1(n19943), .A2(n20348), .ZN(n17966) );
  XNOR2_X1 U8636 ( .A(n16428), .B(n16427), .ZN(n17568) );
  INV_X1 U8638 ( .A(n17568), .ZN(n18095) );
  XNOR2_X1 U8639 ( .A(n17364), .B(n17363), .ZN(n17758) );
  OAI21_X1 U8640 ( .B1(n18115), .B2(n19885), .A(n17968), .ZN(n17460) );
  AND2_X1 U8641 ( .A1(n18033), .A2(n18270), .ZN(n17768) );
  OR2_X1 U8642 ( .A1(n18019), .A2(n18938), .ZN(n17705) );
  XNOR2_X1 U8643 ( .A(n16133), .B(n16132), .ZN(n17063) );
  INV_X1 U8644 ( .A(n17892), .ZN(n16784) );
  OR2_X1 U8645 ( .A1(n17676), .A2(n17078), .ZN(n16314) );
  XNOR2_X1 U8646 ( .A(n15790), .B(n15789), .ZN(n16540) );
  BUF_X1 U8649 ( .A(n17501), .Z(n17504) );
  AOI21_X1 U8650 ( .B1(n17159), .B2(n17158), .A(n17157), .ZN(n17623) );
  AND2_X1 U8651 ( .A1(n20109), .A2(n18097), .ZN(n17164) );
  NOR2_X1 U8655 ( .A1(n20273), .A2(n16673), .ZN(n16636) );
  INV_X1 U8656 ( .A(n19432), .ZN(n19418) );
  OR2_X1 U8657 ( .A1(n18240), .A2(n20128), .ZN(n18247) );
  AND2_X1 U8658 ( .A1(n20003), .A2(n18412), .ZN(n18406) );
  BUF_X1 U8659 ( .A(n17729), .Z(n17640) );
  OR2_X1 U8660 ( .A1(n17476), .A2(n17475), .ZN(n17477) );
  OR2_X1 U8663 ( .A1(n17719), .A2(n17718), .ZN(n17720) );
  OR2_X1 U8665 ( .A1(n18320), .A2(n16155), .ZN(n18321) );
  BUF_X1 U8666 ( .A(n18621), .Z(n18613) );
  OR2_X1 U8667 ( .A1(n19425), .A2(n19409), .ZN(n19428) );
  AND3_X1 U8668 ( .A1(n17789), .A2(n19166), .A3(n17791), .ZN(n17796) );
  INV_X1 U8669 ( .A(Plaintext[71]), .ZN(n3830) );
  XNOR2_X1 U8670 ( .A(n3830), .B(Key[71]), .ZN(n4220) );
  NAND2_X1 U8671 ( .A1(n4223), .A2(n164), .ZN(n3832) );
  INV_X1 U8672 ( .A(Plaintext[70]), .ZN(n3831) );
  XNOR2_X1 U8673 ( .A(Key[66]), .B(Plaintext[66]), .ZN(n4657) );
  AOI21_X1 U8674 ( .B1(n3979), .B2(n4657), .A(n164), .ZN(n3833) );
  INV_X1 U8675 ( .A(n3855), .ZN(n3839) );
  INV_X1 U8677 ( .A(Plaintext[85]), .ZN(n3834) );
  XNOR2_X1 U8678 ( .A(n3834), .B(Key[85]), .ZN(n4663) );
  INV_X1 U8679 ( .A(Plaintext[84]), .ZN(n3835) );
  XNOR2_X1 U8680 ( .A(n3835), .B(Key[84]), .ZN(n4664) );
  INV_X1 U8681 ( .A(n4664), .ZN(n4816) );
  INV_X1 U8682 ( .A(Plaintext[89]), .ZN(n3836) );
  INV_X1 U8683 ( .A(n4410), .ZN(n4411) );
  XNOR2_X1 U8684 ( .A(Key[88]), .B(Plaintext[88]), .ZN(n5071) );
  NAND2_X1 U8685 ( .A1(n4411), .A2(n5071), .ZN(n4814) );
  INV_X1 U8686 ( .A(Plaintext[80]), .ZN(n3840) );
  XNOR2_X1 U8687 ( .A(n3840), .B(Key[80]), .ZN(n3843) );
  INV_X1 U8688 ( .A(n3843), .ZN(n4835) );
  INV_X1 U8689 ( .A(Plaintext[83]), .ZN(n3841) );
  XNOR2_X1 U8690 ( .A(n3841), .B(Key[83]), .ZN(n3846) );
  INV_X1 U8691 ( .A(n3846), .ZN(n4675) );
  INV_X1 U8692 ( .A(n5117), .ZN(n4834) );
  NAND2_X1 U8693 ( .A1(n3842), .A2(n4834), .ZN(n3850) );
  INV_X1 U8694 ( .A(Plaintext[82]), .ZN(n3844) );
  XNOR2_X1 U8695 ( .A(Key[78]), .B(Plaintext[78]), .ZN(n5118) );
  INV_X1 U8696 ( .A(n5118), .ZN(n3845) );
  NAND2_X1 U8697 ( .A1(n3845), .A2(n19508), .ZN(n3847) );
  MUX2_X1 U8698 ( .A(n3848), .B(n3847), .S(n5116), .Z(n3849) );
  INV_X1 U8699 ( .A(n3855), .ZN(n6058) );
  INV_X1 U8700 ( .A(n4670), .ZN(n3854) );
  INV_X1 U8701 ( .A(Plaintext[77]), .ZN(n3851) );
  XNOR2_X1 U8702 ( .A(Key[74]), .B(Plaintext[74]), .ZN(n4669) );
  INV_X1 U8703 ( .A(n4669), .ZN(n4828) );
  INV_X1 U8704 ( .A(n4214), .ZN(n4673) );
  INV_X1 U8705 ( .A(n5258), .ZN(n4668) );
  NOR2_X1 U8706 ( .A1(n4827), .A2(n4829), .ZN(n4213) );
  INV_X1 U8707 ( .A(n4213), .ZN(n3852) );
  OAI211_X1 U8708 ( .C1(n4670), .C2(n4673), .A(n4668), .B(n3852), .ZN(n3853)
         );
  NAND3_X1 U8709 ( .A1(n6058), .A2(n906), .A3(n6057), .ZN(n3866) );
  XNOR2_X1 U8710 ( .A(Key[99]), .B(Plaintext[99]), .ZN(n5081) );
  XNOR2_X1 U8711 ( .A(Key[97]), .B(Plaintext[97]), .ZN(n4719) );
  INV_X1 U8712 ( .A(n4719), .ZN(n5074) );
  XNOR2_X1 U8713 ( .A(Key[96]), .B(Plaintext[96]), .ZN(n5079) );
  XNOR2_X1 U8714 ( .A(Key[100]), .B(Plaintext[100]), .ZN(n5077) );
  INV_X1 U8715 ( .A(n5077), .ZN(n4081) );
  INV_X1 U8718 ( .A(Plaintext[95]), .ZN(n3856) );
  INV_X1 U8719 ( .A(Plaintext[90]), .ZN(n3857) );
  INV_X1 U8721 ( .A(Plaintext[91]), .ZN(n3858) );
  OAI211_X1 U8722 ( .C1(n5093), .C2(n4788), .A(n3859), .B(n2461), .ZN(n3862)
         );
  INV_X1 U8723 ( .A(Plaintext[94]), .ZN(n3860) );
  XNOR2_X1 U8724 ( .A(n3860), .B(Key[94]), .ZN(n5094) );
  INV_X1 U8725 ( .A(n5094), .ZN(n4783) );
  OAI21_X1 U8726 ( .B1(n5098), .B2(n4783), .A(n5092), .ZN(n3861) );
  NAND3_X1 U8728 ( .A1(n6064), .A2(n20670), .A3(n6059), .ZN(n3864) );
  NAND4_X2 U8729 ( .A1(n3865), .A2(n3867), .A3(n3866), .A4(n3864), .ZN(n7201)
         );
  XNOR2_X1 U8730 ( .A(n7201), .B(n2263), .ZN(n3902) );
  INV_X1 U8731 ( .A(Plaintext[32]), .ZN(n3868) );
  XNOR2_X1 U8732 ( .A(n3868), .B(Key[32]), .ZN(n4953) );
  INV_X1 U8733 ( .A(Plaintext[31]), .ZN(n3869) );
  INV_X1 U8735 ( .A(n4474), .ZN(n4913) );
  INV_X1 U8736 ( .A(Plaintext[34]), .ZN(n3870) );
  NAND2_X1 U8738 ( .A1(n3871), .A2(n4952), .ZN(n3873) );
  INV_X1 U8739 ( .A(n4911), .ZN(n4140) );
  OAI21_X1 U8740 ( .B1(n4912), .B2(n4913), .A(n4140), .ZN(n3872) );
  NAND2_X1 U8742 ( .A1(n4021), .A2(n4928), .ZN(n4978) );
  INV_X1 U8743 ( .A(Plaintext[18]), .ZN(n3875) );
  NAND2_X1 U8744 ( .A1(n4131), .A2(n4296), .ZN(n4980) );
  XNOR2_X1 U8745 ( .A(Key[22]), .B(Plaintext[22]), .ZN(n4974) );
  INV_X1 U8746 ( .A(n4297), .ZN(n4932) );
  MUX2_X1 U8747 ( .A(n4974), .B(n4932), .S(n4131), .Z(n3879) );
  INV_X1 U8748 ( .A(n4978), .ZN(n3877) );
  AND2_X1 U8749 ( .A1(n4979), .A2(n4928), .ZN(n3876) );
  INV_X1 U8750 ( .A(n4622), .ZN(n4290) );
  XNOR2_X1 U8751 ( .A(Key[4]), .B(Plaintext[4]), .ZN(n4285) );
  INV_X1 U8752 ( .A(n4285), .ZN(n3882) );
  INV_X1 U8753 ( .A(Plaintext[0]), .ZN(n3880) );
  INV_X1 U8754 ( .A(n4169), .ZN(n4621) );
  AOI21_X1 U8755 ( .B1(n4630), .B2(n4621), .A(n4623), .ZN(n3886) );
  INV_X1 U8756 ( .A(Plaintext[2]), .ZN(n3881) );
  NAND2_X1 U8757 ( .A1(n4290), .A2(n4171), .ZN(n3884) );
  XNOR2_X1 U8758 ( .A(Key[1]), .B(Plaintext[1]), .ZN(n4626) );
  INV_X1 U8759 ( .A(n4626), .ZN(n4170) );
  NAND2_X1 U8760 ( .A1(n4170), .A2(n4623), .ZN(n3883) );
  AOI21_X1 U8761 ( .B1(n3884), .B2(n3883), .A(n3882), .ZN(n3885) );
  XNOR2_X1 U8762 ( .A(Key[7]), .B(Plaintext[7]), .ZN(n4324) );
  INV_X1 U8763 ( .A(n4324), .ZN(n4647) );
  XNOR2_X1 U8764 ( .A(Key[6]), .B(Plaintext[6]), .ZN(n4318) );
  INV_X1 U8765 ( .A(n4318), .ZN(n4646) );
  NAND2_X1 U8766 ( .A1(n4647), .A2(n4646), .ZN(n3888) );
  XNOR2_X2 U8767 ( .A(Key[8]), .B(Plaintext[8]), .ZN(n4640) );
  INV_X1 U8768 ( .A(n4640), .ZN(n4648) );
  INV_X1 U8769 ( .A(Plaintext[11]), .ZN(n3887) );
  XNOR2_X1 U8770 ( .A(n3887), .B(Key[11]), .ZN(n4317) );
  MUX2_X1 U8771 ( .A(n3888), .B(n4648), .S(n4325), .Z(n3891) );
  INV_X1 U8773 ( .A(n4125), .ZN(n4641) );
  NAND2_X1 U8774 ( .A1(n4319), .A2(n4324), .ZN(n4323) );
  INV_X1 U8775 ( .A(n4323), .ZN(n3889) );
  OAI21_X1 U8776 ( .B1(n4641), .B2(n4325), .A(n3889), .ZN(n3890) );
  XNOR2_X1 U8777 ( .A(Key[24]), .B(Plaintext[24]), .ZN(n4114) );
  INV_X1 U8778 ( .A(n4114), .ZN(n4470) );
  INV_X1 U8779 ( .A(n4118), .ZN(n4941) );
  INV_X1 U8780 ( .A(n4945), .ZN(n4467) );
  INV_X1 U8781 ( .A(n4940), .ZN(n4117) );
  INV_X1 U8782 ( .A(Plaintext[28]), .ZN(n3893) );
  XNOR2_X1 U8783 ( .A(n3893), .B(Key[28]), .ZN(n4946) );
  NAND3_X1 U8784 ( .A1(n4946), .A2(n4945), .A3(n4947), .ZN(n3894) );
  OAI211_X1 U8785 ( .C1(n3896), .C2(n4947), .A(n3895), .B(n3894), .ZN(n5795)
         );
  XNOR2_X1 U8786 ( .A(Key[15]), .B(Plaintext[15]), .ZN(n3897) );
  NAND2_X1 U8788 ( .A1(n4988), .A2(n4982), .ZN(n4005) );
  INV_X1 U8789 ( .A(n3897), .ZN(n4983) );
  XNOR2_X1 U8790 ( .A(Key[13]), .B(Plaintext[13]), .ZN(n4618) );
  NAND2_X1 U8791 ( .A1(n4983), .A2(n4618), .ZN(n3898) );
  INV_X1 U8793 ( .A(n4306), .ZN(n4003) );
  XNOR2_X1 U8794 ( .A(Key[16]), .B(Plaintext[16]), .ZN(n4305) );
  NAND2_X1 U8795 ( .A1(n4003), .A2(n4305), .ZN(n3900) );
  NAND2_X1 U8796 ( .A1(n4988), .A2(n4306), .ZN(n3899) );
  INV_X1 U8797 ( .A(n5017), .ZN(n5014) );
  INV_X1 U8799 ( .A(n5018), .ZN(n4736) );
  XNOR2_X1 U8800 ( .A(Key[139]), .B(Plaintext[139]), .ZN(n4277) );
  INV_X1 U8801 ( .A(n4277), .ZN(n5012) );
  NAND2_X1 U8802 ( .A1(n5012), .A2(n4734), .ZN(n3903) );
  INV_X1 U8804 ( .A(n4734), .ZN(n3904) );
  XNOR2_X1 U8805 ( .A(Key[138]), .B(Plaintext[138]), .ZN(n4110) );
  INV_X1 U8806 ( .A(n4110), .ZN(n4554) );
  INV_X1 U8807 ( .A(Plaintext[161]), .ZN(n3906) );
  XNOR2_X2 U8808 ( .A(n3906), .B(Key[161]), .ZN(n4370) );
  INV_X1 U8809 ( .A(n4576), .ZN(n4570) );
  XNOR2_X1 U8811 ( .A(Key[157]), .B(Plaintext[157]), .ZN(n4507) );
  NAND2_X1 U8812 ( .A1(n4507), .A2(n4575), .ZN(n4510) );
  NAND3_X1 U8813 ( .A1(n4510), .A2(n4576), .A3(n3907), .ZN(n3910) );
  INV_X1 U8814 ( .A(n4370), .ZN(n4511) );
  INV_X1 U8815 ( .A(Plaintext[156]), .ZN(n3908) );
  INV_X1 U8816 ( .A(n4571), .ZN(n4573) );
  NAND3_X1 U8817 ( .A1(n4511), .A2(n4372), .A3(n4573), .ZN(n3909) );
  INV_X1 U8818 ( .A(n6048), .ZN(n5139) );
  NAND2_X1 U8819 ( .A1(n5328), .A2(n5139), .ZN(n3920) );
  INV_X1 U8820 ( .A(Plaintext[149]), .ZN(n3911) );
  XNOR2_X1 U8821 ( .A(n3911), .B(Key[149]), .ZN(n5005) );
  INV_X1 U8822 ( .A(n5005), .ZN(n4746) );
  INV_X1 U8823 ( .A(n5010), .ZN(n3912) );
  NAND2_X1 U8824 ( .A1(n4746), .A2(n3912), .ZN(n4557) );
  INV_X1 U8826 ( .A(n4206), .ZN(n4561) );
  NAND2_X1 U8828 ( .A1(n4746), .A2(n4745), .ZN(n3913) );
  NAND2_X1 U8829 ( .A1(n4561), .A2(n3913), .ZN(n3915) );
  NAND2_X1 U8830 ( .A1(n4248), .A2(n4744), .ZN(n3914) );
  INV_X1 U8831 ( .A(n6049), .ZN(n5557) );
  XNOR2_X2 U8832 ( .A(Key[153]), .B(Plaintext[153]), .ZN(n4504) );
  MUX2_X1 U8833 ( .A(n4756), .B(n4504), .S(n4752), .Z(n3918) );
  INV_X1 U8834 ( .A(n4504), .ZN(n4563) );
  XNOR2_X1 U8835 ( .A(Key[151]), .B(Plaintext[151]), .ZN(n4565) );
  INV_X1 U8836 ( .A(n4565), .ZN(n4755) );
  INV_X1 U8837 ( .A(Plaintext[150]), .ZN(n3916) );
  NAND2_X1 U8838 ( .A1(n4754), .A2(n4504), .ZN(n3917) );
  INV_X1 U8839 ( .A(n4567), .ZN(n4198) );
  AOI21_X1 U8840 ( .B1(n3920), .B2(n3919), .A(n6052), .ZN(n3936) );
  XNOR2_X1 U8841 ( .A(Key[171]), .B(Plaintext[171]), .ZN(n4518) );
  INV_X1 U8842 ( .A(n4518), .ZN(n3922) );
  INV_X1 U8843 ( .A(Plaintext[169]), .ZN(n3921) );
  NAND2_X1 U8844 ( .A1(n3922), .A2(n4517), .ZN(n4340) );
  INV_X1 U8845 ( .A(n4340), .ZN(n3924) );
  INV_X1 U8847 ( .A(Plaintext[170]), .ZN(n3923) );
  OAI21_X1 U8848 ( .B1(n3924), .B2(n4522), .A(n4343), .ZN(n3928) );
  INV_X1 U8849 ( .A(n4517), .ZN(n4520) );
  INV_X1 U8850 ( .A(Plaintext[172]), .ZN(n3926) );
  XNOR2_X1 U8851 ( .A(n3926), .B(Key[172]), .ZN(n4342) );
  NAND2_X1 U8852 ( .A1(n3943), .A2(n4342), .ZN(n3927) );
  AND2_X2 U8853 ( .A1(n3928), .A2(n3927), .ZN(n5559) );
  NAND2_X1 U8854 ( .A1(n3929), .A2(n6048), .ZN(n4995) );
  INV_X1 U8856 ( .A(n3948), .ZN(n4542) );
  NAND2_X1 U8858 ( .A1(n4539), .A2(n4350), .ZN(n3931) );
  INV_X1 U8859 ( .A(Plaintext[164]), .ZN(n3930) );
  OAI211_X1 U8860 ( .C1(n4542), .C2(n4539), .A(n3931), .B(n4347), .ZN(n3933)
         );
  NAND2_X1 U8861 ( .A1(n5559), .A2(n6050), .ZN(n3934) );
  OAI22_X1 U8862 ( .A1(n6054), .A2(n4995), .B1(n3934), .B2(n3351), .ZN(n3935)
         );
  XNOR2_X1 U8863 ( .A(Key[175]), .B(Plaintext[175]), .ZN(n4532) );
  XNOR2_X1 U8864 ( .A(Key[174]), .B(Plaintext[174]), .ZN(n4528) );
  NAND2_X1 U8865 ( .A1(n19524), .A2(n4529), .ZN(n3938) );
  INV_X1 U8866 ( .A(Plaintext[179]), .ZN(n3937) );
  XNOR2_X2 U8867 ( .A(n3937), .B(Key[179]), .ZN(n4633) );
  OAI211_X1 U8868 ( .C1(n19524), .C2(n4532), .A(n3938), .B(n4633), .ZN(n5576)
         );
  INV_X1 U8869 ( .A(n4633), .ZN(n4337) );
  INV_X1 U8870 ( .A(Plaintext[178]), .ZN(n3939) );
  NAND2_X2 U8872 ( .A1(n5575), .A2(n5576), .ZN(n5408) );
  NAND2_X1 U8873 ( .A1(n4343), .A2(n4516), .ZN(n3942) );
  AND2_X1 U8875 ( .A1(n4520), .A2(n4523), .ZN(n3941) );
  INV_X1 U8876 ( .A(n4342), .ZN(n4160) );
  INV_X1 U8878 ( .A(n5581), .ZN(n5404) );
  INV_X1 U8879 ( .A(Plaintext[182]), .ZN(n3944) );
  INV_X1 U8880 ( .A(Plaintext[181]), .ZN(n3945) );
  INV_X1 U8881 ( .A(n4313), .ZN(n4603) );
  INV_X1 U8882 ( .A(Plaintext[183]), .ZN(n3946) );
  XNOR2_X1 U8883 ( .A(n3946), .B(Key[183]), .ZN(n4152) );
  INV_X1 U8884 ( .A(Plaintext[180]), .ZN(n3947) );
  INV_X1 U8885 ( .A(n4548), .ZN(n4353) );
  XNOR2_X1 U8886 ( .A(Key[185]), .B(Plaintext[185]), .ZN(n4602) );
  XNOR2_X1 U8887 ( .A(Key[184]), .B(Plaintext[184]), .ZN(n4601) );
  NAND2_X1 U8888 ( .A1(n4355), .A2(n4601), .ZN(n4312) );
  INV_X1 U8889 ( .A(n4602), .ZN(n4607) );
  OAI211_X1 U8890 ( .C1(n4541), .C2(n4349), .A(n4542), .B(n4539), .ZN(n3950)
         );
  NAND2_X1 U8891 ( .A1(n3950), .A2(n3949), .ZN(n3951) );
  XNOR2_X1 U8892 ( .A(Key[189]), .B(Plaintext[189]), .ZN(n4176) );
  INV_X1 U8893 ( .A(n4176), .ZN(n4011) );
  INV_X1 U8894 ( .A(Plaintext[186]), .ZN(n3952) );
  XNOR2_X1 U8895 ( .A(n3952), .B(Key[186]), .ZN(n4611) );
  NAND2_X1 U8896 ( .A1(n4011), .A2(n4611), .ZN(n4010) );
  INV_X1 U8897 ( .A(Plaintext[187]), .ZN(n3953) );
  INV_X1 U8898 ( .A(n4611), .ZN(n4364) );
  XNOR2_X1 U8899 ( .A(Key[190]), .B(Plaintext[190]), .ZN(n4013) );
  NAND2_X1 U8900 ( .A1(n1537), .A2(n748), .ZN(n3954) );
  INV_X1 U8901 ( .A(n4365), .ZN(n4609) );
  OR2_X1 U8902 ( .A1(n4010), .A2(n748), .ZN(n5574) );
  NAND2_X1 U8903 ( .A1(n5573), .A2(n5574), .ZN(n5405) );
  AND2_X1 U8904 ( .A1(n4169), .A2(n4623), .ZN(n4291) );
  OAI21_X1 U8905 ( .B1(n4170), .B2(n4621), .A(n4171), .ZN(n3956) );
  INV_X1 U8907 ( .A(n4171), .ZN(n4631) );
  AOI21_X1 U8908 ( .B1(n4018), .B2(n4627), .A(n4285), .ZN(n3957) );
  XNOR2_X1 U8910 ( .A(n6693), .B(n7304), .ZN(n3962) );
  XNOR2_X1 U8911 ( .A(n3963), .B(n3962), .ZN(n4065) );
  INV_X1 U8913 ( .A(n4968), .ZN(n3965) );
  INV_X1 U8914 ( .A(Plaintext[42]), .ZN(n3964) );
  XNOR2_X1 U8915 ( .A(n3964), .B(Key[42]), .ZN(n4970) );
  NAND2_X1 U8916 ( .A1(n3965), .A2(n4970), .ZN(n4967) );
  AND2_X1 U8917 ( .A1(n4969), .A2(n4968), .ZN(n4483) );
  NAND2_X1 U8919 ( .A1(n4965), .A2(n4479), .ZN(n3966) );
  NAND2_X1 U8920 ( .A1(n4483), .A2(n3966), .ZN(n3968) );
  OAI211_X1 U8922 ( .C1(n4967), .C2(n3967), .A(n3968), .B(n4966), .ZN(n5978)
         );
  INV_X1 U8923 ( .A(Plaintext[41]), .ZN(n3969) );
  XNOR2_X2 U8924 ( .A(n3969), .B(Key[41]), .ZN(n4899) );
  NAND2_X1 U8925 ( .A1(n4377), .A2(n4899), .ZN(n3973) );
  INV_X1 U8926 ( .A(Plaintext[37]), .ZN(n3970) );
  XNOR2_X1 U8928 ( .A(Key[39]), .B(Plaintext[39]), .ZN(n4894) );
  NAND2_X1 U8929 ( .A1(n4960), .A2(n4894), .ZN(n3972) );
  INV_X1 U8930 ( .A(Plaintext[40]), .ZN(n3971) );
  AOI21_X1 U8931 ( .B1(n3973), .B2(n3972), .A(n4962), .ZN(n3976) );
  AOI21_X1 U8932 ( .B1(n3974), .B2(n4136), .A(n3231), .ZN(n3975) );
  NOR2_X1 U8933 ( .A1(n5978), .A2(n6072), .ZN(n3993) );
  NOR2_X1 U8934 ( .A1(n4840), .A2(n4657), .ZN(n4421) );
  INV_X1 U8935 ( .A(Plaintext[65]), .ZN(n3982) );
  NAND2_X1 U8937 ( .A1(n289), .A2(n4652), .ZN(n3986) );
  INV_X1 U8938 ( .A(Plaintext[60]), .ZN(n3983) );
  XNOR2_X1 U8939 ( .A(n3983), .B(Key[60]), .ZN(n4867) );
  INV_X1 U8940 ( .A(Plaintext[62]), .ZN(n3984) );
  NOR2_X1 U8941 ( .A1(n6069), .A2(n5320), .ZN(n3992) );
  INV_X1 U8942 ( .A(Plaintext[49]), .ZN(n3987) );
  XNOR2_X1 U8943 ( .A(n3987), .B(Key[49]), .ZN(n4232) );
  INV_X1 U8944 ( .A(Plaintext[48]), .ZN(n3988) );
  XNOR2_X1 U8945 ( .A(n3988), .B(Key[48]), .ZN(n4497) );
  INV_X1 U8946 ( .A(n4907), .ZN(n4493) );
  XNOR2_X1 U8947 ( .A(Key[52]), .B(Plaintext[52]), .ZN(n4855) );
  NAND2_X1 U8948 ( .A1(n4493), .A2(n4855), .ZN(n3989) );
  INV_X1 U8951 ( .A(n3996), .ZN(n4853) );
  INV_X1 U8952 ( .A(n176), .ZN(n4485) );
  XNOR2_X1 U8953 ( .A(Key[55]), .B(Plaintext[55]), .ZN(n4685) );
  MUX2_X1 U8954 ( .A(n4851), .B(n4682), .S(n4685), .Z(n3998) );
  INV_X1 U8955 ( .A(Plaintext[58]), .ZN(n3994) );
  XNOR2_X1 U8957 ( .A(Key[54]), .B(Plaintext[54]), .ZN(n4391) );
  NAND2_X1 U8958 ( .A1(n178), .A2(n4391), .ZN(n4224) );
  NAND2_X1 U8960 ( .A1(n6068), .A2(n209), .ZN(n4000) );
  OAI21_X1 U8961 ( .B1(n4118), .B2(n4940), .A(n4470), .ZN(n4002) );
  INV_X1 U8962 ( .A(n4305), .ZN(n4989) );
  MUX2_X1 U8963 ( .A(n4005), .B(n4004), .S(n19822), .Z(n4009) );
  INV_X1 U8964 ( .A(n4618), .ZN(n4006) );
  NAND2_X1 U8965 ( .A1(n4988), .A2(n4618), .ZN(n4985) );
  NAND2_X1 U8966 ( .A1(n4007), .A2(n4985), .ZN(n4008) );
  INV_X1 U8967 ( .A(n5395), .ZN(n5367) );
  NAND2_X1 U8968 ( .A1(n1537), .A2(n4615), .ZN(n4366) );
  NAND2_X1 U8970 ( .A1(n4012), .A2(n4011), .ZN(n4014) );
  INV_X1 U8971 ( .A(n4614), .ZN(n4177) );
  NAND2_X1 U8973 ( .A1(n4640), .A2(n4319), .ZN(n4015) );
  OAI21_X1 U8974 ( .B1(n4641), .B2(n4640), .A(n4015), .ZN(n4016) );
  INV_X1 U8975 ( .A(n4317), .ZN(n4642) );
  NAND2_X1 U8976 ( .A1(n5368), .A2(n5322), .ZN(n4019) );
  INV_X1 U8977 ( .A(n4296), .ZN(n4927) );
  INV_X1 U8978 ( .A(n4928), .ZN(n4298) );
  OAI211_X1 U8979 ( .C1(n4927), .C2(n4297), .A(n4020), .B(n4298), .ZN(n4024)
         );
  NAND3_X1 U8980 ( .A1(n4975), .A2(n4928), .A3(n4131), .ZN(n4023) );
  NAND3_X1 U8981 ( .A1(n4932), .A2(n4296), .A3(n4976), .ZN(n4022) );
  NAND3_X1 U8982 ( .A1(n4282), .A2(n5323), .A3(n5398), .ZN(n4025) );
  XNOR2_X1 U8983 ( .A(n7264), .B(n6745), .ZN(n4063) );
  NAND2_X1 U8984 ( .A1(n4796), .A2(n5045), .ZN(n4027) );
  NAND2_X1 U8986 ( .A1(n5042), .A2(n5046), .ZN(n4026) );
  XNOR2_X1 U8987 ( .A(Key[115]), .B(Plaintext[115]), .ZN(n4440) );
  INV_X1 U8988 ( .A(n4439), .ZN(n5048) );
  INV_X1 U8989 ( .A(Plaintext[114]), .ZN(n4028) );
  XNOR2_X1 U8990 ( .A(Key[119]), .B(Plaintext[119]), .ZN(n4088) );
  INV_X1 U8991 ( .A(n4088), .ZN(n4698) );
  INV_X1 U8992 ( .A(n6044), .ZN(n5144) );
  NAND2_X1 U8994 ( .A1(n5087), .A2(n5086), .ZN(n4032) );
  INV_X1 U8996 ( .A(n5086), .ZN(n4802) );
  INV_X1 U8997 ( .A(Plaintext[113]), .ZN(n4030) );
  INV_X1 U8999 ( .A(n4701), .ZN(n4807) );
  OAI21_X1 U9000 ( .B1(n4032), .B2(n5083), .A(n4031), .ZN(n4034) );
  AOI21_X1 U9001 ( .B1(n4032), .B2(n5090), .A(n4807), .ZN(n4033) );
  INV_X1 U9002 ( .A(Plaintext[132]), .ZN(n4035) );
  XNOR2_X1 U9003 ( .A(Key[137]), .B(Plaintext[137]), .ZN(n4268) );
  INV_X1 U9004 ( .A(n4268), .ZN(n5026) );
  INV_X1 U9005 ( .A(Plaintext[134]), .ZN(n4036) );
  XNOR2_X1 U9006 ( .A(n4036), .B(Key[134]), .ZN(n4094) );
  INV_X1 U9007 ( .A(n4094), .ZN(n4761) );
  NAND2_X1 U9008 ( .A1(n4765), .A2(n4269), .ZN(n4037) );
  AOI21_X1 U9009 ( .B1(n4037), .B2(n4095), .A(n4761), .ZN(n4038) );
  INV_X1 U9010 ( .A(Plaintext[125]), .ZN(n4039) );
  XNOR2_X1 U9011 ( .A(n4039), .B(Key[125]), .ZN(n4041) );
  INV_X1 U9012 ( .A(n4041), .ZN(n5035) );
  INV_X1 U9013 ( .A(Plaintext[120]), .ZN(n4040) );
  XNOR2_X1 U9014 ( .A(Key[123]), .B(Plaintext[123]), .ZN(n4107) );
  INV_X1 U9015 ( .A(n5031), .ZN(n4707) );
  NAND2_X1 U9016 ( .A1(n4709), .A2(n4707), .ZN(n4042) );
  AND2_X1 U9017 ( .A1(n4107), .A2(n4769), .ZN(n5037) );
  INV_X1 U9018 ( .A(n4769), .ZN(n4452) );
  XNOR2_X1 U9019 ( .A(Key[105]), .B(Plaintext[105]), .ZN(n4048) );
  INV_X1 U9020 ( .A(Plaintext[104]), .ZN(n4044) );
  XNOR2_X1 U9021 ( .A(n4044), .B(Key[104]), .ZN(n5106) );
  INV_X1 U9022 ( .A(Plaintext[106]), .ZN(n4045) );
  INV_X1 U9024 ( .A(n5101), .ZN(n4077) );
  MUX2_X1 U9025 ( .A(n5105), .B(n5102), .S(n4077), .Z(n4051) );
  INV_X1 U9026 ( .A(Plaintext[107]), .ZN(n4046) );
  XNOR2_X2 U9027 ( .A(n4046), .B(Key[107]), .ZN(n5107) );
  XNOR2_X1 U9028 ( .A(Key[103]), .B(Plaintext[103]), .ZN(n5100) );
  INV_X1 U9029 ( .A(n5100), .ZN(n4793) );
  INV_X1 U9030 ( .A(Plaintext[102]), .ZN(n4047) );
  XNOR2_X1 U9031 ( .A(n4047), .B(Key[102]), .ZN(n5108) );
  INV_X1 U9032 ( .A(n5108), .ZN(n5099) );
  INV_X1 U9033 ( .A(n4048), .ZN(n4693) );
  MUX2_X1 U9034 ( .A(n4049), .B(n5099), .S(n4693), .Z(n4050) );
  INV_X1 U9035 ( .A(Plaintext[129]), .ZN(n4053) );
  XNOR2_X1 U9036 ( .A(Key[131]), .B(Plaintext[131]), .ZN(n4056) );
  INV_X1 U9037 ( .A(n4056), .ZN(n5055) );
  XNOR2_X1 U9038 ( .A(Key[126]), .B(Plaintext[126]), .ZN(n4058) );
  INV_X1 U9039 ( .A(Plaintext[130]), .ZN(n4054) );
  XNOR2_X1 U9040 ( .A(n4054), .B(Key[130]), .ZN(n4445) );
  INV_X1 U9041 ( .A(Plaintext[128]), .ZN(n4055) );
  XNOR2_X1 U9042 ( .A(n4055), .B(Key[128]), .ZN(n4060) );
  INV_X1 U9043 ( .A(n4060), .ZN(n5059) );
  NAND3_X1 U9044 ( .A1(n4585), .A2(n5059), .A3(n5058), .ZN(n4057) );
  INV_X1 U9045 ( .A(n4058), .ZN(n5056) );
  INV_X1 U9046 ( .A(Plaintext[127]), .ZN(n4059) );
  INV_X1 U9047 ( .A(n5052), .ZN(n4739) );
  NAND2_X1 U9048 ( .A1(n6046), .A2(n5309), .ZN(n4061) );
  NOR2_X1 U9049 ( .A1(n4061), .A2(n6044), .ZN(n4062) );
  XNOR2_X1 U9050 ( .A(n4063), .B(n7345), .ZN(n4064) );
  XNOR2_X1 U9051 ( .A(n4065), .B(n4064), .ZN(n8061) );
  INV_X1 U9052 ( .A(n4418), .ZN(n4066) );
  INV_X1 U9053 ( .A(n5093), .ZN(n4715) );
  INV_X1 U9054 ( .A(n4405), .ZN(n4713) );
  NAND3_X1 U9055 ( .A1(n4788), .A2(n4715), .A3(n2460), .ZN(n4069) );
  OAI21_X1 U9057 ( .B1(n4214), .B2(n4827), .A(n4824), .ZN(n4072) );
  INV_X1 U9058 ( .A(n4824), .ZN(n4426) );
  NAND2_X1 U9059 ( .A1(n4426), .A2(n4829), .ZN(n4071) );
  AND2_X1 U9060 ( .A1(n4072), .A2(n4071), .ZN(n4075) );
  NAND2_X1 U9061 ( .A1(n4426), .A2(n4214), .ZN(n4073) );
  AOI21_X1 U9062 ( .B1(n4425), .B2(n4073), .A(n4668), .ZN(n4074) );
  INV_X1 U9063 ( .A(n5434), .ZN(n5995) );
  AOI21_X1 U9064 ( .B1(n5998), .B2(n5997), .A(n5995), .ZN(n4087) );
  AOI21_X1 U9065 ( .B1(n4076), .B2(n5108), .A(n5102), .ZN(n4079) );
  NAND2_X1 U9066 ( .A1(n4793), .A2(n5108), .ZN(n4449) );
  NAND2_X1 U9067 ( .A1(n5998), .A2(n5434), .ZN(n4080) );
  NAND2_X1 U9069 ( .A1(n4081), .A2(n5075), .ZN(n4082) );
  MUX2_X1 U9070 ( .A(n4083), .B(n4082), .S(n5080), .Z(n4086) );
  NAND2_X1 U9071 ( .A1(n4084), .A2(n4457), .ZN(n4085) );
  INV_X1 U9072 ( .A(n6000), .ZN(n6002) );
  NAND2_X1 U9073 ( .A1(n4088), .A2(n5045), .ZN(n4089) );
  NAND2_X1 U9074 ( .A1(n4698), .A2(n5046), .ZN(n4798) );
  INV_X1 U9075 ( .A(n5990), .ZN(n5708) );
  MUX2_X1 U9076 ( .A(n20202), .B(n5086), .S(n5087), .Z(n4093) );
  NAND2_X1 U9077 ( .A1(n4090), .A2(n19776), .ZN(n4092) );
  NOR2_X1 U9078 ( .A1(n4801), .A2(n5083), .ZN(n4091) );
  AOI21_X1 U9079 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n5711) );
  NAND2_X1 U9080 ( .A1(n4765), .A2(n4095), .ZN(n4098) );
  INV_X1 U9081 ( .A(n4095), .ZN(n4764) );
  NAND3_X1 U9083 ( .A1(n5025), .A2(n4761), .A3(n5024), .ZN(n4097) );
  NAND2_X1 U9084 ( .A1(n20461), .A2(n5059), .ZN(n4099) );
  AOI21_X1 U9085 ( .B1(n5054), .B2(n4099), .A(n5058), .ZN(n4104) );
  INV_X1 U9086 ( .A(n4100), .ZN(n5057) );
  NAND3_X1 U9087 ( .A1(n5057), .A2(n5058), .A3(n873), .ZN(n4101) );
  NAND2_X1 U9088 ( .A1(n4102), .A2(n4101), .ZN(n4103) );
  NAND2_X1 U9089 ( .A1(n4708), .A2(n4107), .ZN(n4105) );
  OAI21_X1 U9090 ( .B1(n4107), .B2(n4769), .A(n4105), .ZN(n4106) );
  NAND2_X1 U9091 ( .A1(n4106), .A2(n5032), .ZN(n4109) );
  NAND2_X1 U9092 ( .A1(n303), .A2(n153), .ZN(n4108) );
  INV_X1 U9093 ( .A(n5815), .ZN(n5709) );
  OAI21_X1 U9094 ( .B1(n4734), .B2(n4277), .A(n4554), .ZN(n4111) );
  INV_X1 U9095 ( .A(n5276), .ZN(n5986) );
  NAND2_X1 U9096 ( .A1(n5986), .A2(n5989), .ZN(n4112) );
  XNOR2_X1 U9097 ( .A(n6711), .B(n7390), .ZN(n7016) );
  AND2_X1 U9098 ( .A1(n4887), .A2(n4946), .ZN(n4471) );
  NAND2_X1 U9099 ( .A1(n4114), .A2(n4118), .ZN(n4943) );
  INV_X1 U9100 ( .A(n4943), .ZN(n4115) );
  AOI22_X1 U9101 ( .A1(n4467), .A2(n4471), .B1(n4115), .B2(n4947), .ZN(n4121)
         );
  OAI21_X1 U9102 ( .B1(n4467), .B2(n4117), .A(n4116), .ZN(n4119) );
  INV_X1 U9104 ( .A(n4886), .ZN(n4888) );
  NAND2_X1 U9105 ( .A1(n4119), .A2(n4888), .ZN(n4120) );
  NAND2_X1 U9106 ( .A1(n4003), .A2(n19822), .ZN(n4122) );
  NAND2_X1 U9107 ( .A1(n4620), .A2(n4122), .ZN(n4123) );
  NAND2_X1 U9108 ( .A1(n4125), .A2(n4640), .ZN(n4126) );
  NAND2_X1 U9109 ( .A1(n4647), .A2(n4125), .ZN(n4128) );
  MUX2_X1 U9110 ( .A(n4128), .B(n4318), .S(n4127), .Z(n4129) );
  OAI21_X1 U9111 ( .B1(n4130), .B2(n4642), .A(n4129), .ZN(n5968) );
  INV_X1 U9112 ( .A(n5968), .ZN(n5525) );
  NAND2_X1 U9114 ( .A1(n4298), .A2(n4975), .ZN(n4133) );
  NAND2_X1 U9115 ( .A1(n4296), .A2(n4297), .ZN(n4132) );
  MUX2_X1 U9116 ( .A(n4133), .B(n4132), .S(n4976), .Z(n4134) );
  OAI21_X2 U9117 ( .B1(n4135), .B2(n4297), .A(n4134), .ZN(n5697) );
  INV_X1 U9118 ( .A(n5697), .ZN(n5294) );
  NAND2_X1 U9120 ( .A1(n4899), .A2(n4892), .ZN(n4137) );
  INV_X1 U9121 ( .A(n4912), .ZN(n4914) );
  NAND2_X1 U9124 ( .A1(n4474), .A2(n4911), .ZN(n4141) );
  NAND2_X1 U9126 ( .A1(n4952), .A2(n4954), .ZN(n4142) );
  INV_X1 U9127 ( .A(n4953), .ZN(n4950) );
  OR2_X1 U9128 ( .A1(n4144), .A2(n4954), .ZN(n5522) );
  AOI21_X1 U9129 ( .B1(n4146), .B2(n4646), .A(n4640), .ZN(n4150) );
  NAND3_X1 U9131 ( .A1(n4641), .A2(n4325), .A3(n4640), .ZN(n4147) );
  NAND2_X1 U9133 ( .A1(n4354), .A2(n4547), .ZN(n4151) );
  NAND2_X1 U9135 ( .A1(n19524), .A2(n4532), .ZN(n4158) );
  NAND2_X1 U9136 ( .A1(n4186), .A2(n4637), .ZN(n4157) );
  NAND2_X1 U9137 ( .A1(n4516), .A2(n4342), .ZN(n4527) );
  AOI21_X1 U9138 ( .B1(n4527), .B2(n4522), .A(n4523), .ZN(n4164) );
  NAND3_X1 U9139 ( .A1(n4343), .A2(n4516), .A3(n4160), .ZN(n4162) );
  NAND2_X1 U9140 ( .A1(n4162), .A2(n4161), .ZN(n4163) );
  OAI21_X1 U9142 ( .B1(n5645), .B2(n5443), .A(n4165), .ZN(n4777) );
  INV_X1 U9143 ( .A(n4623), .ZN(n4166) );
  AOI21_X1 U9144 ( .B1(n4166), .B2(n4169), .A(n20143), .ZN(n4175) );
  NAND2_X1 U9145 ( .A1(n4288), .A2(n4167), .ZN(n4174) );
  INV_X1 U9146 ( .A(n4291), .ZN(n4168) );
  OAI21_X1 U9147 ( .B1(n4170), .B2(n4169), .A(n4168), .ZN(n4172) );
  NAND3_X1 U9148 ( .A1(n4613), .A2(n4364), .A3(n748), .ZN(n4178) );
  NAND2_X1 U9149 ( .A1(n4179), .A2(n5442), .ZN(n4180) );
  AOI22_X1 U9150 ( .A1(n4777), .A2(n5649), .B1(n4180), .B2(n5443), .ZN(n6352)
         );
  INV_X1 U9151 ( .A(n6352), .ZN(n7298) );
  XNOR2_X1 U9152 ( .A(n7298), .B(n7196), .ZN(n6858) );
  XNOR2_X1 U9153 ( .A(n7016), .B(n6858), .ZN(n4247) );
  NAND2_X1 U9154 ( .A1(n5798), .A2(n5428), .ZN(n5301) );
  INV_X1 U9155 ( .A(n5795), .ZN(n5791) );
  AOI21_X1 U9156 ( .B1(n4182), .B2(n4181), .A(n5300), .ZN(n4183) );
  INV_X1 U9157 ( .A(n4187), .ZN(n4339) );
  NAND2_X1 U9158 ( .A1(n4516), .A2(n4339), .ZN(n4191) );
  NAND2_X1 U9159 ( .A1(n4517), .A2(n4187), .ZN(n4188) );
  OAI211_X1 U9160 ( .C1(n4523), .C2(n4522), .A(n4188), .B(n4343), .ZN(n4190)
         );
  NAND2_X1 U9161 ( .A1(n4575), .A2(n4576), .ZN(n4257) );
  NAND2_X1 U9162 ( .A1(n4570), .A2(n4574), .ZN(n4192) );
  AND2_X1 U9163 ( .A1(n4257), .A2(n4192), .ZN(n4195) );
  NAND2_X1 U9164 ( .A1(n20190), .A2(n4575), .ZN(n4193) );
  OAI21_X1 U9165 ( .B1(n4372), .B2(n4507), .A(n4193), .ZN(n4194) );
  INV_X1 U9166 ( .A(n5424), .ZN(n5675) );
  NAND2_X1 U9167 ( .A1(n4567), .A2(n4756), .ZN(n4196) );
  NAND2_X1 U9168 ( .A1(n4196), .A2(n4504), .ZN(n4197) );
  NAND2_X1 U9169 ( .A1(n4198), .A2(n4752), .ZN(n4758) );
  NAND2_X1 U9170 ( .A1(n4347), .A2(n4199), .ZN(n4201) );
  MUX2_X1 U9171 ( .A(n4201), .B(n4200), .S(n4541), .Z(n4202) );
  NAND3_X1 U9172 ( .A1(n5424), .A2(n5669), .A3(n5670), .ZN(n4211) );
  INV_X1 U9173 ( .A(n4204), .ZN(n5003) );
  NAND2_X1 U9174 ( .A1(n4744), .A2(n4745), .ZN(n4207) );
  NAND2_X1 U9175 ( .A1(n4207), .A2(n4248), .ZN(n4208) );
  NAND2_X1 U9176 ( .A1(n5424), .A2(n5279), .ZN(n4210) );
  XNOR2_X1 U9177 ( .A(n6708), .B(n6489), .ZN(n4245) );
  NAND2_X1 U9178 ( .A1(n4213), .A2(n4214), .ZN(n4219) );
  AND2_X1 U9179 ( .A1(n4214), .A2(n4669), .ZN(n4823) );
  NAND2_X1 U9180 ( .A1(n4823), .A2(n19688), .ZN(n4218) );
  INV_X1 U9181 ( .A(n4829), .ZN(n4215) );
  OAI21_X1 U9182 ( .B1(n4824), .B2(n4827), .A(n4215), .ZN(n4216) );
  NAND2_X1 U9183 ( .A1(n4216), .A2(n4828), .ZN(n4217) );
  INV_X1 U9184 ( .A(n4220), .ZN(n4841) );
  NAND3_X1 U9185 ( .A1(n4659), .A2(n2601), .A3(n4221), .ZN(n4222) );
  AND2_X1 U9186 ( .A1(n6016), .A2(n6022), .ZN(n5124) );
  INV_X1 U9187 ( .A(n4685), .ZN(n4484) );
  OAI211_X1 U9188 ( .C1(n4484), .C2(n177), .A(n4224), .B(n4853), .ZN(n4225) );
  INV_X1 U9189 ( .A(n5825), .ZN(n5824) );
  NAND2_X1 U9190 ( .A1(n5124), .A2(n5824), .ZN(n4243) );
  NAND2_X1 U9191 ( .A1(n4381), .A2(n4651), .ZN(n4228) );
  INV_X1 U9192 ( .A(n4228), .ZN(n4231) );
  OAI21_X1 U9193 ( .B1(n4652), .B2(n4865), .A(n20356), .ZN(n4230) );
  MUX2_X1 U9194 ( .A(n4228), .B(n4227), .S(n896), .Z(n4229) );
  INV_X1 U9195 ( .A(n4232), .ZN(n4492) );
  INV_X1 U9196 ( .A(n4497), .ZN(n4901) );
  OAI21_X1 U9197 ( .B1(n4492), .B2(n4901), .A(n4378), .ZN(n4905) );
  NAND2_X1 U9198 ( .A1(n4493), .A2(n4499), .ZN(n4236) );
  NAND2_X1 U9199 ( .A1(n4492), .A2(n4856), .ZN(n4857) );
  INV_X1 U9200 ( .A(n4857), .ZN(n4235) );
  NAND2_X1 U9201 ( .A1(n4855), .A2(n4860), .ZN(n4234) );
  NAND3_X1 U9202 ( .A1(n5823), .A2(n5825), .A3(n3569), .ZN(n4242) );
  INV_X1 U9203 ( .A(n4965), .ZN(n4383) );
  INV_X1 U9204 ( .A(n4482), .ZN(n4919) );
  INV_X1 U9205 ( .A(n4969), .ZN(n4921) );
  OAI211_X1 U9206 ( .C1(n4965), .C2(n4479), .A(n4921), .B(n19507), .ZN(n4238)
         );
  OAI21_X1 U9207 ( .B1(n4383), .B2(n4968), .A(n4969), .ZN(n4237) );
  INV_X1 U9208 ( .A(n6017), .ZN(n5827) );
  NAND2_X1 U9209 ( .A1(n5827), .A2(n5825), .ZN(n4241) );
  NAND3_X1 U9210 ( .A1(n3569), .A2(n6017), .A3(n6022), .ZN(n4240) );
  NAND4_X2 U9211 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n7013)
         );
  XNOR2_X1 U9212 ( .A(n7013), .B(n20682), .ZN(n4244) );
  XNOR2_X1 U9213 ( .A(n4245), .B(n4244), .ZN(n4246) );
  INV_X1 U9214 ( .A(n4750), .ZN(n5007) );
  NAND2_X1 U9215 ( .A1(n4248), .A2(n5007), .ZN(n4253) );
  INV_X1 U9216 ( .A(n4744), .ZN(n5006) );
  NAND3_X1 U9217 ( .A1(n4559), .A2(n5006), .A3(n4746), .ZN(n4251) );
  INV_X1 U9218 ( .A(n4350), .ZN(n4537) );
  INV_X1 U9220 ( .A(n4539), .ZN(n4255) );
  OAI21_X1 U9221 ( .B1(n4370), .B2(n4372), .A(n20190), .ZN(n4263) );
  INV_X1 U9222 ( .A(n4257), .ZN(n4262) );
  OAI21_X1 U9223 ( .B1(n4370), .B2(n4574), .A(n4576), .ZN(n4260) );
  NAND2_X1 U9226 ( .A1(n4260), .A2(n4259), .ZN(n4261) );
  OAI21_X1 U9227 ( .B1(n4263), .B2(n4262), .A(n4261), .ZN(n6131) );
  NAND2_X1 U9228 ( .A1(n4563), .A2(n4752), .ZN(n4264) );
  MUX2_X1 U9229 ( .A(n4758), .B(n4264), .S(n4565), .Z(n4267) );
  INV_X1 U9230 ( .A(n4756), .ZN(n4566) );
  INV_X1 U9231 ( .A(n4752), .ZN(n4564) );
  NAND2_X1 U9232 ( .A1(n4566), .A2(n4564), .ZN(n4265) );
  NOR2_X1 U9233 ( .A1(n6129), .A2(n5691), .ZN(n4274) );
  NOR2_X1 U9234 ( .A1(n5025), .A2(n5022), .ZN(n4270) );
  NAND2_X1 U9235 ( .A1(n4094), .A2(n4271), .ZN(n4763) );
  NOR2_X1 U9236 ( .A1(n4763), .A2(n5024), .ZN(n4272) );
  AOI22_X2 U9237 ( .A1(n4275), .A2(n6131), .B1(n4274), .B2(n5621), .ZN(n6496)
         );
  INV_X1 U9238 ( .A(n4276), .ZN(n4279) );
  INV_X1 U9240 ( .A(n5691), .ZN(n6132) );
  AOI21_X1 U9241 ( .B1(n5623), .B2(n6132), .A(n6133), .ZN(n4280) );
  NAND2_X1 U9242 ( .A1(n4280), .A2(n5694), .ZN(n6500) );
  NAND2_X1 U9243 ( .A1(n6496), .A2(n6500), .ZN(n6362) );
  INV_X1 U9244 ( .A(n5322), .ZN(n5394) );
  NAND2_X1 U9245 ( .A1(n5250), .A2(n5322), .ZN(n4281) );
  NAND3_X1 U9246 ( .A1(n5395), .A2(n5368), .A3(n5323), .ZN(n4283) );
  OAI211_X2 U9247 ( .C1(n5251), .C2(n5373), .A(n4284), .B(n4283), .ZN(n7211)
         );
  XNOR2_X1 U9248 ( .A(n6362), .B(n7211), .ZN(n4336) );
  NAND3_X1 U9249 ( .A1(n20143), .A2(n4171), .A3(n4285), .ZN(n4287) );
  NAND2_X1 U9250 ( .A1(n4290), .A2(n4626), .ZN(n4286) );
  NAND2_X1 U9252 ( .A1(n4291), .A2(n4290), .ZN(n4292) );
  INV_X1 U9253 ( .A(n4979), .ZN(n4293) );
  NAND2_X1 U9254 ( .A1(n4293), .A2(n4296), .ZN(n4294) );
  NAND2_X1 U9255 ( .A1(n4294), .A2(n4978), .ZN(n4295) );
  NAND2_X1 U9256 ( .A1(n4295), .A2(n4975), .ZN(n4301) );
  OAI21_X1 U9257 ( .B1(n4297), .B2(n4979), .A(n4296), .ZN(n4299) );
  NAND2_X1 U9258 ( .A1(n4299), .A2(n4298), .ZN(n4300) );
  AND2_X1 U9259 ( .A1(n5628), .A2(n5363), .ZN(n5360) );
  NAND2_X1 U9260 ( .A1(n4983), .A2(n19822), .ZN(n4304) );
  NAND2_X1 U9261 ( .A1(n4003), .A2(n4618), .ZN(n4303) );
  OAI21_X1 U9263 ( .B1(n4983), .B2(n4982), .A(n4003), .ZN(n4308) );
  AND2_X1 U9264 ( .A1(n4306), .A2(n4305), .ZN(n4987) );
  INV_X1 U9265 ( .A(n4987), .ZN(n4307) );
  INV_X1 U9266 ( .A(n4601), .ZN(n4358) );
  AOI21_X1 U9267 ( .B1(n4312), .B2(n4311), .A(n4361), .ZN(n4316) );
  NAND2_X1 U9268 ( .A1(n4152), .A2(n4548), .ZN(n4362) );
  OAI21_X1 U9270 ( .B1(n4640), .B2(n4125), .A(n4317), .ZN(n4322) );
  NAND2_X1 U9271 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  NAND2_X1 U9272 ( .A1(n4320), .A2(n4642), .ZN(n4321) );
  NAND2_X1 U9273 ( .A1(n4322), .A2(n4321), .ZN(n4327) );
  OAI211_X1 U9274 ( .C1(n4325), .C2(n4324), .A(n4323), .B(n4640), .ZN(n4326)
         );
  AND2_X2 U9275 ( .A1(n4327), .A2(n4326), .ZN(n5364) );
  INV_X1 U9276 ( .A(n5364), .ZN(n5630) );
  NOR2_X1 U9277 ( .A1(n5633), .A2(n5630), .ZN(n4328) );
  INV_X1 U9278 ( .A(n5363), .ZN(n5463) );
  AOI22_X1 U9279 ( .A1(n5360), .A2(n4598), .B1(n4328), .B2(n5463), .ZN(n4334)
         );
  AND2_X1 U9280 ( .A1(n4013), .A2(n3717), .ZN(n4331) );
  NAND2_X1 U9281 ( .A1(n4611), .A2(n4614), .ZN(n4367) );
  MUX2_X1 U9282 ( .A(n4367), .B(n4365), .S(n4615), .Z(n4329) );
  NAND2_X1 U9283 ( .A1(n5631), .A2(n5363), .ZN(n4332) );
  OAI21_X1 U9284 ( .B1(n5364), .B2(n5631), .A(n4332), .ZN(n4333) );
  XNOR2_X1 U9285 ( .A(n6165), .B(n2248), .ZN(n4335) );
  XNOR2_X1 U9286 ( .A(n4336), .B(n4335), .ZN(n4466) );
  NAND2_X1 U9287 ( .A1(n3551), .A2(n20487), .ZN(n4338) );
  NAND2_X1 U9288 ( .A1(n4518), .A2(n4339), .ZN(n4341) );
  AOI21_X1 U9289 ( .B1(n4341), .B2(n4340), .A(n4524), .ZN(n4346) );
  NAND2_X1 U9290 ( .A1(n4343), .A2(n4342), .ZN(n4345) );
  NAND2_X1 U9291 ( .A1(n5605), .A2(n5719), .ZN(n5242) );
  NAND3_X1 U9295 ( .A1(n4603), .A2(n4355), .A3(n4353), .ZN(n4357) );
  NAND3_X1 U9296 ( .A1(n4355), .A2(n4548), .A3(n4354), .ZN(n4356) );
  AND2_X1 U9297 ( .A1(n4357), .A2(n4356), .ZN(n4360) );
  OR2_X1 U9298 ( .A1(n4367), .A2(n4013), .ZN(n4369) );
  INV_X1 U9299 ( .A(n4507), .ZN(n4577) );
  NAND2_X1 U9300 ( .A1(n4371), .A2(n4370), .ZN(n4572) );
  AOI21_X1 U9301 ( .B1(n4572), .B2(n4573), .A(n4372), .ZN(n4373) );
  INV_X1 U9302 ( .A(n5715), .ZN(n5346) );
  INV_X1 U9303 ( .A(n4962), .ZN(n4893) );
  INV_X1 U9304 ( .A(n4855), .ZN(n4904) );
  AOI21_X1 U9305 ( .B1(n4493), .B2(n4904), .A(n4860), .ZN(n4380) );
  OAI21_X1 U9306 ( .B1(n4493), .B2(n4902), .A(n4378), .ZN(n4379) );
  NOR2_X1 U9307 ( .A1(n5611), .A2(n5349), .ZN(n5856) );
  INV_X1 U9308 ( .A(n4864), .ZN(n4381) );
  NAND2_X1 U9309 ( .A1(n4921), .A2(n4482), .ZN(n4384) );
  NAND2_X1 U9312 ( .A1(n4385), .A2(n4968), .ZN(n4386) );
  INV_X1 U9313 ( .A(n6150), .ZN(n6152) );
  OAI21_X1 U9314 ( .B1(n6151), .B2(n6155), .A(n6152), .ZN(n4404) );
  NAND2_X1 U9315 ( .A1(n6150), .A2(n6155), .ZN(n5855) );
  INV_X1 U9316 ( .A(n4684), .ZN(n4848) );
  OAI21_X1 U9317 ( .B1(n4853), .B2(n4848), .A(n4687), .ZN(n4390) );
  NAND2_X1 U9318 ( .A1(n4685), .A2(n4391), .ZN(n4388) );
  NAND2_X1 U9319 ( .A1(n4388), .A2(n4387), .ZN(n4389) );
  INV_X1 U9321 ( .A(n4391), .ZN(n4486) );
  AND2_X1 U9323 ( .A1(n4475), .A2(n4912), .ZN(n4397) );
  INV_X1 U9324 ( .A(n4474), .ZN(n4395) );
  AND2_X1 U9325 ( .A1(n4395), .A2(n4912), .ZN(n4958) );
  INV_X1 U9326 ( .A(n4958), .ZN(n4396) );
  OAI21_X1 U9327 ( .B1(n4398), .B2(n4397), .A(n4396), .ZN(n4401) );
  NOR2_X1 U9328 ( .A1(n4912), .A2(n4475), .ZN(n4399) );
  INV_X1 U9329 ( .A(n4954), .ZN(n4916) );
  INV_X1 U9330 ( .A(n6153), .ZN(n6149) );
  NAND3_X1 U9331 ( .A1(n6149), .A2(n20405), .A3(n6156), .ZN(n4402) );
  AOI21_X1 U9332 ( .B1(n5096), .B2(n5095), .A(n5092), .ZN(n4408) );
  NAND2_X1 U9333 ( .A1(n5098), .A2(n5092), .ZN(n4786) );
  NAND2_X1 U9334 ( .A1(n5095), .A2(n4405), .ZN(n4406) );
  AOI21_X1 U9335 ( .B1(n4786), .B2(n4406), .A(n4783), .ZN(n4407) );
  OAI21_X1 U9336 ( .B1(n5069), .B2(n5073), .A(n2632), .ZN(n4416) );
  INV_X1 U9337 ( .A(n4409), .ZN(n4415) );
  OAI21_X1 U9338 ( .B1(n5069), .B2(n5071), .A(n4410), .ZN(n4413) );
  NAND2_X1 U9339 ( .A1(n4816), .A2(n291), .ZN(n4412) );
  AND2_X1 U9340 ( .A1(n6123), .A2(n5873), .ZN(n5387) );
  NAND3_X1 U9341 ( .A1(n19508), .A2(n1916), .A3(n169), .ZN(n4419) );
  INV_X1 U9342 ( .A(n4420), .ZN(n4844) );
  AND2_X1 U9343 ( .A1(n4841), .A2(n4844), .ZN(n4424) );
  NAND2_X1 U9344 ( .A1(n4840), .A2(n164), .ZN(n4423) );
  INV_X1 U9345 ( .A(n6119), .ZN(n5869) );
  NAND2_X1 U9346 ( .A1(n4824), .A2(n4669), .ZN(n4826) );
  AND2_X1 U9347 ( .A1(n4425), .A2(n4826), .ZN(n5257) );
  NAND2_X1 U9348 ( .A1(n4824), .A2(n4829), .ZN(n4667) );
  NAND3_X1 U9349 ( .A1(n6124), .A2(n5873), .A3(n6119), .ZN(n4434) );
  INV_X2 U9350 ( .A(n5873), .ZN(n6128) );
  NAND2_X1 U9351 ( .A1(n20459), .A2(n20356), .ZN(n4654) );
  NAND2_X1 U9353 ( .A1(n19523), .A2(n896), .ZN(n4428) );
  AOI21_X1 U9354 ( .B1(n4654), .B2(n4428), .A(n4652), .ZN(n4432) );
  NAND2_X1 U9355 ( .A1(n20357), .A2(n4652), .ZN(n4430) );
  AOI21_X1 U9356 ( .B1(n4430), .B2(n3560), .A(n896), .ZN(n4431) );
  OR2_X1 U9357 ( .A1(n4432), .A2(n4431), .ZN(n6118) );
  AND2_X1 U9358 ( .A1(n4433), .A2(n4434), .ZN(n4435) );
  NAND2_X1 U9359 ( .A1(n4436), .A2(n4435), .ZN(n6738) );
  INV_X1 U9360 ( .A(n5083), .ZN(n4804) );
  NAND3_X1 U9361 ( .A1(n19776), .A2(n20016), .A3(n5087), .ZN(n4437) );
  INV_X1 U9362 ( .A(n4697), .ZN(n5047) );
  NAND3_X1 U9363 ( .A1(n20464), .A2(n5042), .A3(n5047), .ZN(n4443) );
  INV_X1 U9364 ( .A(n6138), .ZN(n5342) );
  NAND2_X1 U9365 ( .A1(n5056), .A2(n20461), .ZN(n4743) );
  INV_X1 U9366 ( .A(n4445), .ZN(n4738) );
  AOI21_X1 U9367 ( .B1(n4743), .B2(n4741), .A(n4738), .ZN(n4448) );
  NAND2_X1 U9368 ( .A1(n4100), .A2(n20461), .ZN(n4446) );
  AOI21_X1 U9369 ( .B1(n4446), .B2(n2929), .A(n5059), .ZN(n4447) );
  INV_X1 U9370 ( .A(n5860), .ZN(n6141) );
  NAND3_X1 U9371 ( .A1(n4450), .A2(n3167), .A3(n5105), .ZN(n4451) );
  MUX2_X1 U9373 ( .A(n303), .B(n4452), .S(n4771), .Z(n4456) );
  NAND2_X1 U9374 ( .A1(n303), .A2(n4708), .ZN(n4454) );
  MUX2_X1 U9375 ( .A(n4454), .B(n4453), .S(n5035), .Z(n4455) );
  OAI21_X1 U9377 ( .B1(n5080), .B2(n5077), .A(n5079), .ZN(n4460) );
  MUX2_X1 U9378 ( .A(n4462), .B(n4461), .S(n6141), .Z(n4463) );
  OAI21_X2 U9379 ( .B1(n4464), .B2(n6143), .A(n4463), .ZN(n7363) );
  XNOR2_X1 U9380 ( .A(n7363), .B(n6738), .ZN(n7036) );
  XNOR2_X1 U9381 ( .A(n6881), .B(n7036), .ZN(n4465) );
  NOR2_X1 U9383 ( .A1(n4941), .A2(n4940), .ZN(n4469) );
  INV_X1 U9384 ( .A(n4946), .ZN(n4468) );
  OAI21_X1 U9385 ( .B1(n4889), .B2(n4469), .A(n4468), .ZN(n4473) );
  OAI21_X1 U9386 ( .B1(n4471), .B2(n4470), .A(n4941), .ZN(n4472) );
  NAND2_X1 U9387 ( .A1(n4474), .A2(n4954), .ZN(n4951) );
  NAND2_X1 U9388 ( .A1(n4954), .A2(n4475), .ZN(n4476) );
  AOI21_X1 U9390 ( .B1(n4854), .B2(n4851), .A(n4848), .ZN(n4489) );
  AOI21_X1 U9391 ( .B1(n4487), .B2(n4486), .A(n4687), .ZN(n4488) );
  MUX2_X1 U9392 ( .A(n4960), .B(n20205), .S(n4894), .Z(n4491) );
  MUX2_X1 U9393 ( .A(n4962), .B(n292), .S(n4892), .Z(n4490) );
  OAI21_X1 U9394 ( .B1(n4499), .B2(n4855), .A(n4907), .ZN(n4496) );
  NAND2_X1 U9395 ( .A1(n4494), .A2(n4493), .ZN(n4495) );
  AOI21_X1 U9396 ( .B1(n6202), .B2(n6206), .A(n6204), .ZN(n4502) );
  MUX2_X1 U9397 ( .A(n4504), .B(n4752), .S(n4756), .Z(n4506) );
  OAI21_X1 U9398 ( .B1(n4566), .B2(n4565), .A(n4504), .ZN(n4503) );
  OAI21_X1 U9399 ( .B1(n4754), .B2(n4504), .A(n4503), .ZN(n4505) );
  OAI21_X1 U9400 ( .B1(n4507), .B2(n4573), .A(n4511), .ZN(n4508) );
  NAND2_X1 U9401 ( .A1(n4574), .A2(n4511), .ZN(n4512) );
  NAND2_X1 U9402 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  NAND3_X1 U9404 ( .A1(n4524), .A2(n4523), .A3(n4522), .ZN(n4525) );
  MUX2_X1 U9405 ( .A(n5545), .B(n5734), .S(n5765), .Z(n4552) );
  INV_X1 U9406 ( .A(n4528), .ZN(n4529) );
  OAI21_X1 U9408 ( .B1(n4529), .B2(n4532), .A(n20369), .ZN(n4533) );
  NAND2_X1 U9409 ( .A1(n4636), .A2(n4533), .ZN(n4534) );
  OAI21_X1 U9410 ( .B1(n4636), .B2(n3753), .A(n4534), .ZN(n5539) );
  NAND2_X1 U9411 ( .A1(n4535), .A2(n4185), .ZN(n5540) );
  NAND2_X1 U9412 ( .A1(n5539), .A2(n5540), .ZN(n5763) );
  OAI22_X1 U9413 ( .A1(n4538), .A2(n4537), .B1(n4536), .B2(n4540), .ZN(n5537)
         );
  INV_X1 U9414 ( .A(n5765), .ZN(n5546) );
  NAND2_X1 U9415 ( .A1(n4313), .A2(n4548), .ZN(n4608) );
  NAND2_X1 U9416 ( .A1(n4546), .A2(n4313), .ZN(n4549) );
  AOI21_X1 U9417 ( .B1(n4549), .B2(n4548), .A(n4547), .ZN(n4550) );
  INV_X1 U9418 ( .A(n5768), .ZN(n5735) );
  MUX2_X2 U9419 ( .A(n4552), .B(n4551), .S(n5735), .Z(n7288) );
  NAND2_X1 U9420 ( .A1(n4734), .A2(n20229), .ZN(n4553) );
  INV_X1 U9421 ( .A(n4555), .ZN(n5016) );
  OAI211_X1 U9422 ( .C1(n5018), .C2(n20229), .A(n4553), .B(n5016), .ZN(n4556)
         );
  NAND2_X1 U9423 ( .A1(n4557), .A2(n4744), .ZN(n4562) );
  MUX2_X1 U9424 ( .A(n4559), .B(n4558), .S(n4746), .Z(n4560) );
  OAI21_X2 U9425 ( .B1(n4562), .B2(n4561), .A(n4560), .ZN(n5805) );
  NAND2_X1 U9426 ( .A1(n5378), .A2(n5805), .ZN(n6191) );
  OAI21_X1 U9427 ( .B1(n4754), .B2(n4565), .A(n4564), .ZN(n4569) );
  NAND2_X1 U9428 ( .A1(n4566), .A2(n4752), .ZN(n4568) );
  NAND2_X1 U9429 ( .A1(n5803), .A2(n5802), .ZN(n6195) );
  MUX2_X1 U9430 ( .A(n4572), .B(n20190), .S(n4570), .Z(n4580) );
  OAI22_X1 U9431 ( .A1(n4576), .A2(n4575), .B1(n4574), .B2(n4573), .ZN(n4578)
         );
  NAND2_X1 U9432 ( .A1(n4578), .A2(n4577), .ZN(n4579) );
  NAND3_X1 U9433 ( .A1(n6191), .A2(n6195), .A3(n5382), .ZN(n4596) );
  AND2_X1 U9434 ( .A1(n5805), .A2(n6189), .ZN(n5379) );
  INV_X1 U9435 ( .A(n5379), .ZN(n4594) );
  INV_X1 U9436 ( .A(n5805), .ZN(n6193) );
  NAND3_X1 U9437 ( .A1(n5060), .A2(n5055), .A3(n4585), .ZN(n4587) );
  NAND2_X1 U9438 ( .A1(n5057), .A2(n4738), .ZN(n4586) );
  AOI22_X1 U9439 ( .A1(n4587), .A2(n4586), .B1(n4739), .B2(n4738), .ZN(n4592)
         );
  NAND3_X1 U9440 ( .A1(n4588), .A2(n5055), .A3(n4738), .ZN(n4589) );
  NAND2_X1 U9441 ( .A1(n4590), .A2(n4589), .ZN(n4591) );
  NOR2_X2 U9442 ( .A1(n4592), .A2(n4591), .ZN(n6192) );
  INV_X1 U9443 ( .A(n6192), .ZN(n5804) );
  XNOR2_X1 U9445 ( .A(n6477), .B(n19180), .ZN(n4597) );
  XNOR2_X1 U9446 ( .A(n6864), .B(n4597), .ZN(n4729) );
  MUX2_X1 U9447 ( .A(n5631), .B(n5633), .S(n5364), .Z(n4599) );
  MUX2_X1 U9448 ( .A(n4599), .B(n5465), .S(n5463), .Z(n4600) );
  NAND2_X1 U9449 ( .A1(n4602), .A2(n4601), .ZN(n4604) );
  INV_X1 U9450 ( .A(n4982), .ZN(n4617) );
  OAI21_X1 U9451 ( .B1(n4988), .B2(n4618), .A(n4617), .ZN(n4619) );
  AOI22_X1 U9452 ( .A1(n4620), .A2(n4989), .B1(n4003), .B2(n4619), .ZN(n4882)
         );
  NAND2_X1 U9453 ( .A1(n4631), .A2(n4626), .ZN(n4625) );
  MUX2_X1 U9454 ( .A(n4625), .B(n4624), .S(n4623), .Z(n4629) );
  OAI211_X1 U9455 ( .C1(n4631), .C2(n4630), .A(n4629), .B(n4628), .ZN(n5744)
         );
  INV_X1 U9456 ( .A(n5744), .ZN(n4632) );
  NAND2_X1 U9457 ( .A1(n3551), .A2(n19524), .ZN(n4635) );
  NAND2_X1 U9458 ( .A1(n4633), .A2(n4185), .ZN(n4634) );
  NAND2_X1 U9459 ( .A1(n4185), .A2(n19524), .ZN(n4639) );
  NAND2_X1 U9460 ( .A1(n4127), .A2(n4646), .ZN(n4644) );
  NAND2_X1 U9461 ( .A1(n4641), .A2(n4640), .ZN(n4643) );
  NOR2_X1 U9462 ( .A1(n5201), .A2(n5747), .ZN(n5496) );
  INV_X1 U9463 ( .A(n6719), .ZN(n4650) );
  XNOR2_X1 U9464 ( .A(n4650), .B(n20203), .ZN(n4727) );
  AND2_X1 U9465 ( .A1(n4651), .A2(n896), .ZN(n4653) );
  NAND2_X1 U9466 ( .A1(n4659), .A2(n4658), .ZN(n4660) );
  AOI21_X1 U9467 ( .B1(n4662), .B2(n2632), .A(n4410), .ZN(n4666) );
  NAND2_X1 U9468 ( .A1(n4664), .A2(n4663), .ZN(n5070) );
  INV_X1 U9469 ( .A(n6171), .ZN(n4691) );
  MUX2_X1 U9470 ( .A(n4675), .B(n4835), .S(n19508), .Z(n4680) );
  NAND2_X1 U9471 ( .A1(n5115), .A2(n4675), .ZN(n4678) );
  NAND2_X1 U9472 ( .A1(n2042), .A2(n169), .ZN(n4677) );
  MUX2_X1 U9473 ( .A(n4678), .B(n4677), .S(n4676), .Z(n4679) );
  NAND2_X1 U9474 ( .A1(n1867), .A2(n6166), .ZN(n4689) );
  OAI21_X1 U9475 ( .B1(n4682), .B2(n4684), .A(n4681), .ZN(n4683) );
  NAND2_X1 U9476 ( .A1(n4683), .A2(n4391), .ZN(n5219) );
  NAND2_X1 U9477 ( .A1(n4684), .A2(n177), .ZN(n5217) );
  AND2_X1 U9478 ( .A1(n178), .A2(n4685), .ZN(n4850) );
  OAI21_X1 U9479 ( .B1(n3996), .B2(n4687), .A(n4850), .ZN(n5218) );
  OAI21_X2 U9480 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(n7216) );
  MUX2_X1 U9481 ( .A(n5101), .B(n4693), .S(n5102), .Z(n4695) );
  NAND2_X1 U9482 ( .A1(n4693), .A2(n5100), .ZN(n4790) );
  AND2_X1 U9483 ( .A1(n4790), .A2(n4792), .ZN(n4694) );
  NOR2_X1 U9484 ( .A1(n6183), .A2(n5847), .ZN(n6182) );
  AND2_X1 U9485 ( .A1(n4699), .A2(n4700), .ZN(n4704) );
  NAND2_X1 U9486 ( .A1(n4804), .A2(n19777), .ZN(n5091) );
  NAND2_X1 U9487 ( .A1(n4801), .A2(n5086), .ZN(n4702) );
  MUX2_X1 U9488 ( .A(n5091), .B(n4702), .S(n5088), .Z(n4703) );
  NOR2_X1 U9489 ( .A1(n5846), .A2(n5730), .ZN(n4705) );
  NOR2_X1 U9490 ( .A1(n6182), .A2(n4705), .ZN(n6382) );
  INV_X1 U9491 ( .A(n6382), .ZN(n4725) );
  AOI22_X1 U9492 ( .A1(n303), .A2(n4707), .B1(n4706), .B2(n4708), .ZN(n4711)
         );
  MUX2_X1 U9493 ( .A(n4709), .B(n4708), .S(n4707), .Z(n4710) );
  OAI211_X1 U9494 ( .C1(n5093), .C2(n4713), .A(n4712), .B(n4783), .ZN(n4718)
         );
  NAND2_X1 U9495 ( .A1(n4714), .A2(n5094), .ZN(n4717) );
  NOR2_X1 U9496 ( .A1(n4788), .A2(n4715), .ZN(n4716) );
  AND2_X1 U9498 ( .A1(n5080), .A2(n5077), .ZN(n4722) );
  NAND2_X1 U9499 ( .A1(n5081), .A2(n4719), .ZN(n5076) );
  NAND2_X1 U9500 ( .A1(n4720), .A2(n5078), .ZN(n4721) );
  INV_X1 U9501 ( .A(n5383), .ZN(n4723) );
  OAI211_X1 U9502 ( .C1(n19476), .C2(n6379), .A(n4723), .B(n6184), .ZN(n4724)
         );
  OAI21_X1 U9503 ( .B1(n4725), .B2(n6184), .A(n4724), .ZN(n4726) );
  XNOR2_X1 U9504 ( .A(n7216), .B(n4726), .ZN(n6562) );
  XNOR2_X1 U9505 ( .A(n4727), .B(n6562), .ZN(n4728) );
  MUX2_X1 U9507 ( .A(n7461), .B(n4730), .S(n8190), .Z(n5137) );
  OAI21_X1 U9508 ( .B1(n5012), .B2(n5014), .A(n4731), .ZN(n4733) );
  NAND2_X1 U9509 ( .A1(n5058), .A2(n4738), .ZN(n4740) );
  NAND3_X1 U9510 ( .A1(n4740), .A2(n4739), .A3(n5057), .ZN(n4742) );
  INV_X1 U9511 ( .A(n6104), .ZN(n5659) );
  INV_X1 U9512 ( .A(n4745), .ZN(n5004) );
  NAND2_X1 U9513 ( .A1(n4750), .A2(n5010), .ZN(n4747) );
  MUX2_X1 U9514 ( .A(n4748), .B(n4747), .S(n5006), .Z(n4749) );
  AOI21_X1 U9515 ( .B1(n4753), .B2(n4754), .A(n4752), .ZN(n4760) );
  NAND2_X1 U9516 ( .A1(n4755), .A2(n4754), .ZN(n4757) );
  AOI21_X1 U9517 ( .B1(n4758), .B2(n4757), .A(n4756), .ZN(n4759) );
  NOR2_X1 U9518 ( .A1(n5172), .A2(n6109), .ZN(n4776) );
  NAND2_X1 U9519 ( .A1(n4761), .A2(n19788), .ZN(n4762) );
  NAND2_X1 U9520 ( .A1(n4763), .A2(n4762), .ZN(n4768) );
  NAND2_X1 U9521 ( .A1(n4765), .A2(n5022), .ZN(n4766) );
  NAND2_X1 U9522 ( .A1(n5027), .A2(n4766), .ZN(n4767) );
  MUX2_X2 U9523 ( .A(n4768), .B(n4767), .S(n5026), .Z(n6105) );
  OAI22_X1 U9524 ( .A1(n153), .A2(n5035), .B1(n303), .B2(n4769), .ZN(n4770) );
  NAND3_X1 U9525 ( .A1(n5038), .A2(n303), .A3(n4772), .ZN(n4773) );
  INV_X1 U9526 ( .A(n6107), .ZN(n5656) );
  NAND3_X1 U9527 ( .A1(n5657), .A2(n6104), .A3(n5656), .ZN(n4775) );
  XNOR2_X1 U9528 ( .A(n7384), .B(n2122), .ZN(n4781) );
  NOR2_X1 U9529 ( .A1(n5649), .A2(n5643), .ZN(n4779) );
  NAND2_X1 U9531 ( .A1(n4777), .A2(n5648), .ZN(n4778) );
  INV_X1 U9532 ( .A(n7336), .ZN(n4780) );
  INV_X1 U9533 ( .A(n4782), .ZN(n4785) );
  NAND2_X1 U9534 ( .A1(n2460), .A2(n4783), .ZN(n4784) );
  NAND2_X1 U9535 ( .A1(n4785), .A2(n4784), .ZN(n4787) );
  OAI211_X1 U9536 ( .C1(n4789), .C2(n4788), .A(n4787), .B(n4786), .ZN(n5952)
         );
  NAND2_X1 U9537 ( .A1(n5101), .A2(n5107), .ZN(n4791) );
  MUX2_X1 U9538 ( .A(n4791), .B(n4790), .S(n5102), .Z(n4794) );
  INV_X1 U9539 ( .A(n4795), .ZN(n4797) );
  NAND2_X1 U9540 ( .A1(n4799), .A2(n4798), .ZN(n4800) );
  NAND2_X1 U9541 ( .A1(n4801), .A2(n20016), .ZN(n4808) );
  NAND2_X1 U9542 ( .A1(n4802), .A2(n20202), .ZN(n4803) );
  NAND3_X1 U9543 ( .A1(n4808), .A2(n5090), .A3(n4803), .ZN(n4806) );
  OAI211_X1 U9544 ( .C1(n4808), .C2(n4807), .A(n4806), .B(n4805), .ZN(n5949)
         );
  NOR2_X1 U9545 ( .A1(n6101), .A2(n5949), .ZN(n4822) );
  NAND2_X1 U9546 ( .A1(n20431), .A2(n5075), .ZN(n4811) );
  OAI21_X1 U9547 ( .B1(n5075), .B2(n5077), .A(n4811), .ZN(n4812) );
  INV_X1 U9548 ( .A(n6097), .ZN(n5662) );
  INV_X1 U9549 ( .A(n4814), .ZN(n4815) );
  NAND2_X1 U9550 ( .A1(n4815), .A2(n5069), .ZN(n4820) );
  OAI21_X1 U9551 ( .B1(n2971), .B2(n291), .A(n5073), .ZN(n4817) );
  NAND2_X1 U9552 ( .A1(n4818), .A2(n4817), .ZN(n4819) );
  NAND2_X1 U9553 ( .A1(n5950), .A2(n5664), .ZN(n4821) );
  INV_X1 U9554 ( .A(n4823), .ZN(n4833) );
  NAND2_X1 U9555 ( .A1(n4828), .A2(n4827), .ZN(n4830) );
  MUX2_X1 U9556 ( .A(n4831), .B(n4830), .S(n4829), .Z(n4832) );
  OAI21_X1 U9557 ( .B1(n19688), .B2(n4833), .A(n4832), .ZN(n5200) );
  AOI21_X1 U9558 ( .B1(n20256), .B2(n4834), .A(n169), .ZN(n4836) );
  OR2_X1 U9559 ( .A1(n4836), .A2(n4835), .ZN(n4837) );
  INV_X1 U9560 ( .A(n6092), .ZN(n5912) );
  INV_X1 U9561 ( .A(n4839), .ZN(n4843) );
  NOR2_X1 U9562 ( .A1(n4841), .A2(n4840), .ZN(n4842) );
  NOR2_X1 U9563 ( .A1(n4846), .A2(n4845), .ZN(n5902) );
  INV_X1 U9564 ( .A(n5902), .ZN(n4847) );
  INV_X1 U9566 ( .A(n6090), .ZN(n5493) );
  NAND2_X1 U9567 ( .A1(n4850), .A2(n4849), .ZN(n4852) );
  OAI211_X1 U9568 ( .C1(n4854), .C2(n4853), .A(n4852), .B(n4851), .ZN(n6087)
         );
  INV_X1 U9569 ( .A(n6087), .ZN(n5176) );
  NAND2_X1 U9570 ( .A1(n5493), .A2(n5176), .ZN(n4876) );
  INV_X1 U9572 ( .A(n4856), .ZN(n4903) );
  NAND2_X1 U9573 ( .A1(n4903), .A2(n4901), .ZN(n4858) );
  NAND2_X1 U9574 ( .A1(n4858), .A2(n4857), .ZN(n4859) );
  INV_X1 U9575 ( .A(n5901), .ZN(n4862) );
  NAND3_X1 U9576 ( .A1(n20357), .A2(n4867), .A3(n896), .ZN(n4869) );
  NAND3_X1 U9577 ( .A1(n4871), .A2(n4870), .A3(n4869), .ZN(n4872) );
  NAND2_X1 U9578 ( .A1(n890), .A2(n5899), .ZN(n4874) );
  XNOR2_X1 U9579 ( .A(n7184), .B(n6918), .ZN(n7040) );
  INV_X1 U9580 ( .A(n5670), .ZN(n5185) );
  NAND2_X1 U9581 ( .A1(n5185), .A2(n5425), .ZN(n4880) );
  NAND2_X1 U9582 ( .A1(n5675), .A2(n5668), .ZN(n5677) );
  INV_X1 U9583 ( .A(n5669), .ZN(n5676) );
  OAI21_X1 U9584 ( .B1(n3397), .B2(n5670), .A(n5676), .ZN(n4878) );
  OAI21_X1 U9585 ( .B1(n5279), .B2(n5668), .A(n5669), .ZN(n4877) );
  NAND2_X1 U9586 ( .A1(n4878), .A2(n4877), .ZN(n4879) );
  NOR2_X1 U9587 ( .A1(n20509), .A2(n5745), .ZN(n5497) );
  NAND2_X1 U9588 ( .A1(n5201), .A2(n5741), .ZN(n4881) );
  NAND2_X1 U9589 ( .A1(n5497), .A2(n4881), .ZN(n4884) );
  INV_X1 U9590 ( .A(n4882), .ZN(n5749) );
  NAND3_X1 U9591 ( .A1(n5741), .A2(n5743), .A3(n5745), .ZN(n4883) );
  XNOR2_X1 U9592 ( .A(n7188), .B(n7337), .ZN(n4938) );
  INV_X1 U9593 ( .A(n4885), .ZN(n4891) );
  OAI21_X1 U9594 ( .B1(n4946), .B2(n4887), .A(n4886), .ZN(n4890) );
  OAI21_X1 U9596 ( .B1(n4892), .B2(n4893), .A(n4899), .ZN(n4897) );
  AOI21_X1 U9598 ( .B1(n4903), .B2(n4902), .A(n4901), .ZN(n4908) );
  NAND2_X1 U9599 ( .A1(n4905), .A2(n4904), .ZN(n4906) );
  NAND2_X1 U9600 ( .A1(n4912), .A2(n4911), .ZN(n4955) );
  NAND3_X1 U9602 ( .A1(n4955), .A2(n4916), .A3(n4915), .ZN(n4917) );
  NAND2_X1 U9603 ( .A1(n5684), .A2(n5476), .ZN(n5680) );
  NAND2_X1 U9604 ( .A1(n4968), .A2(n19507), .ZN(n4920) );
  OAI211_X1 U9605 ( .C1(n4921), .C2(n19507), .A(n4920), .B(n4919), .ZN(n4923)
         );
  OAI21_X1 U9606 ( .B1(n3967), .B2(n4965), .A(n4482), .ZN(n4922) );
  NAND2_X1 U9607 ( .A1(n4923), .A2(n4922), .ZN(n4924) );
  OAI21_X1 U9608 ( .B1(n4926), .B2(n19507), .A(n4924), .ZN(n6083) );
  INV_X1 U9609 ( .A(n6083), .ZN(n5411) );
  AOI22_X1 U9610 ( .A1(n5686), .A2(n5680), .B1(n5411), .B2(n3529), .ZN(n4936)
         );
  NAND2_X1 U9611 ( .A1(n4928), .A2(n4974), .ZN(n4929) );
  AOI22_X1 U9612 ( .A1(n4931), .A2(n4930), .B1(n4929), .B2(n4976), .ZN(n4934)
         );
  NOR2_X1 U9613 ( .A1(n4932), .A2(n4974), .ZN(n4933) );
  OR2_X1 U9614 ( .A1(n5683), .A2(n5410), .ZN(n5412) );
  NOR2_X1 U9615 ( .A1(n5412), .A2(n5684), .ZN(n4935) );
  OR2_X1 U9616 ( .A1(n4936), .A2(n4935), .ZN(n7383) );
  INV_X1 U9617 ( .A(n7383), .ZN(n4937) );
  XNOR2_X1 U9618 ( .A(n4938), .B(n4937), .ZN(n6877) );
  XNOR2_X1 U9619 ( .A(n4939), .B(n6877), .ZN(n8185) );
  INV_X1 U9620 ( .A(n8062), .ZN(n7606) );
  NAND2_X1 U9623 ( .A1(n4945), .A2(n4118), .ZN(n4944) );
  OAI21_X1 U9624 ( .B1(n4946), .B2(n4945), .A(n4944), .ZN(n4948) );
  NAND2_X1 U9625 ( .A1(n4951), .A2(n4950), .ZN(n4959) );
  NAND2_X1 U9626 ( .A1(n292), .A2(n20205), .ZN(n4964) );
  NAND2_X1 U9627 ( .A1(n4962), .A2(n4892), .ZN(n4963) );
  AOI21_X1 U9628 ( .B1(n4967), .B2(n4966), .A(n4965), .ZN(n4973) );
  AOI21_X1 U9629 ( .B1(n4971), .B2(n4970), .A(n4482), .ZN(n4972) );
  INV_X1 U9630 ( .A(n6036), .ZN(n5564) );
  INV_X1 U9631 ( .A(n5531), .ZN(n4981) );
  INV_X1 U9632 ( .A(n4974), .ZN(n4975) );
  NAND3_X1 U9633 ( .A1(n6033), .A2(n4981), .A3(n20241), .ZN(n4992) );
  NAND2_X1 U9634 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  NAND2_X1 U9635 ( .A1(n4985), .A2(n4984), .ZN(n4986) );
  NAND2_X1 U9636 ( .A1(n4989), .A2(n4988), .ZN(n4990) );
  AND2_X1 U9637 ( .A1(n4992), .A2(n5471), .ZN(n4993) );
  NAND2_X1 U9638 ( .A1(n5328), .A2(n6048), .ZN(n4999) );
  NOR2_X1 U9639 ( .A1(n5559), .A2(n6050), .ZN(n4994) );
  NAND2_X1 U9640 ( .A1(n3351), .A2(n4994), .ZN(n4998) );
  NAND3_X1 U9642 ( .A1(n5139), .A2(n5138), .A3(n6049), .ZN(n4996) );
  XNOR2_X1 U9644 ( .A(n7318), .B(n7371), .ZN(n6889) );
  AOI21_X1 U9645 ( .B1(n5405), .B2(n3959), .A(n5148), .ZN(n5002) );
  NOR2_X1 U9646 ( .A1(n5408), .A2(n5580), .ZN(n5318) );
  OAI21_X1 U9647 ( .B1(n5318), .B2(n5000), .A(n946), .ZN(n5001) );
  AOI22_X1 U9648 ( .A1(n5007), .A2(n5004), .B1(n5003), .B2(n5006), .ZN(n5011)
         );
  NAND2_X1 U9649 ( .A1(n4248), .A2(n5004), .ZN(n5008) );
  NAND3_X1 U9651 ( .A1(n5015), .A2(n5014), .A3(n5013), .ZN(n5020) );
  NAND3_X1 U9652 ( .A1(n5018), .A2(n20229), .A3(n5016), .ZN(n5019) );
  NAND2_X1 U9653 ( .A1(n5030), .A2(n5927), .ZN(n5066) );
  INV_X1 U9654 ( .A(n6027), .ZN(n5192) );
  NAND2_X1 U9655 ( .A1(n5032), .A2(n153), .ZN(n5033) );
  NAND2_X1 U9656 ( .A1(n5034), .A2(n5033), .ZN(n5039) );
  INV_X1 U9657 ( .A(n6025), .ZN(n5520) );
  NAND3_X1 U9658 ( .A1(n6026), .A2(n5192), .A3(n5520), .ZN(n5065) );
  NAND2_X1 U9659 ( .A1(n5040), .A2(n5045), .ZN(n5041) );
  OAI211_X1 U9660 ( .C1(n5044), .C2(n5043), .A(n5042), .B(n5041), .ZN(n5051)
         );
  AND2_X1 U9661 ( .A1(n5046), .A2(n5045), .ZN(n5049) );
  OAI211_X1 U9662 ( .C1(n5049), .C2(n20464), .A(n5048), .B(n5047), .ZN(n5050)
         );
  NAND2_X1 U9663 ( .A1(n5927), .A2(n5926), .ZN(n5064) );
  NAND3_X1 U9664 ( .A1(n5057), .A2(n5056), .A3(n5055), .ZN(n5062) );
  NAND3_X1 U9665 ( .A1(n5060), .A2(n5059), .A3(n5058), .ZN(n5061) );
  NAND3_X1 U9666 ( .A1(n5192), .A2(n19789), .A3(n5930), .ZN(n5063) );
  INV_X1 U9667 ( .A(n7373), .ZN(n5067) );
  XNOR2_X1 U9668 ( .A(n7088), .B(n5067), .ZN(n5068) );
  XNOR2_X1 U9669 ( .A(n5068), .B(n6889), .ZN(n5134) );
  OR2_X1 U9670 ( .A1(n5070), .A2(n5069), .ZN(n5504) );
  AND3_X1 U9671 ( .A1(n5080), .A2(n3451), .A3(n5079), .ZN(n5508) );
  OAI21_X1 U9673 ( .B1(n5083), .B2(n5086), .A(n20016), .ZN(n5085) );
  OR3_X1 U9674 ( .A1(n5088), .A2(n5087), .A3(n5086), .ZN(n5089) );
  INV_X1 U9675 ( .A(n19979), .ZN(n5921) );
  OAI22_X1 U9676 ( .A1(n6007), .A2(n5914), .B1(n5921), .B2(n861), .ZN(n5111)
         );
  MUX2_X1 U9678 ( .A(n5107), .B(n5106), .S(n4048), .Z(n5109) );
  NAND2_X1 U9679 ( .A1(n5109), .A2(n5108), .ZN(n5110) );
  NAND2_X1 U9680 ( .A1(n5111), .A2(n5590), .ZN(n5123) );
  NAND2_X1 U9681 ( .A1(n20256), .A2(n19508), .ZN(n5113) );
  AOI21_X1 U9682 ( .B1(n5114), .B2(n5113), .A(n5115), .ZN(n5121) );
  NAND2_X1 U9683 ( .A1(n5116), .A2(n5115), .ZN(n5119) );
  AOI21_X1 U9684 ( .B1(n5119), .B2(n169), .A(n19508), .ZN(n5120) );
  INV_X1 U9685 ( .A(n5823), .ZN(n5828) );
  NAND3_X1 U9686 ( .A1(n5828), .A2(n5447), .A3(n3569), .ZN(n5127) );
  NAND2_X1 U9687 ( .A1(n5124), .A2(n5823), .ZN(n5126) );
  NAND3_X1 U9688 ( .A1(n5447), .A2(n5825), .A3(n6016), .ZN(n5125) );
  XNOR2_X1 U9689 ( .A(n7046), .B(n7179), .ZN(n6579) );
  NAND2_X1 U9690 ( .A1(n5647), .A2(n5641), .ZN(n5128) );
  AOI21_X1 U9691 ( .B1(n5128), .B2(n5648), .A(n5649), .ZN(n5131) );
  NAND2_X1 U9692 ( .A1(n5442), .A2(n5444), .ZN(n5291) );
  NAND3_X1 U9693 ( .A1(n5649), .A2(n5444), .A3(n5643), .ZN(n5129) );
  NAND2_X1 U9694 ( .A1(n5291), .A2(n5129), .ZN(n5130) );
  XNOR2_X1 U9695 ( .A(n7144), .B(n1840), .ZN(n5132) );
  XNOR2_X1 U9696 ( .A(n6579), .B(n5132), .ZN(n5133) );
  AOI21_X1 U9697 ( .B1(n20465), .B2(n8184), .A(n8060), .ZN(n5135) );
  AND2_X1 U9698 ( .A1(n8182), .A2(n5135), .ZN(n5136) );
  INV_X1 U9699 ( .A(n5559), .ZN(n6051) );
  AND2_X1 U9702 ( .A1(n5559), .A2(n6049), .ZN(n5329) );
  NOR3_X1 U9703 ( .A1(n5329), .A2(n3351), .A3(n5330), .ZN(n5142) );
  NAND2_X1 U9704 ( .A1(n6044), .A2(n5888), .ZN(n5781) );
  INV_X1 U9705 ( .A(n6041), .ZN(n5776) );
  NAND3_X1 U9706 ( .A1(n135), .A2(n5776), .A3(n5309), .ZN(n5145) );
  XNOR2_X1 U9707 ( .A(n6674), .B(n6494), .ZN(n7228) );
  NAND3_X1 U9708 ( .A1(n5571), .A2(n5580), .A3(n5582), .ZN(n5151) );
  NAND2_X1 U9709 ( .A1(n5408), .A2(n3959), .ZN(n5317) );
  NAND3_X2 U9710 ( .A1(n5152), .A2(n5151), .A3(n5150), .ZN(n7212) );
  OAI21_X1 U9711 ( .B1(n6068), .B2(n5978), .A(n6069), .ZN(n5155) );
  INV_X1 U9712 ( .A(n5978), .ZN(n6075) );
  NOR2_X1 U9713 ( .A1(n6067), .A2(n6072), .ZN(n5880) );
  XNOR2_X1 U9714 ( .A(n7212), .B(n7232), .ZN(n6801) );
  XNOR2_X1 U9715 ( .A(n6801), .B(n7228), .ZN(n5166) );
  INV_X1 U9716 ( .A(n5796), .ZN(n5792) );
  XNOR2_X1 U9717 ( .A(n7364), .B(n7211), .ZN(n5164) );
  INV_X1 U9718 ( .A(n6057), .ZN(n6056) );
  NAND3_X1 U9719 ( .A1(n6064), .A2(n6056), .A3(n5891), .ZN(n5162) );
  NAND3_X1 U9720 ( .A1(n6064), .A2(n6057), .A3(n6055), .ZN(n5161) );
  INV_X1 U9721 ( .A(n5782), .ZN(n5895) );
  NAND3_X1 U9722 ( .A1(n6058), .A2(n20670), .A3(n5895), .ZN(n5160) );
  NAND3_X1 U9723 ( .A1(n906), .A2(n5891), .A3(n6059), .ZN(n5159) );
  XNOR2_X1 U9724 ( .A(n7365), .B(n2096), .ZN(n5163) );
  XNOR2_X1 U9725 ( .A(n5164), .B(n5163), .ZN(n5165) );
  NAND2_X1 U9726 ( .A1(n5663), .A2(n5953), .ZN(n5167) );
  NAND2_X1 U9727 ( .A1(n5661), .A2(n5167), .ZN(n5171) );
  OAI21_X1 U9728 ( .B1(n6097), .B2(n5949), .A(n6101), .ZN(n5170) );
  INV_X1 U9729 ( .A(n5949), .ZN(n5168) );
  NOR2_X1 U9730 ( .A1(n5663), .A2(n5168), .ZN(n5169) );
  AOI21_X2 U9731 ( .B1(n5171), .B2(n5170), .A(n5169), .ZN(n6679) );
  INV_X1 U9732 ( .A(n6105), .ZN(n5955) );
  NAND3_X1 U9733 ( .A1(n5955), .A2(n5957), .A3(n6109), .ZN(n5175) );
  NAND3_X1 U9734 ( .A1(n5172), .A2(n6108), .A3(n6109), .ZN(n5174) );
  NAND3_X1 U9735 ( .A1(n6113), .A2(n5957), .A3(n6104), .ZN(n5173) );
  XNOR2_X1 U9736 ( .A(n6679), .B(n6634), .ZN(n7279) );
  INV_X1 U9737 ( .A(n7279), .ZN(n6926) );
  OAI21_X1 U9738 ( .B1(n5199), .B2(n890), .A(n20149), .ZN(n5177) );
  INV_X1 U9739 ( .A(n5200), .ZN(n5494) );
  NAND3_X1 U9740 ( .A1(n5742), .A2(n5201), .A3(n5749), .ZN(n5178) );
  XNOR2_X1 U9741 ( .A(n6926), .B(n7377), .ZN(n5191) );
  INV_X1 U9742 ( .A(n5682), .ZN(n6084) );
  INV_X1 U9743 ( .A(n5476), .ZN(n6082) );
  OAI21_X1 U9744 ( .B1(n6082), .B2(n6083), .A(n5684), .ZN(n5182) );
  AND2_X1 U9745 ( .A1(n5682), .A2(n6083), .ZN(n5181) );
  INV_X1 U9746 ( .A(n5425), .ZN(n5184) );
  NAND2_X1 U9747 ( .A1(n5668), .A2(n5184), .ZN(n5188) );
  NAND3_X1 U9748 ( .A1(n5669), .A2(n5185), .A3(n5184), .ZN(n5186) );
  XNOR2_X1 U9749 ( .A(n7144), .B(n19205), .ZN(n5189) );
  XNOR2_X1 U9750 ( .A(n6838), .B(n5189), .ZN(n5190) );
  INV_X1 U9751 ( .A(n5926), .ZN(n5931) );
  OR2_X1 U9752 ( .A1(n5931), .A2(n6025), .ZN(n6030) );
  AOI21_X1 U9753 ( .B1(n6028), .B2(n6030), .A(n5192), .ZN(n5195) );
  AOI21_X1 U9755 ( .B1(n5193), .B2(n5926), .A(n5929), .ZN(n5194) );
  NAND2_X1 U9756 ( .A1(n5736), .A2(n5768), .ZN(n5224) );
  INV_X1 U9758 ( .A(n5763), .ZN(n5769) );
  AOI21_X1 U9759 ( .B1(n5224), .B2(n5225), .A(n5769), .ZN(n5198) );
  NAND2_X1 U9760 ( .A1(n5765), .A2(n5767), .ZN(n5196) );
  AOI21_X1 U9761 ( .B1(n5766), .B2(n5196), .A(n5736), .ZN(n5197) );
  NAND2_X1 U9762 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  NAND2_X1 U9763 ( .A1(n5204), .A2(n5745), .ZN(n5206) );
  NAND2_X1 U9764 ( .A1(n5742), .A2(n5746), .ZN(n5205) );
  XNOR2_X1 U9766 ( .A(n7238), .B(n6824), .ZN(n5214) );
  INV_X1 U9767 ( .A(n6007), .ZN(n5207) );
  INV_X1 U9768 ( .A(n5917), .ZN(n6013) );
  AOI21_X1 U9769 ( .B1(n5916), .B2(n5207), .A(n6013), .ZN(n5210) );
  NAND2_X1 U9770 ( .A1(n5208), .A2(n6010), .ZN(n5209) );
  XNOR2_X1 U9771 ( .A(n7392), .B(n6854), .ZN(n5212) );
  INV_X1 U9772 ( .A(n20672), .ZN(n18660) );
  XNOR2_X1 U9773 ( .A(n7196), .B(n18660), .ZN(n5211) );
  XNOR2_X1 U9774 ( .A(n5212), .B(n5211), .ZN(n5213) );
  NOR2_X1 U9775 ( .A1(n8304), .A2(n8301), .ZN(n5272) );
  AOI21_X1 U9777 ( .B1(n5631), .B2(n5633), .A(n5363), .ZN(n5216) );
  INV_X1 U9778 ( .A(n6808), .ZN(n5222) );
  INV_X1 U9779 ( .A(n6167), .ZN(n6176) );
  AND2_X1 U9780 ( .A1(n5218), .A2(n5217), .ZN(n5220) );
  NAND2_X1 U9782 ( .A1(n6176), .A2(n5945), .ZN(n5943) );
  NAND2_X1 U9783 ( .A1(n6172), .A2(n6168), .ZN(n6175) );
  INV_X1 U9784 ( .A(n6171), .ZN(n5842) );
  OAI211_X1 U9785 ( .C1(n6166), .C2(n6172), .A(n170), .B(n5842), .ZN(n5221) );
  XNOR2_X1 U9786 ( .A(n5222), .B(n6873), .ZN(n7381) );
  INV_X1 U9787 ( .A(n7381), .ZN(n6464) );
  OAI211_X1 U9788 ( .C1(n5763), .C2(n5768), .A(n5546), .B(n5734), .ZN(n5223)
         );
  INV_X1 U9790 ( .A(n5839), .ZN(n6203) );
  NOR2_X1 U9792 ( .A1(n6204), .A2(n19968), .ZN(n5230) );
  NAND3_X1 U9793 ( .A1(n6218), .A2(n6205), .A3(n19492), .ZN(n5227) );
  OAI21_X1 U9794 ( .B1(n5226), .B2(n6218), .A(n5227), .ZN(n5228) );
  INV_X1 U9795 ( .A(n5228), .ZN(n5229) );
  XNOR2_X1 U9796 ( .A(n7187), .B(n7249), .ZN(n6810) );
  XNOR2_X1 U9797 ( .A(n6810), .B(n6464), .ZN(n5239) );
  NAND2_X1 U9798 ( .A1(n5382), .A2(n6189), .ZN(n5234) );
  INV_X1 U9799 ( .A(n6190), .ZN(n5232) );
  NOR2_X1 U9800 ( .A1(n5805), .A2(n6189), .ZN(n5231) );
  OAI22_X1 U9801 ( .A1(n5232), .A2(n5231), .B1(n6194), .B2(n5803), .ZN(n5233)
         );
  INV_X1 U9802 ( .A(n6919), .ZN(n6513) );
  NOR2_X1 U9803 ( .A1(n6184), .A2(n5845), .ZN(n5235) );
  INV_X1 U9804 ( .A(n5728), .ZN(n6380) );
  XNOR2_X1 U9805 ( .A(n6513), .B(n7248), .ZN(n5237) );
  XNOR2_X1 U9806 ( .A(n7188), .B(n2221), .ZN(n5236) );
  XNOR2_X1 U9807 ( .A(n5237), .B(n5236), .ZN(n5238) );
  NOR2_X1 U9808 ( .A1(n8046), .A2(n8044), .ZN(n5271) );
  INV_X1 U9809 ( .A(n5240), .ZN(n5241) );
  OAI211_X1 U9810 ( .C1(n5346), .C2(n5605), .A(n5243), .B(n5720), .ZN(n5244)
         );
  NAND2_X1 U9811 ( .A1(n6150), .A2(n5612), .ZN(n5246) );
  XNOR2_X1 U9813 ( .A(n7254), .B(n5249), .ZN(n6590) );
  INV_X1 U9814 ( .A(n6590), .ZN(n6818) );
  NAND2_X1 U9815 ( .A1(n5401), .A2(n5251), .ZN(n5252) );
  INV_X1 U9816 ( .A(n6123), .ZN(n5338) );
  NAND2_X1 U9817 ( .A1(n6128), .A2(n5338), .ZN(n5870) );
  OAI21_X1 U9818 ( .B1(n6128), .B2(n6119), .A(n5386), .ZN(n5260) );
  NAND2_X1 U9819 ( .A1(n5255), .A2(n19688), .ZN(n5256) );
  OAI211_X1 U9820 ( .C1(n19688), .C2(n5257), .A(n6128), .B(n5256), .ZN(n5259)
         );
  OAI211_X1 U9821 ( .C1(n6117), .C2(n6128), .A(n5260), .B(n5259), .ZN(n5261)
         );
  XNOR2_X1 U9822 ( .A(n6818), .B(n7353), .ZN(n5270) );
  XNOR2_X1 U9823 ( .A(n20203), .B(n2296), .ZN(n5268) );
  MUX2_X1 U9824 ( .A(n6129), .B(n6131), .S(n6133), .Z(n5263) );
  NAND2_X1 U9826 ( .A1(n6139), .A2(n6138), .ZN(n5265) );
  MUX2_X1 U9827 ( .A(n5267), .B(n5266), .S(n5860), .Z(n6285) );
  XNOR2_X1 U9828 ( .A(n6285), .B(n6520), .ZN(n7256) );
  XNOR2_X1 U9829 ( .A(n7256), .B(n5268), .ZN(n5269) );
  AND2_X1 U9830 ( .A1(n5704), .A2(n5997), .ZN(n5433) );
  NAND2_X1 U9831 ( .A1(n5433), .A2(n5434), .ZN(n5274) );
  NAND3_X1 U9832 ( .A1(n19562), .A2(n5996), .A3(n6002), .ZN(n5273) );
  XNOR2_X1 U9833 ( .A(n6850), .B(n19222), .ZN(n5278) );
  NAND2_X1 U9834 ( .A1(n5711), .A2(n5985), .ZN(n5993) );
  INV_X1 U9835 ( .A(n5711), .ZN(n5817) );
  NAND2_X1 U9836 ( .A1(n5818), .A2(n5989), .ZN(n5277) );
  XNOR2_X1 U9837 ( .A(n5278), .B(n6947), .ZN(n5284) );
  NAND2_X1 U9838 ( .A1(n3397), .A2(n5425), .ZN(n5282) );
  NOR2_X1 U9839 ( .A1(n5670), .A2(n5279), .ZN(n5280) );
  XNOR2_X1 U9840 ( .A(n7202), .B(n6945), .ZN(n5283) );
  XNOR2_X1 U9841 ( .A(n5284), .B(n5283), .ZN(n5297) );
  NOR2_X1 U9842 ( .A1(n3569), .A2(n6017), .ZN(n5286) );
  NOR2_X1 U9843 ( .A1(n5823), .A2(n5827), .ZN(n5285) );
  OAI21_X1 U9844 ( .B1(n5286), .B2(n5285), .A(n5825), .ZN(n5288) );
  NAND3_X1 U9845 ( .A1(n5824), .A2(n5826), .A3(n6022), .ZN(n5287) );
  INV_X1 U9846 ( .A(n5442), .ZN(n5646) );
  NAND2_X1 U9847 ( .A1(n5646), .A2(n5641), .ZN(n5289) );
  INV_X1 U9848 ( .A(n5443), .ZN(n5642) );
  NAND3_X1 U9849 ( .A1(n5645), .A2(n5649), .A3(n5642), .ZN(n5290) );
  XNOR2_X1 U9850 ( .A(n7006), .B(n7266), .ZN(n5296) );
  MUX2_X1 U9851 ( .A(n5699), .B(n5971), .S(n5968), .Z(n5295) );
  INV_X1 U9852 ( .A(n5524), .ZN(n5967) );
  NOR2_X1 U9853 ( .A1(n5697), .A2(n5967), .ZN(n5450) );
  NAND2_X1 U9854 ( .A1(n5450), .A2(n5973), .ZN(n5293) );
  NAND2_X1 U9855 ( .A1(n957), .A2(n5971), .ZN(n5292) );
  OAI211_X1 U9856 ( .C1(n5295), .C2(n5294), .A(n5293), .B(n5292), .ZN(n6348)
         );
  INV_X1 U9857 ( .A(n6348), .ZN(n7344) );
  XNOR2_X1 U9858 ( .A(n7344), .B(n5296), .ZN(n6835) );
  NAND3_X1 U9859 ( .A1(n20001), .A2(n8301), .A3(n8303), .ZN(n5298) );
  NAND2_X1 U9860 ( .A1(n5792), .A2(n5300), .ZN(n5303) );
  NOR2_X1 U9861 ( .A1(n5798), .A2(n19912), .ZN(n5302) );
  INV_X1 U9862 ( .A(n5300), .ZN(n5790) );
  OAI211_X1 U9863 ( .C1(n5304), .C2(n6059), .A(n5895), .B(n6057), .ZN(n5307)
         );
  INV_X1 U9864 ( .A(n6061), .ZN(n5306) );
  XNOR2_X1 U9865 ( .A(n6687), .B(n7338), .ZN(n5315) );
  OAI21_X1 U9866 ( .B1(n6044), .B2(n5309), .A(n5308), .ZN(n6047) );
  NOR2_X1 U9867 ( .A1(n6046), .A2(n5888), .ZN(n5310) );
  NOR2_X1 U9868 ( .A1(n5311), .A2(n5310), .ZN(n5313) );
  INV_X1 U9869 ( .A(n5311), .ZN(n5312) );
  INV_X1 U9870 ( .A(n6728), .ZN(n5314) );
  XNOR2_X1 U9871 ( .A(n5315), .B(n5314), .ZN(n6630) );
  OAI21_X1 U9872 ( .B1(n5582), .B2(n5581), .A(n5317), .ZN(n5406) );
  INV_X1 U9873 ( .A(n5318), .ZN(n5319) );
  INV_X1 U9874 ( .A(n6782), .ZN(n5321) );
  XNOR2_X1 U9875 ( .A(n5321), .B(n7134), .ZN(n5690) );
  NOR2_X1 U9876 ( .A1(n1838), .A2(n5398), .ZN(n5327) );
  NAND2_X1 U9877 ( .A1(n5397), .A2(n5323), .ZN(n5324) );
  XNOR2_X1 U9878 ( .A(n7041), .B(n18691), .ZN(n5335) );
  NAND2_X1 U9879 ( .A1(n5329), .A2(n5328), .ZN(n5334) );
  NAND2_X1 U9880 ( .A1(n6052), .A2(n6051), .ZN(n5333) );
  NAND2_X1 U9881 ( .A1(n5330), .A2(n6050), .ZN(n5332) );
  NAND2_X1 U9882 ( .A1(n5330), .A2(n6051), .ZN(n5331) );
  NAND4_X1 U9883 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n6573)
         );
  INV_X1 U9884 ( .A(n6573), .ZN(n6038) );
  XNOR2_X1 U9885 ( .A(n5335), .B(n6038), .ZN(n5336) );
  XNOR2_X1 U9886 ( .A(n5690), .B(n5336), .ZN(n5337) );
  NAND3_X1 U9888 ( .A1(n5868), .A2(n5338), .A3(n6119), .ZN(n5339) );
  NAND2_X1 U9889 ( .A1(n5386), .A2(n6118), .ZN(n6127) );
  AND2_X1 U9890 ( .A1(n6127), .A2(n5339), .ZN(n5340) );
  OAI21_X2 U9891 ( .B1(n6128), .B2(n5341), .A(n5340), .ZN(n7087) );
  INV_X1 U9892 ( .A(n6140), .ZN(n5866) );
  NAND2_X1 U9893 ( .A1(n5866), .A2(n5860), .ZN(n5345) );
  OAI21_X1 U9894 ( .B1(n20334), .B2(n6140), .A(n5342), .ZN(n5344) );
  INV_X1 U9895 ( .A(n6724), .ZN(n6633) );
  XNOR2_X1 U9896 ( .A(n6633), .B(n7087), .ZN(n6237) );
  INV_X1 U9897 ( .A(n6237), .ZN(n5354) );
  MUX2_X1 U9898 ( .A(n5604), .B(n5605), .S(n5716), .Z(n5348) );
  NAND2_X1 U9899 ( .A1(n5605), .A2(n5346), .ZN(n5347) );
  OR2_X1 U9900 ( .A1(n5610), .A2(n1277), .ZN(n5352) );
  NAND2_X1 U9901 ( .A1(n6153), .A2(n5349), .ZN(n5351) );
  NAND3_X1 U9902 ( .A1(n5611), .A2(n6156), .A3(n6159), .ZN(n5350) );
  XNOR2_X1 U9903 ( .A(n5354), .B(n6506), .ZN(n5377) );
  NAND2_X1 U9904 ( .A1(n5356), .A2(n5623), .ZN(n5355) );
  AOI21_X1 U9905 ( .B1(n5355), .B2(n5692), .A(n6131), .ZN(n5359) );
  NAND2_X1 U9906 ( .A1(n5691), .A2(n6131), .ZN(n5357) );
  AOI21_X1 U9907 ( .B1(n5621), .B2(n5357), .A(n5356), .ZN(n5358) );
  INV_X1 U9908 ( .A(n7142), .ZN(n6469) );
  INV_X1 U9909 ( .A(n5360), .ZN(n5362) );
  NAND2_X1 U9910 ( .A1(n5631), .A2(n5364), .ZN(n5361) );
  AOI21_X1 U9911 ( .B1(n5362), .B2(n5361), .A(n4598), .ZN(n5366) );
  NAND2_X1 U9912 ( .A1(n4598), .A2(n5363), .ZN(n5629) );
  INV_X1 U9913 ( .A(n5633), .ZN(n5466) );
  AOI21_X1 U9914 ( .B1(n5629), .B2(n5466), .A(n5364), .ZN(n5365) );
  NOR2_X1 U9915 ( .A1(n5366), .A2(n5365), .ZN(n7048) );
  INV_X1 U9916 ( .A(n7048), .ZN(n6680) );
  XNOR2_X1 U9917 ( .A(n6469), .B(n6680), .ZN(n5375) );
  NAND2_X1 U9918 ( .A1(n5392), .A2(n5367), .ZN(n5372) );
  OAI21_X1 U9919 ( .B1(n5394), .B2(n5398), .A(n5395), .ZN(n5370) );
  NAND2_X1 U9920 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  XNOR2_X1 U9921 ( .A(n7316), .B(n2123), .ZN(n5374) );
  XNOR2_X1 U9922 ( .A(n5375), .B(n5374), .ZN(n5376) );
  OAI21_X1 U9923 ( .B1(n5379), .B2(n6192), .A(n5802), .ZN(n5381) );
  OAI211_X1 U9924 ( .C1(n5733), .C2(n5382), .A(n5381), .B(n5380), .ZN(n6714)
         );
  NAND2_X1 U9925 ( .A1(n5728), .A2(n5845), .ZN(n5385) );
  NAND3_X1 U9926 ( .A1(n6183), .A2(n5845), .A3(n6184), .ZN(n5384) );
  XNOR2_X1 U9927 ( .A(n7065), .B(n6714), .ZN(n6640) );
  INV_X1 U9928 ( .A(n6640), .ZN(n5403) );
  NAND3_X1 U9929 ( .A1(n6120), .A2(n5386), .A3(n6119), .ZN(n5391) );
  AND2_X1 U9930 ( .A1(n6118), .A2(n6119), .ZN(n5867) );
  NAND2_X1 U9931 ( .A1(n5867), .A2(n6123), .ZN(n5389) );
  NAND2_X1 U9932 ( .A1(n5387), .A2(n6124), .ZN(n5388) );
  INV_X1 U9933 ( .A(n5392), .ZN(n5402) );
  OAI21_X1 U9934 ( .B1(n5395), .B2(n5394), .A(n5393), .ZN(n5396) );
  NAND2_X1 U9935 ( .A1(n5396), .A2(n5401), .ZN(n5400) );
  OAI211_X2 U9936 ( .C1(n5402), .C2(n5401), .A(n5400), .B(n5399), .ZN(n6777)
         );
  XNOR2_X1 U9937 ( .A(n7128), .B(n6777), .ZN(n6488) );
  XNOR2_X1 U9938 ( .A(n5403), .B(n6488), .ZN(n5423) );
  NAND2_X1 U9939 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  OR2_X1 U9940 ( .A1(n5410), .A2(n5682), .ZN(n6081) );
  INV_X1 U9941 ( .A(n5683), .ZN(n5479) );
  AOI21_X1 U9942 ( .B1(n6081), .B2(n5479), .A(n5476), .ZN(n5414) );
  AOI21_X1 U9943 ( .B1(n5412), .B2(n5680), .A(n5411), .ZN(n5413) );
  INV_X1 U9944 ( .A(n7014), .ZN(n5415) );
  XNOR2_X1 U9945 ( .A(n19855), .B(n5415), .ZN(n5421) );
  NAND2_X1 U9946 ( .A1(n6204), .A2(n19968), .ZN(n5419) );
  INV_X1 U9947 ( .A(n19492), .ZN(n5416) );
  OAI21_X1 U9948 ( .B1(n19522), .B2(n5416), .A(n6205), .ZN(n5417) );
  NAND3_X1 U9949 ( .A1(n6205), .A2(n19492), .A3(n3640), .ZN(n5418) );
  XNOR2_X1 U9950 ( .A(n7296), .B(n2376), .ZN(n5420) );
  XNOR2_X1 U9951 ( .A(n5421), .B(n5420), .ZN(n5422) );
  MUX2_X1 U9952 ( .A(n5670), .B(n5425), .S(n5424), .Z(n5427) );
  MUX2_X1 U9953 ( .A(n19912), .B(n5796), .S(n5428), .Z(n5430) );
  MUX2_X2 U9954 ( .A(n5431), .B(n5430), .S(n5429), .Z(n7253) );
  XNOR2_X1 U9955 ( .A(n7116), .B(n7253), .ZN(n5441) );
  INV_X1 U9956 ( .A(n5998), .ZN(n5432) );
  NAND2_X1 U9957 ( .A1(n5437), .A2(n5436), .ZN(n7081) );
  MUX2_X1 U9958 ( .A(n5711), .B(n5990), .S(n5985), .Z(n5440) );
  NOR2_X1 U9959 ( .A1(n5815), .A2(n5989), .ZN(n5988) );
  NOR2_X1 U9960 ( .A1(n5988), .A2(n5438), .ZN(n5439) );
  MUX2_X2 U9961 ( .A(n5440), .B(n5439), .S(n5818), .Z(n7122) );
  XNOR2_X1 U9962 ( .A(n5441), .B(n6621), .ZN(n5454) );
  MUX2_X1 U9963 ( .A(n5442), .B(n5641), .S(n5444), .Z(n5446) );
  MUX2_X1 U9964 ( .A(n5444), .B(n5649), .S(n5443), .Z(n5445) );
  MUX2_X1 U9965 ( .A(n5825), .B(n6017), .S(n6016), .Z(n5448) );
  XNOR2_X1 U9966 ( .A(n7257), .B(n7121), .ZN(n5599) );
  NAND3_X1 U9968 ( .A1(n5973), .A2(n19804), .A3(n20673), .ZN(n5451) );
  XNOR2_X1 U9969 ( .A(n7289), .B(n2455), .ZN(n5452) );
  XNOR2_X1 U9970 ( .A(n5599), .B(n5452), .ZN(n5453) );
  AOI21_X1 U9971 ( .B1(n6107), .B2(n6104), .A(n6105), .ZN(n5455) );
  NAND2_X1 U9972 ( .A1(n5663), .A2(n6101), .ZN(n5456) );
  OAI21_X1 U9973 ( .B1(n5662), .B2(n5663), .A(n5456), .ZN(n5457) );
  NAND2_X1 U9974 ( .A1(n5457), .A2(n283), .ZN(n5459) );
  INV_X1 U9975 ( .A(n6225), .ZN(n6646) );
  INV_X1 U9976 ( .A(n5945), .ZN(n6173) );
  NAND3_X1 U9977 ( .A1(n1867), .A2(n170), .A3(n6173), .ZN(n5460) );
  NAND2_X1 U9978 ( .A1(n5463), .A2(n4598), .ZN(n5470) );
  NAND3_X1 U9979 ( .A1(n5467), .A2(n5466), .A3(n31), .ZN(n5468) );
  XNOR2_X1 U9980 ( .A(n7160), .B(n7263), .ZN(n6484) );
  XNOR2_X1 U9981 ( .A(n6646), .B(n6484), .ZN(n5491) );
  INV_X1 U9982 ( .A(n5532), .ZN(n5529) );
  OAI21_X1 U9983 ( .B1(n5562), .B2(n2940), .A(n5529), .ZN(n5474) );
  NOR2_X1 U9984 ( .A1(n5532), .A2(n6036), .ZN(n5565) );
  INV_X1 U9985 ( .A(n5565), .ZN(n5473) );
  INV_X1 U9986 ( .A(n5566), .ZN(n6034) );
  NAND2_X1 U9987 ( .A1(n5476), .A2(n6083), .ZN(n5478) );
  MUX2_X1 U9988 ( .A(n5478), .B(n5477), .S(n5684), .Z(n5482) );
  NAND2_X1 U9989 ( .A1(n5682), .A2(n5479), .ZN(n6080) );
  OAI21_X1 U9990 ( .B1(n5681), .B2(n5479), .A(n6080), .ZN(n5480) );
  NAND2_X1 U9991 ( .A1(n5480), .A2(n6082), .ZN(n5481) );
  XNOR2_X1 U9992 ( .A(n7267), .B(n7306), .ZN(n5489) );
  NOR2_X1 U9993 ( .A1(n5719), .A2(n5715), .ZN(n5603) );
  NAND2_X1 U9994 ( .A1(n5603), .A2(n5717), .ZN(n5487) );
  NAND3_X1 U9995 ( .A1(n5605), .A2(n5715), .A3(n5720), .ZN(n5486) );
  AND2_X1 U9996 ( .A1(n5719), .A2(n5483), .ZN(n5602) );
  NAND3_X1 U9997 ( .A1(n5718), .A2(n5604), .A3(n5715), .ZN(n5484) );
  XNOR2_X1 U9998 ( .A(n7163), .B(n2395), .ZN(n5488) );
  XNOR2_X1 U9999 ( .A(n5489), .B(n5488), .ZN(n5490) );
  INV_X1 U10000 ( .A(n8034), .ZN(n7603) );
  INV_X1 U10001 ( .A(n5492), .ZN(n5900) );
  INV_X1 U10003 ( .A(n5497), .ZN(n5498) );
  NAND3_X1 U10004 ( .A1(n4632), .A2(n5741), .A3(n5746), .ZN(n5499) );
  INV_X1 U10007 ( .A(n862), .ZN(n5919) );
  NAND2_X1 U10008 ( .A1(n5502), .A2(n5919), .ZN(n5515) );
  INV_X1 U10009 ( .A(n5503), .ZN(n5513) );
  INV_X1 U10010 ( .A(n5504), .ZN(n5507) );
  INV_X1 U10011 ( .A(n5505), .ZN(n5506) );
  NOR2_X1 U10012 ( .A1(n5507), .A2(n5506), .ZN(n5512) );
  INV_X1 U10013 ( .A(n5508), .ZN(n5509) );
  AND2_X1 U10014 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  NAND4_X1 U10015 ( .A1(n5513), .A2(n862), .A3(n5512), .A4(n5511), .ZN(n5514)
         );
  NAND3_X1 U10016 ( .A1(n6014), .A2(n5515), .A3(n5514), .ZN(n5517) );
  NAND2_X1 U10017 ( .A1(n5517), .A2(n5516), .ZN(n6420) );
  NAND2_X1 U10018 ( .A1(n5927), .A2(n6025), .ZN(n5518) );
  NOR2_X1 U10019 ( .A1(n5926), .A2(n6031), .ZN(n5519) );
  XNOR2_X1 U10020 ( .A(n6420), .B(n6736), .ZN(n6626) );
  XNOR2_X1 U10021 ( .A(n6495), .B(n6626), .ZN(n5553) );
  NAND3_X1 U10022 ( .A1(n5528), .A2(n5967), .A3(n5523), .ZN(n5527) );
  NAND3_X1 U10023 ( .A1(n5700), .A2(n5525), .A3(n19804), .ZN(n5526) );
  OAI211_X1 U10024 ( .C1(n5700), .C2(n5528), .A(n5527), .B(n5526), .ZN(n7035)
         );
  NAND2_X1 U10025 ( .A1(n6036), .A2(n20241), .ZN(n5530) );
  NAND2_X1 U10026 ( .A1(n5531), .A2(n6036), .ZN(n5533) );
  OAI22_X1 U10027 ( .A1(n5534), .A2(n5569), .B1(n5533), .B2(n5532), .ZN(n5535)
         );
  NOR2_X1 U10028 ( .A1(n5536), .A2(n5535), .ZN(n6293) );
  INV_X1 U10029 ( .A(n6293), .ZN(n7326) );
  XNOR2_X1 U10030 ( .A(n7326), .B(n7035), .ZN(n5551) );
  NAND2_X1 U10031 ( .A1(n5736), .A2(n5734), .ZN(n5544) );
  INV_X1 U10032 ( .A(n5537), .ZN(n5542) );
  INV_X1 U10033 ( .A(n5538), .ZN(n5541) );
  NAND4_X1 U10034 ( .A1(n5542), .A2(n5541), .A3(n5540), .A4(n5539), .ZN(n5543)
         );
  NAND3_X1 U10035 ( .A1(n5544), .A2(n5768), .A3(n5543), .ZN(n5549) );
  NAND3_X1 U10036 ( .A1(n5736), .A2(n5734), .A3(n5765), .ZN(n5548) );
  NAND3_X1 U10037 ( .A1(n5546), .A2(n5735), .A3(n5545), .ZN(n5547) );
  XNOR2_X1 U10039 ( .A(n7155), .B(n2222), .ZN(n5550) );
  XNOR2_X1 U10040 ( .A(n5551), .B(n5550), .ZN(n5552) );
  XNOR2_X1 U10041 ( .A(n5553), .B(n5552), .ZN(n8033) );
  OAI21_X1 U10042 ( .B1(n7600), .B2(n8033), .A(n7445), .ZN(n5554) );
  INV_X1 U10043 ( .A(n8286), .ZN(n7444) );
  NAND2_X1 U10044 ( .A1(n5554), .A2(n7444), .ZN(n5555) );
  OAI21_X1 U10045 ( .B1(n7796), .B2(n8034), .A(n5555), .ZN(n5556) );
  NAND2_X1 U10047 ( .A1(n5562), .A2(n6036), .ZN(n5570) );
  OAI21_X1 U10048 ( .B1(n5564), .B2(n20241), .A(n5569), .ZN(n5567) );
  MUX2_X1 U10049 ( .A(n5567), .B(n5566), .S(n5565), .Z(n5568) );
  XNOR2_X1 U10050 ( .A(n7080), .B(n7287), .ZN(n6759) );
  NAND2_X1 U10051 ( .A1(n5572), .A2(n5571), .ZN(n5586) );
  INV_X1 U10052 ( .A(n5573), .ZN(n5578) );
  NAND3_X1 U10053 ( .A1(n5576), .A2(n5575), .A3(n5574), .ZN(n5577) );
  OAI21_X1 U10054 ( .B1(n5578), .B2(n5577), .A(n5580), .ZN(n5579) );
  OAI21_X1 U10055 ( .B1(n5581), .B2(n5580), .A(n5579), .ZN(n5585) );
  XNOR2_X1 U10056 ( .A(n5884), .B(n19158), .ZN(n5587) );
  XNOR2_X1 U10057 ( .A(n6759), .B(n5587), .ZN(n5601) );
  NAND2_X1 U10059 ( .A1(n20368), .A2(n5588), .ZN(n5594) );
  NOR2_X1 U10060 ( .A1(n5920), .A2(n19980), .ZN(n5593) );
  NAND3_X1 U10061 ( .A1(n5916), .A2(n6007), .A3(n19980), .ZN(n5592) );
  INV_X1 U10062 ( .A(n7115), .ZN(n5598) );
  INV_X1 U10063 ( .A(n5927), .ZN(n5595) );
  XNOR2_X1 U10064 ( .A(n5598), .B(n6819), .ZN(n7285) );
  XNOR2_X1 U10065 ( .A(n7285), .B(n5599), .ZN(n5600) );
  XNOR2_X1 U10066 ( .A(n5600), .B(n5601), .ZN(n7420) );
  NAND2_X1 U10067 ( .A1(n5602), .A2(n5720), .ZN(n5609) );
  INV_X1 U10068 ( .A(n5603), .ZN(n5608) );
  NAND3_X1 U10069 ( .A1(n20034), .A2(n5715), .A3(n5483), .ZN(n5606) );
  XNOR2_X1 U10072 ( .A(n6558), .B(n7297), .ZN(n6526) );
  INV_X1 U10073 ( .A(n6526), .ZN(n6774) );
  NAND2_X1 U10075 ( .A1(n5615), .A2(n6140), .ZN(n5619) );
  NAND2_X1 U10076 ( .A1(n6138), .A2(n5859), .ZN(n5616) );
  NAND2_X1 U10077 ( .A1(n5617), .A2(n6143), .ZN(n5618) );
  INV_X1 U10078 ( .A(n6133), .ZN(n6130) );
  AOI22_X1 U10079 ( .A1(n5623), .A2(n5622), .B1(n6130), .B2(n5691), .ZN(n5693)
         );
  INV_X1 U10080 ( .A(n6131), .ZN(n5626) );
  OAI21_X1 U10081 ( .B1(n5624), .B2(n5621), .A(n6133), .ZN(n5625) );
  OAI21_X1 U10082 ( .B1(n5693), .B2(n5626), .A(n5625), .ZN(n6855) );
  XNOR2_X1 U10083 ( .A(n6855), .B(n6713), .ZN(n7295) );
  XNOR2_X1 U10084 ( .A(n6774), .B(n7295), .ZN(n5639) );
  NAND3_X1 U10085 ( .A1(n5631), .A2(n4598), .A3(n5633), .ZN(n5627) );
  OAI21_X1 U10086 ( .B1(n5629), .B2(n5628), .A(n5627), .ZN(n5636) );
  AOI21_X1 U10087 ( .B1(n5634), .B2(n5633), .A(n5632), .ZN(n5635) );
  INV_X1 U10088 ( .A(n6301), .ZN(n6936) );
  XNOR2_X1 U10089 ( .A(n6936), .B(n404), .ZN(n5637) );
  XNOR2_X1 U10090 ( .A(n6488), .B(n5637), .ZN(n5638) );
  INV_X1 U10091 ( .A(n5640), .ZN(n5654) );
  INV_X1 U10092 ( .A(n5641), .ZN(n5644) );
  OAI21_X1 U10093 ( .B1(n5644), .B2(n5643), .A(n5642), .ZN(n5653) );
  NAND3_X1 U10094 ( .A1(n5647), .A2(n5646), .A3(n5645), .ZN(n5652) );
  NAND2_X1 U10096 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  XNOR2_X1 U10098 ( .A(n6912), .B(n18203), .ZN(n5655) );
  XNOR2_X1 U10099 ( .A(n6495), .B(n5655), .ZN(n5689) );
  OAI21_X1 U10100 ( .B1(n284), .B2(n6101), .A(n5662), .ZN(n5666) );
  NAND2_X1 U10101 ( .A1(n6097), .A2(n5949), .ZN(n6096) );
  XNOR2_X1 U10103 ( .A(n6966), .B(n6735), .ZN(n7323) );
  NOR2_X1 U10104 ( .A1(n5424), .A2(n5669), .ZN(n5671) );
  OAI22_X1 U10106 ( .A1(n5677), .A2(n5676), .B1(n3127), .B2(n5674), .ZN(n5678)
         );
  OAI21_X1 U10108 ( .B1(n5681), .B2(n6082), .A(n5680), .ZN(n5687) );
  NAND3_X1 U10109 ( .A1(n5684), .A2(n6082), .A3(n6083), .ZN(n5685) );
  XNOR2_X1 U10110 ( .A(n19765), .B(n19698), .ZN(n6752) );
  XNOR2_X1 U10111 ( .A(n7323), .B(n6752), .ZN(n5688) );
  XNOR2_X1 U10112 ( .A(n5689), .B(n5688), .ZN(n5762) );
  NOR2_X1 U10113 ( .A1(n5691), .A2(n6131), .ZN(n5695) );
  NAND2_X1 U10114 ( .A1(n5698), .A2(n5970), .ZN(n5702) );
  INV_X1 U10115 ( .A(n5699), .ZN(n5972) );
  OAI211_X1 U10116 ( .C1(n5973), .C2(n5967), .A(n5972), .B(n5700), .ZN(n5701)
         );
  INV_X1 U10117 ( .A(n7332), .ZN(n5703) );
  XNOR2_X1 U10118 ( .A(n5703), .B(n7097), .ZN(n6534) );
  INV_X1 U10119 ( .A(n5813), .ZN(n5706) );
  AOI22_X1 U10120 ( .A1(n5707), .A2(n6003), .B1(n5706), .B2(n5705), .ZN(n7133)
         );
  INV_X1 U10121 ( .A(n7133), .ZN(n6512) );
  NAND2_X1 U10122 ( .A1(n5708), .A2(n5989), .ZN(n5713) );
  OAI21_X1 U10123 ( .B1(n5985), .B2(n5990), .A(n3468), .ZN(n5710) );
  NAND3_X1 U10124 ( .A1(n5276), .A2(n5711), .A3(n5990), .ZN(n5712) );
  INV_X1 U10125 ( .A(n6872), .ZN(n6811) );
  NAND3_X1 U10126 ( .A1(n5718), .A2(n5717), .A3(n5720), .ZN(n5723) );
  NAND2_X1 U10127 ( .A1(n5719), .A2(n5720), .ZN(n5721) );
  XNOR2_X1 U10128 ( .A(n6917), .B(n17637), .ZN(n5725) );
  XNOR2_X1 U10129 ( .A(n7334), .B(n5725), .ZN(n5726) );
  NOR2_X1 U10130 ( .A1(n8205), .A2(n8204), .ZN(n5760) );
  MUX2_X1 U10131 ( .A(n6379), .B(n5728), .S(n19475), .Z(n5729) );
  NOR2_X1 U10132 ( .A1(n5729), .A2(n6183), .ZN(n5731) );
  NAND2_X1 U10133 ( .A1(n6192), .A2(n6189), .ZN(n5732) );
  INV_X1 U10134 ( .A(n5736), .ZN(n5770) );
  AND2_X1 U10136 ( .A1(n5765), .A2(n5768), .ZN(n5764) );
  NAND2_X1 U10137 ( .A1(n5764), .A2(n5766), .ZN(n5739) );
  XNOR2_X1 U10139 ( .A(n6767), .B(n17089), .ZN(n5754) );
  NAND2_X1 U10140 ( .A1(n5742), .A2(n5741), .ZN(n5753) );
  NAND2_X1 U10141 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  MUX2_X1 U10142 ( .A(n5226), .B(n6204), .S(n6206), .Z(n5757) );
  NOR2_X1 U10143 ( .A1(n6202), .A2(n19492), .ZN(n5756) );
  NAND2_X1 U10144 ( .A1(n6218), .A2(n19968), .ZN(n5758) );
  INV_X1 U10145 ( .A(n5762), .ZN(n7871) );
  NAND2_X1 U10146 ( .A1(n5764), .A2(n5763), .ZN(n5774) );
  NAND2_X1 U10147 ( .A1(n5766), .A2(n5765), .ZN(n5773) );
  NAND3_X1 U10148 ( .A1(n5769), .A2(n5546), .A3(n5767), .ZN(n5772) );
  NAND3_X1 U10149 ( .A1(n5770), .A2(n5769), .A3(n5768), .ZN(n5771) );
  XNOR2_X1 U10150 ( .A(n6927), .B(n19140), .ZN(n5775) );
  XNOR2_X1 U10151 ( .A(n6506), .B(n5775), .ZN(n5812) );
  NAND2_X1 U10152 ( .A1(n6041), .A2(n6042), .ZN(n5778) );
  NAND3_X1 U10153 ( .A1(n6046), .A2(n6041), .A3(n5888), .ZN(n5780) );
  NAND2_X1 U10154 ( .A1(n6059), .A2(n5782), .ZN(n5783) );
  OAI21_X1 U10155 ( .B1(n6064), .B2(n6059), .A(n5783), .ZN(n5784) );
  NAND2_X1 U10156 ( .A1(n5784), .A2(n5891), .ZN(n5789) );
  NOR2_X1 U10157 ( .A1(n6057), .A2(n6055), .ZN(n5787) );
  INV_X1 U10158 ( .A(n6059), .ZN(n5786) );
  AOI22_X1 U10159 ( .A1(n5787), .A2(n5786), .B1(n5785), .B2(n6055), .ZN(n5788)
         );
  NAND2_X1 U10160 ( .A1(n5789), .A2(n5788), .ZN(n6723) );
  XNOR2_X1 U10161 ( .A(n6839), .B(n6723), .ZN(n7313) );
  AND2_X1 U10162 ( .A1(n5794), .A2(n5793), .ZN(n5801) );
  MUX2_X1 U10163 ( .A(n5797), .B(n5796), .S(n19912), .Z(n5799) );
  NAND2_X1 U10164 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  NAND2_X1 U10165 ( .A1(n5801), .A2(n5800), .ZN(n7317) );
  INV_X1 U10166 ( .A(n5803), .ZN(n5806) );
  NOR2_X1 U10167 ( .A1(n5806), .A2(n5805), .ZN(n5810) );
  OAI21_X1 U10168 ( .B1(n5803), .B2(n5802), .A(n6194), .ZN(n5809) );
  NAND3_X1 U10169 ( .A1(n6193), .A2(n5806), .A3(n6189), .ZN(n5807) );
  OAI211_X2 U10170 ( .C1(n5809), .C2(n5810), .A(n5808), .B(n5807), .ZN(n7091)
         );
  XNOR2_X1 U10171 ( .A(n7317), .B(n7091), .ZN(n6790) );
  XNOR2_X1 U10172 ( .A(n6790), .B(n7313), .ZN(n5811) );
  XNOR2_X1 U10173 ( .A(n5812), .B(n5811), .ZN(n7615) );
  INV_X1 U10174 ( .A(n5997), .ZN(n5999) );
  NAND2_X1 U10175 ( .A1(n5816), .A2(n5986), .ZN(n5821) );
  NAND3_X1 U10176 ( .A1(n5818), .A2(n285), .A3(n5817), .ZN(n5819) );
  OAI211_X1 U10177 ( .C1(n5988), .C2(n5821), .A(n5820), .B(n5819), .ZN(n6754)
         );
  XNOR2_X1 U10178 ( .A(n7231), .B(n6754), .ZN(n6268) );
  INV_X1 U10179 ( .A(n6268), .ZN(n6603) );
  XNOR2_X1 U10180 ( .A(n19765), .B(n7364), .ZN(n5822) );
  XNOR2_X1 U10181 ( .A(n6603), .B(n5822), .ZN(n5834) );
  NOR2_X1 U10182 ( .A1(n3569), .A2(n5823), .ZN(n6018) );
  AND2_X1 U10183 ( .A1(n5825), .A2(n6016), .ZN(n6020) );
  NAND2_X1 U10184 ( .A1(n6020), .A2(n6022), .ZN(n5830) );
  XNOR2_X1 U10185 ( .A(n6912), .B(n7154), .ZN(n6676) );
  XNOR2_X1 U10186 ( .A(n7035), .B(n2284), .ZN(n5832) );
  XNOR2_X1 U10187 ( .A(n6676), .B(n5832), .ZN(n5833) );
  XNOR2_X1 U10188 ( .A(n5833), .B(n5834), .ZN(n7453) );
  OAI21_X1 U10189 ( .B1(n5226), .B2(n19968), .A(n6204), .ZN(n5837) );
  OAI21_X1 U10190 ( .B1(n5839), .B2(n5838), .A(n5837), .ZN(n5840) );
  OAI21_X1 U10191 ( .B1(n5846), .B2(n5845), .A(n6184), .ZN(n5849) );
  XNOR2_X1 U10192 ( .A(n6680), .B(n7091), .ZN(n5852) );
  XNOR2_X1 U10193 ( .A(n6985), .B(n19243), .ZN(n5851) );
  XNOR2_X1 U10194 ( .A(n5852), .B(n5851), .ZN(n5853) );
  NAND2_X1 U10195 ( .A1(n7453), .A2(n8040), .ZN(n7788) );
  INV_X1 U10197 ( .A(n5856), .ZN(n5857) );
  XNOR2_X1 U10198 ( .A(n19780), .B(n6917), .ZN(n6686) );
  XNOR2_X1 U10199 ( .A(n7097), .B(n6808), .ZN(n5858) );
  XNOR2_X1 U10200 ( .A(n6686), .B(n5858), .ZN(n5878) );
  NAND2_X1 U10201 ( .A1(n6143), .A2(n5860), .ZN(n5863) );
  NAND2_X1 U10202 ( .A1(n5861), .A2(n6141), .ZN(n5862) );
  OAI21_X1 U10203 ( .B1(n5864), .B2(n5863), .A(n5862), .ZN(n5865) );
  INV_X1 U10204 ( .A(n5867), .ZN(n5874) );
  NAND3_X1 U10205 ( .A1(n5870), .A2(n5869), .A3(n5868), .ZN(n5872) );
  NAND2_X1 U10206 ( .A1(n6124), .A2(n5873), .ZN(n5871) );
  XNOR2_X1 U10207 ( .A(n6249), .B(n6786), .ZN(n6598) );
  INV_X1 U10208 ( .A(n2306), .ZN(n5875) );
  XNOR2_X1 U10209 ( .A(n7041), .B(n5875), .ZN(n5876) );
  XNOR2_X1 U10210 ( .A(n6598), .B(n5876), .ZN(n5877) );
  XNOR2_X1 U10211 ( .A(n5878), .B(n5877), .ZN(n8041) );
  INV_X1 U10212 ( .A(n8041), .ZN(n8298) );
  NOR2_X1 U10213 ( .A1(n6068), .A2(n6067), .ZN(n5881) );
  NOR2_X2 U10214 ( .A1(n5883), .A2(n5882), .ZN(n7118) );
  NAND3_X1 U10215 ( .A1(n6044), .A2(n1007), .A3(n5885), .ZN(n5886) );
  OAI21_X1 U10216 ( .B1(n6041), .B2(n6044), .A(n5886), .ZN(n5887) );
  INV_X1 U10217 ( .A(n5887), .ZN(n5890) );
  XNOR2_X1 U10219 ( .A(n6761), .B(n7258), .ZN(n6588) );
  XNOR2_X1 U10220 ( .A(n7080), .B(n7253), .ZN(n5897) );
  XNOR2_X1 U10221 ( .A(n6977), .B(n2347), .ZN(n5896) );
  XNOR2_X1 U10222 ( .A(n5897), .B(n5896), .ZN(n5898) );
  INV_X1 U10223 ( .A(n6942), .ZN(n5913) );
  NAND2_X1 U10224 ( .A1(n5900), .A2(n5899), .ZN(n6091) );
  NOR2_X1 U10225 ( .A1(n5902), .A2(n5901), .ZN(n5906) );
  NAND4_X1 U10226 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n5907)
         );
  OAI21_X1 U10227 ( .B1(n5199), .B2(n6087), .A(n5907), .ZN(n5909) );
  NAND2_X1 U10228 ( .A1(n5909), .A2(n5908), .ZN(n5911) );
  NAND3_X1 U10229 ( .A1(n20149), .A2(n5199), .A3(n890), .ZN(n5910) );
  OAI211_X1 U10230 ( .C1(n5912), .C2(n6091), .A(n5911), .B(n5910), .ZN(n7164)
         );
  XNOR2_X1 U10231 ( .A(n5913), .B(n7164), .ZN(n6692) );
  OAI21_X1 U10233 ( .B1(n5914), .B2(n861), .A(n5915), .ZN(n5918) );
  NAND2_X1 U10234 ( .A1(n5918), .A2(n5917), .ZN(n5925) );
  NAND3_X1 U10235 ( .A1(n5919), .A2(n6007), .A3(n6013), .ZN(n5923) );
  NAND3_X1 U10236 ( .A1(n5921), .A2(n6010), .A3(n862), .ZN(n5922) );
  AND2_X1 U10237 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  NAND2_X1 U10238 ( .A1(n5925), .A2(n5924), .ZN(n6946) );
  OAI21_X1 U10239 ( .B1(n5595), .B2(n19790), .A(n5926), .ZN(n5935) );
  NOR2_X1 U10240 ( .A1(n5927), .A2(n5930), .ZN(n5934) );
  XNOR2_X1 U10241 ( .A(n6946), .B(n6768), .ZN(n6611) );
  INV_X1 U10242 ( .A(n6611), .ZN(n5936) );
  XNOR2_X1 U10243 ( .A(n6692), .B(n5936), .ZN(n5940) );
  XNOR2_X1 U10244 ( .A(n6348), .B(n7267), .ZN(n5938) );
  XNOR2_X1 U10245 ( .A(n20225), .B(n17686), .ZN(n5937) );
  XNOR2_X1 U10246 ( .A(n5938), .B(n5937), .ZN(n5939) );
  INV_X1 U10247 ( .A(n7787), .ZN(n5963) );
  INV_X1 U10248 ( .A(n6166), .ZN(n5942) );
  AOI21_X1 U10249 ( .B1(n5943), .B2(n6175), .A(n5942), .ZN(n5947) );
  NAND2_X1 U10250 ( .A1(n6176), .A2(n6171), .ZN(n5944) );
  AOI21_X1 U10251 ( .B1(n5945), .B2(n5944), .A(n6168), .ZN(n5946) );
  XNOR2_X1 U10252 ( .A(n7127), .B(n6936), .ZN(n6665) );
  INV_X1 U10253 ( .A(n5948), .ZN(n5951) );
  XNOR2_X1 U10254 ( .A(n7240), .B(n941), .ZN(n6606) );
  XNOR2_X1 U10255 ( .A(n6665), .B(n6606), .ZN(n5962) );
  INV_X1 U10256 ( .A(n7392), .ZN(n5958) );
  XNOR2_X1 U10257 ( .A(n7014), .B(n5958), .ZN(n5960) );
  XNOR2_X1 U10258 ( .A(n6558), .B(n2401), .ZN(n5959) );
  XNOR2_X1 U10259 ( .A(n5960), .B(n5959), .ZN(n5961) );
  AND2_X1 U10262 ( .A1(n5967), .A2(n5971), .ZN(n5969) );
  INV_X1 U10263 ( .A(n5973), .ZN(n5974) );
  NAND2_X1 U10264 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  XNOR2_X1 U10265 ( .A(n7372), .B(n7142), .ZN(n6721) );
  INV_X1 U10266 ( .A(n6721), .ZN(n5983) );
  NAND2_X1 U10267 ( .A1(n209), .A2(n5978), .ZN(n5979) );
  AOI22_X1 U10268 ( .A1(n5980), .A2(n6069), .B1(n6072), .B2(n6067), .ZN(n5981)
         );
  XNOR2_X1 U10269 ( .A(n7047), .B(n7088), .ZN(n7315) );
  XNOR2_X1 U10270 ( .A(n7315), .B(n5983), .ZN(n6006) );
  XNOR2_X1 U10271 ( .A(n7272), .B(n2410), .ZN(n6004) );
  AND2_X1 U10272 ( .A1(n5985), .A2(n5989), .ZN(n5987) );
  OAI21_X1 U10273 ( .B1(n5988), .B2(n5987), .A(n5986), .ZN(n5994) );
  INV_X1 U10274 ( .A(n5989), .ZN(n5991) );
  NAND3_X1 U10275 ( .A1(n5991), .A2(n285), .A3(n5990), .ZN(n5992) );
  NAND3_X1 U10276 ( .A1(n6000), .A2(n5999), .A3(n5998), .ZN(n6001) );
  INV_X1 U10277 ( .A(n6328), .ZN(n7177) );
  XNOR2_X1 U10278 ( .A(n7177), .B(n6004), .ZN(n6005) );
  OAI211_X1 U10279 ( .C1(n6010), .C2(n19980), .A(n20368), .B(n6007), .ZN(n6012) );
  INV_X1 U10280 ( .A(n2349), .ZN(n6015) );
  XNOR2_X1 U10281 ( .A(n6990), .B(n6015), .ZN(n6024) );
  AOI21_X1 U10282 ( .B1(n3569), .B2(n6017), .A(n6016), .ZN(n6021) );
  INV_X1 U10283 ( .A(n6021), .ZN(n6023) );
  OAI211_X1 U10285 ( .C1(n6027), .C2(n19789), .A(n5595), .B(n6025), .ZN(n6029)
         );
  XNOR2_X1 U10286 ( .A(n6782), .B(n7042), .ZN(n6032) );
  XNOR2_X1 U10287 ( .A(n7382), .B(n7336), .ZN(n6039) );
  XNOR2_X1 U10288 ( .A(n6039), .B(n6038), .ZN(n6732) );
  NAND2_X1 U10289 ( .A1(n6043), .A2(n6042), .ZN(n6045) );
  AOI22_X2 U10290 ( .A1(n6047), .A2(n6046), .B1(n6045), .B2(n6044), .ZN(n6997)
         );
  XNOR2_X1 U10292 ( .A(n6997), .B(n7018), .ZN(n7193) );
  INV_X1 U10293 ( .A(n7193), .ZN(n6066) );
  AOI21_X1 U10294 ( .B1(n6056), .B2(n5782), .A(n6058), .ZN(n6063) );
  NOR2_X1 U10295 ( .A1(n6058), .A2(n6057), .ZN(n6060) );
  XNOR2_X1 U10296 ( .A(n7017), .B(n6708), .ZN(n7294) );
  INV_X1 U10297 ( .A(n7294), .ZN(n6065) );
  XNOR2_X1 U10298 ( .A(n6065), .B(n6066), .ZN(n6079) );
  XNOR2_X1 U10299 ( .A(n6707), .B(n7391), .ZN(n6077) );
  XNOR2_X1 U10300 ( .A(n6777), .B(n1148), .ZN(n6076) );
  XNOR2_X1 U10301 ( .A(n6077), .B(n6076), .ZN(n6078) );
  NAND2_X1 U10302 ( .A1(n6081), .A2(n6080), .ZN(n6086) );
  MUX2_X1 U10303 ( .A(n6084), .B(n6083), .S(n6082), .Z(n6085) );
  NAND2_X1 U10305 ( .A1(n890), .A2(n6087), .ZN(n6088) );
  NAND3_X1 U10306 ( .A1(n6093), .A2(n6092), .A3(n6091), .ZN(n6094) );
  XNOR2_X1 U10307 ( .A(n6095), .B(n6718), .ZN(n6116) );
  OAI21_X1 U10308 ( .B1(n6098), .B2(n6097), .A(n6096), .ZN(n6103) );
  NAND2_X1 U10309 ( .A1(n6100), .A2(n6099), .ZN(n6102) );
  MUX2_X1 U10310 ( .A(n6105), .B(n6104), .S(n6109), .Z(n6106) );
  INV_X1 U10311 ( .A(n6106), .ZN(n6112) );
  XNOR2_X1 U10312 ( .A(n7218), .B(n7221), .ZN(n6337) );
  XNOR2_X1 U10313 ( .A(n7257), .B(n2368), .ZN(n6114) );
  XNOR2_X1 U10314 ( .A(n6337), .B(n6114), .ZN(n6115) );
  NAND2_X1 U10315 ( .A1(n8196), .A2(n20198), .ZN(n7628) );
  NOR2_X1 U10316 ( .A1(n6119), .A2(n6118), .ZN(n6121) );
  OAI21_X1 U10317 ( .B1(n6122), .B2(n6121), .A(n6120), .ZN(n6126) );
  NAND3_X1 U10318 ( .A1(n6124), .A2(n6128), .A3(n6123), .ZN(n6125) );
  OAI211_X1 U10319 ( .C1(n6128), .C2(n6127), .A(n6126), .B(n6125), .ZN(n7009)
         );
  XNOR2_X1 U10320 ( .A(n7009), .B(n6745), .ZN(n7308) );
  MUX2_X1 U10321 ( .A(n6130), .B(n6132), .S(n6129), .Z(n6137) );
  NAND2_X1 U10322 ( .A1(n6132), .A2(n6131), .ZN(n6135) );
  MUX2_X1 U10323 ( .A(n6135), .B(n6134), .S(n6133), .Z(n6136) );
  OAI21_X2 U10324 ( .B1(n6137), .B2(n5621), .A(n6136), .ZN(n7007) );
  MUX2_X1 U10325 ( .A(n6139), .B(n6141), .S(n6138), .Z(n6147) );
  NAND2_X1 U10326 ( .A1(n6141), .A2(n6140), .ZN(n6145) );
  NAND2_X1 U10327 ( .A1(n6148), .A2(n20334), .ZN(n6144) );
  MUX2_X1 U10328 ( .A(n6145), .B(n6144), .S(n6143), .Z(n6146) );
  XNOR2_X1 U10329 ( .A(n7007), .B(n7206), .ZN(n6349) );
  XNOR2_X1 U10330 ( .A(n6349), .B(n7308), .ZN(n6164) );
  NAND3_X1 U10331 ( .A1(n6151), .A2(n6150), .A3(n6149), .ZN(n6158) );
  OAI211_X1 U10332 ( .C1(n6156), .C2(n6155), .A(n6154), .B(n6153), .ZN(n6157)
         );
  INV_X1 U10334 ( .A(n2445), .ZN(n6161) );
  XNOR2_X1 U10335 ( .A(n7263), .B(n6161), .ZN(n6162) );
  XNOR2_X1 U10336 ( .A(n6744), .B(n6162), .ZN(n6163) );
  XNOR2_X1 U10337 ( .A(n6164), .B(n6163), .ZN(n8192) );
  INV_X1 U10338 ( .A(n6165), .ZN(n6180) );
  NAND2_X1 U10339 ( .A1(n6167), .A2(n6171), .ZN(n6169) );
  MUX2_X1 U10340 ( .A(n6170), .B(n6169), .S(n6168), .Z(n6179) );
  NOR2_X1 U10341 ( .A1(n6172), .A2(n6171), .ZN(n6174) );
  NAND2_X1 U10342 ( .A1(n6174), .A2(n6173), .ZN(n6178) );
  XNOR2_X1 U10343 ( .A(n6180), .B(n7032), .ZN(n7324) );
  INV_X1 U10344 ( .A(n7324), .ZN(n6546) );
  NOR2_X1 U10345 ( .A1(n6379), .A2(n288), .ZN(n6181) );
  OAI21_X1 U10346 ( .B1(n6380), .B2(n6184), .A(n6183), .ZN(n6185) );
  NOR2_X1 U10347 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  MUX2_X1 U10349 ( .A(n6191), .B(n6190), .S(n6189), .Z(n6198) );
  NAND2_X1 U10350 ( .A1(n6193), .A2(n6192), .ZN(n6196) );
  XNOR2_X1 U10352 ( .A(n19778), .B(n7031), .ZN(n6199) );
  XNOR2_X1 U10353 ( .A(n6546), .B(n6199), .ZN(n6210) );
  XNOR2_X1 U10354 ( .A(n7230), .B(n484), .ZN(n6209) );
  NAND2_X1 U10355 ( .A1(n6218), .A2(n19492), .ZN(n6201) );
  NAND2_X1 U10356 ( .A1(n6220), .A2(n6204), .ZN(n6208) );
  NOR2_X1 U10357 ( .A1(n6206), .A2(n6205), .ZN(n6219) );
  NAND2_X1 U10358 ( .A1(n6219), .A2(n6218), .ZN(n6207) );
  XNOR2_X1 U10359 ( .A(n6970), .B(n7155), .ZN(n6737) );
  NAND3_X1 U10361 ( .A1(n9238), .A2(n9233), .A3(n8708), .ZN(n6213) );
  XNOR2_X1 U10362 ( .A(n9819), .B(n17791), .ZN(n6658) );
  XNOR2_X1 U10363 ( .A(n7151), .B(n19840), .ZN(n6911) );
  XNOR2_X1 U10364 ( .A(n6165), .B(n17791), .ZN(n6216) );
  XNOR2_X1 U10365 ( .A(n6911), .B(n6216), .ZN(n6224) );
  XNOR2_X1 U10366 ( .A(n6736), .B(n7360), .ZN(n6222) );
  XNOR2_X1 U10367 ( .A(n6420), .B(n19764), .ZN(n7058) );
  XNOR2_X1 U10368 ( .A(n7058), .B(n6222), .ZN(n6223) );
  XNOR2_X1 U10369 ( .A(n20224), .B(n6745), .ZN(n7073) );
  XNOR2_X1 U10370 ( .A(n6225), .B(n7073), .ZN(n6228) );
  INV_X1 U10371 ( .A(n7160), .ZN(n6226) );
  XNOR2_X1 U10372 ( .A(n6228), .B(n6227), .ZN(n7931) );
  XNOR2_X1 U10373 ( .A(n7080), .B(n7354), .ZN(n6565) );
  XNOR2_X1 U10374 ( .A(n6565), .B(n19847), .ZN(n6233) );
  XNOR2_X1 U10375 ( .A(n6719), .B(n7121), .ZN(n6231) );
  XNOR2_X1 U10376 ( .A(n7258), .B(n18006), .ZN(n6230) );
  XNOR2_X1 U10377 ( .A(n6231), .B(n6230), .ZN(n6232) );
  INV_X1 U10378 ( .A(n7372), .ZN(n6234) );
  XNOR2_X1 U10379 ( .A(n7088), .B(n6234), .ZN(n6236) );
  XNOR2_X1 U10380 ( .A(n7091), .B(n17932), .ZN(n6235) );
  XNOR2_X1 U10381 ( .A(n6236), .B(n6235), .ZN(n6239) );
  XNOR2_X1 U10382 ( .A(n7146), .B(n7274), .ZN(n6925) );
  XNOR2_X1 U10383 ( .A(n6237), .B(n6925), .ZN(n6238) );
  INV_X1 U10384 ( .A(n7936), .ZN(n7933) );
  XNOR2_X1 U10385 ( .A(n7240), .B(n7128), .ZN(n6935) );
  XNOR2_X1 U10386 ( .A(n6935), .B(n6640), .ZN(n6243) );
  XNOR2_X1 U10387 ( .A(n6558), .B(n6708), .ZN(n7066) );
  INV_X1 U10388 ( .A(n7066), .ZN(n6241) );
  XNOR2_X1 U10389 ( .A(n7391), .B(n18304), .ZN(n6240) );
  XNOR2_X1 U10390 ( .A(n6241), .B(n6240), .ZN(n6242) );
  XNOR2_X1 U10391 ( .A(n6687), .B(n649), .ZN(n6246) );
  INV_X1 U10392 ( .A(n7097), .ZN(n6783) );
  XNOR2_X1 U10393 ( .A(n6246), .B(n6783), .ZN(n6248) );
  XNOR2_X1 U10394 ( .A(n6728), .B(n7382), .ZN(n6247) );
  XNOR2_X1 U10395 ( .A(n6248), .B(n6247), .ZN(n6252) );
  XNOR2_X1 U10396 ( .A(n943), .B(n7336), .ZN(n6250) );
  XNOR2_X1 U10397 ( .A(n6250), .B(n7134), .ZN(n6251) );
  XNOR2_X1 U10398 ( .A(n6252), .B(n6251), .ZN(n7763) );
  NOR2_X1 U10399 ( .A1(n7930), .A2(n1063), .ZN(n6438) );
  INV_X1 U10400 ( .A(n7297), .ZN(n6253) );
  XNOR2_X1 U10401 ( .A(n941), .B(n6253), .ZN(n6255) );
  XNOR2_X1 U10403 ( .A(n6777), .B(n16788), .ZN(n6254) );
  XNOR2_X1 U10404 ( .A(n6255), .B(n6254), .ZN(n6258) );
  XNOR2_X1 U10405 ( .A(n7240), .B(n6641), .ZN(n6256) );
  XNOR2_X1 U10406 ( .A(n7127), .B(n6854), .ZN(n6398) );
  XNOR2_X1 U10407 ( .A(n6256), .B(n6398), .ZN(n6257) );
  XNOR2_X2 U10408 ( .A(n6257), .B(n6258), .ZN(n7903) );
  XNOR2_X1 U10409 ( .A(n6611), .B(n7305), .ZN(n6262) );
  XNOR2_X1 U10410 ( .A(n7263), .B(Key[63]), .ZN(n6259) );
  XNOR2_X1 U10411 ( .A(n6259), .B(n6945), .ZN(n6260) );
  XNOR2_X1 U10412 ( .A(n7164), .B(n6850), .ZN(n6393) );
  XNOR2_X1 U10413 ( .A(n6260), .B(n6393), .ZN(n6261) );
  XNOR2_X1 U10414 ( .A(n6261), .B(n6262), .ZN(n7530) );
  XNOR2_X1 U10415 ( .A(n7332), .B(n2216), .ZN(n6263) );
  XNOR2_X1 U10416 ( .A(n6263), .B(n6598), .ZN(n6266) );
  XNOR2_X1 U10417 ( .A(n6782), .B(n6919), .ZN(n7247) );
  XNOR2_X1 U10418 ( .A(n6873), .B(n7137), .ZN(n6368) );
  INV_X1 U10419 ( .A(n6368), .ZN(n6264) );
  XNOR2_X1 U10420 ( .A(n6264), .B(n7247), .ZN(n6265) );
  XNOR2_X1 U10421 ( .A(n6265), .B(n6266), .ZN(n6904) );
  INV_X1 U10422 ( .A(n6904), .ZN(n7902) );
  INV_X1 U10423 ( .A(n6494), .ZN(n6545) );
  XNOR2_X1 U10424 ( .A(n6545), .B(n7230), .ZN(n6267) );
  XNOR2_X1 U10425 ( .A(n6268), .B(n6267), .ZN(n6271) );
  XNOR2_X1 U10426 ( .A(n19699), .B(n18338), .ZN(n6269) );
  XNOR2_X1 U10427 ( .A(n7154), .B(n7365), .ZN(n6364) );
  XNOR2_X1 U10428 ( .A(n6269), .B(n6364), .ZN(n6270) );
  XNOR2_X1 U10429 ( .A(n6271), .B(n6270), .ZN(n7002) );
  BUF_X2 U10430 ( .A(n7002), .Z(n7909) );
  NOR2_X1 U10431 ( .A1(n7902), .A2(n7909), .ZN(n6272) );
  XNOR2_X1 U10432 ( .A(n7272), .B(n7317), .ZN(n6274) );
  XNOR2_X1 U10433 ( .A(n6634), .B(n18011), .ZN(n6273) );
  XNOR2_X1 U10434 ( .A(n6274), .B(n6273), .ZN(n6276) );
  XNOR2_X1 U10435 ( .A(n6593), .B(n6374), .ZN(n6275) );
  XNOR2_X1 U10436 ( .A(n6276), .B(n6275), .ZN(n7908) );
  INV_X1 U10437 ( .A(n7118), .ZN(n6384) );
  XNOR2_X1 U10438 ( .A(n6384), .B(n6520), .ZN(n6277) );
  XNOR2_X1 U10439 ( .A(n6277), .B(n6588), .ZN(n6282) );
  INV_X1 U10440 ( .A(n7257), .ZN(n6278) );
  XNOR2_X1 U10441 ( .A(n6278), .B(n1053), .ZN(n6280) );
  XNOR2_X1 U10442 ( .A(n19730), .B(n17587), .ZN(n6279) );
  XNOR2_X1 U10443 ( .A(n6280), .B(n6279), .ZN(n6281) );
  NAND2_X1 U10444 ( .A1(n7754), .A2(n7903), .ZN(n6283) );
  XNOR2_X1 U10445 ( .A(n5884), .B(n6477), .ZN(n7356) );
  XNOR2_X1 U10446 ( .A(n7254), .B(n7289), .ZN(n7078) );
  XNOR2_X1 U10447 ( .A(n7356), .B(n7078), .ZN(n6289) );
  INV_X1 U10448 ( .A(n6285), .ZN(n6661) );
  XNOR2_X1 U10449 ( .A(n6661), .B(n7216), .ZN(n6287) );
  XNOR2_X1 U10450 ( .A(n19730), .B(n2423), .ZN(n6286) );
  XNOR2_X1 U10451 ( .A(n6287), .B(n6286), .ZN(n6288) );
  XNOR2_X1 U10452 ( .A(n6289), .B(n6288), .ZN(n7919) );
  XNOR2_X1 U10454 ( .A(n6942), .B(n6693), .ZN(n7346) );
  XNOR2_X1 U10455 ( .A(n6850), .B(n6947), .ZN(n6446) );
  XNOR2_X1 U10456 ( .A(n7346), .B(n6446), .ZN(n6292) );
  XNOR2_X1 U10457 ( .A(n7201), .B(n7266), .ZN(n6346) );
  XNOR2_X1 U10458 ( .A(n7306), .B(n2375), .ZN(n6290) );
  XNOR2_X1 U10459 ( .A(n6346), .B(n6290), .ZN(n6291) );
  XNOR2_X1 U10460 ( .A(n6362), .B(n6912), .ZN(n7361) );
  INV_X1 U10461 ( .A(n7057), .ZN(n6294) );
  XNOR2_X1 U10462 ( .A(n6294), .B(n7361), .ZN(n6298) );
  XNOR2_X1 U10463 ( .A(n6674), .B(n6738), .ZN(n6296) );
  XNOR2_X1 U10464 ( .A(n7365), .B(n16035), .ZN(n6295) );
  XNOR2_X1 U10465 ( .A(n6296), .B(n6295), .ZN(n6297) );
  INV_X1 U10466 ( .A(n7978), .ZN(n6299) );
  XNOR2_X1 U10467 ( .A(n6711), .B(n6300), .ZN(n6355) );
  XNOR2_X1 U10468 ( .A(n6301), .B(n6489), .ZN(n7395) );
  XNOR2_X1 U10469 ( .A(n7395), .B(n6355), .ZN(n6305) );
  XNOR2_X1 U10470 ( .A(n6776), .B(n6854), .ZN(n6303) );
  XNOR2_X1 U10471 ( .A(n7296), .B(n1911), .ZN(n6302) );
  XNOR2_X1 U10472 ( .A(n6303), .B(n6302), .ZN(n6304) );
  INV_X1 U10474 ( .A(n6679), .ZN(n6307) );
  XNOR2_X1 U10475 ( .A(n6927), .B(n645), .ZN(n6308) );
  XNOR2_X1 U10476 ( .A(n6309), .B(n6308), .ZN(n6311) );
  XNOR2_X1 U10477 ( .A(n7316), .B(n7373), .ZN(n6505) );
  XNOR2_X1 U10478 ( .A(n7273), .B(n7179), .ZN(n6327) );
  XNOR2_X1 U10479 ( .A(n6505), .B(n6327), .ZN(n6310) );
  NAND2_X1 U10480 ( .A1(n7982), .A2(n7984), .ZN(n7110) );
  XNOR2_X1 U10481 ( .A(n7249), .B(n7184), .ZN(n6334) );
  INV_X1 U10482 ( .A(n7338), .ZN(n6313) );
  XNOR2_X1 U10483 ( .A(n7384), .B(n6313), .ZN(n6514) );
  XNOR2_X1 U10484 ( .A(n6514), .B(n6334), .ZN(n6317) );
  XNOR2_X1 U10485 ( .A(n6873), .B(n6917), .ZN(n6315) );
  XNOR2_X1 U10486 ( .A(n7248), .B(n2341), .ZN(n6314) );
  XNOR2_X1 U10487 ( .A(n6314), .B(n6315), .ZN(n6316) );
  NAND2_X1 U10489 ( .A1(n7110), .A2(n6318), .ZN(n6319) );
  NAND2_X1 U10491 ( .A1(n8470), .A2(n20010), .ZN(n6442) );
  XNOR2_X1 U10492 ( .A(n7325), .B(n1904), .ZN(n6321) );
  XNOR2_X1 U10493 ( .A(n6321), .B(n6735), .ZN(n6323) );
  XNOR2_X1 U10494 ( .A(n7232), .B(n7364), .ZN(n6322) );
  XNOR2_X1 U10495 ( .A(n6323), .B(n6322), .ZN(n6326) );
  XNOR2_X1 U10496 ( .A(n6738), .B(n7031), .ZN(n6325) );
  INV_X1 U10497 ( .A(n19778), .ZN(n6324) );
  XNOR2_X1 U10498 ( .A(n6325), .B(n6324), .ZN(n7214) );
  XNOR2_X1 U10499 ( .A(n7214), .B(n6326), .ZN(n6344) );
  INV_X1 U10500 ( .A(n6344), .ZN(n8355) );
  XNOR2_X1 U10501 ( .A(n6328), .B(n6327), .ZN(n6332) );
  XNOR2_X1 U10502 ( .A(n6723), .B(n7318), .ZN(n6330) );
  XNOR2_X1 U10503 ( .A(n6985), .B(n2392), .ZN(n6329) );
  XNOR2_X1 U10504 ( .A(n6330), .B(n6329), .ZN(n6331) );
  NAND2_X1 U10505 ( .A1(n8355), .A2(n7739), .ZN(n7501) );
  INV_X1 U10506 ( .A(n7501), .ZN(n6343) );
  XNOR2_X1 U10507 ( .A(n899), .B(n2257), .ZN(n6333) );
  XNOR2_X1 U10508 ( .A(n7042), .B(n6990), .ZN(n7185) );
  XNOR2_X1 U10509 ( .A(n7185), .B(n6333), .ZN(n6336) );
  XNOR2_X1 U10510 ( .A(n6808), .B(n7337), .ZN(n6992) );
  XNOR2_X1 U10511 ( .A(n6334), .B(n6992), .ZN(n6335) );
  NOR2_X1 U10512 ( .A1(n8354), .A2(n7739), .ZN(n6342) );
  XNOR2_X1 U10513 ( .A(n6478), .B(n7216), .ZN(n6717) );
  XNOR2_X1 U10514 ( .A(n6717), .B(n6337), .ZN(n6341) );
  XNOR2_X1 U10515 ( .A(n7254), .B(n7288), .ZN(n6339) );
  XNOR2_X1 U10516 ( .A(n6977), .B(n2100), .ZN(n6338) );
  XNOR2_X1 U10517 ( .A(n6339), .B(n6338), .ZN(n6340) );
  XNOR2_X1 U10518 ( .A(n6341), .B(n6340), .ZN(n6345) );
  OAI21_X1 U10519 ( .B1(n6343), .B2(n6342), .A(n7743), .ZN(n6361) );
  NAND2_X1 U10520 ( .A1(n8359), .A2(n7739), .ZN(n6359) );
  XNOR2_X1 U10521 ( .A(n6743), .B(n2420), .ZN(n6347) );
  XNOR2_X1 U10522 ( .A(n6346), .B(n6347), .ZN(n6351) );
  XNOR2_X1 U10524 ( .A(n6961), .B(n6349), .ZN(n6350) );
  XNOR2_X1 U10525 ( .A(n6350), .B(n6351), .ZN(n7741) );
  NAND2_X1 U10526 ( .A1(n7504), .A2(n7741), .ZN(n6358) );
  XNOR2_X1 U10527 ( .A(n7392), .B(n6352), .ZN(n6995) );
  INV_X1 U10528 ( .A(n6995), .ZN(n6354) );
  XNOR2_X1 U10529 ( .A(n6713), .B(n1996), .ZN(n6353) );
  XNOR2_X1 U10530 ( .A(n6354), .B(n6353), .ZN(n6357) );
  XNOR2_X1 U10531 ( .A(n7193), .B(n6355), .ZN(n6356) );
  MUX2_X1 U10532 ( .A(n6359), .B(n6358), .S(n8358), .Z(n6360) );
  NOR2_X1 U10533 ( .A1(n8128), .A2(n8884), .ZN(n9089) );
  XNOR2_X1 U10534 ( .A(n6967), .B(n7363), .ZN(n6363) );
  XNOR2_X1 U10535 ( .A(n6362), .B(n7035), .ZN(n6672) );
  XNOR2_X1 U10536 ( .A(n6672), .B(n6363), .ZN(n6367) );
  XNOR2_X1 U10537 ( .A(n7212), .B(n1857), .ZN(n6365) );
  XNOR2_X1 U10538 ( .A(n6365), .B(n6364), .ZN(n6366) );
  XNOR2_X1 U10539 ( .A(n6367), .B(n6366), .ZN(n6951) );
  INV_X1 U10540 ( .A(n6951), .ZN(n8361) );
  XNOR2_X1 U10541 ( .A(n7041), .B(n7384), .ZN(n6689) );
  XNOR2_X1 U10542 ( .A(n6368), .B(n6689), .ZN(n6372) );
  XNOR2_X1 U10543 ( .A(n6918), .B(n19944), .ZN(n6370) );
  XNOR2_X1 U10544 ( .A(n6990), .B(n19216), .ZN(n6369) );
  XNOR2_X1 U10545 ( .A(n6370), .B(n6369), .ZN(n6371) );
  INV_X1 U10546 ( .A(n7709), .ZN(n8360) );
  XNOR2_X1 U10547 ( .A(n6982), .B(n6680), .ZN(n6373) );
  XNOR2_X1 U10548 ( .A(n6374), .B(n6373), .ZN(n6378) );
  XNOR2_X1 U10549 ( .A(n7046), .B(n7373), .ZN(n6376) );
  XNOR2_X1 U10550 ( .A(n6376), .B(n6375), .ZN(n6377) );
  XNOR2_X1 U10551 ( .A(n6378), .B(n6377), .ZN(n7673) );
  OAI21_X1 U10552 ( .B1(n8361), .B2(n8360), .A(n7673), .ZN(n6390) );
  MUX2_X1 U10553 ( .A(n19476), .B(n6380), .S(n6379), .Z(n6383) );
  XNOR2_X1 U10554 ( .A(n6384), .B(n7355), .ZN(n6385) );
  XNOR2_X1 U10556 ( .A(n6385), .B(n6660), .ZN(n6389) );
  XNOR2_X1 U10557 ( .A(n6867), .B(n7218), .ZN(n6387) );
  XNOR2_X1 U10558 ( .A(n6386), .B(n6387), .ZN(n6388) );
  XNOR2_X2 U10559 ( .A(n6389), .B(n6388), .ZN(n7675) );
  NAND2_X1 U10560 ( .A1(n6390), .A2(n7675), .ZN(n6402) );
  AND2_X1 U10561 ( .A1(n7709), .A2(n7673), .ZN(n8364) );
  XNOR2_X1 U10562 ( .A(n7006), .B(n18284), .ZN(n6391) );
  XNOR2_X1 U10563 ( .A(n6391), .B(n7206), .ZN(n6392) );
  XNOR2_X1 U10564 ( .A(n6693), .B(n7267), .ZN(n6612) );
  XNOR2_X1 U10565 ( .A(n6392), .B(n6612), .ZN(n6395) );
  XNOR2_X1 U10566 ( .A(n7345), .B(n6393), .ZN(n6394) );
  NAND2_X1 U10567 ( .A1(n8364), .A2(n7674), .ZN(n6401) );
  XNOR2_X1 U10568 ( .A(n6997), .B(n632), .ZN(n6397) );
  XNOR2_X1 U10569 ( .A(n7195), .B(n7390), .ZN(n6396) );
  XNOR2_X1 U10570 ( .A(n6397), .B(n6396), .ZN(n6400) );
  XNOR2_X1 U10571 ( .A(n6489), .B(n7014), .ZN(n6666) );
  XNOR2_X1 U10572 ( .A(n6666), .B(n6398), .ZN(n6399) );
  NOR2_X1 U10573 ( .A1(n9453), .A2(n6438), .ZN(n6403) );
  NAND2_X1 U10574 ( .A1(n9089), .A2(n6403), .ZN(n6441) );
  XNOR2_X1 U10575 ( .A(n6404), .B(n7196), .ZN(n7126) );
  INV_X1 U10576 ( .A(n7126), .ZN(n6557) );
  XNOR2_X1 U10577 ( .A(n6557), .B(n7295), .ZN(n6407) );
  XNOR2_X1 U10578 ( .A(n7017), .B(n7065), .ZN(n6773) );
  XNOR2_X1 U10579 ( .A(n7013), .B(n2424), .ZN(n6405) );
  XNOR2_X1 U10580 ( .A(n6773), .B(n6405), .ZN(n6406) );
  XNOR2_X2 U10581 ( .A(n6407), .B(n6406), .ZN(n7749) );
  INV_X1 U10582 ( .A(n7116), .ZN(n6409) );
  XNOR2_X1 U10583 ( .A(n7115), .B(n17170), .ZN(n6408) );
  XNOR2_X1 U10584 ( .A(n6408), .B(n6409), .ZN(n6412) );
  XNOR2_X1 U10585 ( .A(n6410), .B(n7081), .ZN(n6411) );
  XNOR2_X1 U10586 ( .A(n6412), .B(n6411), .ZN(n6415) );
  XNOR2_X1 U10587 ( .A(n7026), .B(n6819), .ZN(n6413) );
  XNOR2_X1 U10588 ( .A(n6413), .B(n20203), .ZN(n6414) );
  XNOR2_X1 U10589 ( .A(n7070), .B(n7202), .ZN(n6416) );
  XNOR2_X1 U10590 ( .A(n7303), .B(n6416), .ZN(n6419) );
  XNOR2_X1 U10591 ( .A(n7163), .B(n7264), .ZN(n6443) );
  XNOR2_X1 U10592 ( .A(n179), .B(n2344), .ZN(n6417) );
  XNOR2_X1 U10593 ( .A(n6443), .B(n6417), .ZN(n6418) );
  XNOR2_X1 U10594 ( .A(n6419), .B(n6418), .ZN(n7914) );
  INV_X1 U10595 ( .A(n7914), .ZN(n7746) );
  INV_X1 U10596 ( .A(n6420), .ZN(n6675) );
  XNOR2_X1 U10597 ( .A(n6675), .B(n7032), .ZN(n6422) );
  XNOR2_X1 U10598 ( .A(n7155), .B(n18090), .ZN(n6421) );
  XNOR2_X1 U10599 ( .A(n6422), .B(n6421), .ZN(n6425) );
  XNOR2_X1 U10600 ( .A(n6883), .B(n6423), .ZN(n6424) );
  XNOR2_X1 U10601 ( .A(n7383), .B(n7333), .ZN(n6426) );
  XNOR2_X1 U10602 ( .A(n7334), .B(n6426), .ZN(n6431) );
  XNOR2_X1 U10603 ( .A(n6427), .B(n6573), .ZN(n7135) );
  INV_X1 U10604 ( .A(n7135), .ZN(n6429) );
  XNOR2_X1 U10605 ( .A(n6687), .B(n875), .ZN(n6428) );
  XNOR2_X1 U10606 ( .A(n6429), .B(n6428), .ZN(n6430) );
  XNOR2_X1 U10607 ( .A(n6431), .B(n6430), .ZN(n7508) );
  INV_X1 U10608 ( .A(n7087), .ZN(n6432) );
  XNOR2_X1 U10609 ( .A(n7047), .B(n6432), .ZN(n6433) );
  XNOR2_X1 U10610 ( .A(n7313), .B(n6433), .ZN(n6437) );
  XNOR2_X1 U10611 ( .A(n7371), .B(n6469), .ZN(n6435) );
  XNOR2_X1 U10612 ( .A(n7144), .B(n17999), .ZN(n6434) );
  XNOR2_X1 U10613 ( .A(n6435), .B(n6434), .ZN(n6436) );
  INV_X1 U10614 ( .A(n6438), .ZN(n8126) );
  INV_X1 U10615 ( .A(n6443), .ZN(n6445) );
  XNOR2_X1 U10616 ( .A(n7007), .B(n17851), .ZN(n6444) );
  XNOR2_X1 U10617 ( .A(n6445), .B(n6444), .ZN(n6448) );
  XNOR2_X1 U10618 ( .A(n6446), .B(n6961), .ZN(n6447) );
  XNOR2_X1 U10619 ( .A(n7116), .B(n7221), .ZN(n6449) );
  XNOR2_X1 U10620 ( .A(n6864), .B(n6449), .ZN(n6452) );
  XNOR2_X1 U10621 ( .A(n6661), .B(n610), .ZN(n6450) );
  XNOR2_X1 U10622 ( .A(n7353), .B(n6450), .ZN(n6451) );
  XNOR2_X1 U10623 ( .A(n6452), .B(n6451), .ZN(n6467) );
  XNOR2_X1 U10624 ( .A(n6707), .B(n2023), .ZN(n6453) );
  XNOR2_X1 U10625 ( .A(n6776), .B(n7018), .ZN(n6669) );
  XNOR2_X1 U10626 ( .A(n6453), .B(n6669), .ZN(n6455) );
  XNOR2_X1 U10627 ( .A(n7013), .B(n6854), .ZN(n7397) );
  XNOR2_X1 U10628 ( .A(n7397), .B(n6995), .ZN(n6454) );
  XNOR2_X1 U10629 ( .A(n7364), .B(n7031), .ZN(n6456) );
  XNOR2_X1 U10630 ( .A(n6881), .B(n6456), .ZN(n6460) );
  XNOR2_X1 U10631 ( .A(n6674), .B(n7155), .ZN(n6458) );
  XNOR2_X1 U10632 ( .A(n7365), .B(n18478), .ZN(n6457) );
  XNOR2_X1 U10633 ( .A(n6458), .B(n6457), .ZN(n6459) );
  XNOR2_X1 U10634 ( .A(n7383), .B(n6573), .ZN(n6463) );
  INV_X1 U10635 ( .A(n20593), .ZN(n6461) );
  XNOR2_X1 U10636 ( .A(n7337), .B(n6461), .ZN(n6462) );
  XNOR2_X1 U10637 ( .A(n6463), .B(n6462), .ZN(n6466) );
  XNOR2_X1 U10638 ( .A(n7248), .B(n7042), .ZN(n6685) );
  XNOR2_X1 U10639 ( .A(n6464), .B(n6685), .ZN(n6465) );
  XNOR2_X1 U10640 ( .A(n6466), .B(n6465), .ZN(n7644) );
  NAND2_X1 U10641 ( .A1(n8219), .A2(n7644), .ZN(n7646) );
  INV_X1 U10642 ( .A(n6467), .ZN(n8079) );
  NAND3_X1 U10643 ( .A1(n7646), .A2(n8079), .A3(n6468), .ZN(n6475) );
  INV_X1 U10644 ( .A(n8076), .ZN(n7645) );
  XNOR2_X1 U10645 ( .A(n7377), .B(n6889), .ZN(n6473) );
  XNOR2_X1 U10646 ( .A(n6679), .B(n6469), .ZN(n6471) );
  XNOR2_X1 U10647 ( .A(n7050), .B(n19052), .ZN(n6470) );
  XNOR2_X1 U10648 ( .A(n6471), .B(n6470), .ZN(n6472) );
  NAND3_X1 U10649 ( .A1(n8220), .A2(n7645), .A3(n8219), .ZN(n6474) );
  XNOR2_X1 U10650 ( .A(n7289), .B(n6520), .ZN(n6619) );
  XNOR2_X1 U10651 ( .A(n6761), .B(n20227), .ZN(n6476) );
  XNOR2_X1 U10652 ( .A(n6619), .B(n6476), .ZN(n6482) );
  XNOR2_X1 U10653 ( .A(n6477), .B(n7257), .ZN(n6480) );
  XNOR2_X1 U10654 ( .A(n6478), .B(n2151), .ZN(n6479) );
  XNOR2_X1 U10655 ( .A(n6480), .B(n6479), .ZN(n6481) );
  XNOR2_X1 U10656 ( .A(n6743), .B(n6693), .ZN(n6483) );
  XNOR2_X1 U10657 ( .A(n6768), .B(n7306), .ZN(n7074) );
  XNOR2_X1 U10658 ( .A(n7074), .B(n6483), .ZN(n6487) );
  XNOR2_X1 U10659 ( .A(n6945), .B(n2446), .ZN(n6485) );
  XNOR2_X1 U10660 ( .A(n6485), .B(n6484), .ZN(n6486) );
  XNOR2_X1 U10661 ( .A(n6487), .B(n6486), .ZN(n8113) );
  XNOR2_X1 U10662 ( .A(n7064), .B(n6488), .ZN(n6493) );
  XNOR2_X1 U10663 ( .A(n6489), .B(n6641), .ZN(n6491) );
  INV_X1 U10664 ( .A(n2305), .ZN(n18389) );
  XNOR2_X1 U10665 ( .A(n6713), .B(n18389), .ZN(n6490) );
  XNOR2_X1 U10666 ( .A(n6491), .B(n6490), .ZN(n6492) );
  NAND3_X1 U10667 ( .A1(n8253), .A2(n7844), .A3(n8114), .ZN(n6519) );
  AND2_X1 U10668 ( .A1(n6702), .A2(n8113), .ZN(n8254) );
  XNOR2_X1 U10669 ( .A(n6495), .B(n6625), .ZN(n6504) );
  XNOR2_X1 U10670 ( .A(n6735), .B(n19850), .ZN(n6502) );
  NAND3_X1 U10671 ( .A1(n6496), .A2(n641), .A3(n6500), .ZN(n6499) );
  INV_X1 U10672 ( .A(n6496), .ZN(n6497) );
  INV_X1 U10673 ( .A(n641), .ZN(n18379) );
  NAND2_X1 U10674 ( .A1(n6497), .A2(n18379), .ZN(n6498) );
  OAI211_X1 U10675 ( .C1(n641), .C2(n6500), .A(n6499), .B(n6498), .ZN(n6501)
         );
  XNOR2_X1 U10676 ( .A(n6502), .B(n6501), .ZN(n6503) );
  XNOR2_X1 U10677 ( .A(n6504), .B(n6503), .ZN(n6510) );
  NAND2_X1 U10678 ( .A1(n8254), .A2(n7560), .ZN(n6518) );
  XNOR2_X1 U10679 ( .A(n6723), .B(n6793), .ZN(n6508) );
  XNOR2_X1 U10680 ( .A(n6634), .B(n18863), .ZN(n6507) );
  XNOR2_X1 U10681 ( .A(n6508), .B(n6507), .ZN(n6509) );
  NAND2_X1 U10682 ( .A1(n7560), .A2(n8245), .ZN(n6517) );
  XNOR2_X1 U10683 ( .A(n6512), .B(n6511), .ZN(n6730) );
  XNOR2_X1 U10684 ( .A(n6513), .B(n16651), .ZN(n6515) );
  NAND3_X1 U10685 ( .A1(n8248), .A2(n8251), .A3(n7844), .ZN(n6516) );
  NAND4_X1 U10686 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n8713)
         );
  XNOR2_X1 U10687 ( .A(n7286), .B(n6759), .ZN(n6524) );
  XNOR2_X1 U10688 ( .A(n6520), .B(n7218), .ZN(n6522) );
  XNOR2_X1 U10689 ( .A(n7122), .B(n18984), .ZN(n6521) );
  XNOR2_X1 U10690 ( .A(n6522), .B(n6521), .ZN(n6523) );
  INV_X1 U10691 ( .A(n6997), .ZN(n6525) );
  XNOR2_X1 U10692 ( .A(n6525), .B(n6714), .ZN(n6856) );
  XNOR2_X1 U10693 ( .A(n6526), .B(n6856), .ZN(n6529) );
  XNOR2_X1 U10694 ( .A(n6641), .B(n2035), .ZN(n6527) );
  XNOR2_X1 U10695 ( .A(n7294), .B(n6527), .ZN(n6528) );
  XNOR2_X1 U10696 ( .A(n6529), .B(n6528), .ZN(n8087) );
  XNOR2_X1 U10697 ( .A(n6982), .B(n6633), .ZN(n6887) );
  XNOR2_X1 U10698 ( .A(n20455), .B(n7315), .ZN(n6533) );
  INV_X1 U10699 ( .A(n17060), .ZN(n6530) );
  XNOR2_X1 U10700 ( .A(n6634), .B(n6530), .ZN(n6531) );
  XNOR2_X1 U10701 ( .A(n6790), .B(n6531), .ZN(n6532) );
  XNOR2_X1 U10702 ( .A(n6533), .B(n6532), .ZN(n8085) );
  XNOR2_X1 U10703 ( .A(n6728), .B(n6990), .ZN(n6876) );
  XNOR2_X1 U10704 ( .A(n6534), .B(n6876), .ZN(n6538) );
  XNOR2_X1 U10705 ( .A(n7333), .B(n6919), .ZN(n6536) );
  XNOR2_X1 U10706 ( .A(n7336), .B(n18396), .ZN(n6535) );
  XNOR2_X1 U10707 ( .A(n6536), .B(n6535), .ZN(n6537) );
  XNOR2_X1 U10708 ( .A(n6538), .B(n6537), .ZN(n8086) );
  AOI22_X1 U10709 ( .A1(n19826), .A2(n20254), .B1(n8085), .B2(n8086), .ZN(
        n7556) );
  INV_X1 U10710 ( .A(n8087), .ZN(n6539) );
  XNOR2_X1 U10711 ( .A(n6742), .B(n7206), .ZN(n6849) );
  XNOR2_X1 U10712 ( .A(n6767), .B(n18997), .ZN(n6540) );
  XNOR2_X1 U10713 ( .A(n6540), .B(n6945), .ZN(n6541) );
  XNOR2_X1 U10714 ( .A(n6541), .B(n6849), .ZN(n6544) );
  INV_X1 U10715 ( .A(n7308), .ZN(n6542) );
  XNOR2_X1 U10716 ( .A(n7305), .B(n6542), .ZN(n6543) );
  XNOR2_X1 U10717 ( .A(n6545), .B(n2382), .ZN(n6547) );
  XNOR2_X1 U10718 ( .A(n6546), .B(n6547), .ZN(n6549) );
  XNOR2_X1 U10719 ( .A(n19778), .B(n6736), .ZN(n6879) );
  XNOR2_X1 U10720 ( .A(n6879), .B(n6752), .ZN(n6548) );
  INV_X1 U10722 ( .A(n8086), .ZN(n8230) );
  OAI211_X1 U10723 ( .C1(n20254), .C2(n8232), .A(n20108), .B(n8230), .ZN(n6550) );
  XNOR2_X1 U10724 ( .A(n7201), .B(n18084), .ZN(n6551) );
  XNOR2_X1 U10725 ( .A(n7202), .B(n6551), .ZN(n6553) );
  XNOR2_X1 U10726 ( .A(n6552), .B(n6553), .ZN(n6556) );
  XNOR2_X1 U10727 ( .A(n7345), .B(n6554), .ZN(n6555) );
  XNOR2_X2 U10728 ( .A(n6556), .B(n6555), .ZN(n8241) );
  XNOR2_X1 U10729 ( .A(n6855), .B(n7391), .ZN(n6996) );
  XNOR2_X1 U10730 ( .A(n6557), .B(n6996), .ZN(n6561) );
  XNOR2_X1 U10731 ( .A(n6558), .B(n347), .ZN(n6559) );
  XNOR2_X1 U10732 ( .A(n7016), .B(n6559), .ZN(n6560) );
  XNOR2_X1 U10733 ( .A(n7116), .B(n20203), .ZN(n6563) );
  XNOR2_X1 U10734 ( .A(n6562), .B(n6563), .ZN(n6567) );
  XNOR2_X1 U10735 ( .A(n6819), .B(n18208), .ZN(n6564) );
  XNOR2_X1 U10736 ( .A(n6565), .B(n6564), .ZN(n6566) );
  XNOR2_X1 U10737 ( .A(n6567), .B(n6566), .ZN(n7862) );
  XNOR2_X1 U10738 ( .A(n6883), .B(n7036), .ZN(n6571) );
  XNOR2_X1 U10739 ( .A(n19764), .B(n18433), .ZN(n6569) );
  XNOR2_X1 U10740 ( .A(n6569), .B(n6737), .ZN(n6570) );
  XNOR2_X1 U10741 ( .A(n6570), .B(n6571), .ZN(n6578) );
  NOR2_X1 U10742 ( .A1(n8239), .A2(n8100), .ZN(n6572) );
  NAND2_X1 U10743 ( .A1(n6572), .A2(n7862), .ZN(n6586) );
  XNOR2_X1 U10744 ( .A(n7097), .B(n6573), .ZN(n6574) );
  XNOR2_X1 U10745 ( .A(n7040), .B(n6574), .ZN(n6577) );
  XNOR2_X1 U10746 ( .A(n7382), .B(n6872), .ZN(n6993) );
  XNOR2_X1 U10747 ( .A(n7188), .B(n2280), .ZN(n6575) );
  XNOR2_X1 U10748 ( .A(n6993), .B(n6575), .ZN(n6576) );
  XNOR2_X1 U10749 ( .A(n6577), .B(n6576), .ZN(n8098) );
  INV_X1 U10750 ( .A(n6578), .ZN(n8099) );
  OAI21_X1 U10751 ( .B1(n20493), .B2(n8238), .A(n8099), .ZN(n6585) );
  XNOR2_X1 U10752 ( .A(n6721), .B(n6579), .ZN(n6583) );
  XNOR2_X1 U10753 ( .A(n6839), .B(n7091), .ZN(n6581) );
  XNOR2_X1 U10754 ( .A(n7144), .B(n19018), .ZN(n6580) );
  XNOR2_X1 U10755 ( .A(n6581), .B(n6580), .ZN(n6582) );
  OAI21_X1 U10756 ( .B1(n8112), .B2(n8111), .A(n8239), .ZN(n6584) );
  OAI21_X1 U10757 ( .B1(n8628), .B2(n8713), .A(n6587), .ZN(n6655) );
  XNOR2_X1 U10758 ( .A(n6588), .B(n6660), .ZN(n6592) );
  XNOR2_X1 U10759 ( .A(n7288), .B(n17535), .ZN(n6589) );
  XNOR2_X1 U10760 ( .A(n6590), .B(n6589), .ZN(n6591) );
  XNOR2_X2 U10761 ( .A(n6592), .B(n6591), .ZN(n8095) );
  XNOR2_X1 U10762 ( .A(n6593), .B(n6838), .ZN(n6597) );
  XNOR2_X1 U10763 ( .A(n6680), .B(n7318), .ZN(n6595) );
  XNOR2_X1 U10764 ( .A(n7373), .B(n1386), .ZN(n6594) );
  XNOR2_X1 U10765 ( .A(n6595), .B(n6594), .ZN(n6596) );
  XNOR2_X1 U10766 ( .A(n6597), .B(n6596), .ZN(n8090) );
  XNOR2_X1 U10768 ( .A(n6810), .B(n6598), .ZN(n6601) );
  INV_X1 U10769 ( .A(n2369), .ZN(n18503) );
  XNOR2_X1 U10770 ( .A(n7337), .B(n18503), .ZN(n6599) );
  XNOR2_X1 U10771 ( .A(n6689), .B(n6599), .ZN(n6600) );
  NAND2_X1 U10772 ( .A1(n20511), .A2(n8211), .ZN(n6618) );
  XNOR2_X1 U10773 ( .A(n883), .B(n2307), .ZN(n6602) );
  XOR2_X1 U10774 ( .A(n6801), .B(n6602), .Z(n6605) );
  XNOR2_X1 U10775 ( .A(n6672), .B(n6603), .ZN(n6604) );
  XNOR2_X1 U10776 ( .A(n6824), .B(n6606), .ZN(n6609) );
  XNOR2_X1 U10777 ( .A(n7298), .B(n2954), .ZN(n6607) );
  XNOR2_X1 U10778 ( .A(n6666), .B(n6607), .ZN(n6608) );
  NAND2_X1 U10779 ( .A1(n8094), .A2(n8212), .ZN(n7898) );
  OAI21_X1 U10780 ( .B1(n8095), .B2(n8094), .A(n7898), .ZN(n6610) );
  XNOR2_X1 U10781 ( .A(n6611), .B(n6612), .ZN(n6616) );
  XNOR2_X1 U10782 ( .A(n7304), .B(n7266), .ZN(n6614) );
  XNOR2_X1 U10783 ( .A(n7006), .B(n19102), .ZN(n6613) );
  XNOR2_X1 U10784 ( .A(n6614), .B(n6613), .ZN(n6615) );
  XNOR2_X1 U10785 ( .A(n6616), .B(n6615), .ZN(n7631) );
  NAND3_X1 U10786 ( .A1(n8095), .A2(n7631), .A3(n8209), .ZN(n6617) );
  XNOR2_X1 U10787 ( .A(n6659), .B(n6619), .ZN(n6623) );
  INV_X1 U10789 ( .A(n8175), .ZN(n8067) );
  XNOR2_X1 U10790 ( .A(n7212), .B(n2233), .ZN(n6624) );
  XNOR2_X1 U10791 ( .A(n6676), .B(n6624), .ZN(n6629) );
  INV_X1 U10792 ( .A(n6625), .ZN(n6627) );
  XNOR2_X1 U10793 ( .A(n6627), .B(n6626), .ZN(n6628) );
  XNOR2_X1 U10794 ( .A(n7187), .B(n538), .ZN(n6631) );
  XNOR2_X1 U10795 ( .A(n20250), .B(n6631), .ZN(n6632) );
  NAND3_X1 U10796 ( .A1(n8067), .A2(n8178), .A3(n8068), .ZN(n6639) );
  XNOR2_X1 U10797 ( .A(n6633), .B(n7178), .ZN(n6636) );
  INV_X1 U10798 ( .A(n2385), .ZN(n19123) );
  XNOR2_X1 U10799 ( .A(n6634), .B(n19123), .ZN(n6635) );
  XNOR2_X1 U10800 ( .A(n6636), .B(n6635), .ZN(n6637) );
  OR2_X1 U10801 ( .A1(n19901), .A2(n8066), .ZN(n7417) );
  NAND2_X1 U10802 ( .A1(n6639), .A2(n7417), .ZN(n6654) );
  XNOR2_X1 U10803 ( .A(n6665), .B(n6640), .ZN(n6645) );
  XNOR2_X1 U10804 ( .A(n6641), .B(n7195), .ZN(n6643) );
  XNOR2_X1 U10805 ( .A(n7296), .B(n2337), .ZN(n6642) );
  XNOR2_X1 U10806 ( .A(n6643), .B(n6642), .ZN(n6644) );
  XNOR2_X2 U10807 ( .A(n6645), .B(n6644), .ZN(n8179) );
  NAND2_X1 U10808 ( .A1(n8068), .A2(n923), .ZN(n6652) );
  INV_X1 U10809 ( .A(n6692), .ZN(n6647) );
  XNOR2_X1 U10810 ( .A(n6647), .B(n6646), .ZN(n6651) );
  XNOR2_X1 U10811 ( .A(n7306), .B(n6945), .ZN(n6649) );
  XNOR2_X1 U10812 ( .A(n7006), .B(n2079), .ZN(n6648) );
  XNOR2_X1 U10813 ( .A(n6649), .B(n6648), .ZN(n6650) );
  XNOR2_X1 U10814 ( .A(n6651), .B(n6650), .ZN(n7621) );
  AOI21_X1 U10815 ( .B1(n7887), .B2(n6652), .A(n8069), .ZN(n6653) );
  XNOR2_X1 U10817 ( .A(n6659), .B(n6660), .ZN(n6664) );
  XNOR2_X1 U10818 ( .A(n6661), .B(n7081), .ZN(n6760) );
  XNOR2_X1 U10819 ( .A(n7221), .B(n18848), .ZN(n6662) );
  XNOR2_X1 U10820 ( .A(n6760), .B(n6662), .ZN(n6663) );
  XNOR2_X2 U10821 ( .A(n6664), .B(n6663), .ZN(n8262) );
  INV_X1 U10822 ( .A(n6665), .ZN(n6667) );
  XNOR2_X1 U10823 ( .A(n7065), .B(n621), .ZN(n6668) );
  XNOR2_X1 U10824 ( .A(n6669), .B(n6668), .ZN(n6670) );
  XNOR2_X1 U10825 ( .A(n7031), .B(n15479), .ZN(n6673) );
  XNOR2_X1 U10826 ( .A(n6672), .B(n6673), .ZN(n6678) );
  XNOR2_X1 U10827 ( .A(n6675), .B(n6674), .ZN(n6751) );
  XNOR2_X1 U10828 ( .A(n6751), .B(n6676), .ZN(n6677) );
  XNOR2_X1 U10829 ( .A(n6678), .B(n6677), .ZN(n7571) );
  INV_X1 U10830 ( .A(n7571), .ZN(n8264) );
  XNOR2_X1 U10831 ( .A(n6679), .B(n7087), .ZN(n6794) );
  XNOR2_X1 U10832 ( .A(n7050), .B(n18830), .ZN(n6682) );
  XNOR2_X1 U10833 ( .A(n6680), .B(n7373), .ZN(n6681) );
  XNOR2_X1 U10834 ( .A(n6682), .B(n6681), .ZN(n6683) );
  XNOR2_X1 U10836 ( .A(n6686), .B(n6685), .ZN(n6691) );
  XNOR2_X1 U10837 ( .A(n6687), .B(n19467), .ZN(n6688) );
  XNOR2_X1 U10838 ( .A(n6689), .B(n6688), .ZN(n6690) );
  XNOR2_X1 U10839 ( .A(n6690), .B(n6691), .ZN(n8150) );
  NAND2_X1 U10840 ( .A1(n8261), .A2(n8150), .ZN(n6699) );
  XNOR2_X1 U10841 ( .A(n6692), .B(n6770), .ZN(n6697) );
  XNOR2_X1 U10842 ( .A(n6693), .B(n7007), .ZN(n6695) );
  XNOR2_X1 U10843 ( .A(n7267), .B(n18308), .ZN(n6694) );
  XNOR2_X1 U10844 ( .A(n6695), .B(n6694), .ZN(n6696) );
  XNOR2_X1 U10845 ( .A(n6697), .B(n6696), .ZN(n8153) );
  INV_X1 U10846 ( .A(n6702), .ZN(n8246) );
  NOR2_X1 U10847 ( .A1(n8253), .A2(n8246), .ZN(n8252) );
  NAND3_X1 U10849 ( .A1(n8253), .A2(n7560), .A3(n8251), .ZN(n6705) );
  AND2_X1 U10850 ( .A1(n9313), .A2(n9305), .ZN(n6896) );
  INV_X1 U10851 ( .A(n941), .ZN(n6706) );
  XNOR2_X1 U10852 ( .A(n19855), .B(n6706), .ZN(n6710) );
  XNOR2_X1 U10853 ( .A(n6708), .B(n2323), .ZN(n6709) );
  XNOR2_X1 U10854 ( .A(n6710), .B(n6709), .ZN(n6716) );
  INV_X1 U10855 ( .A(n6711), .ZN(n6712) );
  XNOR2_X1 U10856 ( .A(n6712), .B(n7391), .ZN(n7194) );
  XNOR2_X1 U10857 ( .A(n6713), .B(n6714), .ZN(n7125) );
  XNOR2_X1 U10858 ( .A(n7194), .B(n7125), .ZN(n6715) );
  XNOR2_X1 U10859 ( .A(n6716), .B(n6715), .ZN(n6734) );
  XNOR2_X1 U10860 ( .A(n7122), .B(n18716), .ZN(n6720) );
  XNOR2_X1 U10861 ( .A(n6722), .B(n6721), .ZN(n6727) );
  XNOR2_X1 U10862 ( .A(n6724), .B(n6723), .ZN(n7148) );
  XNOR2_X1 U10863 ( .A(n7179), .B(n2317), .ZN(n6725) );
  XNOR2_X1 U10864 ( .A(n7148), .B(n6725), .ZN(n6726) );
  XNOR2_X1 U10865 ( .A(n6727), .B(n6726), .ZN(n7671) );
  INV_X1 U10866 ( .A(n7671), .ZN(n8375) );
  XNOR2_X1 U10867 ( .A(n6729), .B(n7184), .ZN(n6731) );
  INV_X1 U10868 ( .A(n6734), .ZN(n8377) );
  XNOR2_X1 U10870 ( .A(n6736), .B(n6735), .ZN(n7152) );
  XNOR2_X1 U10871 ( .A(n7152), .B(n6737), .ZN(n6741) );
  XNOR2_X1 U10872 ( .A(n6738), .B(n19321), .ZN(n6739) );
  XNOR2_X1 U10873 ( .A(n6754), .B(n6165), .ZN(n7060) );
  XNOR2_X1 U10874 ( .A(n6739), .B(n7060), .ZN(n6740) );
  XNOR2_X1 U10876 ( .A(n6743), .B(n6742), .ZN(n7162) );
  XNOR2_X1 U10877 ( .A(n6744), .B(n7162), .ZN(n6749) );
  XNOR2_X1 U10878 ( .A(n6768), .B(n6745), .ZN(n6747) );
  XNOR2_X1 U10879 ( .A(n7201), .B(n2381), .ZN(n6746) );
  XNOR2_X1 U10880 ( .A(n6747), .B(n6746), .ZN(n6748) );
  XNOR2_X1 U10881 ( .A(n6749), .B(n6748), .ZN(n7542) );
  NAND2_X1 U10882 ( .A1(n7542), .A2(n6734), .ZN(n8142) );
  INV_X1 U10883 ( .A(n6751), .ZN(n6753) );
  XNOR2_X1 U10884 ( .A(n6753), .B(n6752), .ZN(n6758) );
  XNOR2_X1 U10885 ( .A(n7230), .B(n7032), .ZN(n6756) );
  XNOR2_X1 U10886 ( .A(n19850), .B(n16366), .ZN(n6755) );
  XNOR2_X1 U10887 ( .A(n6756), .B(n6755), .ZN(n6757) );
  XNOR2_X1 U10889 ( .A(n6759), .B(n6760), .ZN(n6765) );
  XNOR2_X1 U10890 ( .A(n6761), .B(n7257), .ZN(n6763) );
  XNOR2_X1 U10891 ( .A(n7026), .B(n17466), .ZN(n6762) );
  XNOR2_X1 U10892 ( .A(n6763), .B(n6762), .ZN(n6764) );
  XNOR2_X1 U10893 ( .A(n6765), .B(n6764), .ZN(n8380) );
  XNOR2_X1 U10894 ( .A(n179), .B(n7263), .ZN(n6766) );
  XNOR2_X1 U10895 ( .A(n7305), .B(n6766), .ZN(n6772) );
  XNOR2_X1 U10896 ( .A(n20225), .B(n18075), .ZN(n6769) );
  XNOR2_X1 U10897 ( .A(n6769), .B(n6768), .ZN(n6771) );
  MUX2_X1 U10898 ( .A(n8387), .B(n163), .S(n19925), .Z(n6800) );
  INV_X1 U10899 ( .A(n6773), .ZN(n6775) );
  XNOR2_X1 U10900 ( .A(n6775), .B(n6774), .ZN(n6781) );
  XNOR2_X1 U10901 ( .A(n941), .B(n6776), .ZN(n6779) );
  XNOR2_X1 U10902 ( .A(n6777), .B(n573), .ZN(n6778) );
  XNOR2_X1 U10903 ( .A(n6779), .B(n6778), .ZN(n6780) );
  INV_X1 U10904 ( .A(n7684), .ZN(n8385) );
  XNOR2_X1 U10905 ( .A(n6782), .B(n7332), .ZN(n6785) );
  XNOR2_X1 U10906 ( .A(n6783), .B(n7333), .ZN(n6784) );
  XNOR2_X1 U10907 ( .A(n6784), .B(n6785), .ZN(n6789) );
  XNOR2_X1 U10908 ( .A(n7248), .B(n16242), .ZN(n6787) );
  XNOR2_X1 U10909 ( .A(n7098), .B(n6787), .ZN(n6788) );
  NAND3_X1 U10910 ( .A1(n19925), .A2(n8387), .A3(n7497), .ZN(n6799) );
  XNOR2_X1 U10911 ( .A(n7272), .B(n17989), .ZN(n6792) );
  XNOR2_X1 U10913 ( .A(n19852), .B(n6792), .ZN(n6798) );
  XNOR2_X1 U10914 ( .A(n7047), .B(n6793), .ZN(n6796) );
  INV_X1 U10915 ( .A(n6794), .ZN(n6795) );
  XNOR2_X1 U10916 ( .A(n6795), .B(n6796), .ZN(n6797) );
  XNOR2_X1 U10918 ( .A(n6966), .B(n7031), .ZN(n6803) );
  INV_X1 U10919 ( .A(n6801), .ZN(n6802) );
  XNOR2_X1 U10920 ( .A(n6802), .B(n6803), .ZN(n6807) );
  XNOR2_X1 U10921 ( .A(n7364), .B(n19457), .ZN(n6805) );
  XNOR2_X1 U10922 ( .A(n7363), .B(n19840), .ZN(n6804) );
  XNOR2_X1 U10923 ( .A(n6805), .B(n6804), .ZN(n6806) );
  XNOR2_X1 U10924 ( .A(n6808), .B(n7042), .ZN(n6809) );
  XNOR2_X1 U10925 ( .A(n6810), .B(n6809), .ZN(n6815) );
  XNOR2_X1 U10926 ( .A(n6918), .B(n6811), .ZN(n6813) );
  XNOR2_X1 U10927 ( .A(n943), .B(n620), .ZN(n6812) );
  XNOR2_X1 U10928 ( .A(n6813), .B(n6812), .ZN(n6814) );
  XNOR2_X1 U10929 ( .A(n6815), .B(n6814), .ZN(n6830) );
  INV_X1 U10930 ( .A(n7221), .ZN(n6816) );
  XNOR2_X1 U10931 ( .A(n7355), .B(n6816), .ZN(n6817) );
  XNOR2_X1 U10932 ( .A(n6818), .B(n6817), .ZN(n6823) );
  XNOR2_X1 U10933 ( .A(n6977), .B(n6819), .ZN(n6821) );
  XNOR2_X1 U10934 ( .A(n7258), .B(n2055), .ZN(n6820) );
  XNOR2_X1 U10935 ( .A(n6821), .B(n6820), .ZN(n6822) );
  XNOR2_X1 U10936 ( .A(n7240), .B(n6855), .ZN(n6825) );
  XNOR2_X1 U10937 ( .A(n6824), .B(n6825), .ZN(n6829) );
  XNOR2_X1 U10938 ( .A(n7392), .B(n7390), .ZN(n6827) );
  XNOR2_X1 U10939 ( .A(n7018), .B(n457), .ZN(n6826) );
  XOR2_X1 U10940 ( .A(n6827), .B(n6826), .Z(n6828) );
  NAND2_X1 U10941 ( .A1(n7852), .A2(n282), .ZN(n6831) );
  XNOR2_X1 U10942 ( .A(n6832), .B(n7345), .ZN(n6834) );
  XNOR2_X1 U10943 ( .A(n6946), .B(n7007), .ZN(n6833) );
  XNOR2_X1 U10944 ( .A(n6834), .B(n6833), .ZN(n6836) );
  XNOR2_X1 U10945 ( .A(n6836), .B(n6835), .ZN(n8162) );
  INV_X1 U10946 ( .A(n8162), .ZN(n7856) );
  INV_X1 U10947 ( .A(n8159), .ZN(n7851) );
  NAND3_X1 U10948 ( .A1(n7856), .A2(n7724), .A3(n7851), .ZN(n6846) );
  INV_X1 U10949 ( .A(n6838), .ZN(n6841) );
  XNOR2_X1 U10950 ( .A(n7274), .B(n6839), .ZN(n6840) );
  XNOR2_X1 U10951 ( .A(n7050), .B(n18801), .ZN(n6843) );
  XNOR2_X1 U10952 ( .A(n6985), .B(n7046), .ZN(n6842) );
  INV_X1 U10953 ( .A(n8157), .ZN(n6844) );
  OAI21_X1 U10954 ( .B1(n1751), .B2(n20011), .A(n8824), .ZN(n6895) );
  INV_X1 U10955 ( .A(n16424), .ZN(n18792) );
  XNOR2_X1 U10956 ( .A(n6849), .B(n6848), .ZN(n6853) );
  XNOR2_X1 U10957 ( .A(n6850), .B(n7264), .ZN(n7350) );
  XNOR2_X1 U10958 ( .A(n7202), .B(n7304), .ZN(n6851) );
  XNOR2_X1 U10959 ( .A(n7350), .B(n6851), .ZN(n6852) );
  XNOR2_X1 U10960 ( .A(n6853), .B(n6852), .ZN(n8350) );
  XNOR2_X1 U10961 ( .A(n6855), .B(n6854), .ZN(n6857) );
  INV_X1 U10962 ( .A(n6858), .ZN(n6860) );
  XNOR2_X1 U10963 ( .A(n7013), .B(n2275), .ZN(n6859) );
  XNOR2_X1 U10964 ( .A(n6860), .B(n6859), .ZN(n6861) );
  NAND2_X1 U10967 ( .A1(n8350), .A2(n8140), .ZN(n7722) );
  INV_X1 U10968 ( .A(n7122), .ZN(n6863) );
  XNOR2_X1 U10969 ( .A(n20203), .B(n6863), .ZN(n6866) );
  XNOR2_X1 U10971 ( .A(n19741), .B(n6866), .ZN(n6870) );
  XNOR2_X1 U10972 ( .A(n6819), .B(n7218), .ZN(n6976) );
  XNOR2_X1 U10973 ( .A(n19730), .B(n17787), .ZN(n6868) );
  XNOR2_X1 U10974 ( .A(n6976), .B(n6868), .ZN(n6869) );
  XNOR2_X1 U10976 ( .A(n6874), .B(n6873), .ZN(n6875) );
  XNOR2_X1 U10977 ( .A(n6875), .B(n6876), .ZN(n6878) );
  XNOR2_X1 U10978 ( .A(n6878), .B(n6877), .ZN(n8348) );
  NAND2_X1 U10980 ( .A1(n19914), .A2(n8272), .ZN(n6886) );
  INV_X1 U10981 ( .A(n6879), .ZN(n6880) );
  XNOR2_X1 U10982 ( .A(n6880), .B(n6881), .ZN(n6885) );
  XNOR2_X1 U10983 ( .A(n7365), .B(n2298), .ZN(n6882) );
  XNOR2_X1 U10984 ( .A(n6883), .B(n6882), .ZN(n6884) );
  OAI211_X1 U10985 ( .C1(n8352), .C2(n8272), .A(n6886), .B(n8349), .ZN(n6894)
         );
  INV_X1 U10986 ( .A(n6887), .ZN(n6888) );
  XNOR2_X1 U10987 ( .A(n6888), .B(n6889), .ZN(n6893) );
  XNOR2_X1 U10988 ( .A(n7144), .B(n18278), .ZN(n6890) );
  XNOR2_X1 U10989 ( .A(n6891), .B(n6890), .ZN(n6892) );
  INV_X1 U10990 ( .A(n20200), .ZN(n8141) );
  MUX2_X1 U10991 ( .A(n6896), .B(n6895), .S(n9228), .Z(n6898) );
  INV_X1 U10992 ( .A(n9307), .ZN(n9309) );
  AND3_X1 U10993 ( .A1(n20011), .A2(n9309), .A3(n9053), .ZN(n6897) );
  NOR2_X1 U10996 ( .A1(n7500), .A2(n7739), .ZN(n6900) );
  OAI211_X1 U10997 ( .C1(n7931), .C2(n20360), .A(n1063), .B(n20195), .ZN(n6903) );
  INV_X1 U10998 ( .A(n9162), .ZN(n8696) );
  NAND2_X1 U10999 ( .A1(n7904), .A2(n7908), .ZN(n6905) );
  INV_X1 U11001 ( .A(n20166), .ZN(n7755) );
  NOR2_X1 U11002 ( .A1(n7914), .A2(n7750), .ZN(n6907) );
  NOR2_X1 U11003 ( .A1(n7748), .A2(n7507), .ZN(n6906) );
  MUX2_X1 U11004 ( .A(n6907), .B(n6906), .S(n7749), .Z(n6910) );
  XNOR2_X1 U11005 ( .A(n7228), .B(n6911), .ZN(n6916) );
  XNOR2_X1 U11006 ( .A(n7326), .B(n7363), .ZN(n6914) );
  XNOR2_X1 U11007 ( .A(n6912), .B(n2356), .ZN(n6913) );
  XNOR2_X1 U11008 ( .A(n6914), .B(n6913), .ZN(n6915) );
  XNOR2_X1 U11009 ( .A(n7338), .B(Key[60]), .ZN(n6920) );
  XNOR2_X1 U11010 ( .A(n6920), .B(n20250), .ZN(n6921) );
  XNOR2_X1 U11011 ( .A(n7380), .B(n6921), .ZN(n6924) );
  XNOR2_X1 U11012 ( .A(n7248), .B(n943), .ZN(n6922) );
  XNOR2_X1 U11013 ( .A(n6922), .B(n7134), .ZN(n6923) );
  XNOR2_X1 U11014 ( .A(n6924), .B(n6923), .ZN(n7728) );
  XNOR2_X1 U11015 ( .A(n6926), .B(n6925), .ZN(n6930) );
  XNOR2_X1 U11016 ( .A(n6927), .B(n7046), .ZN(n7376) );
  XNOR2_X1 U11017 ( .A(n7316), .B(n18146), .ZN(n6928) );
  XNOR2_X1 U11018 ( .A(n7376), .B(n6928), .ZN(n6929) );
  XNOR2_X1 U11020 ( .A(n5884), .B(n7355), .ZN(n6931) );
  XNOR2_X1 U11021 ( .A(n6931), .B(n7256), .ZN(n6934) );
  XNOR2_X1 U11022 ( .A(n7258), .B(n7121), .ZN(n6933) );
  XNOR2_X1 U11023 ( .A(n6935), .B(n7238), .ZN(n6940) );
  XNOR2_X1 U11024 ( .A(n7390), .B(n7296), .ZN(n6938) );
  INV_X1 U11025 ( .A(n20064), .ZN(n17683) );
  XNOR2_X1 U11026 ( .A(n6936), .B(n17683), .ZN(n6937) );
  XNOR2_X1 U11027 ( .A(n6938), .B(n6937), .ZN(n6939) );
  XNOR2_X1 U11028 ( .A(n6940), .B(n6939), .ZN(n7493) );
  OAI22_X1 U11029 ( .A1(n8166), .A2(n7679), .B1(n8165), .B2(n7728), .ZN(n7729)
         );
  INV_X1 U11030 ( .A(n17024), .ZN(n18670) );
  XNOR2_X1 U11031 ( .A(n7160), .B(n18670), .ZN(n6941) );
  XNOR2_X1 U11032 ( .A(n7345), .B(n6941), .ZN(n6944) );
  XNOR2_X1 U11033 ( .A(n6942), .B(n7306), .ZN(n6943) );
  XNOR2_X1 U11034 ( .A(n6944), .B(n6943), .ZN(n6949) );
  XNOR2_X1 U11035 ( .A(n6948), .B(n6947), .ZN(n7270) );
  NAND2_X1 U11036 ( .A1(n7729), .A2(n8341), .ZN(n6950) );
  NAND2_X1 U11037 ( .A1(n6951), .A2(n7673), .ZN(n7711) );
  NAND2_X1 U11038 ( .A1(n6952), .A2(n8365), .ZN(n6957) );
  INV_X1 U11039 ( .A(n7673), .ZN(n6953) );
  NAND2_X1 U11040 ( .A1(n7709), .A2(n6953), .ZN(n6954) );
  NAND3_X1 U11041 ( .A1(n7711), .A2(n7675), .A3(n6954), .ZN(n6956) );
  INV_X1 U11042 ( .A(n7675), .ZN(n8366) );
  INV_X1 U11043 ( .A(n8365), .ZN(n8363) );
  NAND3_X1 U11044 ( .A1(n1994), .A2(n8363), .A3(n7674), .ZN(n6955) );
  INV_X1 U11045 ( .A(n9163), .ZN(n9161) );
  NAND3_X1 U11046 ( .A1(n8611), .A2(n8609), .A3(n9161), .ZN(n6959) );
  NAND3_X1 U11047 ( .A1(n9164), .A2(n9158), .A3(n1230), .ZN(n6958) );
  XNOR2_X1 U11048 ( .A(n6961), .B(n6960), .ZN(n6965) );
  XNOR2_X1 U11049 ( .A(n7009), .B(n18439), .ZN(n6963) );
  XNOR2_X1 U11050 ( .A(n6963), .B(n6962), .ZN(n6964) );
  XNOR2_X1 U11052 ( .A(n6966), .B(n6967), .ZN(n6969) );
  XNOR2_X1 U11053 ( .A(n7151), .B(n7032), .ZN(n6968) );
  XNOR2_X1 U11054 ( .A(n6969), .B(n6968), .ZN(n6974) );
  XNOR2_X1 U11055 ( .A(n6970), .B(n7364), .ZN(n6972) );
  XNOR2_X1 U11056 ( .A(n883), .B(n18065), .ZN(n6971) );
  XNOR2_X1 U11057 ( .A(n6972), .B(n6971), .ZN(n6973) );
  XNOR2_X2 U11058 ( .A(n6974), .B(n6973), .ZN(n7967) );
  XNOR2_X1 U11059 ( .A(n7354), .B(n7288), .ZN(n6975) );
  XNOR2_X1 U11060 ( .A(n20209), .B(n6975), .ZN(n6981) );
  XNOR2_X1 U11061 ( .A(n6977), .B(n20227), .ZN(n6979) );
  XNOR2_X1 U11062 ( .A(n7026), .B(n16487), .ZN(n6978) );
  XNOR2_X1 U11063 ( .A(n6979), .B(n6978), .ZN(n6980) );
  XNOR2_X1 U11064 ( .A(n6981), .B(n6980), .ZN(n7487) );
  XNOR2_X1 U11065 ( .A(n6982), .B(n7047), .ZN(n6984) );
  XNOR2_X1 U11066 ( .A(n903), .B(n6839), .ZN(n6983) );
  XNOR2_X1 U11067 ( .A(n6984), .B(n6983), .ZN(n6989) );
  XNOR2_X1 U11068 ( .A(n7146), .B(n7318), .ZN(n6987) );
  XNOR2_X1 U11069 ( .A(n6985), .B(n18420), .ZN(n6986) );
  XNOR2_X1 U11070 ( .A(n6987), .B(n6986), .ZN(n6988) );
  XNOR2_X1 U11071 ( .A(n6989), .B(n6988), .ZN(n7971) );
  XNOR2_X1 U11072 ( .A(n6990), .B(n19027), .ZN(n6991) );
  XNOR2_X1 U11073 ( .A(n6993), .B(n7134), .ZN(n6994) );
  XNOR2_X1 U11074 ( .A(n6995), .B(n6996), .ZN(n7001) );
  XNOR2_X1 U11075 ( .A(n7017), .B(n2417), .ZN(n6999) );
  XNOR2_X1 U11076 ( .A(n6997), .B(n7128), .ZN(n6998) );
  XNOR2_X1 U11077 ( .A(n6999), .B(n6998), .ZN(n7000) );
  INV_X1 U11078 ( .A(n8527), .ZN(n8849) );
  INV_X1 U11079 ( .A(n7002), .ZN(n7753) );
  INV_X1 U11080 ( .A(n9046), .ZN(n8852) );
  XNOR2_X1 U11081 ( .A(n7201), .B(n17733), .ZN(n7005) );
  XNOR2_X1 U11082 ( .A(n7005), .B(n7264), .ZN(n7008) );
  XNOR2_X1 U11083 ( .A(n7006), .B(n7007), .ZN(n7204) );
  XNOR2_X1 U11084 ( .A(n7008), .B(n7204), .ZN(n7012) );
  XNOR2_X1 U11085 ( .A(n179), .B(n7267), .ZN(n7010) );
  XNOR2_X1 U11086 ( .A(n7010), .B(n7345), .ZN(n7011) );
  INV_X1 U11087 ( .A(n20165), .ZN(n7915) );
  INV_X1 U11088 ( .A(n7013), .ZN(n7015) );
  XNOR2_X1 U11089 ( .A(n7015), .B(n7014), .ZN(n7237) );
  XNOR2_X1 U11090 ( .A(n7016), .B(n7237), .ZN(n7022) );
  XNOR2_X1 U11091 ( .A(n7017), .B(n1869), .ZN(n7020) );
  XNOR2_X1 U11092 ( .A(n7195), .B(n7018), .ZN(n7019) );
  XNOR2_X1 U11093 ( .A(n7020), .B(n7019), .ZN(n7021) );
  XNOR2_X2 U11094 ( .A(n7022), .B(n7021), .ZN(n8910) );
  INV_X1 U11095 ( .A(n8910), .ZN(n8906) );
  XNOR2_X1 U11096 ( .A(n7355), .B(n7216), .ZN(n7024) );
  XNOR2_X1 U11097 ( .A(n7253), .B(n7221), .ZN(n7023) );
  XNOR2_X1 U11098 ( .A(n7024), .B(n7023), .ZN(n7030) );
  XNOR2_X1 U11099 ( .A(n7026), .B(n7025), .ZN(n7028) );
  XNOR2_X1 U11100 ( .A(n7028), .B(n7027), .ZN(n7029) );
  INV_X1 U11102 ( .A(n7836), .ZN(n7961) );
  XNOR2_X1 U11103 ( .A(n7212), .B(n7031), .ZN(n7034) );
  XNOR2_X1 U11104 ( .A(n7032), .B(n2384), .ZN(n7033) );
  XNOR2_X1 U11105 ( .A(n7034), .B(n7033), .ZN(n7038) );
  XNOR2_X1 U11106 ( .A(n7036), .B(n7229), .ZN(n7037) );
  XNOR2_X1 U11108 ( .A(n19944), .B(n7333), .ZN(n7039) );
  XNOR2_X1 U11109 ( .A(n7040), .B(n7039), .ZN(n7045) );
  XNOR2_X1 U11110 ( .A(n7041), .B(n7383), .ZN(n7246) );
  XNOR2_X1 U11111 ( .A(n7042), .B(n642), .ZN(n7043) );
  XNOR2_X1 U11112 ( .A(n7246), .B(n7043), .ZN(n7044) );
  XNOR2_X1 U11113 ( .A(n7045), .B(n7044), .ZN(n7956) );
  XNOR2_X1 U11114 ( .A(n7046), .B(n7047), .ZN(n7049) );
  XNOR2_X1 U11115 ( .A(n7048), .B(n7371), .ZN(n7277) );
  XNOR2_X1 U11116 ( .A(n7277), .B(n7049), .ZN(n7054) );
  XNOR2_X1 U11117 ( .A(n7050), .B(n7178), .ZN(n7052) );
  XNOR2_X1 U11118 ( .A(n7179), .B(n2448), .ZN(n7051) );
  XNOR2_X1 U11119 ( .A(n7052), .B(n7051), .ZN(n7053) );
  INV_X1 U11120 ( .A(n7958), .ZN(n7835) );
  NAND3_X1 U11121 ( .A1(n277), .A2(n7835), .A3(n8910), .ZN(n7055) );
  XNOR2_X1 U11122 ( .A(n7057), .B(n7058), .ZN(n7062) );
  XNOR2_X1 U11123 ( .A(n7154), .B(n18887), .ZN(n7059) );
  XNOR2_X1 U11124 ( .A(n7060), .B(n7059), .ZN(n7061) );
  XNOR2_X1 U11125 ( .A(n7062), .B(n7061), .ZN(n7096) );
  INV_X1 U11126 ( .A(n7096), .ZN(n7830) );
  XNOR2_X1 U11127 ( .A(n7127), .B(n7241), .ZN(n7063) );
  XNOR2_X1 U11128 ( .A(n7064), .B(n7063), .ZN(n7069) );
  XNOR2_X1 U11129 ( .A(n7065), .B(n2203), .ZN(n7067) );
  XNOR2_X1 U11130 ( .A(n7066), .B(n7067), .ZN(n7068) );
  XNOR2_X1 U11131 ( .A(n7070), .B(n17365), .ZN(n7072) );
  XNOR2_X1 U11132 ( .A(n7164), .B(n7266), .ZN(n7071) );
  XNOR2_X1 U11133 ( .A(n7072), .B(n7071), .ZN(n7076) );
  XNOR2_X1 U11134 ( .A(n7074), .B(n7073), .ZN(n7075) );
  XNOR2_X1 U11135 ( .A(n7078), .B(n7079), .ZN(n7085) );
  XNOR2_X1 U11136 ( .A(n7118), .B(n7080), .ZN(n7083) );
  XNOR2_X1 U11137 ( .A(n7081), .B(n2413), .ZN(n7082) );
  XNOR2_X1 U11138 ( .A(n7083), .B(n7082), .ZN(n7084) );
  NAND2_X1 U11139 ( .A1(n8014), .A2(n7086), .ZN(n7106) );
  XNOR2_X1 U11140 ( .A(n7087), .B(n7088), .ZN(n7090) );
  XNOR2_X1 U11141 ( .A(n7090), .B(n7089), .ZN(n7095) );
  XNOR2_X1 U11142 ( .A(n7273), .B(n7316), .ZN(n7093) );
  XNOR2_X1 U11143 ( .A(n7091), .B(n18366), .ZN(n7092) );
  XNOR2_X1 U11144 ( .A(n7093), .B(n7092), .ZN(n7094) );
  XNOR2_X1 U11145 ( .A(n7095), .B(n7094), .ZN(n8011) );
  NAND2_X1 U11146 ( .A1(n7830), .A2(n8012), .ZN(n7105) );
  XNOR2_X1 U11147 ( .A(n7097), .B(n19780), .ZN(n7099) );
  XNOR2_X1 U11148 ( .A(n7098), .B(n7099), .ZN(n7103) );
  XNOR2_X1 U11149 ( .A(n7249), .B(n7336), .ZN(n7101) );
  XNOR2_X1 U11150 ( .A(n7338), .B(n2164), .ZN(n7100) );
  XNOR2_X1 U11151 ( .A(n7101), .B(n7100), .ZN(n7102) );
  XNOR2_X1 U11152 ( .A(n7103), .B(n7102), .ZN(n7990) );
  INV_X1 U11153 ( .A(n7990), .ZN(n7829) );
  NAND3_X1 U11154 ( .A1(n7096), .A2(n7829), .A3(n8015), .ZN(n7104) );
  INV_X1 U11155 ( .A(n8851), .ZN(n7656) );
  NAND2_X1 U11156 ( .A1(n7919), .A2(n7768), .ZN(n7113) );
  INV_X1 U11157 ( .A(n7984), .ZN(n7534) );
  NAND2_X1 U11158 ( .A1(n7534), .A2(n7981), .ZN(n7108) );
  NAND3_X1 U11159 ( .A1(n7110), .A2(n19812), .A3(n7108), .ZN(n7112) );
  NAND3_X1 U11160 ( .A1(n505), .A2(n7921), .A3(n7984), .ZN(n7111) );
  OAI211_X1 U11161 ( .C1(n7978), .C2(n7113), .A(n7112), .B(n7111), .ZN(n8848)
         );
  INV_X1 U11162 ( .A(n8848), .ZN(n7659) );
  NOR2_X1 U11163 ( .A1(n9046), .A2(n7659), .ZN(n7114) );
  NAND2_X1 U11164 ( .A1(n7114), .A2(n8849), .ZN(n7173) );
  XNOR2_X1 U11165 ( .A(n6478), .B(n2394), .ZN(n7117) );
  XNOR2_X1 U11167 ( .A(n7118), .B(n1053), .ZN(n7119) );
  XNOR2_X1 U11168 ( .A(n7122), .B(n20227), .ZN(n7123) );
  XNOR2_X1 U11169 ( .A(n7126), .B(n7125), .ZN(n7132) );
  XNOR2_X1 U11170 ( .A(n7127), .B(n19953), .ZN(n7130) );
  XNOR2_X1 U11171 ( .A(n7128), .B(n1782), .ZN(n7129) );
  XNOR2_X1 U11172 ( .A(n7130), .B(n7129), .ZN(n7131) );
  XNOR2_X1 U11173 ( .A(n899), .B(n7134), .ZN(n7136) );
  XNOR2_X1 U11174 ( .A(n7136), .B(n7135), .ZN(n7141) );
  XNOR2_X1 U11175 ( .A(n6728), .B(n2442), .ZN(n7139) );
  XNOR2_X1 U11176 ( .A(n7137), .B(n7332), .ZN(n7138) );
  XNOR2_X1 U11177 ( .A(n7139), .B(n7138), .ZN(n7140) );
  XNOR2_X1 U11178 ( .A(n7141), .B(n7140), .ZN(n7952) );
  XNOR2_X1 U11179 ( .A(n7143), .B(n7142), .ZN(n7145) );
  XNOR2_X1 U11180 ( .A(n7317), .B(n7144), .ZN(n7176) );
  XNOR2_X1 U11181 ( .A(n7176), .B(n7145), .ZN(n7150) );
  XNOR2_X1 U11182 ( .A(n7146), .B(n18078), .ZN(n7147) );
  XNOR2_X1 U11183 ( .A(n7148), .B(n7147), .ZN(n7149) );
  XNOR2_X1 U11184 ( .A(n7149), .B(n7150), .ZN(n7951) );
  XNOR2_X1 U11185 ( .A(n7151), .B(n7211), .ZN(n7153) );
  XNOR2_X1 U11186 ( .A(n7152), .B(n7153), .ZN(n7159) );
  XNOR2_X1 U11187 ( .A(n19699), .B(n7154), .ZN(n7157) );
  XNOR2_X1 U11188 ( .A(n7155), .B(n18988), .ZN(n7156) );
  XNOR2_X1 U11189 ( .A(n7157), .B(n7156), .ZN(n7158) );
  XNOR2_X1 U11190 ( .A(n7159), .B(n7158), .ZN(n7481) );
  INV_X1 U11191 ( .A(n7481), .ZN(n7950) );
  INV_X1 U11193 ( .A(n7814), .ZN(n7169) );
  XNOR2_X1 U11194 ( .A(n7160), .B(n311), .ZN(n7161) );
  XNOR2_X1 U11195 ( .A(n7164), .B(n7163), .ZN(n7165) );
  XNOR2_X1 U11196 ( .A(n7305), .B(n7165), .ZN(n7166) );
  XNOR2_X2 U11197 ( .A(n7167), .B(n7166), .ZN(n7948) );
  NAND2_X1 U11198 ( .A1(n7169), .A2(n7168), .ZN(n7171) );
  INV_X1 U11199 ( .A(n7818), .ZN(n7170) );
  INV_X1 U11201 ( .A(n9039), .ZN(n8529) );
  NAND3_X1 U11202 ( .A1(n8529), .A2(n8527), .A3(n7656), .ZN(n7172) );
  NAND2_X1 U11203 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  XNOR2_X1 U11204 ( .A(n7177), .B(n7176), .ZN(n7183) );
  XNOR2_X1 U11205 ( .A(n903), .B(n7178), .ZN(n7181) );
  XNOR2_X1 U11206 ( .A(n7179), .B(n19336), .ZN(n7180) );
  XNOR2_X1 U11207 ( .A(n7181), .B(n7180), .ZN(n7182) );
  XNOR2_X1 U11208 ( .A(n7183), .B(n7182), .ZN(n7475) );
  XNOR2_X1 U11209 ( .A(n7332), .B(n7184), .ZN(n7186) );
  XNOR2_X1 U11210 ( .A(n7186), .B(n7185), .ZN(n7192) );
  XNOR2_X1 U11211 ( .A(n19944), .B(n7382), .ZN(n7190) );
  XNOR2_X1 U11212 ( .A(n7188), .B(n18779), .ZN(n7189) );
  XNOR2_X1 U11213 ( .A(n7190), .B(n7189), .ZN(n7191) );
  INV_X1 U11215 ( .A(n8315), .ZN(n8003) );
  INV_X1 U11216 ( .A(n7594), .ZN(n7227) );
  XNOR2_X1 U11217 ( .A(n7193), .B(n7194), .ZN(n7200) );
  XNOR2_X1 U11218 ( .A(n7195), .B(n19953), .ZN(n7198) );
  XNOR2_X1 U11219 ( .A(n7196), .B(n2329), .ZN(n7197) );
  XNOR2_X1 U11220 ( .A(n7198), .B(n7197), .ZN(n7199) );
  XNOR2_X1 U11222 ( .A(n7201), .B(n16030), .ZN(n7203) );
  XNOR2_X1 U11223 ( .A(n7203), .B(n7202), .ZN(n7205) );
  XNOR2_X1 U11224 ( .A(n7205), .B(n7204), .ZN(n7209) );
  XNOR2_X1 U11225 ( .A(n7348), .B(n7206), .ZN(n7207) );
  XNOR2_X1 U11226 ( .A(n7305), .B(n7207), .ZN(n7208) );
  XNOR2_X1 U11227 ( .A(n7209), .B(n7208), .ZN(n7591) );
  XNOR2_X1 U11228 ( .A(n7212), .B(n7211), .ZN(n7213) );
  OAI211_X1 U11229 ( .C1(n7592), .C2(n8313), .A(n8004), .B(n8315), .ZN(n7226)
         );
  XNOR2_X1 U11230 ( .A(n7217), .B(n7216), .ZN(n7220) );
  XNOR2_X1 U11231 ( .A(n7218), .B(n7354), .ZN(n7219) );
  XNOR2_X1 U11232 ( .A(n7220), .B(n7219), .ZN(n7224) );
  XNOR2_X1 U11233 ( .A(n1052), .B(n7221), .ZN(n7222) );
  XNOR2_X1 U11234 ( .A(n20203), .B(n7222), .ZN(n7223) );
  XNOR2_X1 U11235 ( .A(n7224), .B(n7223), .ZN(n8316) );
  NAND2_X1 U11237 ( .A1(n19520), .A2(n8313), .ZN(n7225) );
  XNOR2_X1 U11238 ( .A(n7228), .B(n7229), .ZN(n7236) );
  XNOR2_X1 U11239 ( .A(n7230), .B(n18854), .ZN(n7234) );
  XNOR2_X1 U11240 ( .A(n19841), .B(n7232), .ZN(n7233) );
  XNOR2_X1 U11241 ( .A(n7234), .B(n7233), .ZN(n7235) );
  INV_X1 U11242 ( .A(n7237), .ZN(n7239) );
  XNOR2_X1 U11243 ( .A(n7239), .B(n7238), .ZN(n7245) );
  XNOR2_X1 U11244 ( .A(n7240), .B(n7241), .ZN(n7243) );
  XNOR2_X1 U11245 ( .A(n6777), .B(n18055), .ZN(n7242) );
  XNOR2_X1 U11246 ( .A(n7243), .B(n7242), .ZN(n7244) );
  XNOR2_X1 U11247 ( .A(n7249), .B(n7248), .ZN(n7251) );
  XNOR2_X1 U11248 ( .A(n6249), .B(n2108), .ZN(n7250) );
  XNOR2_X1 U11249 ( .A(n7251), .B(n7250), .ZN(n7252) );
  XNOR2_X1 U11250 ( .A(n7254), .B(n7253), .ZN(n7255) );
  XNOR2_X1 U11251 ( .A(n7256), .B(n7255), .ZN(n7262) );
  XNOR2_X1 U11252 ( .A(n7025), .B(n7257), .ZN(n7260) );
  XNOR2_X1 U11253 ( .A(n7258), .B(n2032), .ZN(n7259) );
  XNOR2_X1 U11254 ( .A(n7260), .B(n7259), .ZN(n7261) );
  XNOR2_X1 U11255 ( .A(n7261), .B(n7262), .ZN(n7466) );
  INV_X1 U11256 ( .A(n7963), .ZN(n7283) );
  INV_X1 U11257 ( .A(n2192), .ZN(n17940) );
  XNOR2_X1 U11258 ( .A(n7263), .B(n17940), .ZN(n7265) );
  XNOR2_X1 U11259 ( .A(n7265), .B(n7264), .ZN(n7269) );
  XNOR2_X1 U11260 ( .A(n7266), .B(n7267), .ZN(n7268) );
  XNOR2_X1 U11261 ( .A(n7269), .B(n7268), .ZN(n7271) );
  XNOR2_X1 U11262 ( .A(n7271), .B(n7270), .ZN(n7965) );
  INV_X1 U11263 ( .A(n7965), .ZN(n8018) );
  XNOR2_X1 U11264 ( .A(n7272), .B(n17095), .ZN(n7276) );
  XNOR2_X1 U11265 ( .A(n7273), .B(n7274), .ZN(n7275) );
  XNOR2_X1 U11266 ( .A(n7276), .B(n7275), .ZN(n7281) );
  INV_X1 U11267 ( .A(n7277), .ZN(n7278) );
  XNOR2_X1 U11268 ( .A(n7279), .B(n7278), .ZN(n7280) );
  NOR2_X1 U11271 ( .A1(n20347), .A2(n20490), .ZN(n7282) );
  AOI22_X1 U11272 ( .A1(n7283), .A2(n8018), .B1(n208), .B2(n7282), .ZN(n7284)
         );
  XNOR2_X1 U11273 ( .A(n1052), .B(n7288), .ZN(n7291) );
  XNOR2_X1 U11274 ( .A(n7289), .B(n2310), .ZN(n7290) );
  XNOR2_X1 U11275 ( .A(n7291), .B(n7290), .ZN(n7292) );
  XNOR2_X1 U11276 ( .A(n7295), .B(n7294), .ZN(n7302) );
  XNOR2_X1 U11277 ( .A(n7296), .B(n19953), .ZN(n7300) );
  XNOR2_X1 U11278 ( .A(n7298), .B(n18768), .ZN(n7299) );
  XNOR2_X1 U11279 ( .A(n7300), .B(n7299), .ZN(n7301) );
  XNOR2_X1 U11280 ( .A(n7302), .B(n7301), .ZN(n7312) );
  NAND2_X1 U11281 ( .A1(n1425), .A2(n7312), .ZN(n7343) );
  XNOR2_X1 U11282 ( .A(n7306), .B(n17544), .ZN(n7307) );
  XNOR2_X1 U11283 ( .A(n7308), .B(n7307), .ZN(n7309) );
  XNOR2_X1 U11284 ( .A(n7310), .B(n7309), .ZN(n7311) );
  INV_X1 U11285 ( .A(n7312), .ZN(n8001) );
  INV_X1 U11286 ( .A(n7313), .ZN(n7314) );
  XNOR2_X1 U11287 ( .A(n7314), .B(n7315), .ZN(n7322) );
  XNOR2_X1 U11288 ( .A(n7317), .B(n7316), .ZN(n7320) );
  XNOR2_X1 U11289 ( .A(n7318), .B(n345), .ZN(n7319) );
  XNOR2_X1 U11290 ( .A(n7320), .B(n7319), .ZN(n7321) );
  XNOR2_X1 U11291 ( .A(n7323), .B(n7324), .ZN(n7331) );
  XNOR2_X1 U11292 ( .A(n883), .B(n18726), .ZN(n7329) );
  XNOR2_X1 U11293 ( .A(n7326), .B(n19698), .ZN(n7328) );
  XNOR2_X1 U11294 ( .A(n7328), .B(n7329), .ZN(n7330) );
  XNOR2_X1 U11295 ( .A(n7331), .B(n7330), .ZN(n7585) );
  XNOR2_X1 U11296 ( .A(n7332), .B(n7333), .ZN(n7335) );
  XNOR2_X1 U11297 ( .A(n7335), .B(n7334), .ZN(n7342) );
  XNOR2_X1 U11298 ( .A(n7337), .B(n7336), .ZN(n7340) );
  XNOR2_X1 U11299 ( .A(n7338), .B(n17804), .ZN(n7339) );
  XNOR2_X1 U11300 ( .A(n7340), .B(n7339), .ZN(n7341) );
  MUX2_X1 U11301 ( .A(n8925), .B(n8932), .S(n8928), .Z(n7413) );
  XNOR2_X1 U11302 ( .A(n7345), .B(n7344), .ZN(n7347) );
  XNOR2_X1 U11303 ( .A(n7346), .B(n7347), .ZN(n7351) );
  XNOR2_X1 U11304 ( .A(n7348), .B(n18070), .ZN(n7349) );
  XNOR2_X1 U11305 ( .A(n7025), .B(n2383), .ZN(n7352) );
  XNOR2_X1 U11306 ( .A(n7352), .B(n7353), .ZN(n7359) );
  XNOR2_X1 U11307 ( .A(n7355), .B(n7354), .ZN(n7357) );
  XNOR2_X1 U11308 ( .A(n7357), .B(n7356), .ZN(n7358) );
  XNOR2_X1 U11309 ( .A(n7359), .B(n7358), .ZN(n8025) );
  XNOR2_X1 U11310 ( .A(n7361), .B(n7362), .ZN(n7369) );
  XNOR2_X1 U11311 ( .A(n7364), .B(n7363), .ZN(n7367) );
  XNOR2_X1 U11312 ( .A(n7365), .B(n17993), .ZN(n7366) );
  XNOR2_X1 U11313 ( .A(n7367), .B(n7366), .ZN(n7368) );
  XNOR2_X1 U11314 ( .A(n7368), .B(n7369), .ZN(n7389) );
  INV_X1 U11315 ( .A(n7389), .ZN(n8290) );
  OAI21_X1 U11316 ( .B1(n8293), .B2(n20189), .A(n7370), .ZN(n7401) );
  XNOR2_X1 U11317 ( .A(n7371), .B(n903), .ZN(n7375) );
  XNOR2_X1 U11318 ( .A(n7373), .B(n19436), .ZN(n7374) );
  XNOR2_X1 U11319 ( .A(n7375), .B(n7374), .ZN(n7379) );
  XNOR2_X1 U11320 ( .A(n7377), .B(n7376), .ZN(n7378) );
  XNOR2_X1 U11321 ( .A(n7378), .B(n7379), .ZN(n8288) );
  XNOR2_X1 U11322 ( .A(n7382), .B(n7383), .ZN(n7386) );
  XNOR2_X1 U11323 ( .A(n7384), .B(n18809), .ZN(n7385) );
  XNOR2_X1 U11324 ( .A(n7386), .B(n7385), .ZN(n7387) );
  XNOR2_X1 U11325 ( .A(n7390), .B(n7391), .ZN(n7394) );
  XNOR2_X1 U11326 ( .A(n7392), .B(n18819), .ZN(n7393) );
  XNOR2_X1 U11327 ( .A(n7394), .B(n7393), .ZN(n7399) );
  INV_X1 U11328 ( .A(n7395), .ZN(n7396) );
  XNOR2_X1 U11329 ( .A(n7397), .B(n7396), .ZN(n7398) );
  NAND2_X1 U11330 ( .A1(n8928), .A2(n8932), .ZN(n7662) );
  OAI21_X1 U11331 ( .B1(n7950), .B2(n2326), .A(n7951), .ZN(n7404) );
  NAND2_X1 U11332 ( .A1(n8596), .A2(n8931), .ZN(n7406) );
  OAI21_X1 U11333 ( .B1(n7662), .B2(n8931), .A(n7406), .ZN(n7411) );
  OAI211_X1 U11334 ( .C1(n7826), .C2(n7830), .A(n7407), .B(n8012), .ZN(n7410)
         );
  OAI21_X1 U11335 ( .B1(n7826), .B2(n7829), .A(n8011), .ZN(n7409) );
  NAND2_X1 U11336 ( .A1(n8749), .A2(n8748), .ZN(n8640) );
  NAND2_X1 U11337 ( .A1(n7411), .A2(n8640), .ZN(n7412) );
  OAI21_X1 U11338 ( .B1(n7413), .B2(n8596), .A(n7412), .ZN(n10299) );
  NOR2_X1 U11339 ( .A1(n8178), .A2(n19901), .ZN(n7415) );
  OAI21_X1 U11340 ( .B1(n7416), .B2(n7415), .A(n923), .ZN(n7419) );
  NOR2_X1 U11341 ( .A1(n8069), .A2(n8179), .ZN(n7418) );
  INV_X1 U11342 ( .A(n7420), .ZN(n8201) );
  AOI21_X1 U11344 ( .B1(n7615), .B2(n7422), .A(n8201), .ZN(n7423) );
  NAND2_X1 U11345 ( .A1(n9300), .A2(n9018), .ZN(n7424) );
  INV_X1 U11346 ( .A(n7644), .ZN(n8215) );
  NAND2_X1 U11348 ( .A1(n20108), .A2(n8086), .ZN(n7425) );
  NOR2_X1 U11349 ( .A1(n20107), .A2(n6539), .ZN(n7426) );
  INV_X1 U11350 ( .A(n20108), .ZN(n8084) );
  NAND2_X1 U11351 ( .A1(n8084), .A2(n8085), .ZN(n8236) );
  INV_X1 U11352 ( .A(n8236), .ZN(n7428) );
  NAND2_X1 U11353 ( .A1(n7631), .A2(n8212), .ZN(n7431) );
  NAND2_X1 U11354 ( .A1(n8094), .A2(n8211), .ZN(n7430) );
  MUX2_X1 U11355 ( .A(n7431), .B(n7430), .S(n8095), .Z(n7435) );
  INV_X1 U11357 ( .A(n8211), .ZN(n8093) );
  INV_X1 U11358 ( .A(n8098), .ZN(n7638) );
  INV_X1 U11359 ( .A(n8111), .ZN(n8237) );
  MUX2_X1 U11360 ( .A(n3775), .B(n7436), .S(n20493), .Z(n7437) );
  INV_X1 U11362 ( .A(n9304), .ZN(n8845) );
  MUX2_X1 U11364 ( .A(n8323), .B(n7441), .S(n1425), .Z(n8512) );
  OAI21_X1 U11365 ( .B1(n7590), .B2(n7442), .A(n7584), .ZN(n8513) );
  BUF_X2 U11366 ( .A(n7443), .Z(n8282) );
  NAND3_X1 U11367 ( .A1(n8286), .A2(n7603), .A3(n8282), .ZN(n7449) );
  NAND3_X1 U11368 ( .A1(n7444), .A2(n3660), .A3(n7445), .ZN(n7448) );
  NAND3_X1 U11369 ( .A1(n7444), .A2(n8281), .A3(n7600), .ZN(n7447) );
  INV_X1 U11370 ( .A(n8033), .ZN(n8284) );
  NAND3_X1 U11371 ( .A1(n8284), .A2(n8280), .A3(n7445), .ZN(n7446) );
  AND4_X1 U11372 ( .A1(n7448), .A2(n7449), .A3(n7447), .A4(n7446), .ZN(n9021)
         );
  INV_X1 U11373 ( .A(n7877), .ZN(n8305) );
  INV_X1 U11376 ( .A(n20257), .ZN(n7789) );
  INV_X1 U11378 ( .A(n8040), .ZN(n7581) );
  NAND3_X1 U11379 ( .A1(n8297), .A2(n20243), .A3(n7581), .ZN(n7454) );
  MUX2_X1 U11380 ( .A(n20243), .B(n8297), .S(n8298), .Z(n7455) );
  INV_X1 U11381 ( .A(n8676), .ZN(n8841) );
  NAND2_X1 U11382 ( .A1(n8054), .A2(n8193), .ZN(n7456) );
  NOR2_X1 U11383 ( .A1(n8052), .A2(n8192), .ZN(n7458) );
  AOI22_X1 U11384 ( .A1(n7458), .A2(n19802), .B1(n19474), .B2(n8197), .ZN(
        n7459) );
  INV_X1 U11385 ( .A(n8060), .ZN(n7460) );
  NAND2_X1 U11386 ( .A1(n7460), .A2(n8190), .ZN(n8183) );
  INV_X1 U11387 ( .A(n8185), .ZN(n8059) );
  NAND3_X1 U11388 ( .A1(n7462), .A2(n20465), .A3(n8059), .ZN(n7464) );
  NAND3_X1 U11389 ( .A1(n8185), .A2(n7893), .A3(n8184), .ZN(n7463) );
  XNOR2_X1 U11390 ( .A(n9602), .B(n10482), .ZN(n9984) );
  INV_X1 U11391 ( .A(n8025), .ZN(n8292) );
  INV_X1 U11392 ( .A(n8026), .ZN(n8024) );
  INV_X1 U11393 ( .A(n8288), .ZN(n7468) );
  NAND2_X1 U11394 ( .A1(n8292), .A2(n8026), .ZN(n8031) );
  NAND2_X1 U11395 ( .A1(n8290), .A2(n8289), .ZN(n8029) );
  NAND2_X1 U11396 ( .A1(n7470), .A2(n8024), .ZN(n7471) );
  NAND2_X1 U11397 ( .A1(n7096), .A2(n7990), .ZN(n7994) );
  NAND3_X1 U11398 ( .A1(n7096), .A2(n8011), .A3(n20154), .ZN(n7472) );
  NAND2_X1 U11399 ( .A1(n8316), .A2(n7591), .ZN(n8007) );
  INV_X1 U11400 ( .A(n8007), .ZN(n7474) );
  NOR2_X1 U11401 ( .A1(n8004), .A2(n7591), .ZN(n7473) );
  OAI21_X1 U11402 ( .B1(n7474), .B2(n7473), .A(n8313), .ZN(n7478) );
  INV_X1 U11404 ( .A(n8004), .ZN(n7476) );
  OAI21_X1 U11405 ( .B1(n8811), .B2(n8810), .A(n8815), .ZN(n7486) );
  NAND3_X1 U11407 ( .A1(n7479), .A2(n20013), .A3(n7948), .ZN(n7484) );
  NOR2_X1 U11408 ( .A1(n7952), .A2(n7951), .ZN(n7480) );
  INV_X1 U11409 ( .A(n7951), .ZN(n7815) );
  NAND3_X1 U11410 ( .A1(n7949), .A2(n7951), .A3(n7953), .ZN(n7482) );
  AND2_X1 U11411 ( .A1(n8812), .A2(n8815), .ZN(n7485) );
  INV_X1 U11412 ( .A(n8811), .ZN(n9119) );
  AOI22_X1 U11413 ( .A1(n8818), .A2(n7486), .B1(n7485), .B2(n9119), .ZN(n7492)
         );
  NAND2_X1 U11414 ( .A1(n7487), .A2(n7974), .ZN(n7970) );
  INV_X1 U11415 ( .A(n7972), .ZN(n7927) );
  OAI22_X1 U11416 ( .A1(n7970), .A2(n7927), .B1(n278), .B2(n7968), .ZN(n7490)
         );
  INV_X1 U11417 ( .A(n7487), .ZN(n7973) );
  NAND2_X1 U11418 ( .A1(n7973), .A2(n7967), .ZN(n7489) );
  NAND2_X1 U11419 ( .A1(n7972), .A2(n278), .ZN(n7488) );
  NOR2_X1 U11420 ( .A1(n8550), .A2(n9122), .ZN(n9120) );
  NAND2_X1 U11421 ( .A1(n9120), .A2(n8812), .ZN(n7491) );
  INV_X1 U11422 ( .A(n7493), .ZN(n8344) );
  MUX2_X1 U11423 ( .A(n8166), .B(n8344), .S(n8342), .Z(n7495) );
  NOR2_X1 U11424 ( .A1(n8340), .A2(n8343), .ZN(n7494) );
  AND3_X1 U11426 ( .A1(n8340), .A2(n8341), .A3(n7679), .ZN(n9048) );
  INV_X1 U11427 ( .A(n9289), .ZN(n9577) );
  INV_X1 U11428 ( .A(n8387), .ZN(n7496) );
  AOI21_X1 U11429 ( .B1(n7497), .B2(n7496), .A(n20177), .ZN(n7499) );
  INV_X1 U11430 ( .A(n7686), .ZN(n8382) );
  NAND2_X1 U11431 ( .A1(n8359), .A2(n8354), .ZN(n7740) );
  NAND3_X1 U11432 ( .A1(n7501), .A2(n7740), .A3(n7500), .ZN(n7503) );
  NAND3_X1 U11433 ( .A1(n8355), .A2(n8358), .A3(n7504), .ZN(n7502) );
  AOI22_X1 U11435 ( .A1(n2031), .A2(n20360), .B1(n20195), .B2(n7763), .ZN(
        n7505) );
  NAND2_X1 U11436 ( .A1(n2540), .A2(n7936), .ZN(n7506) );
  OAI211_X1 U11437 ( .C1(n7746), .C2(n7749), .A(n7911), .B(n7910), .ZN(n7509)
         );
  NAND2_X1 U11438 ( .A1(n7510), .A2(n7675), .ZN(n7511) );
  NAND3_X1 U11439 ( .A1(n8366), .A2(n7709), .A3(n8365), .ZN(n7514) );
  NAND2_X1 U11440 ( .A1(n9049), .A2(n9576), .ZN(n7515) );
  AOI21_X1 U11441 ( .B1(n9287), .B2(n7515), .A(n19896), .ZN(n7516) );
  AOI21_X2 U11442 ( .B1(n9577), .B2(n20196), .A(n7516), .ZN(n9983) );
  XNOR2_X1 U11443 ( .A(n10028), .B(n9983), .ZN(n7517) );
  XNOR2_X1 U11444 ( .A(n9984), .B(n7517), .ZN(n7580) );
  INV_X1 U11445 ( .A(n7956), .ZN(n7834) );
  MUX2_X1 U11446 ( .A(n277), .B(n7834), .S(n7958), .Z(n8907) );
  AOI21_X1 U11449 ( .B1(n7760), .B2(n7519), .A(n2030), .ZN(n8908) );
  AND2_X1 U11450 ( .A1(n7520), .A2(n2031), .ZN(n8909) );
  NAND2_X1 U11451 ( .A1(n8923), .A2(n8917), .ZN(n7533) );
  INV_X1 U11452 ( .A(n7974), .ZN(n7820) );
  NAND2_X1 U11454 ( .A1(n7523), .A2(n7970), .ZN(n8733) );
  INV_X1 U11455 ( .A(n7948), .ZN(n7819) );
  OAI21_X1 U11456 ( .B1(n7819), .B2(n20013), .A(n7815), .ZN(n7524) );
  NAND2_X1 U11457 ( .A1(n7524), .A2(n7949), .ZN(n7526) );
  NAND3_X1 U11458 ( .A1(n7819), .A2(n7950), .A3(n7952), .ZN(n7525) );
  OAI211_X1 U11459 ( .C1(n7818), .C2(n7948), .A(n7526), .B(n7525), .ZN(n8735)
         );
  NAND2_X1 U11460 ( .A1(n7909), .A2(n7903), .ZN(n7527) );
  OAI21_X1 U11461 ( .B1(n7909), .B2(n7754), .A(n7527), .ZN(n7529) );
  NOR2_X1 U11462 ( .A1(n7754), .A2(n7902), .ZN(n7528) );
  AND3_X1 U11463 ( .A1(n7754), .A2(n19521), .A3(n7530), .ZN(n7531) );
  INV_X1 U11464 ( .A(n7981), .ZN(n7766) );
  NAND3_X1 U11465 ( .A1(n7920), .A2(n7536), .A3(n7921), .ZN(n7535) );
  AOI21_X1 U11466 ( .B1(n9158), .B2(n8696), .A(n9159), .ZN(n7540) );
  INV_X1 U11467 ( .A(n9164), .ZN(n7537) );
  NOR2_X1 U11468 ( .A1(n7537), .A2(n9163), .ZN(n9157) );
  NAND2_X1 U11469 ( .A1(n9157), .A2(n8611), .ZN(n7539) );
  NAND3_X1 U11470 ( .A1(n1230), .A2(n8696), .A3(n9161), .ZN(n7538) );
  XNOR2_X1 U11472 ( .A(n10620), .B(n9947), .ZN(n9416) );
  NOR2_X1 U11474 ( .A1(n7541), .A2(n8372), .ZN(n7546) );
  INV_X1 U11475 ( .A(n8376), .ZN(n7703) );
  NAND3_X1 U11476 ( .A1(n8372), .A2(n20252), .A3(n8377), .ZN(n7543) );
  NAND3_X1 U11477 ( .A1(n7544), .A2(n7543), .A3(n8369), .ZN(n7545) );
  INV_X1 U11478 ( .A(n8352), .ZN(n7717) );
  OAI22_X1 U11479 ( .A1(n7717), .A2(n8140), .B1(n19914), .B2(n8347), .ZN(n8351) );
  INV_X1 U11480 ( .A(n8270), .ZN(n7549) );
  NOR2_X1 U11481 ( .A1(n8349), .A2(n8348), .ZN(n7548) );
  INV_X1 U11482 ( .A(n8350), .ZN(n8268) );
  NAND2_X1 U11483 ( .A1(n8268), .A2(n8140), .ZN(n7547) );
  NAND2_X1 U11484 ( .A1(n7724), .A2(n282), .ZN(n7551) );
  NAND2_X1 U11485 ( .A1(n7552), .A2(n7855), .ZN(n7555) );
  NAND3_X1 U11486 ( .A1(n7856), .A2(n7851), .A3(n7852), .ZN(n7553) );
  NAND2_X1 U11488 ( .A1(n7559), .A2(n9364), .ZN(n7567) );
  AND2_X1 U11489 ( .A1(n7560), .A2(n8114), .ZN(n7843) );
  NOR2_X1 U11490 ( .A1(n7560), .A2(n6704), .ZN(n7561) );
  OAI21_X1 U11491 ( .B1(n7843), .B2(n7561), .A(n8245), .ZN(n7566) );
  NOR2_X1 U11493 ( .A1(n7844), .A2(n8114), .ZN(n7563) );
  AOI22_X1 U11494 ( .A1(n7564), .A2(n20251), .B1(n7563), .B2(n6704), .ZN(n7565) );
  NAND2_X1 U11495 ( .A1(n7567), .A2(n9362), .ZN(n7577) );
  NOR2_X1 U11496 ( .A1(n8961), .A2(n8960), .ZN(n7575) );
  MUX2_X1 U11497 ( .A(n8264), .B(n8263), .S(n895), .Z(n7569) );
  INV_X1 U11498 ( .A(n8104), .ZN(n7570) );
  NAND2_X1 U11499 ( .A1(n7570), .A2(n8262), .ZN(n7573) );
  AND3_X2 U11500 ( .A1(n7574), .A2(n7573), .A3(n7572), .ZN(n8958) );
  INV_X1 U11501 ( .A(n8958), .ZN(n7653) );
  AOI22_X1 U11502 ( .A1(n7575), .A2(n7653), .B1(n8959), .B2(n8726), .ZN(n7576)
         );
  XNOR2_X1 U11503 ( .A(n9802), .B(n2344), .ZN(n7578) );
  XNOR2_X1 U11504 ( .A(n9416), .B(n7578), .ZN(n7579) );
  XNOR2_X1 U11505 ( .A(n7580), .B(n7579), .ZN(n9492) );
  INV_X1 U11506 ( .A(n9492), .ZN(n11160) );
  MUX2_X2 U11507 ( .A(n7583), .B(n7582), .S(n8299), .Z(n8947) );
  INV_X1 U11509 ( .A(n7585), .ZN(n8322) );
  NAND2_X1 U11510 ( .A1(n8322), .A2(n8001), .ZN(n7586) );
  OAI211_X1 U11511 ( .C1(n1425), .C2(n8322), .A(n7586), .B(n8325), .ZN(n7587)
         );
  INV_X1 U11513 ( .A(n8644), .ZN(n7608) );
  INV_X1 U11514 ( .A(n7591), .ZN(n7592) );
  NAND2_X1 U11515 ( .A1(n7593), .A2(n8316), .ZN(n7596) );
  NAND2_X1 U11516 ( .A1(n7594), .A2(n7592), .ZN(n7595) );
  NAND2_X1 U11517 ( .A1(n7608), .A2(n8937), .ZN(n7613) );
  NAND3_X1 U11518 ( .A1(n8304), .A2(n8046), .A3(n8305), .ZN(n7598) );
  NOR2_X1 U11519 ( .A1(n8286), .A2(n19686), .ZN(n7795) );
  NAND3_X1 U11521 ( .A1(n8033), .A2(n8282), .A3(n8281), .ZN(n7604) );
  NAND3_X1 U11523 ( .A1(n8185), .A2(n20247), .A3(n20465), .ZN(n7607) );
  NAND2_X1 U11525 ( .A1(n7610), .A2(n8730), .ZN(n7611) );
  XNOR2_X1 U11526 ( .A(n10054), .B(n1782), .ZN(n7655) );
  INV_X1 U11527 ( .A(n7615), .ZN(n8203) );
  NAND3_X1 U11528 ( .A1(n8201), .A2(n7421), .A3(n8204), .ZN(n7617) );
  INV_X1 U11529 ( .A(n8743), .ZN(n8949) );
  INV_X1 U11530 ( .A(n7887), .ZN(n7620) );
  NOR2_X1 U11531 ( .A1(n8179), .A2(n923), .ZN(n7619) );
  AOI22_X1 U11532 ( .A1(n7620), .A2(n8068), .B1(n7622), .B2(n7619), .ZN(n7625)
         );
  INV_X1 U11533 ( .A(n7621), .ZN(n8176) );
  NAND2_X1 U11534 ( .A1(n8176), .A2(n8179), .ZN(n7623) );
  INV_X1 U11535 ( .A(n8178), .ZN(n7622) );
  INV_X1 U11536 ( .A(n8197), .ZN(n7879) );
  AOI21_X1 U11537 ( .B1(n7628), .B2(n7627), .A(n8051), .ZN(n7629) );
  NAND2_X1 U11539 ( .A1(n8090), .A2(n7633), .ZN(n7634) );
  NOR2_X1 U11540 ( .A1(n8241), .A2(n8112), .ZN(n7637) );
  NAND2_X1 U11541 ( .A1(n7637), .A2(n3775), .ZN(n7643) );
  INV_X1 U11542 ( .A(n8241), .ZN(n7639) );
  NAND3_X1 U11543 ( .A1(n8239), .A2(n7639), .A3(n7638), .ZN(n7642) );
  NAND3_X1 U11544 ( .A1(n8099), .A2(n8100), .A3(n8241), .ZN(n7641) );
  NAND2_X1 U11545 ( .A1(n8099), .A2(n8237), .ZN(n7640) );
  AND2_X1 U11546 ( .A1(n8603), .A2(n8741), .ZN(n8485) );
  INV_X1 U11547 ( .A(n8485), .ZN(n7650) );
  INV_X1 U11548 ( .A(n8741), .ZN(n8953) );
  OAI22_X1 U11549 ( .A1(n20441), .A2(n7645), .B1(n8220), .B2(n7644), .ZN(n7847) );
  INV_X1 U11550 ( .A(n7646), .ZN(n7647) );
  INV_X1 U11551 ( .A(n8742), .ZN(n8950) );
  NAND2_X1 U11552 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  INV_X1 U11553 ( .A(n9362), .ZN(n7654) );
  XNOR2_X1 U11554 ( .A(n10566), .B(n10456), .ZN(n10017) );
  XNOR2_X1 U11555 ( .A(n7655), .B(n10017), .ZN(n7664) );
  OAI21_X1 U11556 ( .B1(n8527), .B2(n8848), .A(n9046), .ZN(n7657) );
  NAND2_X1 U11557 ( .A1(n8749), .A2(n8747), .ZN(n7661) );
  INV_X1 U11558 ( .A(n8932), .ZN(n8638) );
  NAND3_X1 U11559 ( .A1(n8638), .A2(n8749), .A3(n8925), .ZN(n7660) );
  XNOR2_X1 U11560 ( .A(n9430), .B(n10163), .ZN(n7663) );
  INV_X1 U11561 ( .A(n8499), .ZN(n7666) );
  INV_X1 U11562 ( .A(n8733), .ZN(n8497) );
  NOR2_X1 U11563 ( .A1(n8499), .A2(n8734), .ZN(n8738) );
  MUX2_X1 U11564 ( .A(n7665), .B(n8738), .S(n8736), .Z(n7670) );
  NAND2_X1 U11565 ( .A1(n19518), .A2(n8736), .ZN(n7667) );
  INV_X1 U11566 ( .A(n8736), .ZN(n8916) );
  AOI22_X1 U11567 ( .A1(n7668), .A2(n7667), .B1(n7666), .B2(n8916), .ZN(n7669)
         );
  OAI21_X1 U11569 ( .B1(n8146), .B2(n7671), .A(n8370), .ZN(n7672) );
  MUX2_X1 U11570 ( .A(n7673), .B(n7709), .S(n6951), .Z(n7678) );
  INV_X1 U11571 ( .A(n7674), .ZN(n7708) );
  INV_X1 U11572 ( .A(n8342), .ZN(n8167) );
  MUX2_X1 U11573 ( .A(n2964), .B(n7679), .S(n8343), .Z(n7682) );
  NAND3_X1 U11574 ( .A1(n8167), .A2(n8165), .A3(n7679), .ZN(n7681) );
  NOR2_X1 U11575 ( .A1(n8340), .A2(n7679), .ZN(n7733) );
  NAND2_X1 U11576 ( .A1(n7733), .A2(n8341), .ZN(n7680) );
  INV_X1 U11579 ( .A(n8386), .ZN(n7683) );
  INV_X1 U11580 ( .A(n8380), .ZN(n8133) );
  OAI21_X1 U11581 ( .B1(n8132), .B2(n7683), .A(n8133), .ZN(n7688) );
  INV_X1 U11583 ( .A(n7714), .ZN(n7687) );
  MUX2_X1 U11584 ( .A(n9358), .B(n19941), .S(n9528), .Z(n7702) );
  OAI21_X1 U11585 ( .B1(n7746), .B2(n3445), .A(n7748), .ZN(n7693) );
  NOR2_X1 U11586 ( .A1(n7748), .A2(n7910), .ZN(n7690) );
  OAI21_X1 U11587 ( .B1(n7691), .B2(n7690), .A(n7914), .ZN(n7692) );
  NAND2_X1 U11589 ( .A1(n9354), .A2(n8904), .ZN(n8492) );
  NAND3_X1 U11592 ( .A1(n7696), .A2(n7695), .A3(n8355), .ZN(n7697) );
  AOI21_X2 U11593 ( .B1(n9359), .B2(n7702), .A(n7701), .ZN(n10203) );
  XNOR2_X1 U11594 ( .A(n10200), .B(n10203), .ZN(n10596) );
  NAND2_X1 U11596 ( .A1(n7703), .A2(n7671), .ZN(n7704) );
  MUX2_X1 U11597 ( .A(n7705), .B(n7704), .S(n8373), .Z(n7706) );
  MUX2_X1 U11599 ( .A(n8366), .B(n8361), .S(n7674), .Z(n7712) );
  NAND3_X1 U11600 ( .A1(n8361), .A2(n7709), .A3(n7708), .ZN(n7710) );
  INV_X1 U11601 ( .A(n8879), .ZN(n9255) );
  AOI21_X1 U11602 ( .B1(n8132), .B2(n8381), .A(n8387), .ZN(n7713) );
  OAI22_X1 U11603 ( .A1(n7714), .A2(n7713), .B1(n163), .B2(n8131), .ZN(n7715)
         );
  OAI21_X1 U11604 ( .B1(n20177), .B2(n7716), .A(n7715), .ZN(n9250) );
  NAND2_X1 U11605 ( .A1(n20200), .A2(n8271), .ZN(n7719) );
  NAND2_X1 U11606 ( .A1(n8348), .A2(n8347), .ZN(n7718) );
  NAND3_X1 U11607 ( .A1(n7723), .A2(n7719), .A3(n7718), .ZN(n7721) );
  OAI211_X1 U11608 ( .C1(n7723), .C2(n7722), .A(n7721), .B(n7720), .ZN(n8972)
         );
  AND2_X1 U11609 ( .A1(n9252), .A2(n8972), .ZN(n7727) );
  NAND2_X1 U11610 ( .A1(n8167), .A2(n7728), .ZN(n7732) );
  NOR2_X1 U11611 ( .A1(n8341), .A2(n8344), .ZN(n7731) );
  INV_X1 U11612 ( .A(n7729), .ZN(n7730) );
  OAI21_X1 U11613 ( .B1(n7732), .B2(n7731), .A(n7730), .ZN(n7735) );
  NAND2_X1 U11614 ( .A1(n7733), .A2(n7732), .ZN(n7734) );
  INV_X1 U11615 ( .A(n9249), .ZN(n8971) );
  NOR2_X1 U11619 ( .A1(n7736), .A2(n19516), .ZN(n7737) );
  NAND2_X1 U11620 ( .A1(n7740), .A2(n7739), .ZN(n7744) );
  NAND2_X1 U11621 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  NOR2_X1 U11622 ( .A1(n7747), .A2(n7912), .ZN(n8124) );
  INV_X1 U11623 ( .A(n8125), .ZN(n7751) );
  OAI21_X1 U11624 ( .B1(n7002), .B2(n7908), .A(n7903), .ZN(n7757) );
  NAND3_X1 U11625 ( .A1(n7754), .A2(n7753), .A3(n19521), .ZN(n7756) );
  NAND2_X1 U11626 ( .A1(n7752), .A2(n8657), .ZN(n7759) );
  NAND2_X1 U11627 ( .A1(n8658), .A2(n7759), .ZN(n9003) );
  NOR2_X1 U11628 ( .A1(n7761), .A2(n2540), .ZN(n7762) );
  NAND2_X1 U11629 ( .A1(n7931), .A2(n20359), .ZN(n7765) );
  NAND2_X1 U11630 ( .A1(n8998), .A2(n8657), .ZN(n7776) );
  NAND2_X1 U11631 ( .A1(n8999), .A2(n8998), .ZN(n8443) );
  NAND2_X1 U11632 ( .A1(n7919), .A2(n7921), .ZN(n7980) );
  INV_X1 U11634 ( .A(n8998), .ZN(n8773) );
  NOR2_X1 U11635 ( .A1(n7958), .A2(n7834), .ZN(n7770) );
  NAND3_X1 U11636 ( .A1(n7836), .A2(n20165), .A3(n8906), .ZN(n7771) );
  OAI21_X1 U11637 ( .B1(n8443), .B2(n19517), .A(n7774), .ZN(n7775) );
  XNOR2_X1 U11638 ( .A(n9792), .B(n9667), .ZN(n10603) );
  NAND2_X1 U11639 ( .A1(n19520), .A2(n8315), .ZN(n7779) );
  INV_X1 U11640 ( .A(n8313), .ZN(n8314) );
  NAND3_X1 U11641 ( .A1(n8312), .A2(n8314), .A3(n19942), .ZN(n7777) );
  NAND2_X1 U11642 ( .A1(n7807), .A2(n8288), .ZN(n7780) );
  INV_X1 U11643 ( .A(n7780), .ZN(n7784) );
  OAI21_X1 U11644 ( .B1(n934), .B2(n8289), .A(n8292), .ZN(n7783) );
  NAND2_X1 U11645 ( .A1(n8293), .A2(n20189), .ZN(n7781) );
  MUX2_X1 U11646 ( .A(n7781), .B(n7780), .S(n8026), .Z(n7782) );
  AND2_X1 U11648 ( .A1(n7585), .A2(n8001), .ZN(n8324) );
  NAND2_X1 U11649 ( .A1(n7787), .A2(n8299), .ZN(n8043) );
  NAND3_X1 U11650 ( .A1(n8043), .A2(n8295), .A3(n7788), .ZN(n7792) );
  NAND2_X1 U11651 ( .A1(n8297), .A2(n20257), .ZN(n7791) );
  AND3_X1 U11652 ( .A1(n8297), .A2(n7789), .A3(n20485), .ZN(n7790) );
  NAND2_X1 U11653 ( .A1(n8034), .A2(n8282), .ZN(n8287) );
  NAND2_X1 U11654 ( .A1(n7793), .A2(n8287), .ZN(n7794) );
  OAI21_X1 U11655 ( .B1(n7796), .B2(n7795), .A(n7794), .ZN(n8761) );
  OAI21_X1 U11656 ( .B1(n19827), .B2(n9176), .A(n8760), .ZN(n7805) );
  NAND2_X1 U11657 ( .A1(n3212), .A2(n20490), .ZN(n7800) );
  NAND2_X1 U11658 ( .A1(n20347), .A2(n7801), .ZN(n7799) );
  AOI21_X1 U11659 ( .B1(n8016), .B2(n7801), .A(n20270), .ZN(n7802) );
  OR2_X1 U11660 ( .A1(n7802), .A2(n3212), .ZN(n7803) );
  NAND2_X1 U11661 ( .A1(n8293), .A2(n8026), .ZN(n7808) );
  NAND2_X1 U11662 ( .A1(n8293), .A2(n8290), .ZN(n7810) );
  NAND3_X1 U11664 ( .A1(n7950), .A2(n20013), .A3(n7815), .ZN(n7817) );
  MUX2_X1 U11665 ( .A(n9006), .B(n8890), .S(n8895), .Z(n7842) );
  NAND2_X1 U11666 ( .A1(n7972), .A2(n7820), .ZN(n7825) );
  NAND2_X1 U11667 ( .A1(n7974), .A2(n7967), .ZN(n7821) );
  OAI211_X1 U11668 ( .C1(n7967), .C2(n7968), .A(n7821), .B(n278), .ZN(n7823)
         );
  OAI21_X1 U11669 ( .B1(n7922), .B2(n7968), .A(n7971), .ZN(n7822) );
  NAND2_X1 U11670 ( .A1(n7823), .A2(n7822), .ZN(n7824) );
  OAI21_X1 U11671 ( .B1(n7973), .B2(n7825), .A(n7824), .ZN(n9008) );
  NAND3_X1 U11672 ( .A1(n7828), .A2(n7827), .A3(n20154), .ZN(n7832) );
  MUX2_X1 U11673 ( .A(n9008), .B(n8895), .S(n9007), .Z(n7841) );
  NOR2_X1 U11674 ( .A1(n7836), .A2(n7833), .ZN(n7957) );
  INV_X1 U11675 ( .A(n7957), .ZN(n7840) );
  NAND2_X1 U11676 ( .A1(n7837), .A2(n90), .ZN(n7838) );
  INV_X1 U11677 ( .A(n9009), .ZN(n8623) );
  XNOR2_X1 U11678 ( .A(n9420), .B(n10262), .ZN(n8407) );
  XNOR2_X1 U11679 ( .A(n10603), .B(n8407), .ZN(n7947) );
  INV_X1 U11680 ( .A(n7843), .ZN(n7846) );
  NAND2_X1 U11681 ( .A1(n8248), .A2(n8245), .ZN(n7845) );
  INV_X1 U11682 ( .A(n9271), .ZN(n8984) );
  INV_X1 U11683 ( .A(n8221), .ZN(n8216) );
  NAND2_X1 U11684 ( .A1(n7847), .A2(n8216), .ZN(n7850) );
  INV_X1 U11685 ( .A(n8219), .ZN(n8218) );
  AOI21_X1 U11686 ( .B1(n8215), .B2(n8218), .A(n8220), .ZN(n7848) );
  NOR2_X1 U11688 ( .A1(n8984), .A2(n9265), .ZN(n7870) );
  NAND2_X1 U11689 ( .A1(n8162), .A2(n7851), .ZN(n7854) );
  NAND2_X1 U11690 ( .A1(n7856), .A2(n7855), .ZN(n7853) );
  OAI21_X1 U11691 ( .B1(n7857), .B2(n7856), .A(n8160), .ZN(n7858) );
  MUX2_X1 U11692 ( .A(n20108), .B(n6539), .S(n8086), .Z(n7861) );
  INV_X1 U11695 ( .A(n7866), .ZN(n9267) );
  NAND2_X1 U11696 ( .A1(n8981), .A2(n9267), .ZN(n7869) );
  NAND2_X1 U11697 ( .A1(n8238), .A2(n8111), .ZN(n7863) );
  NOR2_X1 U11698 ( .A1(n8979), .A2(n9265), .ZN(n8652) );
  OAI22_X1 U11699 ( .A1(n8262), .A2(n7864), .B1(n8150), .B2(n8261), .ZN(n8154)
         );
  NOR2_X1 U11700 ( .A1(n8264), .A2(n895), .ZN(n7865) );
  INV_X1 U11701 ( .A(n8153), .ZN(n8107) );
  NAND2_X1 U11702 ( .A1(n8107), .A2(n7864), .ZN(n8266) );
  AOI22_X1 U11703 ( .A1(n8154), .A2(n8106), .B1(n7865), .B2(n8266), .ZN(n8653)
         );
  INV_X1 U11704 ( .A(n8653), .ZN(n9262) );
  AOI22_X1 U11705 ( .A1(n19880), .A2(n8652), .B1(n7867), .B2(n7866), .ZN(n7868) );
  INV_X1 U11706 ( .A(n8200), .ZN(n8071) );
  MUX2_X1 U11707 ( .A(n7873), .B(n7872), .S(n8070), .Z(n7875) );
  NOR2_X1 U11709 ( .A1(n8195), .A2(n20198), .ZN(n7880) );
  AOI22_X1 U11710 ( .A1(n7880), .A2(n7879), .B1(n7878), .B2(n8053), .ZN(n7884)
         );
  AOI21_X1 U11711 ( .B1(n8052), .B2(n8193), .A(n8053), .ZN(n7882) );
  NAND2_X1 U11712 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  NAND2_X1 U11713 ( .A1(n1850), .A2(n923), .ZN(n7886) );
  OAI21_X1 U11714 ( .B1(n8179), .B2(n8176), .A(n7622), .ZN(n7885) );
  MUX2_X1 U11715 ( .A(n7886), .B(n7885), .S(n8181), .Z(n7888) );
  NAND2_X1 U11716 ( .A1(n9275), .A2(n20265), .ZN(n7889) );
  NAND3_X1 U11717 ( .A1(n7897), .A2(n9274), .A3(n7889), .ZN(n7901) );
  NAND2_X1 U11718 ( .A1(n8186), .A2(n7893), .ZN(n7890) );
  INV_X1 U11719 ( .A(n7892), .ZN(n7894) );
  NAND2_X1 U11720 ( .A1(n7894), .A2(n7460), .ZN(n7895) );
  INV_X1 U11721 ( .A(n9274), .ZN(n9277) );
  NAND3_X1 U11722 ( .A1(n19732), .A2(n9277), .A3(n20265), .ZN(n7899) );
  XNOR2_X1 U11723 ( .A(n10528), .B(n10264), .ZN(n9974) );
  INV_X1 U11725 ( .A(n7904), .ZN(n7905) );
  INV_X1 U11726 ( .A(n9149), .ZN(n9144) );
  NAND2_X1 U11727 ( .A1(n7961), .A2(n8906), .ZN(n7916) );
  NAND2_X1 U11729 ( .A1(n9144), .A2(n8337), .ZN(n7944) );
  OAI21_X1 U11730 ( .B1(n7972), .B2(n7973), .A(n7974), .ZN(n7925) );
  NAND2_X1 U11731 ( .A1(n7967), .A2(n278), .ZN(n7924) );
  NAND3_X1 U11732 ( .A1(n7925), .A2(n7924), .A3(n7923), .ZN(n7926) );
  OAI21_X1 U11733 ( .B1(n7927), .B2(n7967), .A(n7926), .ZN(n8790) );
  NAND3_X1 U11734 ( .A1(n7932), .A2(n1452), .A3(n7931), .ZN(n7940) );
  NAND3_X1 U11735 ( .A1(n2031), .A2(n1063), .A3(n7933), .ZN(n7939) );
  NAND3_X1 U11736 ( .A1(n2031), .A2(n7936), .A3(n20195), .ZN(n7938) );
  AOI21_X2 U11738 ( .B1(n7944), .B2(n7943), .A(n7942), .ZN(n9937) );
  XNOR2_X1 U11739 ( .A(n9937), .B(n2341), .ZN(n7945) );
  XNOR2_X1 U11740 ( .A(n9974), .B(n7945), .ZN(n7946) );
  INV_X1 U11741 ( .A(n11161), .ZN(n10650) );
  MUX2_X1 U11742 ( .A(n9555), .B(n10945), .S(n10650), .Z(n8402) );
  MUX2_X1 U11743 ( .A(n7952), .B(n7951), .S(n7950), .Z(n7954) );
  NAND2_X1 U11744 ( .A1(n7957), .A2(n8910), .ZN(n7960) );
  OAI211_X1 U11745 ( .C1(n7962), .C2(n7961), .A(n7960), .B(n7959), .ZN(n9171)
         );
  INV_X1 U11746 ( .A(n9171), .ZN(n9080) );
  OAI21_X1 U11747 ( .B1(n7965), .B2(n8017), .A(n20270), .ZN(n7964) );
  AOI22_X1 U11748 ( .A1(n7966), .A2(n7965), .B1(n8016), .B2(n7964), .ZN(n8568)
         );
  NAND2_X1 U11749 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  NAND2_X1 U11750 ( .A1(n7973), .A2(n7972), .ZN(n7975) );
  NOR2_X1 U11751 ( .A1(n269), .A2(n8569), .ZN(n7988) );
  AOI21_X1 U11752 ( .B1(n7980), .B2(n7979), .A(n7978), .ZN(n7987) );
  NAND2_X1 U11753 ( .A1(n7982), .A2(n7981), .ZN(n7985) );
  AOI21_X1 U11754 ( .B1(n7985), .B2(n7984), .A(n7919), .ZN(n7986) );
  OAI22_X1 U11756 ( .A1(n8014), .A2(n20154), .B1(n8011), .B2(n7990), .ZN(n8010) );
  OAI21_X1 U11757 ( .B1(n7995), .B2(n7994), .A(n7993), .ZN(n9168) );
  NOR2_X2 U11758 ( .A1(n7997), .A2(n7996), .ZN(n10150) );
  NOR2_X1 U11759 ( .A1(n7998), .A2(n8322), .ZN(n8000) );
  NOR2_X1 U11761 ( .A1(n1425), .A2(n8001), .ZN(n8002) );
  NAND2_X1 U11762 ( .A1(n19520), .A2(n8004), .ZN(n8006) );
  AND2_X1 U11763 ( .A1(n8006), .A2(n8007), .ZN(n8008) );
  MUX2_X1 U11765 ( .A(n3212), .B(n8017), .S(n8016), .Z(n8023) );
  MUX2_X1 U11766 ( .A(n8020), .B(n8019), .S(n3212), .Z(n8021) );
  OAI21_X1 U11767 ( .B1(n8023), .B2(n20270), .A(n8021), .ZN(n9062) );
  INV_X1 U11768 ( .A(n8677), .ZN(n8037) );
  NAND3_X1 U11769 ( .A1(n8290), .A2(n8024), .A3(n7468), .ZN(n8030) );
  OAI21_X1 U11770 ( .B1(n8026), .B2(n8289), .A(n20189), .ZN(n8027) );
  INV_X1 U11771 ( .A(n8027), .ZN(n8028) );
  NAND2_X1 U11772 ( .A1(n8034), .A2(n8280), .ZN(n8035) );
  OAI21_X1 U11773 ( .B1(n8034), .B2(n8282), .A(n8281), .ZN(n8032) );
  NOR3_X1 U11774 ( .A1(n9029), .A2(n9060), .A3(n8833), .ZN(n8036) );
  AOI21_X1 U11775 ( .B1(n8037), .B2(n8831), .A(n8036), .ZN(n8039) );
  NAND3_X1 U11776 ( .A1(n9031), .A2(n8829), .A3(n9060), .ZN(n8038) );
  XNOR2_X1 U11777 ( .A(n10270), .B(n10150), .ZN(n8524) );
  OAI21_X1 U11778 ( .B1(n8297), .B2(n8298), .A(n8040), .ZN(n8042) );
  AND2_X1 U11779 ( .A1(n8040), .A2(n20485), .ZN(n8296) );
  INV_X1 U11780 ( .A(n8303), .ZN(n8309) );
  NAND3_X1 U11781 ( .A1(n20001), .A2(n8045), .A3(n8044), .ZN(n8049) );
  OAI211_X1 U11782 ( .C1(n20057), .C2(n20001), .A(n8047), .B(n8304), .ZN(n8048) );
  NAND2_X1 U11783 ( .A1(n9836), .A2(n9066), .ZN(n9069) );
  NAND2_X1 U11784 ( .A1(n8054), .A2(n8197), .ZN(n8056) );
  NAND2_X1 U11785 ( .A1(n8056), .A2(n20198), .ZN(n8057) );
  NOR2_X1 U11786 ( .A1(n20247), .A2(n8060), .ZN(n8064) );
  NOR2_X1 U11787 ( .A1(n8185), .A2(n20465), .ZN(n8063) );
  INV_X1 U11789 ( .A(n8066), .ZN(n8177) );
  NOR2_X1 U11791 ( .A1(n7421), .A2(n8070), .ZN(n8073) );
  NOR2_X1 U11793 ( .A1(n3795), .A2(n8219), .ZN(n8078) );
  NOR2_X1 U11794 ( .A1(n8079), .A2(n8215), .ZN(n8080) );
  NOR3_X1 U11795 ( .A1(n19809), .A2(n20441), .A3(n3795), .ZN(n8081) );
  MUX2_X1 U11796 ( .A(n8086), .B(n8085), .S(n20107), .Z(n8088) );
  AND2_X1 U11797 ( .A1(n8093), .A2(n8090), .ZN(n8210) );
  AOI21_X1 U11798 ( .B1(n8094), .B2(n8093), .A(n20511), .ZN(n8096) );
  OR2_X1 U11799 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  NAND2_X1 U11800 ( .A1(n9333), .A2(n9328), .ZN(n8869) );
  MUX2_X1 U11801 ( .A(n8100), .B(n8099), .S(n8098), .Z(n8102) );
  NAND2_X1 U11802 ( .A1(n8241), .A2(n8100), .ZN(n8244) );
  INV_X1 U11803 ( .A(n8244), .ZN(n8101) );
  MUX2_X1 U11804 ( .A(n8102), .B(n8101), .S(n3775), .Z(n8463) );
  INV_X1 U11805 ( .A(n8463), .ZN(n8119) );
  AND2_X1 U11807 ( .A1(n8104), .A2(n8261), .ZN(n8110) );
  NAND2_X1 U11808 ( .A1(n8151), .A2(n895), .ZN(n8105) );
  NAND2_X1 U11809 ( .A1(n8106), .A2(n8105), .ZN(n8108) );
  NAND2_X1 U11810 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  INV_X1 U11811 ( .A(n9330), .ZN(n9074) );
  AND3_X1 U11812 ( .A1(n8112), .A2(n8239), .A3(n8111), .ZN(n8462) );
  INV_X1 U11813 ( .A(n8462), .ZN(n8118) );
  NAND4_X1 U11814 ( .A1(n8119), .A2(n20008), .A3(n9074), .A4(n8118), .ZN(n8123) );
  NAND2_X1 U11815 ( .A1(n8245), .A2(n8246), .ZN(n8117) );
  OAI21_X1 U11816 ( .B1(n8114), .B2(n8113), .A(n8248), .ZN(n8116) );
  MUX2_X1 U11817 ( .A(n8117), .B(n8116), .S(n20251), .Z(n8120) );
  NAND4_X1 U11818 ( .A1(n8119), .A2(n900), .A3(n8120), .A4(n8118), .ZN(n8121)
         );
  XNOR2_X1 U11819 ( .A(n10552), .B(n10271), .ZN(n9998) );
  XNOR2_X1 U11820 ( .A(n9998), .B(n8524), .ZN(n8173) );
  OR2_X1 U11821 ( .A1(n7752), .A2(n8657), .ZN(n8660) );
  XNOR2_X1 U11822 ( .A(n9635), .B(n17587), .ZN(n8171) );
  INV_X1 U11823 ( .A(n8470), .ZN(n9091) );
  NAND2_X1 U11824 ( .A1(n8884), .A2(n9453), .ZN(n8889) );
  NAND2_X1 U11825 ( .A1(n8387), .A2(n8132), .ZN(n8137) );
  NAND2_X1 U11826 ( .A1(n8133), .A2(n8381), .ZN(n8134) );
  MUX2_X1 U11827 ( .A(n20200), .B(n8272), .S(n8348), .Z(n8139) );
  OAI21_X1 U11828 ( .B1(n8370), .B2(n8377), .A(n8142), .ZN(n8144) );
  NAND2_X1 U11829 ( .A1(n20294), .A2(n20252), .ZN(n8143) );
  NAND2_X1 U11830 ( .A1(n8144), .A2(n8143), .ZN(n8148) );
  INV_X1 U11831 ( .A(n8261), .ZN(n8149) );
  OAI21_X1 U11832 ( .B1(n7571), .B2(n8150), .A(n8149), .ZN(n8152) );
  INV_X1 U11833 ( .A(n8156), .ZN(n9341) );
  NAND2_X1 U11834 ( .A1(n9341), .A2(n9346), .ZN(n8701) );
  NOR2_X1 U11835 ( .A1(n8157), .A2(n6830), .ZN(n8158) );
  NOR2_X1 U11836 ( .A1(n8159), .A2(n8158), .ZN(n8161) );
  NOR2_X1 U11837 ( .A1(n9341), .A2(n9563), .ZN(n9191) );
  NAND2_X1 U11838 ( .A1(n9191), .A2(n9564), .ZN(n8168) );
  XNOR2_X1 U11839 ( .A(n9999), .B(n918), .ZN(n10584) );
  XNOR2_X1 U11840 ( .A(n10584), .B(n8171), .ZN(n8172) );
  INV_X1 U11841 ( .A(n10945), .ZN(n8174) );
  NAND2_X1 U11842 ( .A1(n8174), .A2(n11158), .ZN(n8399) );
  NOR2_X1 U11843 ( .A1(n8178), .A2(n8177), .ZN(n8180) );
  AND2_X1 U11844 ( .A1(n8182), .A2(n8184), .ZN(n8191) );
  INV_X1 U11845 ( .A(n8183), .ZN(n8188) );
  OAI21_X1 U11846 ( .B1(n8188), .B2(n8187), .A(n8186), .ZN(n8189) );
  NAND2_X1 U11847 ( .A1(n9218), .A2(n908), .ZN(n8228) );
  OAI21_X1 U11848 ( .B1(n8196), .B2(n8195), .A(n8194), .ZN(n8198) );
  NAND2_X1 U11849 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  INV_X1 U11850 ( .A(n9221), .ZN(n8795) );
  NAND3_X1 U11851 ( .A1(n8205), .A2(n819), .A3(n8203), .ZN(n8206) );
  NAND2_X1 U11852 ( .A1(n8210), .A2(n8209), .ZN(n8214) );
  OAI211_X1 U11853 ( .C1(n7631), .C2(n8212), .A(n7633), .B(n8211), .ZN(n8213)
         );
  NOR2_X1 U11854 ( .A1(n9114), .A2(n9113), .ZN(n8225) );
  NAND2_X1 U11855 ( .A1(n8218), .A2(n20180), .ZN(n8222) );
  OAI22_X1 U11856 ( .A1(n8222), .A2(n19809), .B1(n8219), .B2(n20174), .ZN(
        n8223) );
  AND2_X1 U11857 ( .A1(n8797), .A2(n9113), .ZN(n8428) );
  AOI22_X1 U11858 ( .A1(n8226), .A2(n8225), .B1(n8428), .B2(n8795), .ZN(n8227)
         );
  NAND2_X1 U11859 ( .A1(n8228), .A2(n8227), .ZN(n9769) );
  MUX2_X1 U11860 ( .A(n20107), .B(n8230), .S(n20495), .Z(n8235) );
  AND2_X1 U11861 ( .A1(n6539), .A2(n8232), .ZN(n8234) );
  OAI21_X1 U11862 ( .B1(n8239), .B2(n8098), .A(n8237), .ZN(n8240) );
  NAND2_X1 U11863 ( .A1(n8240), .A2(n3775), .ZN(n8243) );
  NOR3_X1 U11864 ( .A1(n8435), .A2(n8434), .A3(n9201), .ZN(n8279) );
  NAND2_X1 U11865 ( .A1(n8247), .A2(n8246), .ZN(n8249) );
  OR2_X1 U11866 ( .A1(n8256), .A2(n7724), .ZN(n8257) );
  NOR2_X1 U11868 ( .A1(n8349), .A2(n19914), .ZN(n8269) );
  OAI21_X1 U11869 ( .B1(n8270), .B2(n8269), .A(n8268), .ZN(n8275) );
  NAND2_X1 U11870 ( .A1(n8273), .A2(n20200), .ZN(n8274) );
  NAND2_X1 U11871 ( .A1(n9129), .A2(n8276), .ZN(n8432) );
  OR2_X1 U11872 ( .A1(n8432), .A2(n9201), .ZN(n8277) );
  XNOR2_X1 U11874 ( .A(n9769), .B(n10431), .ZN(n9996) );
  NOR2_X1 U11875 ( .A1(n20012), .A2(n8282), .ZN(n8285) );
  NOR2_X1 U11876 ( .A1(n8287), .A2(n8286), .ZN(n8421) );
  OAI21_X1 U11877 ( .B1(n8290), .B2(n8289), .A(n934), .ZN(n8291) );
  OAI211_X1 U11878 ( .C1(n8300), .C2(n8299), .A(n8298), .B(n8297), .ZN(n9099)
         );
  OAI21_X1 U11879 ( .B1(n8303), .B2(n20001), .A(n8301), .ZN(n8308) );
  NAND2_X1 U11880 ( .A1(n20057), .A2(n8304), .ZN(n8307) );
  NAND2_X1 U11882 ( .A1(n7592), .A2(n8314), .ZN(n8318) );
  NAND2_X1 U11883 ( .A1(n19942), .A2(n8315), .ZN(n8317) );
  MUX2_X1 U11884 ( .A(n8318), .B(n8317), .S(n8316), .Z(n8319) );
  NAND2_X1 U11885 ( .A1(n8872), .A2(n9106), .ZN(n8559) );
  NAND3_X1 U11886 ( .A1(n8559), .A2(n9107), .A3(n20000), .ZN(n8326) );
  INV_X1 U11888 ( .A(n9120), .ZN(n8331) );
  INV_X1 U11889 ( .A(n9122), .ZN(n8814) );
  NAND2_X1 U11890 ( .A1(n8815), .A2(n9122), .ZN(n8328) );
  XNOR2_X1 U11891 ( .A(n9861), .B(n19990), .ZN(n8469) );
  XNOR2_X1 U11892 ( .A(n8469), .B(n9996), .ZN(n8398) );
  AND2_X1 U11893 ( .A1(n8332), .A2(n8734), .ZN(n8335) );
  INV_X1 U11894 ( .A(n9648), .ZN(n8339) );
  INV_X1 U11895 ( .A(n9143), .ZN(n8338) );
  MUX2_X1 U11896 ( .A(n8341), .B(n3121), .S(n8340), .Z(n8346) );
  MUX2_X1 U11897 ( .A(n20274), .B(n8343), .S(n8342), .Z(n8345) );
  AOI21_X1 U11898 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(n8353) );
  NAND2_X1 U11899 ( .A1(n8355), .A2(n8354), .ZN(n8356) );
  NAND2_X1 U11900 ( .A1(n8364), .A2(n8363), .ZN(n8368) );
  NAND2_X1 U11901 ( .A1(n1994), .A2(n8365), .ZN(n8367) );
  NAND3_X1 U11902 ( .A1(n20294), .A2(n8373), .A3(n8372), .ZN(n8379) );
  NAND3_X1 U11903 ( .A1(n8377), .A2(n20252), .A3(n8375), .ZN(n8378) );
  INV_X1 U11904 ( .A(n8389), .ZN(n8392) );
  NAND2_X1 U11907 ( .A1(n8386), .A2(n8385), .ZN(n8388) );
  MUX2_X1 U11908 ( .A(n8389), .B(n8388), .S(n8387), .Z(n8390) );
  NAND3_X1 U11909 ( .A1(n9212), .A2(n9211), .A3(n8420), .ZN(n8393) );
  XNOR2_X1 U11910 ( .A(n10236), .B(n2448), .ZN(n8395) );
  XNOR2_X1 U11911 ( .A(n8396), .B(n8395), .ZN(n8397) );
  AOI21_X1 U11913 ( .B1(n8400), .B2(n8399), .A(n11159), .ZN(n8401) );
  MUX2_X1 U11914 ( .A(n8569), .B(n9171), .S(n9167), .Z(n8404) );
  MUX2_X1 U11915 ( .A(n9163), .B(n9160), .S(n8611), .Z(n8406) );
  MUX2_X1 U11916 ( .A(n9159), .B(n9162), .S(n9158), .Z(n8405) );
  XNOR2_X1 U11917 ( .A(n9794), .B(n10472), .ZN(n8408) );
  XNOR2_X1 U11918 ( .A(n8408), .B(n8407), .ZN(n8418) );
  MUX2_X1 U11919 ( .A(n8713), .B(n9241), .S(n9240), .Z(n8410) );
  MUX2_X1 U11920 ( .A(n9240), .B(n9242), .S(n6587), .Z(n8409) );
  MUX2_X1 U11921 ( .A(n8410), .B(n8409), .S(n266), .Z(n10526) );
  XNOR2_X1 U11925 ( .A(n10425), .B(n10526), .ZN(n9459) );
  NAND2_X1 U11926 ( .A1(n9564), .A2(n9338), .ZN(n8413) );
  MUX2_X1 U11927 ( .A(n8699), .B(n8413), .S(n9567), .Z(n8414) );
  OAI21_X2 U11928 ( .B1(n8415), .B2(n9338), .A(n8414), .ZN(n10265) );
  XNOR2_X1 U11929 ( .A(n10265), .B(n2257), .ZN(n8416) );
  XNOR2_X1 U11930 ( .A(n9459), .B(n8416), .ZN(n8417) );
  XNOR2_X1 U11931 ( .A(n8418), .B(n8417), .ZN(n10756) );
  NOR2_X1 U11932 ( .A1(n9111), .A2(n9106), .ZN(n8424) );
  OAI21_X1 U11933 ( .B1(n8555), .B2(n9105), .A(n9111), .ZN(n8425) );
  XNOR2_X1 U11934 ( .A(n10620), .B(n18075), .ZN(n8426) );
  XNOR2_X1 U11935 ( .A(n8427), .B(n8426), .ZN(n8441) );
  NOR2_X1 U11936 ( .A1(n9219), .A2(n9112), .ZN(n8431) );
  NAND2_X1 U11937 ( .A1(n8428), .A2(n9217), .ZN(n8430) );
  AND2_X1 U11938 ( .A1(n8433), .A2(n8432), .ZN(n8437) );
  AOI21_X1 U11939 ( .B1(n9130), .B2(n8276), .A(n8805), .ZN(n8436) );
  OAI22_X1 U11940 ( .A1(n8437), .A2(n9780), .B1(n9204), .B2(n8436), .ZN(n9535)
         );
  XNOR2_X1 U11941 ( .A(n10072), .B(n9535), .ZN(n10543) );
  NAND2_X1 U11942 ( .A1(n9151), .A2(n9143), .ZN(n8438) );
  NAND2_X1 U11943 ( .A1(n9151), .A2(n8790), .ZN(n8789) );
  XNOR2_X1 U11944 ( .A(n10028), .B(n8769), .ZN(n10480) );
  XNOR2_X1 U11945 ( .A(n10480), .B(n10543), .ZN(n8440) );
  OAI21_X1 U11946 ( .B1(n8995), .B2(n8443), .A(n8442), .ZN(n9923) );
  NOR2_X1 U11947 ( .A1(n9209), .A2(n8445), .ZN(n8446) );
  XNOR2_X1 U11948 ( .A(n10303), .B(n9923), .ZN(n9738) );
  OAI21_X1 U11949 ( .B1(n9275), .B2(n9274), .A(n8650), .ZN(n8449) );
  XNOR2_X1 U11950 ( .A(n8450), .B(n10114), .ZN(n8451) );
  XNOR2_X1 U11951 ( .A(n9738), .B(n8451), .ZN(n8461) );
  OAI21_X1 U11952 ( .B1(n8979), .B2(n2118), .A(n9267), .ZN(n8453) );
  NOR2_X1 U11953 ( .A1(n8979), .A2(n19710), .ZN(n8452) );
  INV_X1 U11954 ( .A(n8550), .ZN(n9128) );
  NAND3_X1 U11956 ( .A1(n9119), .A2(n8552), .A3(n8810), .ZN(n8455) );
  OAI211_X2 U11957 ( .C1(n9128), .C2(n8457), .A(n8456), .B(n8455), .ZN(n10572)
         );
  XNOR2_X1 U11958 ( .A(n10570), .B(n10572), .ZN(n8459) );
  XNOR2_X1 U11959 ( .A(n10054), .B(n2067), .ZN(n8458) );
  XNOR2_X1 U11960 ( .A(n8459), .B(n8458), .ZN(n8460) );
  XNOR2_X1 U11961 ( .A(n8461), .B(n8460), .ZN(n11526) );
  INV_X1 U11962 ( .A(n9331), .ZN(n9073) );
  NOR2_X1 U11963 ( .A1(n9836), .A2(n9066), .ZN(n8545) );
  INV_X1 U11964 ( .A(n9834), .ZN(n9317) );
  XNOR2_X1 U11965 ( .A(n9647), .B(n10557), .ZN(n9470) );
  XNOR2_X1 U11966 ( .A(n9470), .B(n8469), .ZN(n8481) );
  NAND2_X1 U11967 ( .A1(n9451), .A2(n9453), .ZN(n8474) );
  NAND3_X1 U11968 ( .A1(n1576), .A2(n9090), .A3(n9091), .ZN(n8473) );
  NAND3_X1 U11969 ( .A1(n8474), .A2(n8473), .A3(n8472), .ZN(n9812) );
  OAI21_X1 U11971 ( .B1(n670), .B2(n8972), .A(n8971), .ZN(n8476) );
  NAND3_X1 U11972 ( .A1(n9249), .A2(n9256), .A3(n8879), .ZN(n8475) );
  XNOR2_X1 U11973 ( .A(n10281), .B(n9812), .ZN(n9722) );
  INV_X1 U11974 ( .A(n9007), .ZN(n9004) );
  NAND2_X1 U11975 ( .A1(n9004), .A2(n19490), .ZN(n8477) );
  INV_X1 U11976 ( .A(n8895), .ZN(n8891) );
  OAI211_X1 U11977 ( .C1(n19490), .C2(n9008), .A(n8891), .B(n9005), .ZN(n8478)
         );
  XNOR2_X1 U11978 ( .A(n10497), .B(n17999), .ZN(n8479) );
  XNOR2_X1 U11979 ( .A(n9722), .B(n8479), .ZN(n8480) );
  NOR2_X1 U11981 ( .A1(n10756), .A2(n11527), .ZN(n10635) );
  MUX2_X1 U11983 ( .A(n8485), .B(n8483), .S(n9368), .Z(n8487) );
  NOR2_X1 U11984 ( .A1(n8603), .A2(n8742), .ZN(n8484) );
  MUX2_X1 U11985 ( .A(n8945), .B(n8941), .S(n8729), .Z(n8489) );
  NOR2_X1 U11986 ( .A1(n8944), .A2(n8939), .ZN(n8490) );
  XNOR2_X1 U11988 ( .A(n10442), .B(n10402), .ZN(n9445) );
  INV_X1 U11989 ( .A(n8492), .ZN(n8496) );
  OAI21_X1 U11990 ( .B1(n8904), .B2(n8720), .A(n9358), .ZN(n8495) );
  NAND2_X1 U11991 ( .A1(n8722), .A2(n9528), .ZN(n8493) );
  MUX2_X1 U11992 ( .A(n8493), .B(n8492), .S(n9359), .Z(n8494) );
  XNOR2_X1 U11994 ( .A(n10506), .B(n9817), .ZN(n8507) );
  NAND2_X1 U11995 ( .A1(n9361), .A2(n207), .ZN(n8505) );
  NAND2_X1 U11996 ( .A1(n9363), .A2(n9362), .ZN(n8501) );
  MUX2_X1 U11997 ( .A(n8502), .B(n8501), .S(n8961), .Z(n8504) );
  NAND3_X1 U11998 ( .A1(n8958), .A2(n8726), .A3(n207), .ZN(n8503) );
  XNOR2_X1 U11999 ( .A(n19785), .B(n2356), .ZN(n8506) );
  XNOR2_X1 U12000 ( .A(n8507), .B(n8506), .ZN(n8508) );
  INV_X1 U12001 ( .A(n11527), .ZN(n10919) );
  INV_X1 U12002 ( .A(n11521), .ZN(n11530) );
  NOR2_X1 U12003 ( .A1(n8676), .A2(n9023), .ZN(n9022) );
  INV_X1 U12006 ( .A(n8512), .ZN(n8517) );
  NAND3_X1 U12007 ( .A1(n8517), .A2(n8516), .A3(n8515), .ZN(n8518) );
  NOR2_X1 U12008 ( .A1(n8846), .A2(n9300), .ZN(n8523) );
  NOR2_X1 U12009 ( .A1(n9018), .A2(n9295), .ZN(n8842) );
  AOI22_X1 U12010 ( .A1(n9304), .A2(n8842), .B1(n8520), .B2(n8846), .ZN(n8521)
         );
  XNOR2_X1 U12011 ( .A(n10551), .B(n10461), .ZN(n9476) );
  XNOR2_X1 U12012 ( .A(n9476), .B(n8524), .ZN(n8536) );
  NOR2_X1 U12013 ( .A1(n8527), .A2(n9039), .ZN(n8526) );
  NOR2_X1 U12014 ( .A1(n9046), .A2(n8851), .ZN(n8525) );
  NAND3_X1 U12015 ( .A1(n8527), .A2(n9046), .A3(n8848), .ZN(n8528) );
  OAI21_X1 U12016 ( .B1(n9037), .B2(n8529), .A(n8528), .ZN(n8530) );
  NOR2_X2 U12017 ( .A1(n8531), .A2(n8530), .ZN(n10491) );
  NOR2_X1 U12018 ( .A1(n9291), .A2(n9576), .ZN(n8532) );
  XNOR2_X1 U12019 ( .A(n9824), .B(n10491), .ZN(n8534) );
  NAND2_X1 U12020 ( .A1(n8823), .A2(n9307), .ZN(n9054) );
  XNOR2_X1 U12021 ( .A(n10274), .B(n2218), .ZN(n8533) );
  XNOR2_X1 U12022 ( .A(n8534), .B(n8533), .ZN(n8535) );
  NOR2_X1 U12024 ( .A1(n9331), .A2(n9326), .ZN(n8538) );
  AOI22_X1 U12025 ( .A1(n8539), .A2(n9333), .B1(n8538), .B2(n9329), .ZN(n8540)
         );
  NOR2_X1 U12027 ( .A1(n8543), .A2(n8542), .ZN(n8547) );
  XNOR2_X1 U12028 ( .A(n872), .B(n10604), .ZN(n9503) );
  INV_X1 U12030 ( .A(n9420), .ZN(n10173) );
  XNOR2_X1 U12031 ( .A(n10173), .B(n2442), .ZN(n8548) );
  NOR2_X1 U12033 ( .A1(n8550), .A2(n8813), .ZN(n8551) );
  AOI21_X1 U12034 ( .B1(n8552), .B2(n8818), .A(n8551), .ZN(n8554) );
  INV_X1 U12035 ( .A(n9107), .ZN(n8871) );
  OAI21_X1 U12036 ( .B1(n8871), .B2(n9111), .A(n9106), .ZN(n8558) );
  INV_X1 U12037 ( .A(n8555), .ZN(n8557) );
  INV_X1 U12038 ( .A(n8780), .ZN(n8556) );
  INV_X1 U12039 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U12040 ( .A1(n9111), .A2(n8560), .ZN(n8561) );
  XNOR2_X1 U12041 ( .A(n10171), .B(n10421), .ZN(n9208) );
  INV_X1 U12042 ( .A(n9087), .ZN(n8562) );
  OAI211_X1 U12043 ( .C1(n9451), .C2(n8884), .A(n8563), .B(n1576), .ZN(n8564)
         );
  OAI21_X1 U12044 ( .B1(n1576), .B2(n9454), .A(n8564), .ZN(n9500) );
  XNOR2_X1 U12045 ( .A(n9500), .B(n19767), .ZN(n9750) );
  XNOR2_X1 U12046 ( .A(n9208), .B(n9750), .ZN(n8566) );
  NOR3_X1 U12048 ( .A1(n9167), .A2(n9080), .A3(n9166), .ZN(n8570) );
  INV_X1 U12049 ( .A(n8833), .ZN(n9059) );
  INV_X1 U12050 ( .A(n9029), .ZN(n8571) );
  MUX2_X1 U12051 ( .A(n8829), .B(n8571), .S(n9060), .Z(n8575) );
  MUX2_X1 U12053 ( .A(n8573), .B(n8572), .S(n8829), .Z(n8574) );
  XNOR2_X1 U12054 ( .A(n10254), .B(n10186), .ZN(n9325) );
  NAND2_X1 U12055 ( .A1(n9579), .A2(n19896), .ZN(n8581) );
  NAND3_X1 U12056 ( .A1(n8577), .A2(n19519), .A3(n19715), .ZN(n8580) );
  AND2_X1 U12057 ( .A1(n9291), .A2(n9576), .ZN(n9290) );
  NOR2_X1 U12058 ( .A1(n19896), .A2(n9576), .ZN(n8578) );
  OAI21_X1 U12059 ( .B1(n9290), .B2(n8578), .A(n9287), .ZN(n8579) );
  OAI211_X1 U12060 ( .C1(n9289), .C2(n8581), .A(n8580), .B(n8579), .ZN(n9844)
         );
  XNOR2_X1 U12061 ( .A(n9844), .B(n10252), .ZN(n9773) );
  XNOR2_X1 U12062 ( .A(n9325), .B(n9773), .ZN(n8591) );
  MUX2_X1 U12063 ( .A(n891), .B(n8846), .S(n2984), .Z(n8585) );
  NAND2_X1 U12064 ( .A1(n9304), .A2(n9296), .ZN(n8583) );
  INV_X1 U12065 ( .A(n8671), .ZN(n8588) );
  INV_X1 U12066 ( .A(n9023), .ZN(n8836) );
  INV_X1 U12067 ( .A(n9021), .ZN(n8837) );
  NAND2_X1 U12068 ( .A1(n8672), .A2(n8837), .ZN(n8586) );
  XNOR2_X1 U12069 ( .A(n10612), .B(n10367), .ZN(n9512) );
  XNOR2_X1 U12070 ( .A(n9842), .B(n2384), .ZN(n8589) );
  XNOR2_X1 U12071 ( .A(n9512), .B(n8589), .ZN(n8590) );
  XNOR2_X1 U12072 ( .A(n9754), .B(n8593), .ZN(n10182) );
  NAND2_X1 U12073 ( .A1(n8947), .A2(n8937), .ZN(n8728) );
  OAI21_X1 U12074 ( .B1(n8939), .B2(n8945), .A(n8728), .ZN(n8648) );
  AOI21_X2 U12075 ( .B1(n8644), .B2(n8648), .A(n8594), .ZN(n10320) );
  XNOR2_X1 U12076 ( .A(n10320), .B(n2375), .ZN(n8595) );
  XNOR2_X1 U12077 ( .A(n10182), .B(n8595), .ZN(n8608) );
  INV_X1 U12078 ( .A(n8928), .ZN(n8752) );
  INV_X1 U12079 ( .A(n8925), .ZN(n8639) );
  OAI22_X1 U12081 ( .A1(n8752), .A2(n8639), .B1(n8933), .B2(n8931), .ZN(n8643)
         );
  INV_X1 U12082 ( .A(n8749), .ZN(n8929) );
  NAND2_X1 U12083 ( .A1(n8932), .A2(n8925), .ZN(n8597) );
  NAND2_X1 U12085 ( .A1(n9037), .A2(n9045), .ZN(n8601) );
  NAND2_X1 U12086 ( .A1(n9039), .A2(n9038), .ZN(n8599) );
  AOI21_X1 U12087 ( .B1(n8599), .B2(n8851), .A(n8849), .ZN(n8600) );
  AOI21_X1 U12088 ( .B1(n8601), .B2(n8848), .A(n8600), .ZN(n9402) );
  XNOR2_X1 U12089 ( .A(n9402), .B(n10179), .ZN(n9232) );
  INV_X1 U12090 ( .A(n9232), .ZN(n8606) );
  NAND2_X1 U12091 ( .A1(n9372), .A2(n9367), .ZN(n8605) );
  OAI21_X1 U12092 ( .B1(n8953), .B2(n8742), .A(n8603), .ZN(n8604) );
  AOI22_X1 U12093 ( .A1(n8605), .A2(n8743), .B1(n8956), .B2(n8604), .ZN(n9537)
         );
  INV_X1 U12094 ( .A(n9537), .ZN(n10286) );
  INV_X1 U12096 ( .A(n9756), .ZN(n10619) );
  XNOR2_X1 U12097 ( .A(n10619), .B(n8606), .ZN(n8607) );
  OAI21_X1 U12098 ( .B1(n11544), .B2(n11545), .A(n11550), .ZN(n8692) );
  NAND3_X1 U12100 ( .A1(n9160), .A2(n8609), .A3(n9159), .ZN(n8612) );
  INV_X1 U12101 ( .A(n9879), .ZN(n8615) );
  XNOR2_X1 U12102 ( .A(n8615), .B(n10150), .ZN(n8627) );
  NOR2_X1 U12103 ( .A1(n9172), .A2(n8761), .ZN(n8616) );
  NAND2_X1 U12105 ( .A1(n9172), .A2(n9177), .ZN(n8619) );
  INV_X1 U12106 ( .A(n9176), .ZN(n8617) );
  NAND3_X1 U12107 ( .A1(n9005), .A2(n8895), .A3(n9007), .ZN(n8625) );
  NAND3_X1 U12108 ( .A1(n8623), .A2(n8891), .A3(n8622), .ZN(n8624) );
  INV_X1 U12110 ( .A(n8713), .ZN(n9239) );
  NAND3_X1 U12111 ( .A1(n266), .A2(n9239), .A3(n9186), .ZN(n8629) );
  OAI21_X1 U12112 ( .B1(n9233), .B2(n1041), .A(n19716), .ZN(n8634) );
  XNOR2_X1 U12113 ( .A(n10359), .B(n10582), .ZN(n9508) );
  XNOR2_X1 U12114 ( .A(n917), .B(n16487), .ZN(n8635) );
  NAND2_X1 U12117 ( .A1(n8933), .A2(n8747), .ZN(n8642) );
  AND3_X1 U12118 ( .A1(n8640), .A2(n8639), .A3(n8638), .ZN(n8641) );
  NAND2_X1 U12120 ( .A1(n111), .A2(n8937), .ZN(n8647) );
  OAI211_X1 U12121 ( .C1(n8644), .C2(n8937), .A(n8941), .B(n8945), .ZN(n8645)
         );
  INV_X1 U12122 ( .A(n8645), .ZN(n8646) );
  AOI21_X2 U12123 ( .B1(n8648), .B2(n8647), .A(n8646), .ZN(n10157) );
  XNOR2_X1 U12124 ( .A(n10157), .B(n10240), .ZN(n9360) );
  INV_X1 U12125 ( .A(n8649), .ZN(n9273) );
  OAI211_X1 U12126 ( .C1(n9273), .C2(n20265), .A(n9277), .B(n9275), .ZN(n8651)
         );
  NAND2_X1 U12127 ( .A1(n8771), .A2(n19710), .ZN(n8654) );
  XNOR2_X1 U12129 ( .A(n10351), .B(n10589), .ZN(n9523) );
  INV_X1 U12130 ( .A(n9523), .ZN(n8656) );
  XNOR2_X1 U12131 ( .A(n8656), .B(n9360), .ZN(n8664) );
  NOR2_X1 U12132 ( .A1(n8998), .A2(n19517), .ZN(n8659) );
  XNOR2_X1 U12133 ( .A(n9861), .B(n9862), .ZN(n8662) );
  XNOR2_X1 U12134 ( .A(n10236), .B(n18366), .ZN(n8661) );
  XNOR2_X1 U12135 ( .A(n8662), .B(n8661), .ZN(n8663) );
  XNOR2_X1 U12136 ( .A(n8664), .B(n8663), .ZN(n10760) );
  INV_X1 U12137 ( .A(n10760), .ZN(n11549) );
  INV_X1 U12138 ( .A(n10928), .ZN(n8689) );
  NOR2_X1 U12140 ( .A1(n20146), .A2(n8805), .ZN(n9781) );
  NAND3_X1 U12143 ( .A1(n9217), .A2(n1428), .A3(n9114), .ZN(n8668) );
  XNOR2_X1 U12144 ( .A(n10595), .B(n20161), .ZN(n9518) );
  OAI21_X1 U12145 ( .B1(n19857), .B2(n8672), .A(n8671), .ZN(n8673) );
  NAND2_X1 U12147 ( .A1(n8831), .A2(n9029), .ZN(n9032) );
  OAI21_X1 U12148 ( .B1(n9031), .B2(n9060), .A(n9032), .ZN(n8679) );
  INV_X1 U12149 ( .A(n9062), .ZN(n8830) );
  NAND2_X1 U12150 ( .A1(n8677), .A2(n9059), .ZN(n8678) );
  XNOR2_X1 U12152 ( .A(n10567), .B(n19806), .ZN(n9294) );
  XNOR2_X1 U12153 ( .A(n8680), .B(n9518), .ZN(n8687) );
  XNOR2_X1 U12154 ( .A(n10163), .B(n10203), .ZN(n8685) );
  NOR2_X1 U12155 ( .A1(n8338), .A2(n8786), .ZN(n8682) );
  XNOR2_X1 U12156 ( .A(n9777), .B(n18819), .ZN(n8684) );
  XNOR2_X1 U12157 ( .A(n8685), .B(n8684), .ZN(n8686) );
  XNOR2_X1 U12158 ( .A(n8687), .B(n8686), .ZN(n11548) );
  NAND2_X1 U12160 ( .A1(n647), .A2(n11546), .ZN(n8688) );
  NAND2_X1 U12161 ( .A1(n8689), .A2(n8688), .ZN(n8691) );
  NOR2_X1 U12162 ( .A1(n10926), .A2(n11546), .ZN(n8690) );
  NAND2_X1 U12164 ( .A1(n8987), .A2(n8761), .ZN(n8695) );
  OAI21_X1 U12165 ( .B1(n19827), .B2(n8695), .A(n8694), .ZN(n10043) );
  INV_X1 U12166 ( .A(n10497), .ZN(n9589) );
  XNOR2_X1 U12167 ( .A(n10043), .B(n9589), .ZN(n9524) );
  OAI21_X1 U12168 ( .B1(n9159), .B2(n9162), .A(n8609), .ZN(n8697) );
  INV_X1 U12169 ( .A(n8699), .ZN(n8704) );
  OAI21_X1 U12170 ( .B1(n19590), .B2(n9340), .A(n8700), .ZN(n9072) );
  NAND2_X1 U12171 ( .A1(n9072), .A2(n8701), .ZN(n8702) );
  OAI21_X1 U12172 ( .B1(n8704), .B2(n8703), .A(n8702), .ZN(n9685) );
  XNOR2_X1 U12173 ( .A(n10280), .B(n9685), .ZN(n9651) );
  XNOR2_X1 U12174 ( .A(n9524), .B(n9651), .ZN(n8719) );
  NAND2_X1 U12175 ( .A1(n269), .A2(n9168), .ZN(n9081) );
  INV_X1 U12176 ( .A(n9168), .ZN(n8706) );
  OAI211_X1 U12177 ( .C1(n9171), .C2(n9166), .A(n264), .B(n8706), .ZN(n8707)
         );
  NAND3_X1 U12178 ( .A1(n2097), .A2(n8411), .A3(n1041), .ZN(n8710) );
  OAI211_X1 U12179 ( .C1(n8712), .C2(n8711), .A(n8710), .B(n9236), .ZN(n10088)
         );
  XNOR2_X1 U12180 ( .A(n9908), .B(n10088), .ZN(n8717) );
  XNOR2_X1 U12181 ( .A(n8717), .B(n8716), .ZN(n8718) );
  OAI22_X1 U12182 ( .A1(n8721), .A2(n8720), .B1(n8905), .B2(n9358), .ZN(n8725)
         );
  NOR2_X1 U12183 ( .A1(n19941), .A2(n8904), .ZN(n8723) );
  XNOR2_X1 U12184 ( .A(n10273), .B(n10126), .ZN(n9632) );
  NOR2_X1 U12185 ( .A1(n8729), .A2(n8937), .ZN(n8732) );
  NOR3_X1 U12186 ( .A1(n8917), .A2(n8736), .A3(n8735), .ZN(n8737) );
  AOI21_X1 U12187 ( .B1(n8738), .B2(n3645), .A(n8737), .ZN(n8739) );
  XNOR2_X1 U12188 ( .A(n9632), .B(n8740), .ZN(n8757) );
  NOR2_X1 U12189 ( .A1(n8741), .A2(n8950), .ZN(n9371) );
  NAND2_X1 U12190 ( .A1(n8482), .A2(n8743), .ZN(n8744) );
  XNOR2_X1 U12192 ( .A(n10213), .B(n2151), .ZN(n8755) );
  NOR2_X1 U12193 ( .A1(n8932), .A2(n8747), .ZN(n8751) );
  NOR2_X1 U12194 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  XNOR2_X1 U12196 ( .A(n9952), .B(n10491), .ZN(n9507) );
  XNOR2_X1 U12197 ( .A(n8755), .B(n9507), .ZN(n8756) );
  INV_X1 U12199 ( .A(n9172), .ZN(n8765) );
  INV_X1 U12200 ( .A(n8761), .ZN(n9178) );
  NOR2_X1 U12201 ( .A1(n19827), .A2(n9178), .ZN(n8762) );
  OAI21_X1 U12202 ( .B1(n8763), .B2(n8762), .A(n9177), .ZN(n8764) );
  OAI21_X1 U12203 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n10071) );
  XNOR2_X1 U12204 ( .A(n9894), .B(n10071), .ZN(n8770) );
  AOI22_X1 U12205 ( .A1(n8768), .A2(n9008), .B1(n8767), .B2(n9004), .ZN(n9710)
         );
  XNOR2_X1 U12206 ( .A(n9600), .B(n9710), .ZN(n9538) );
  XNOR2_X1 U12207 ( .A(n8770), .B(n9538), .ZN(n8778) );
  OAI21_X1 U12208 ( .B1(n8773), .B2(n8772), .A(n8997), .ZN(n8774) );
  NAND2_X1 U12209 ( .A1(n8774), .A2(n3518), .ZN(n8775) );
  XNOR2_X1 U12211 ( .A(n8777), .B(n8778), .ZN(n10640) );
  NOR2_X1 U12212 ( .A1(n9107), .A2(n9105), .ZN(n8784) );
  OAI21_X1 U12213 ( .B1(n8779), .B2(n20000), .A(n9111), .ZN(n8783) );
  INV_X1 U12214 ( .A(n8872), .ZN(n8781) );
  NAND3_X1 U12215 ( .A1(n1960), .A2(n8781), .A3(n9106), .ZN(n8782) );
  INV_X1 U12217 ( .A(n8790), .ZN(n9148) );
  INV_X1 U12218 ( .A(n8789), .ZN(n8792) );
  NOR2_X1 U12219 ( .A1(n9145), .A2(n8790), .ZN(n8791) );
  XNOR2_X1 U12220 ( .A(n20211), .B(n9771), .ZN(n8802) );
  INV_X1 U12221 ( .A(n8793), .ZN(n8794) );
  AND3_X1 U12222 ( .A1(n1603), .A2(n8794), .A3(n9217), .ZN(n8800) );
  INV_X1 U12223 ( .A(n8796), .ZN(n8799) );
  AND2_X1 U12224 ( .A1(n9114), .A2(n8797), .ZN(n8798) );
  XNOR2_X1 U12225 ( .A(n10247), .B(n2382), .ZN(n8801) );
  XNOR2_X1 U12226 ( .A(n8802), .B(n8801), .ZN(n8822) );
  NAND2_X1 U12227 ( .A1(n8803), .A2(n9135), .ZN(n8804) );
  NAND2_X1 U12228 ( .A1(n9204), .A2(n8665), .ZN(n8809) );
  NOR2_X1 U12229 ( .A1(n9129), .A2(n8276), .ZN(n8806) );
  OAI21_X1 U12230 ( .B1(n9202), .B2(n8806), .A(n3542), .ZN(n8808) );
  NAND2_X1 U12231 ( .A1(n9782), .A2(n9129), .ZN(n8807) );
  OAI211_X1 U12232 ( .C1(n9780), .C2(n8809), .A(n8808), .B(n8807), .ZN(n9691)
         );
  XNOR2_X1 U12233 ( .A(n9691), .B(n10296), .ZN(n8820) );
  MUX2_X1 U12234 ( .A(n8811), .B(n8810), .S(n8815), .Z(n8819) );
  NAND2_X1 U12235 ( .A1(n9122), .A2(n8812), .ZN(n8817) );
  NAND3_X1 U12236 ( .A1(n8815), .A2(n8814), .A3(n8813), .ZN(n8816) );
  XNOR2_X1 U12237 ( .A(n10506), .B(n10404), .ZN(n9514) );
  XNOR2_X1 U12238 ( .A(n9514), .B(n8820), .ZN(n8821) );
  MUX2_X1 U12239 ( .A(n8823), .B(n9228), .S(n9313), .Z(n8827) );
  NAND2_X1 U12240 ( .A1(n9305), .A2(n9228), .ZN(n8825) );
  OAI21_X1 U12241 ( .B1(n9307), .B2(n8827), .A(n8826), .ZN(n9668) );
  XNOR2_X1 U12242 ( .A(n10261), .B(n9668), .ZN(n9625) );
  INV_X1 U12243 ( .A(n9031), .ZN(n9061) );
  NAND3_X1 U12244 ( .A1(n9061), .A2(n9060), .A3(n9029), .ZN(n8835) );
  INV_X1 U12245 ( .A(n9060), .ZN(n9028) );
  NAND2_X1 U12246 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  NAND3_X1 U12247 ( .A1(n8833), .A2(n9029), .A3(n9028), .ZN(n8834) );
  XNOR2_X1 U12248 ( .A(n9934), .B(n10472), .ZN(n9499) );
  XNOR2_X1 U12249 ( .A(n9625), .B(n9499), .ZN(n8859) );
  MUX2_X1 U12250 ( .A(n8839), .B(n8838), .S(n19857), .Z(n8840) );
  NAND2_X1 U12251 ( .A1(n2984), .A2(n9018), .ZN(n8844) );
  INV_X1 U12252 ( .A(n8842), .ZN(n8843) );
  OAI22_X1 U12253 ( .A1(n8845), .A2(n8844), .B1(n8843), .B2(n20472), .ZN(n8847) );
  XNOR2_X1 U12255 ( .A(n9623), .B(n10422), .ZN(n9407) );
  NOR2_X1 U12256 ( .A1(n9046), .A2(n8848), .ZN(n9040) );
  NOR2_X1 U12257 ( .A1(n9046), .A2(n9038), .ZN(n8850) );
  MUX2_X1 U12258 ( .A(n9040), .B(n8850), .S(n8849), .Z(n8856) );
  NOR2_X1 U12259 ( .A1(n8852), .A2(n8851), .ZN(n8854) );
  NOR2_X1 U12260 ( .A1(n1933), .A2(n9039), .ZN(n8853) );
  XNOR2_X1 U12262 ( .A(n20483), .B(n19467), .ZN(n8857) );
  XNOR2_X1 U12263 ( .A(n9407), .B(n8857), .ZN(n8858) );
  XNOR2_X1 U12264 ( .A(n8858), .B(n8859), .ZN(n10638) );
  INV_X1 U12265 ( .A(n9066), .ZN(n9321) );
  NOR2_X1 U12266 ( .A1(n9837), .A2(n9065), .ZN(n8862) );
  OR2_X1 U12267 ( .A1(n9317), .A2(n9066), .ZN(n8861) );
  AOI22_X1 U12268 ( .A1(n8862), .A2(n9069), .B1(n8861), .B2(n9065), .ZN(n8863)
         );
  INV_X1 U12269 ( .A(n8866), .ZN(n9327) );
  OAI21_X1 U12270 ( .B1(n8866), .B2(n9326), .A(n9074), .ZN(n8865) );
  NAND2_X1 U12271 ( .A1(n8865), .A2(n9329), .ZN(n8868) );
  OAI211_X2 U12273 ( .C1(n8869), .C2(n9327), .A(n8868), .B(n8867), .ZN(n10204)
         );
  XNOR2_X1 U12274 ( .A(n10594), .B(n10204), .ZN(n8878) );
  NAND2_X1 U12276 ( .A1(n8872), .A2(n19515), .ZN(n8876) );
  OAI21_X1 U12277 ( .B1(n8872), .B2(n9106), .A(n9105), .ZN(n8870) );
  NAND2_X1 U12278 ( .A1(n8871), .A2(n8870), .ZN(n8875) );
  NOR2_X1 U12279 ( .A1(n8781), .A2(n20000), .ZN(n8873) );
  OAI211_X2 U12280 ( .C1(n1960), .C2(n8876), .A(n8875), .B(n8874), .ZN(n10388)
         );
  INV_X1 U12281 ( .A(n10572), .ZN(n8877) );
  XNOR2_X1 U12282 ( .A(n8877), .B(n10388), .ZN(n9520) );
  XNOR2_X1 U12283 ( .A(n8878), .B(n9520), .ZN(n8900) );
  INV_X1 U12284 ( .A(n8972), .ZN(n9251) );
  NAND2_X1 U12285 ( .A1(n19516), .A2(n9249), .ZN(n8883) );
  NAND2_X1 U12286 ( .A1(n8974), .A2(n8879), .ZN(n8882) );
  OAI21_X1 U12287 ( .B1(n9252), .B2(n8972), .A(n670), .ZN(n8881) );
  INV_X1 U12288 ( .A(n8884), .ZN(n9452) );
  AND3_X1 U12289 ( .A1(n8887), .A2(n8886), .A3(n8885), .ZN(n8888) );
  XNOR2_X1 U12290 ( .A(n9429), .B(n9922), .ZN(n8898) );
  INV_X1 U12291 ( .A(n9008), .ZN(n8896) );
  OAI21_X1 U12292 ( .B1(n9004), .B2(n9008), .A(n19490), .ZN(n8893) );
  NAND2_X1 U12293 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  OAI21_X1 U12294 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n9926) );
  XNOR2_X1 U12295 ( .A(n9926), .B(n2323), .ZN(n8897) );
  XNOR2_X1 U12296 ( .A(n8898), .B(n8897), .ZN(n8899) );
  NAND2_X1 U12297 ( .A1(n11538), .A2(n11532), .ZN(n8901) );
  MUX2_X1 U12298 ( .A(n8902), .B(n8901), .S(n11534), .Z(n8903) );
  NAND2_X1 U12299 ( .A1(n8907), .A2(n8906), .ZN(n8915) );
  INV_X1 U12300 ( .A(n8908), .ZN(n8914) );
  INV_X1 U12301 ( .A(n8909), .ZN(n8913) );
  NAND2_X1 U12302 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  NAND4_X1 U12303 ( .A1(n8915), .A2(n8914), .A3(n8913), .A4(n8912), .ZN(n8919)
         );
  NAND4_X1 U12304 ( .A1(n8921), .A2(n8920), .A3(n8919), .A4(n8918), .ZN(n8922)
         );
  NOR2_X1 U12305 ( .A1(n8932), .A2(n8931), .ZN(n8927) );
  INV_X1 U12306 ( .A(n8924), .ZN(n8926) );
  NAND2_X1 U12309 ( .A1(n8932), .A2(n8931), .ZN(n8934) );
  XNOR2_X1 U12310 ( .A(n9624), .B(n20484), .ZN(n9456) );
  XNOR2_X1 U12311 ( .A(n8936), .B(n9456), .ZN(n8969) );
  NAND2_X1 U12313 ( .A1(n8953), .A2(n904), .ZN(n8955) );
  NAND3_X1 U12314 ( .A1(n8953), .A2(n8952), .A3(n8482), .ZN(n8954) );
  OAI21_X1 U12315 ( .B1(n8956), .B2(n8955), .A(n8954), .ZN(n8957) );
  XNOR2_X1 U12316 ( .A(n10527), .B(n9670), .ZN(n9421) );
  NOR2_X1 U12317 ( .A1(n9362), .A2(n8961), .ZN(n8962) );
  NAND2_X1 U12318 ( .A1(n8962), .A2(n9363), .ZN(n8963) );
  NAND2_X1 U12319 ( .A1(n8964), .A2(n8963), .ZN(n8967) );
  NOR2_X1 U12320 ( .A1(n8965), .A2(n8726), .ZN(n8966) );
  NOR2_X2 U12321 ( .A1(n8967), .A2(n8966), .ZN(n9869) );
  XNOR2_X1 U12322 ( .A(n9421), .B(n9869), .ZN(n8968) );
  XNOR2_X1 U12323 ( .A(n8969), .B(n8968), .ZN(n9017) );
  NOR2_X1 U12324 ( .A1(n9256), .A2(n9255), .ZN(n8973) );
  AND2_X1 U12325 ( .A1(n8973), .A2(n8974), .ZN(n8975) );
  AND2_X1 U12326 ( .A1(n8979), .A2(n19710), .ZN(n8980) );
  NAND2_X1 U12327 ( .A1(n8984), .A2(n8980), .ZN(n8982) );
  OAI211_X1 U12328 ( .C1(n8984), .C2(n8983), .A(n8982), .B(n3797), .ZN(n9398)
         );
  INV_X1 U12329 ( .A(n9398), .ZN(n10094) );
  XNOR2_X1 U12330 ( .A(n9692), .B(n10094), .ZN(n8994) );
  NAND2_X1 U12331 ( .A1(n9177), .A2(n8987), .ZN(n8989) );
  OAI21_X1 U12332 ( .B1(n265), .B2(n9178), .A(n9172), .ZN(n8986) );
  NAND2_X1 U12333 ( .A1(n265), .A2(n9176), .ZN(n9175) );
  MUX2_X1 U12334 ( .A(n8987), .B(n8986), .S(n9175), .Z(n8988) );
  OAI21_X1 U12335 ( .B1(n9172), .B2(n8989), .A(n8988), .ZN(n10613) );
  XNOR2_X1 U12336 ( .A(n10441), .B(n10613), .ZN(n10257) );
  XNOR2_X1 U12337 ( .A(n10257), .B(n8994), .ZN(n9016) );
  MUX2_X1 U12338 ( .A(n19517), .B(n8998), .S(n8997), .Z(n9001) );
  NAND3_X1 U12339 ( .A1(n8999), .A2(n8998), .A3(n8997), .ZN(n9000) );
  OAI21_X1 U12340 ( .B1(n9001), .B2(n8657), .A(n9000), .ZN(n9002) );
  XNOR2_X1 U12341 ( .A(n10026), .B(n2248), .ZN(n9014) );
  INV_X1 U12342 ( .A(n9010), .ZN(n9013) );
  OAI21_X1 U12343 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n9012) );
  XNOR2_X1 U12344 ( .A(n10008), .B(n9771), .ZN(n9446) );
  XNOR2_X1 U12345 ( .A(n9446), .B(n9014), .ZN(n9015) );
  XNOR2_X1 U12346 ( .A(n9016), .B(n9015), .ZN(n11553) );
  NOR2_X1 U12348 ( .A1(n9304), .A2(n9018), .ZN(n9020) );
  AND2_X1 U12349 ( .A1(n19857), .A2(n9021), .ZN(n9027) );
  INV_X1 U12350 ( .A(n9022), .ZN(n9026) );
  NOR2_X1 U12351 ( .A1(n9062), .A2(n9029), .ZN(n9030) );
  NOR2_X1 U12352 ( .A1(n9034), .A2(n9030), .ZN(n9036) );
  INV_X1 U12353 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U12354 ( .A1(n9034), .A2(n9033), .ZN(n9035) );
  XNOR2_X1 U12355 ( .A(n9908), .B(n9991), .ZN(n9469) );
  XNOR2_X1 U12356 ( .A(n10242), .B(n9469), .ZN(n9058) );
  INV_X1 U12357 ( .A(n9037), .ZN(n9043) );
  NOR2_X1 U12358 ( .A1(n9039), .A2(n9038), .ZN(n9042) );
  INV_X1 U12359 ( .A(n9040), .ZN(n9041) );
  OAI21_X1 U12360 ( .B1(n9043), .B2(n9042), .A(n9041), .ZN(n9044) );
  NOR2_X1 U12361 ( .A1(n9049), .A2(n9576), .ZN(n9050) );
  XNOR2_X1 U12362 ( .A(n10046), .B(n10350), .ZN(n9056) );
  NAND2_X1 U12363 ( .A1(n1751), .A2(n20011), .ZN(n9226) );
  XNOR2_X1 U12365 ( .A(n10087), .B(n2385), .ZN(n9055) );
  XNOR2_X1 U12366 ( .A(n9056), .B(n9055), .ZN(n9057) );
  XNOR2_X1 U12367 ( .A(n9058), .B(n9057), .ZN(n10913) );
  AOI21_X1 U12368 ( .B1(n9061), .B2(n9060), .A(n9059), .ZN(n9064) );
  OAI21_X1 U12369 ( .B1(n9317), .B2(n9065), .A(n9837), .ZN(n9068) );
  AND3_X1 U12370 ( .A1(n20476), .A2(n9837), .A3(n9066), .ZN(n9067) );
  XNOR2_X1 U12371 ( .A(n865), .B(n10220), .ZN(n9415) );
  INV_X1 U12372 ( .A(n9070), .ZN(n9339) );
  OAI21_X1 U12373 ( .B1(n19590), .B2(n9564), .A(n9563), .ZN(n9071) );
  AOI22_X1 U12374 ( .A1(n9075), .A2(n9329), .B1(n9074), .B2(n9333), .ZN(n9079)
         );
  XNOR2_X1 U12377 ( .A(n9414), .B(n10382), .ZN(n9674) );
  XNOR2_X1 U12378 ( .A(n9415), .B(n9674), .ZN(n9097) );
  AOI21_X1 U12379 ( .B1(n1027), .B2(n9081), .A(n9080), .ZN(n9084) );
  XNOR2_X1 U12381 ( .A(n20134), .B(n9986), .ZN(n9464) );
  NOR2_X1 U12382 ( .A1(n9087), .A2(n20010), .ZN(n9094) );
  NAND2_X1 U12383 ( .A1(n9089), .A2(n9088), .ZN(n9093) );
  NAND3_X1 U12384 ( .A1(n9452), .A2(n9091), .A3(n9090), .ZN(n9092) );
  XNOR2_X1 U12386 ( .A(n10027), .B(n19222), .ZN(n9095) );
  XNOR2_X1 U12387 ( .A(n9464), .B(n9095), .ZN(n9096) );
  AOI21_X1 U12390 ( .B1(n19564), .B2(n10913), .A(n19957), .ZN(n9098) );
  NAND3_X1 U12391 ( .A1(n9107), .A2(n9106), .A3(n9105), .ZN(n9108) );
  OAI211_X1 U12392 ( .C1(n9111), .C2(n9110), .A(n9109), .B(n9108), .ZN(n10578)
         );
  NAND3_X1 U12393 ( .A1(n1056), .A2(n8795), .A3(n9112), .ZN(n9117) );
  XNOR2_X1 U12394 ( .A(n10578), .B(n10154), .ZN(n10210) );
  NAND2_X1 U12395 ( .A1(n9120), .A2(n9119), .ZN(n9126) );
  AOI22_X1 U12396 ( .A1(n9124), .A2(n9128), .B1(n9123), .B2(n9122), .ZN(n9125)
         );
  XNOR2_X1 U12397 ( .A(n10079), .B(n9902), .ZN(n9477) );
  XNOR2_X1 U12398 ( .A(n20491), .B(n9477), .ZN(n9156) );
  NAND2_X1 U12399 ( .A1(n9780), .A2(n3542), .ZN(n9132) );
  INV_X1 U12402 ( .A(n9134), .ZN(n9142) );
  NOR2_X1 U12403 ( .A1(n9211), .A2(n9214), .ZN(n9136) );
  NAND2_X1 U12404 ( .A1(n9213), .A2(n9136), .ZN(n9141) );
  AND2_X1 U12405 ( .A1(n9137), .A2(n9214), .ZN(n9139) );
  AOI22_X1 U12406 ( .A1(n9213), .A2(n9139), .B1(n9138), .B2(n9211), .ZN(n9140)
         );
  XNOR2_X1 U12407 ( .A(n19945), .B(n10358), .ZN(n9154) );
  NOR2_X1 U12408 ( .A1(n9144), .A2(n9143), .ZN(n9152) );
  XNOR2_X1 U12410 ( .A(n10061), .B(n20394), .ZN(n9153) );
  XNOR2_X1 U12411 ( .A(n9154), .B(n9153), .ZN(n9155) );
  NAND2_X1 U12412 ( .A1(n10913), .A2(n11556), .ZN(n10645) );
  OR2_X1 U12413 ( .A1(n10645), .A2(n9017), .ZN(n9200) );
  INV_X1 U12414 ( .A(n11556), .ZN(n11162) );
  AND2_X1 U12415 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  OAI21_X1 U12416 ( .B1(n9167), .B2(n9171), .A(n9166), .ZN(n9170) );
  NAND2_X1 U12417 ( .A1(n264), .A2(n9168), .ZN(n9169) );
  NAND2_X1 U12418 ( .A1(n264), .A2(n9171), .ZN(n10328) );
  XNOR2_X1 U12420 ( .A(n9587), .B(n10052), .ZN(n9179) );
  OAI21_X1 U12421 ( .B1(n9172), .B2(n9177), .A(n2243), .ZN(n9174) );
  INV_X1 U12422 ( .A(n9177), .ZN(n9173) );
  XNOR2_X1 U12423 ( .A(n9926), .B(n9643), .ZN(n9480) );
  XNOR2_X1 U12424 ( .A(n9480), .B(n9179), .ZN(n9198) );
  NAND2_X1 U12425 ( .A1(n9234), .A2(n19716), .ZN(n9180) );
  AOI21_X1 U12426 ( .B1(n9183), .B2(n9182), .A(n9234), .ZN(n9184) );
  NAND2_X1 U12427 ( .A1(n9186), .A2(n9241), .ZN(n9187) );
  AOI21_X1 U12428 ( .B1(n9188), .B2(n9187), .A(n9242), .ZN(n9703) );
  OR2_X1 U12429 ( .A1(n9703), .A2(n9700), .ZN(n10166) );
  XNOR2_X1 U12430 ( .A(n10166), .B(n10571), .ZN(n10201) );
  OAI21_X1 U12431 ( .B1(n9339), .B2(n9563), .A(n9342), .ZN(n9192) );
  NOR2_X1 U12432 ( .A1(n9192), .A2(n9191), .ZN(n9195) );
  AOI21_X1 U12433 ( .B1(n8701), .B2(n9193), .A(n9339), .ZN(n9194) );
  XNOR2_X1 U12434 ( .A(n10107), .B(n2023), .ZN(n9196) );
  XNOR2_X1 U12435 ( .A(n10201), .B(n9196), .ZN(n9197) );
  XNOR2_X1 U12436 ( .A(n9197), .B(n9198), .ZN(n11559) );
  INV_X1 U12437 ( .A(n11559), .ZN(n10914) );
  NAND3_X1 U12438 ( .A1(n19957), .A2(n11162), .A3(n10914), .ZN(n9199) );
  NAND2_X1 U12439 ( .A1(n12354), .A2(n12349), .ZN(n11032) );
  XNOR2_X1 U12440 ( .A(n10229), .B(n18779), .ZN(n9206) );
  XNOR2_X1 U12441 ( .A(n19746), .B(n9206), .ZN(n9207) );
  XNOR2_X1 U12442 ( .A(n9208), .B(n9207), .ZN(n9225) );
  XNOR2_X1 U12443 ( .A(n9977), .B(n9937), .ZN(n10098) );
  NAND2_X1 U12444 ( .A1(n9218), .A2(n1056), .ZN(n9216) );
  OAI21_X1 U12445 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(n9223) );
  NOR2_X1 U12446 ( .A1(n9220), .A2(n9219), .ZN(n9222) );
  XNOR2_X1 U12447 ( .A(n10098), .B(n10473), .ZN(n9224) );
  INV_X1 U12448 ( .A(n9305), .ZN(n9308) );
  AOI21_X1 U12449 ( .B1(n9227), .B2(n9226), .A(n9308), .ZN(n9231) );
  INV_X1 U12450 ( .A(n9228), .ZN(n9306) );
  AOI21_X1 U12451 ( .B1(n9229), .B2(n20011), .A(n9306), .ZN(n9230) );
  XNOR2_X1 U12452 ( .A(n10417), .B(n9232), .ZN(n9248) );
  INV_X1 U12453 ( .A(n9234), .ZN(n9235) );
  XNOR2_X1 U12454 ( .A(n10484), .B(n10027), .ZN(n9246) );
  XNOR2_X1 U12456 ( .A(n9854), .B(n17365), .ZN(n9245) );
  XNOR2_X1 U12457 ( .A(n9246), .B(n9245), .ZN(n9247) );
  XNOR2_X1 U12458 ( .A(n9248), .B(n9247), .ZN(n9351) );
  NAND2_X1 U12459 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  NAND3_X1 U12460 ( .A1(n9260), .A2(n670), .A3(n9253), .ZN(n9258) );
  NAND3_X1 U12461 ( .A1(n19516), .A2(n9256), .A3(n9255), .ZN(n9257) );
  XNOR2_X1 U12462 ( .A(n10462), .B(n9261), .ZN(n9286) );
  INV_X1 U12463 ( .A(n9264), .ZN(n9269) );
  NOR2_X1 U12464 ( .A1(n9266), .A2(n9265), .ZN(n9268) );
  XNOR2_X1 U12466 ( .A(n19718), .B(n10360), .ZN(n9284) );
  XNOR2_X1 U12467 ( .A(n10061), .B(n2383), .ZN(n9283) );
  XNOR2_X1 U12468 ( .A(n9284), .B(n9283), .ZN(n9285) );
  XNOR2_X2 U12469 ( .A(n9286), .B(n9285), .ZN(n11174) );
  NOR2_X1 U12470 ( .A1(n19715), .A2(n9576), .ZN(n9288) );
  AOI22_X1 U12471 ( .A1(n9578), .A2(n9291), .B1(n9577), .B2(n9290), .ZN(n9292)
         );
  NAND2_X1 U12472 ( .A1(n9582), .A2(n9292), .ZN(n9293) );
  XNOR2_X1 U12473 ( .A(n9293), .B(n9430), .ZN(n10453) );
  XNOR2_X1 U12474 ( .A(n9294), .B(n10453), .ZN(n9316) );
  INV_X1 U12475 ( .A(n9299), .ZN(n9301) );
  NAND2_X1 U12476 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  MUX2_X1 U12477 ( .A(n9306), .B(n9307), .S(n9305), .Z(n9314) );
  NAND3_X1 U12478 ( .A1(n9308), .A2(n9307), .A3(n1751), .ZN(n9312) );
  NAND2_X1 U12479 ( .A1(n20011), .A2(n9309), .ZN(n9311) );
  XNOR2_X1 U12480 ( .A(n10205), .B(n2401), .ZN(n9315) );
  NAND2_X1 U12481 ( .A1(n20505), .A2(n9837), .ZN(n9320) );
  NOR2_X1 U12482 ( .A1(n9837), .A2(n9317), .ZN(n9318) );
  NOR2_X1 U12483 ( .A1(n9321), .A2(n9836), .ZN(n9322) );
  XNOR2_X1 U12484 ( .A(n9324), .B(n9325), .ZN(n9350) );
  NAND2_X1 U12485 ( .A1(n9329), .A2(n3800), .ZN(n9335) );
  NOR2_X1 U12486 ( .A1(n9331), .A2(n9330), .ZN(n9332) );
  NAND2_X1 U12487 ( .A1(n9333), .A2(n9332), .ZN(n9334) );
  XNOR2_X1 U12488 ( .A(n10248), .B(n18854), .ZN(n9348) );
  NAND2_X1 U12489 ( .A1(n9339), .A2(n9338), .ZN(n9566) );
  NAND3_X1 U12490 ( .A1(n19590), .A2(n9346), .A3(n9340), .ZN(n9343) );
  NAND3_X1 U12491 ( .A1(n9342), .A2(n9341), .A3(n9563), .ZN(n9568) );
  AND2_X1 U12492 ( .A1(n9343), .A2(n9568), .ZN(n9345) );
  NAND3_X1 U12493 ( .A1(n9564), .A2(n9346), .A3(n9563), .ZN(n9344) );
  OAI211_X1 U12494 ( .C1(n9346), .C2(n9566), .A(n9345), .B(n9344), .ZN(n9347)
         );
  XNOR2_X1 U12495 ( .A(n9957), .B(n9347), .ZN(n10447) );
  XNOR2_X1 U12496 ( .A(n9348), .B(n10447), .ZN(n9349) );
  XNOR2_X1 U12497 ( .A(n9350), .B(n9349), .ZN(n11175) );
  NOR2_X1 U12498 ( .A1(n11175), .A2(n11178), .ZN(n9379) );
  NOR2_X1 U12499 ( .A1(n19941), .A2(n2756), .ZN(n9355) );
  XNOR2_X1 U12500 ( .A(n10436), .B(n9648), .ZN(n10085) );
  XNOR2_X1 U12501 ( .A(n10085), .B(n9360), .ZN(n9377) );
  NOR2_X1 U12502 ( .A1(n9362), .A2(n9361), .ZN(n9365) );
  XNOR2_X1 U12503 ( .A(n10349), .B(n10046), .ZN(n9375) );
  INV_X1 U12504 ( .A(n9367), .ZN(n9369) );
  NAND2_X1 U12505 ( .A1(n9373), .A2(n9372), .ZN(n10498) );
  XNOR2_X1 U12506 ( .A(n10498), .B(n345), .ZN(n9374) );
  XNOR2_X1 U12507 ( .A(n9375), .B(n9374), .ZN(n9376) );
  NOR3_X1 U12508 ( .A1(n12002), .A2(n12001), .A3(n19769), .ZN(n9380) );
  XNOR2_X1 U12509 ( .A(n9383), .B(n10002), .ZN(n9679) );
  XNOR2_X1 U12510 ( .A(n10077), .B(n10273), .ZN(n10409) );
  XNOR2_X1 U12511 ( .A(n10409), .B(n9679), .ZN(n9386) );
  XNOR2_X1 U12512 ( .A(n9824), .B(n10061), .ZN(n9728) );
  XNOR2_X1 U12513 ( .A(n10213), .B(n2347), .ZN(n9384) );
  XNOR2_X1 U12514 ( .A(n9728), .B(n9384), .ZN(n9385) );
  XNOR2_X1 U12515 ( .A(n9386), .B(n9385), .ZN(n11283) );
  INV_X1 U12516 ( .A(n11283), .ZN(n11282) );
  XNOR2_X1 U12517 ( .A(n10240), .B(n10088), .ZN(n10433) );
  XNOR2_X1 U12518 ( .A(n9812), .B(n10046), .ZN(n9387) );
  XNOR2_X1 U12519 ( .A(n10397), .B(n9388), .ZN(n9389) );
  INV_X1 U12520 ( .A(n10199), .ZN(n9392) );
  XNOR2_X1 U12521 ( .A(n10107), .B(n9429), .ZN(n10392) );
  XNOR2_X1 U12522 ( .A(n10392), .B(n10454), .ZN(n9396) );
  XNOR2_X1 U12523 ( .A(n9923), .B(n10204), .ZN(n9394) );
  XNOR2_X1 U12524 ( .A(n10052), .B(n404), .ZN(n9393) );
  XNOR2_X1 U12525 ( .A(n9394), .B(n9393), .ZN(n9395) );
  XNOR2_X1 U12526 ( .A(n9396), .B(n9395), .ZN(n10693) );
  INV_X1 U12527 ( .A(n10693), .ZN(n11281) );
  INV_X1 U12529 ( .A(n20210), .ZN(n9397) );
  XNOR2_X1 U12530 ( .A(n9397), .B(n10254), .ZN(n10444) );
  XNOR2_X1 U12531 ( .A(n10026), .B(n9817), .ZN(n9717) );
  XNOR2_X1 U12532 ( .A(n10444), .B(n9717), .ZN(n9401) );
  XNOR2_X1 U12533 ( .A(n10247), .B(n2222), .ZN(n9399) );
  XNOR2_X1 U12534 ( .A(n10406), .B(n9399), .ZN(n9400) );
  XNOR2_X1 U12535 ( .A(n9401), .B(n9400), .ZN(n9559) );
  XNOR2_X1 U12536 ( .A(n10027), .B(n9799), .ZN(n9713) );
  INV_X1 U12537 ( .A(n9402), .ZN(n10219) );
  XNOR2_X1 U12538 ( .A(n10219), .B(n19818), .ZN(n10416) );
  XNOR2_X1 U12539 ( .A(n20268), .B(n9713), .ZN(n9406) );
  XNOR2_X1 U12540 ( .A(n9894), .B(n10382), .ZN(n9403) );
  XNOR2_X1 U12541 ( .A(n9404), .B(n9403), .ZN(n9405) );
  NAND2_X1 U12542 ( .A1(n9559), .A2(n10995), .ZN(n9411) );
  XNOR2_X1 U12543 ( .A(n9869), .B(n10261), .ZN(n10036) );
  XNOR2_X1 U12544 ( .A(n10036), .B(n9407), .ZN(n9410) );
  XNOR2_X1 U12545 ( .A(n10421), .B(n2221), .ZN(n9408) );
  INV_X1 U12546 ( .A(n9794), .ZN(n9458) );
  XNOR2_X1 U12547 ( .A(n20608), .B(n19746), .ZN(n9733) );
  XNOR2_X1 U12548 ( .A(n9408), .B(n9733), .ZN(n9409) );
  XNOR2_X1 U12549 ( .A(n9415), .B(n10321), .ZN(n9419) );
  XNOR2_X1 U12550 ( .A(n9416), .B(n9417), .ZN(n9418) );
  XNOR2_X2 U12551 ( .A(n9419), .B(n9418), .ZN(n11278) );
  INV_X1 U12552 ( .A(n11278), .ZN(n10688) );
  XNOR2_X1 U12553 ( .A(n9420), .B(n10261), .ZN(n9422) );
  INV_X1 U12554 ( .A(n9421), .ZN(n10233) );
  XNOR2_X1 U12555 ( .A(n9422), .B(n10233), .ZN(n9425) );
  XNOR2_X1 U12556 ( .A(n10229), .B(n9669), .ZN(n10342) );
  XNOR2_X1 U12557 ( .A(n9937), .B(n2164), .ZN(n9423) );
  XNOR2_X1 U12558 ( .A(n10342), .B(n9423), .ZN(n9424) );
  INV_X1 U12559 ( .A(n9861), .ZN(n9426) );
  XNOR2_X1 U12560 ( .A(n9426), .B(n10558), .ZN(n10588) );
  XNOR2_X1 U12561 ( .A(n9648), .B(n10349), .ZN(n9427) );
  XNOR2_X1 U12562 ( .A(n9427), .B(n10350), .ZN(n9944) );
  XNOR2_X1 U12563 ( .A(n9697), .B(n9856), .ZN(n10334) );
  XNOR2_X1 U12564 ( .A(n10334), .B(n10201), .ZN(n9431) );
  XNOR2_X1 U12565 ( .A(n9432), .B(n9431), .ZN(n11413) );
  INV_X1 U12566 ( .A(n11413), .ZN(n9547) );
  INV_X1 U12567 ( .A(n10248), .ZN(n9846) );
  XNOR2_X1 U12568 ( .A(n9846), .B(n9692), .ZN(n10371) );
  XNOR2_X1 U12569 ( .A(n10296), .B(n19760), .ZN(n9661) );
  XNOR2_X1 U12570 ( .A(n9842), .B(n18065), .ZN(n9433) );
  XNOR2_X1 U12571 ( .A(n9661), .B(n9433), .ZN(n9434) );
  XNOR2_X1 U12572 ( .A(n10257), .B(n9434), .ZN(n9435) );
  XNOR2_X1 U12573 ( .A(n9435), .B(n10371), .ZN(n11411) );
  NAND2_X1 U12574 ( .A1(n11276), .A2(n11411), .ZN(n9444) );
  XNOR2_X1 U12575 ( .A(n10210), .B(n10150), .ZN(n9438) );
  INV_X1 U12576 ( .A(n10273), .ZN(n9436) );
  XNOR2_X1 U12577 ( .A(n9436), .B(n2394), .ZN(n9437) );
  XNOR2_X1 U12578 ( .A(n9438), .B(n9437), .ZN(n9441) );
  XNOR2_X1 U12579 ( .A(n928), .B(n9635), .ZN(n9440) );
  INV_X1 U12580 ( .A(n10360), .ZN(n9439) );
  XNOR2_X1 U12581 ( .A(n9441), .B(n926), .ZN(n9545) );
  INV_X1 U12582 ( .A(n9545), .ZN(n11408) );
  OAI21_X1 U12583 ( .B1(n11408), .B2(n11277), .A(n11413), .ZN(n9442) );
  NAND2_X1 U12584 ( .A1(n9442), .A2(n19851), .ZN(n9443) );
  NOR2_X1 U12585 ( .A1(n11841), .A2(n11674), .ZN(n9543) );
  XNOR2_X1 U12586 ( .A(n9691), .B(n9817), .ZN(n10508) );
  XNOR2_X1 U12587 ( .A(n9445), .B(n10508), .ZN(n9450) );
  INV_X1 U12588 ( .A(n9446), .ZN(n9448) );
  XNOR2_X1 U12589 ( .A(n9844), .B(n2307), .ZN(n9447) );
  XNOR2_X1 U12590 ( .A(n9448), .B(n9447), .ZN(n9449) );
  XNOR2_X1 U12591 ( .A(n9450), .B(n9449), .ZN(n11011) );
  XNOR2_X1 U12592 ( .A(n9868), .B(n2280), .ZN(n9457) );
  XNOR2_X1 U12593 ( .A(n9457), .B(n9456), .ZN(n9461) );
  XNOR2_X1 U12594 ( .A(n9458), .B(n9668), .ZN(n10475) );
  XNOR2_X1 U12595 ( .A(n10475), .B(n9459), .ZN(n9460) );
  XNOR2_X1 U12597 ( .A(n10072), .B(n2079), .ZN(n9463) );
  XNOR2_X1 U12598 ( .A(n10481), .B(n9463), .ZN(n9467) );
  XNOR2_X1 U12599 ( .A(n9464), .B(n9465), .ZN(n9466) );
  XNOR2_X1 U12600 ( .A(n9467), .B(n9466), .ZN(n9548) );
  NOR2_X1 U12601 ( .A1(n10953), .A2(n10952), .ZN(n11013) );
  INV_X1 U12602 ( .A(n9812), .ZN(n9468) );
  XNOR2_X1 U12603 ( .A(n9468), .B(n9685), .ZN(n10501) );
  XNOR2_X1 U12604 ( .A(n10501), .B(n9469), .ZN(n9474) );
  INV_X1 U12605 ( .A(n9470), .ZN(n9472) );
  XNOR2_X1 U12606 ( .A(n9862), .B(n17060), .ZN(n9471) );
  XNOR2_X1 U12607 ( .A(n9472), .B(n9471), .ZN(n9473) );
  XNOR2_X1 U12610 ( .A(n9879), .B(n610), .ZN(n9475) );
  XNOR2_X1 U12611 ( .A(n9476), .B(n9475), .ZN(n9478) );
  INV_X1 U12612 ( .A(n9551), .ZN(n11147) );
  XNOR2_X1 U12613 ( .A(n9923), .B(n10114), .ZN(n9479) );
  XNOR2_X1 U12614 ( .A(n9479), .B(n9480), .ZN(n9484) );
  XNOR2_X1 U12615 ( .A(n9922), .B(n10570), .ZN(n9482) );
  INV_X1 U12616 ( .A(n621), .ZN(n18355) );
  XNOR2_X1 U12617 ( .A(n9777), .B(n18355), .ZN(n9481) );
  XNOR2_X1 U12618 ( .A(n9482), .B(n9481), .ZN(n9483) );
  XNOR2_X1 U12619 ( .A(n9484), .B(n9483), .ZN(n11149) );
  INV_X1 U12620 ( .A(n11149), .ZN(n10951) );
  NAND3_X1 U12621 ( .A1(n11016), .A2(n10952), .A3(n10951), .ZN(n9485) );
  NOR2_X1 U12622 ( .A1(n11175), .A2(n9351), .ZN(n10657) );
  INV_X1 U12623 ( .A(n10657), .ZN(n10912) );
  NAND2_X1 U12624 ( .A1(n11174), .A2(n10962), .ZN(n9487) );
  NAND2_X1 U12627 ( .A1(n11175), .A2(n11178), .ZN(n9488) );
  OAI22_X1 U12628 ( .A1(n9488), .A2(n11176), .B1(n11177), .B2(n11174), .ZN(
        n9489) );
  NOR2_X1 U12629 ( .A1(n11161), .A2(n10649), .ZN(n11157) );
  INV_X1 U12630 ( .A(n11157), .ZN(n9495) );
  INV_X1 U12631 ( .A(n11156), .ZN(n9494) );
  NAND2_X1 U12632 ( .A1(n10649), .A2(n11159), .ZN(n9493) );
  NAND3_X1 U12633 ( .A1(n9495), .A2(n9494), .A3(n9493), .ZN(n9497) );
  OAI211_X1 U12634 ( .C1(n11158), .C2(n11160), .A(n11155), .B(n11159), .ZN(
        n9496) );
  INV_X1 U12635 ( .A(n9499), .ZN(n9501) );
  XNOR2_X1 U12636 ( .A(n9500), .B(n10265), .ZN(n10524) );
  XNOR2_X1 U12637 ( .A(n10524), .B(n9501), .ZN(n9505) );
  XNOR2_X1 U12638 ( .A(n9667), .B(n16242), .ZN(n9502) );
  XNOR2_X1 U12639 ( .A(n9503), .B(n9502), .ZN(n9504) );
  INV_X1 U12640 ( .A(n10274), .ZN(n9506) );
  XNOR2_X1 U12641 ( .A(n9879), .B(n9506), .ZN(n10548) );
  XNOR2_X1 U12642 ( .A(n10548), .B(n9507), .ZN(n9511) );
  XNOR2_X1 U12643 ( .A(n9999), .B(n18716), .ZN(n9509) );
  XNOR2_X1 U12644 ( .A(n9509), .B(n9508), .ZN(n9510) );
  NOR2_X1 U12645 ( .A1(n1721), .A2(n20366), .ZN(n9517) );
  XNOR2_X1 U12646 ( .A(n9844), .B(n19786), .ZN(n10535) );
  XNOR2_X1 U12647 ( .A(n10535), .B(n9512), .ZN(n9516) );
  XNOR2_X1 U12648 ( .A(n10249), .B(n2298), .ZN(n9513) );
  XNOR2_X1 U12649 ( .A(n9514), .B(n9513), .ZN(n9515) );
  XNOR2_X1 U12650 ( .A(n9516), .B(n9515), .ZN(n10642) );
  XNOR2_X1 U12651 ( .A(n20176), .B(n1996), .ZN(n9519) );
  XNOR2_X1 U12652 ( .A(n9518), .B(n9519), .ZN(n9522) );
  XNOR2_X1 U12653 ( .A(n10303), .B(n9777), .ZN(n10568) );
  XNOR2_X1 U12654 ( .A(n10568), .B(n9520), .ZN(n9521) );
  XNOR2_X1 U12655 ( .A(n9524), .B(n9523), .ZN(n9525) );
  XNOR2_X1 U12656 ( .A(n9526), .B(n9525), .ZN(n9616) );
  NAND3_X1 U12657 ( .A1(n9527), .A2(n18177), .A3(n9530), .ZN(n9533) );
  INV_X1 U12658 ( .A(n18177), .ZN(n9531) );
  NAND3_X1 U12659 ( .A1(n9529), .A2(n9531), .A3(n9528), .ZN(n9532) );
  XNOR2_X1 U12660 ( .A(n9534), .B(n9983), .ZN(n9536) );
  INV_X1 U12661 ( .A(n9535), .ZN(n10180) );
  XNOR2_X1 U12662 ( .A(n10180), .B(n10320), .ZN(n9711) );
  XNOR2_X1 U12663 ( .A(n9711), .B(n9536), .ZN(n9541) );
  INV_X1 U12664 ( .A(n9538), .ZN(n9539) );
  XNOR2_X1 U12665 ( .A(n10483), .B(n9539), .ZN(n9540) );
  INV_X1 U12666 ( .A(n13042), .ZN(n9544) );
  XNOR2_X1 U12667 ( .A(n9544), .B(n13070), .ZN(n11801) );
  INV_X1 U12669 ( .A(n11000), .ZN(n11005) );
  INV_X1 U12670 ( .A(n11952), .ZN(n11827) );
  INV_X1 U12671 ( .A(n11011), .ZN(n11153) );
  NOR2_X1 U12672 ( .A1(n10953), .A2(n11153), .ZN(n9550) );
  NOR2_X1 U12673 ( .A1(n20470), .A2(n11147), .ZN(n9549) );
  INV_X1 U12674 ( .A(n9548), .ZN(n11009) );
  MUX2_X1 U12675 ( .A(n9550), .B(n9549), .S(n11009), .Z(n9554) );
  NOR2_X1 U12676 ( .A1(n9552), .A2(n11010), .ZN(n9553) );
  NOR2_X1 U12677 ( .A1(n11157), .A2(n9555), .ZN(n9558) );
  NAND2_X1 U12678 ( .A1(n10947), .A2(n10694), .ZN(n11289) );
  INV_X1 U12679 ( .A(n9559), .ZN(n10950) );
  NAND3_X1 U12680 ( .A1(n10995), .A2(n11283), .A3(n11281), .ZN(n9562) );
  INV_X1 U12681 ( .A(n10946), .ZN(n11284) );
  NAND2_X1 U12682 ( .A1(n11284), .A2(n11283), .ZN(n10998) );
  NAND3_X1 U12683 ( .A1(n19817), .A2(n10998), .A3(n9560), .ZN(n9561) );
  XNOR2_X1 U12684 ( .A(n10506), .B(n10186), .ZN(n10533) );
  INV_X1 U12685 ( .A(n9568), .ZN(n9569) );
  XNOR2_X1 U12686 ( .A(n10249), .B(n1857), .ZN(n9571) );
  XNOR2_X1 U12687 ( .A(n9571), .B(n9843), .ZN(n9572) );
  XNOR2_X1 U12688 ( .A(n10533), .B(n9572), .ZN(n9575) );
  XNOR2_X1 U12689 ( .A(n9960), .B(n10445), .ZN(n9573) );
  NAND2_X1 U12693 ( .A1(n9577), .A2(n9576), .ZN(n9581) );
  AOI21_X1 U12694 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9584) );
  XNOR2_X1 U12695 ( .A(n10572), .B(n1911), .ZN(n9585) );
  XNOR2_X1 U12696 ( .A(n9585), .B(n10016), .ZN(n9586) );
  XNOR2_X1 U12697 ( .A(n10567), .B(n10456), .ZN(n10165) );
  XNOR2_X1 U12698 ( .A(n10514), .B(n9587), .ZN(n9588) );
  XNOR2_X1 U12699 ( .A(n10157), .B(n10350), .ZN(n9591) );
  XNOR2_X1 U12700 ( .A(n10498), .B(n9589), .ZN(n9590) );
  XNOR2_X1 U12701 ( .A(n9591), .B(n9590), .ZN(n9595) );
  XNOR2_X1 U12702 ( .A(n9994), .B(n10431), .ZN(n9593) );
  XNOR2_X1 U12703 ( .A(n10436), .B(n17932), .ZN(n9592) );
  XNOR2_X1 U12704 ( .A(n9593), .B(n9592), .ZN(n9594) );
  XNOR2_X1 U12705 ( .A(n9595), .B(n9594), .ZN(n11294) );
  INV_X1 U12706 ( .A(n11406), .ZN(n9612) );
  INV_X1 U12707 ( .A(n10264), .ZN(n9597) );
  XNOR2_X1 U12708 ( .A(n9597), .B(n9667), .ZN(n9598) );
  XNOR2_X1 U12709 ( .A(n9598), .B(n10473), .ZN(n9599) );
  XNOR2_X1 U12710 ( .A(n10179), .B(n9600), .ZN(n9800) );
  INV_X1 U12711 ( .A(n9987), .ZN(n9601) );
  XNOR2_X1 U12712 ( .A(n9601), .B(n10484), .ZN(n9853) );
  XNOR2_X1 U12713 ( .A(n9853), .B(n9800), .ZN(n9604) );
  NOR2_X1 U12714 ( .A1(n11292), .A2(n19506), .ZN(n9610) );
  XNOR2_X1 U12715 ( .A(n9999), .B(n10271), .ZN(n9605) );
  XNOR2_X1 U12716 ( .A(n10358), .B(n2100), .ZN(n9607) );
  XNOR2_X1 U12717 ( .A(n878), .B(n19717), .ZN(n9606) );
  XNOR2_X1 U12718 ( .A(n9607), .B(n9606), .ZN(n9608) );
  INV_X1 U12719 ( .A(n11294), .ZN(n11402) );
  OAI21_X1 U12720 ( .B1(n11403), .B2(n11402), .A(n10980), .ZN(n9609) );
  MUX2_X1 U12722 ( .A(n9613), .B(n981), .S(n11951), .Z(n9622) );
  INV_X1 U12723 ( .A(n10958), .ZN(n9615) );
  NAND2_X1 U12724 ( .A1(n9615), .A2(n9614), .ZN(n9619) );
  NAND2_X1 U12725 ( .A1(n11145), .A2(n11142), .ZN(n9618) );
  INV_X1 U12726 ( .A(n10642), .ZN(n11140) );
  AND3_X1 U12727 ( .A1(n1749), .A2(n11140), .A3(n10701), .ZN(n9617) );
  INV_X1 U12728 ( .A(n11830), .ZN(n11953) );
  OAI21_X1 U12729 ( .B1(n11659), .B2(n11953), .A(n11828), .ZN(n9620) );
  NOR2_X1 U12730 ( .A1(n9620), .A2(n981), .ZN(n9621) );
  INV_X1 U12731 ( .A(n10343), .ZN(n9626) );
  XNOR2_X1 U12732 ( .A(n9626), .B(n9625), .ZN(n9631) );
  INV_X1 U12733 ( .A(n9937), .ZN(n9627) );
  XNOR2_X1 U12734 ( .A(n10265), .B(n9627), .ZN(n9629) );
  XNOR2_X1 U12735 ( .A(n10425), .B(n17804), .ZN(n9628) );
  XNOR2_X1 U12736 ( .A(n9629), .B(n9628), .ZN(n9630) );
  INV_X1 U12738 ( .A(n9632), .ZN(n9634) );
  XNOR2_X1 U12739 ( .A(n10461), .B(n10079), .ZN(n9633) );
  XNOR2_X1 U12740 ( .A(n9634), .B(n9633), .ZN(n9639) );
  XNOR2_X1 U12741 ( .A(n10213), .B(n9635), .ZN(n9637) );
  XNOR2_X1 U12742 ( .A(n10274), .B(n19410), .ZN(n9636) );
  XNOR2_X1 U12743 ( .A(n9637), .B(n9636), .ZN(n9638) );
  XNOR2_X1 U12744 ( .A(n9639), .B(n9638), .ZN(n10685) );
  NOR2_X1 U12745 ( .A1(n20496), .A2(n12101), .ZN(n9660) );
  XNOR2_X1 U12746 ( .A(n10303), .B(n20672), .ZN(n9640) );
  XNOR2_X1 U12747 ( .A(n10304), .B(n9640), .ZN(n9642) );
  XNOR2_X1 U12748 ( .A(n9967), .B(n9922), .ZN(n9641) );
  XNOR2_X1 U12749 ( .A(n9642), .B(n9641), .ZN(n9645) );
  XNOR2_X1 U12750 ( .A(n9644), .B(n10105), .ZN(n10337) );
  XNOR2_X1 U12751 ( .A(n10337), .B(n9645), .ZN(n10683) );
  XNOR2_X1 U12753 ( .A(n20156), .B(n9648), .ZN(n10438) );
  INV_X1 U12754 ( .A(n10438), .ZN(n9649) );
  XNOR2_X1 U12755 ( .A(n10086), .B(n9649), .ZN(n9653) );
  XNOR2_X1 U12756 ( .A(n10281), .B(n2123), .ZN(n9650) );
  XNOR2_X1 U12757 ( .A(n9651), .B(n9650), .ZN(n9652) );
  INV_X1 U12758 ( .A(n10684), .ZN(n10864) );
  INV_X1 U12759 ( .A(n10290), .ZN(n9655) );
  XNOR2_X1 U12760 ( .A(n9947), .B(n2192), .ZN(n9654) );
  XNOR2_X1 U12761 ( .A(n9655), .B(n9654), .ZN(n9658) );
  XNOR2_X1 U12762 ( .A(n9894), .B(n9986), .ZN(n10318) );
  XNOR2_X1 U12763 ( .A(n9656), .B(n10318), .ZN(n9657) );
  XNOR2_X1 U12764 ( .A(n9658), .B(n9657), .ZN(n9666) );
  XNOR2_X1 U12765 ( .A(n10442), .B(n9691), .ZN(n9662) );
  XNOR2_X1 U12766 ( .A(n9662), .B(n9661), .ZN(n9665) );
  XNOR2_X1 U12768 ( .A(n19786), .B(n17993), .ZN(n9663) );
  XNOR2_X1 U12769 ( .A(n929), .B(n9663), .ZN(n9664) );
  XNOR2_X1 U12770 ( .A(n9664), .B(n9665), .ZN(n11380) );
  INV_X1 U12771 ( .A(n11380), .ZN(n11275) );
  NAND2_X1 U12772 ( .A1(n11275), .A2(n11383), .ZN(n12100) );
  INV_X1 U12773 ( .A(n10422), .ZN(n10605) );
  XNOR2_X1 U12774 ( .A(n9869), .B(n10605), .ZN(n10099) );
  XNOR2_X1 U12775 ( .A(n9667), .B(n10421), .ZN(n9975) );
  XNOR2_X1 U12776 ( .A(n10099), .B(n9975), .ZN(n9673) );
  XNOR2_X1 U12777 ( .A(n19853), .B(n9668), .ZN(n10138) );
  INV_X1 U12778 ( .A(n9670), .ZN(n10174) );
  XNOR2_X1 U12779 ( .A(n10174), .B(n642), .ZN(n9671) );
  XNOR2_X1 U12780 ( .A(n10138), .B(n9671), .ZN(n9672) );
  XNOR2_X1 U12781 ( .A(n9673), .B(n9672), .ZN(n11328) );
  XNOR2_X1 U12782 ( .A(n10416), .B(n9674), .ZN(n9678) );
  XNOR2_X1 U12783 ( .A(n10220), .B(n9983), .ZN(n9676) );
  XNOR2_X1 U12784 ( .A(n9462), .B(n2208), .ZN(n9675) );
  XNOR2_X1 U12785 ( .A(n9676), .B(n9675), .ZN(n9677) );
  XNOR2_X1 U12786 ( .A(n9678), .B(n9677), .ZN(n11244) );
  XNOR2_X1 U12787 ( .A(n10077), .B(n10126), .ZN(n9680) );
  INV_X1 U12788 ( .A(n9679), .ZN(n10465) );
  XNOR2_X1 U12789 ( .A(n10465), .B(n9680), .ZN(n9684) );
  XNOR2_X1 U12790 ( .A(n9999), .B(n1057), .ZN(n9682) );
  XNOR2_X1 U12791 ( .A(n928), .B(n2423), .ZN(n9681) );
  XNOR2_X1 U12792 ( .A(n9682), .B(n9681), .ZN(n9683) );
  XNOR2_X2 U12793 ( .A(n9684), .B(n9683), .ZN(n11376) );
  XNOR2_X1 U12794 ( .A(n10350), .B(n9685), .ZN(n10122) );
  INV_X1 U12795 ( .A(n10122), .ZN(n9687) );
  XNOR2_X1 U12796 ( .A(n9994), .B(n18420), .ZN(n9686) );
  XNOR2_X1 U12797 ( .A(n9687), .B(n9686), .ZN(n9690) );
  XNOR2_X1 U12798 ( .A(n10430), .B(n10087), .ZN(n9688) );
  XNOR2_X1 U12799 ( .A(n10433), .B(n9688), .ZN(n9689) );
  MUX2_X1 U12800 ( .A(n11375), .B(n10661), .S(n11329), .Z(n12363) );
  XNOR2_X1 U12801 ( .A(n9692), .B(n9691), .ZN(n10134) );
  XNOR2_X1 U12802 ( .A(n10444), .B(n10134), .ZN(n9696) );
  XNOR2_X1 U12803 ( .A(n10441), .B(n10094), .ZN(n9694) );
  XNOR2_X1 U12804 ( .A(n10249), .B(n18338), .ZN(n9693) );
  XNOR2_X1 U12805 ( .A(n9694), .B(n9693), .ZN(n9695) );
  XNOR2_X1 U12806 ( .A(n9696), .B(n9695), .ZN(n11373) );
  INV_X1 U12807 ( .A(n11373), .ZN(n10856) );
  INV_X1 U12808 ( .A(n11376), .ZN(n11332) );
  XNOR2_X1 U12809 ( .A(n9697), .B(n9922), .ZN(n10118) );
  INV_X1 U12810 ( .A(n10118), .ZN(n9698) );
  XNOR2_X1 U12811 ( .A(n9698), .B(n20176), .ZN(n9708) );
  INV_X1 U12812 ( .A(n9700), .ZN(n9699) );
  NAND2_X1 U12813 ( .A1(n9699), .A2(n2203), .ZN(n9704) );
  INV_X1 U12814 ( .A(n2203), .ZN(n18909) );
  NAND2_X1 U12815 ( .A1(n9703), .A2(n18909), .ZN(n9702) );
  NAND2_X1 U12816 ( .A1(n9700), .A2(n18909), .ZN(n9701) );
  OAI211_X1 U12817 ( .C1(n9704), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9705)
         );
  XNOR2_X1 U12818 ( .A(n9705), .B(n10107), .ZN(n9706) );
  XNOR2_X1 U12819 ( .A(n10454), .B(n9706), .ZN(n9707) );
  NAND2_X1 U12820 ( .A1(n2858), .A2(n11330), .ZN(n9709) );
  MUX2_X1 U12821 ( .A(n10662), .B(n9709), .S(n11244), .Z(n12362) );
  INV_X1 U12822 ( .A(n9710), .ZN(n10031) );
  XNOR2_X1 U12823 ( .A(n10072), .B(n10031), .ZN(n10379) );
  XNOR2_X1 U12824 ( .A(n10379), .B(n9711), .ZN(n9715) );
  XNOR2_X1 U12825 ( .A(n9802), .B(n2263), .ZN(n9712) );
  XNOR2_X1 U12826 ( .A(n9713), .B(n9712), .ZN(n9714) );
  XNOR2_X2 U12827 ( .A(n9715), .B(n9714), .ZN(n11399) );
  INV_X1 U12828 ( .A(n10404), .ZN(n9716) );
  XNOR2_X1 U12829 ( .A(n9716), .B(n10402), .ZN(n10131) );
  XNOR2_X1 U12830 ( .A(n10131), .B(n9717), .ZN(n9721) );
  XNOR2_X1 U12831 ( .A(n10252), .B(n10367), .ZN(n9719) );
  XNOR2_X1 U12832 ( .A(n19785), .B(n484), .ZN(n9718) );
  XNOR2_X1 U12833 ( .A(n9719), .B(n9718), .ZN(n9720) );
  XNOR2_X1 U12834 ( .A(n9721), .B(n9720), .ZN(n11297) );
  XNOR2_X1 U12835 ( .A(n10043), .B(n10557), .ZN(n10396) );
  XNOR2_X1 U12836 ( .A(n10396), .B(n9722), .ZN(n9726) );
  XNOR2_X1 U12837 ( .A(n10236), .B(n1386), .ZN(n9723) );
  XNOR2_X1 U12838 ( .A(n9724), .B(n9723), .ZN(n9725) );
  XNOR2_X1 U12839 ( .A(n9726), .B(n9725), .ZN(n10667) );
  INV_X1 U12840 ( .A(n10667), .ZN(n11394) );
  INV_X1 U12841 ( .A(n9952), .ZN(n9727) );
  XNOR2_X1 U12842 ( .A(n9727), .B(n10551), .ZN(n10125) );
  XNOR2_X1 U12843 ( .A(n10125), .B(n9728), .ZN(n9732) );
  XNOR2_X1 U12844 ( .A(n10359), .B(n917), .ZN(n9730) );
  XNOR2_X1 U12845 ( .A(n10274), .B(n19158), .ZN(n9729) );
  XNOR2_X1 U12846 ( .A(n9730), .B(n9729), .ZN(n9731) );
  NAND2_X1 U12847 ( .A1(n11394), .A2(n11397), .ZN(n9746) );
  XNOR2_X1 U12848 ( .A(n19767), .B(n10339), .ZN(n9734) );
  XNOR2_X1 U12849 ( .A(n9734), .B(n9733), .ZN(n9737) );
  XNOR2_X1 U12850 ( .A(n10037), .B(n10526), .ZN(n10376) );
  XNOR2_X1 U12851 ( .A(n10265), .B(n538), .ZN(n9735) );
  XNOR2_X1 U12852 ( .A(n10376), .B(n9735), .ZN(n9736) );
  XNOR2_X1 U12853 ( .A(n20161), .B(n10052), .ZN(n9739) );
  XNOR2_X1 U12854 ( .A(n9738), .B(n9739), .ZN(n9743) );
  XNOR2_X1 U12855 ( .A(n10388), .B(n10203), .ZN(n9741) );
  XNOR2_X1 U12856 ( .A(n10570), .B(n347), .ZN(n9740) );
  XNOR2_X1 U12857 ( .A(n9741), .B(n9740), .ZN(n9742) );
  XNOR2_X1 U12858 ( .A(n9743), .B(n9742), .ZN(n10986) );
  NAND2_X1 U12859 ( .A1(n10667), .A2(n10986), .ZN(n9744) );
  OAI21_X1 U12860 ( .B1(n11395), .B2(n11399), .A(n9744), .ZN(n10985) );
  NAND2_X1 U12861 ( .A1(n10985), .A2(n11401), .ZN(n9745) );
  INV_X1 U12863 ( .A(n12009), .ZN(n12510) );
  XNOR2_X1 U12864 ( .A(n9748), .B(n620), .ZN(n9749) );
  XNOR2_X1 U12865 ( .A(n20483), .B(n9749), .ZN(n9751) );
  XNOR2_X1 U12866 ( .A(n9750), .B(n9751), .ZN(n9753) );
  XNOR2_X1 U12867 ( .A(n10528), .B(n10262), .ZN(n9752) );
  XNOR2_X1 U12868 ( .A(n10137), .B(n9752), .ZN(n10477) );
  XNOR2_X1 U12869 ( .A(n9753), .B(n10477), .ZN(n11871) );
  XNOR2_X1 U12870 ( .A(n9754), .B(n10482), .ZN(n10540) );
  XNOR2_X1 U12871 ( .A(n9987), .B(n18997), .ZN(n9755) );
  XNOR2_X1 U12872 ( .A(n10540), .B(n9755), .ZN(n9758) );
  XNOR2_X1 U12873 ( .A(n20134), .B(n10028), .ZN(n10287) );
  XNOR2_X1 U12874 ( .A(n9756), .B(n10287), .ZN(n9757) );
  INV_X1 U12876 ( .A(n11303), .ZN(n10862) );
  XNOR2_X1 U12879 ( .A(n9760), .B(n10270), .ZN(n10489) );
  XNOR2_X1 U12881 ( .A(n9761), .B(n9902), .ZN(n9763) );
  XNOR2_X1 U12882 ( .A(n9879), .B(n878), .ZN(n9762) );
  XNOR2_X1 U12883 ( .A(n9763), .B(n9762), .ZN(n9764) );
  XNOR2_X1 U12884 ( .A(n10489), .B(n9764), .ZN(n11389) );
  XNOR2_X1 U12886 ( .A(n10236), .B(n18278), .ZN(n9766) );
  INV_X1 U12887 ( .A(n9908), .ZN(n9765) );
  XNOR2_X1 U12888 ( .A(n9766), .B(n9765), .ZN(n9768) );
  XNOR2_X1 U12889 ( .A(n9862), .B(n10436), .ZN(n9767) );
  XNOR2_X1 U12890 ( .A(n9768), .B(n9767), .ZN(n9770) );
  XNOR2_X1 U12891 ( .A(n10589), .B(n10048), .ZN(n10279) );
  INV_X1 U12892 ( .A(n9769), .ZN(n10561) );
  XNOR2_X1 U12893 ( .A(n10279), .B(n10561), .ZN(n10503) );
  INV_X1 U12895 ( .A(n11866), .ZN(n10990) );
  XNOR2_X1 U12896 ( .A(n9772), .B(n9843), .ZN(n9774) );
  INV_X1 U12897 ( .A(n9819), .ZN(n10401) );
  XNOR2_X1 U12898 ( .A(n10401), .B(n10612), .ZN(n9775) );
  XNOR2_X1 U12899 ( .A(n9775), .B(n19871), .ZN(n10510) );
  NAND2_X1 U12900 ( .A1(n11302), .A2(n19750), .ZN(n10711) );
  INV_X1 U12901 ( .A(n9777), .ZN(n9778) );
  INV_X1 U12902 ( .A(n9779), .ZN(n9785) );
  AOI21_X1 U12904 ( .B1(n19553), .B2(n9782), .A(n9781), .ZN(n9783) );
  OAI21_X1 U12905 ( .B1(n9785), .B2(n19553), .A(n9783), .ZN(n9786) );
  XNOR2_X1 U12906 ( .A(n9786), .B(n10054), .ZN(n10517) );
  XNOR2_X1 U12907 ( .A(n10517), .B(n9860), .ZN(n9790) );
  INV_X1 U12908 ( .A(n10566), .ZN(n10387) );
  INV_X1 U12909 ( .A(n10203), .ZN(n9787) );
  XNOR2_X1 U12910 ( .A(n9926), .B(n573), .ZN(n9788) );
  XNOR2_X1 U12911 ( .A(n9789), .B(n9790), .ZN(n10709) );
  AOI21_X1 U12912 ( .B1(n10711), .B2(n20517), .A(n20601), .ZN(n9791) );
  MUX2_X1 U12913 ( .A(n12008), .B(n12510), .S(n12508), .Z(n9887) );
  XNOR2_X1 U12914 ( .A(n10171), .B(n10472), .ZN(n10525) );
  XNOR2_X1 U12915 ( .A(n10525), .B(n9974), .ZN(n9798) );
  XNOR2_X1 U12918 ( .A(n10229), .B(n18396), .ZN(n9795) );
  XNOR2_X1 U12919 ( .A(n9796), .B(n9795), .ZN(n9797) );
  XNOR2_X1 U12920 ( .A(n10482), .B(n9799), .ZN(n9801) );
  INV_X1 U12921 ( .A(n9800), .ZN(n10541) );
  XNOR2_X1 U12922 ( .A(n10541), .B(n9801), .ZN(n9805) );
  XNOR2_X1 U12923 ( .A(n9854), .B(n9802), .ZN(n10223) );
  XNOR2_X1 U12924 ( .A(n10289), .B(n19102), .ZN(n9803) );
  XNOR2_X1 U12925 ( .A(n9803), .B(n10223), .ZN(n9804) );
  XNOR2_X1 U12926 ( .A(n9805), .B(n9804), .ZN(n10194) );
  INV_X1 U12927 ( .A(n10194), .ZN(n11337) );
  XNOR2_X1 U12928 ( .A(n10203), .B(n9923), .ZN(n9806) );
  XNOR2_X1 U12929 ( .A(n10165), .B(n9806), .ZN(n9810) );
  XNOR2_X1 U12930 ( .A(n10387), .B(n10205), .ZN(n9808) );
  XNOR2_X1 U12931 ( .A(n10572), .B(n457), .ZN(n9807) );
  XNOR2_X1 U12932 ( .A(n9808), .B(n9807), .ZN(n9809) );
  XNOR2_X1 U12933 ( .A(n9809), .B(n9810), .ZN(n10673) );
  XNOR2_X1 U12934 ( .A(n10497), .B(n10157), .ZN(n10559) );
  INV_X1 U12935 ( .A(n9996), .ZN(n9811) );
  XNOR2_X1 U12936 ( .A(n9811), .B(n10559), .ZN(n9816) );
  XNOR2_X1 U12937 ( .A(n9812), .B(n10349), .ZN(n9814) );
  XNOR2_X1 U12938 ( .A(n10236), .B(n18863), .ZN(n9813) );
  XNOR2_X1 U12939 ( .A(n9814), .B(n9813), .ZN(n9815) );
  INV_X1 U12940 ( .A(n9830), .ZN(n11264) );
  XNOR2_X1 U12941 ( .A(n10252), .B(n9817), .ZN(n9818) );
  XNOR2_X1 U12942 ( .A(n10533), .B(n9818), .ZN(n9823) );
  XNOR2_X1 U12943 ( .A(n10248), .B(n18478), .ZN(n9821) );
  INV_X1 U12944 ( .A(n10445), .ZN(n9820) );
  XNOR2_X1 U12945 ( .A(n9819), .B(n9820), .ZN(n10011) );
  XNOR2_X1 U12946 ( .A(n9821), .B(n10011), .ZN(n9822) );
  INV_X1 U12947 ( .A(n11267), .ZN(n11343) );
  XNOR2_X1 U12948 ( .A(n9998), .B(n10549), .ZN(n9829) );
  XNOR2_X1 U12949 ( .A(n9824), .B(n10360), .ZN(n9827) );
  XNOR2_X1 U12950 ( .A(n918), .B(n18208), .ZN(n9826) );
  XNOR2_X1 U12951 ( .A(n9827), .B(n9826), .ZN(n9828) );
  MUX2_X1 U12952 ( .A(n20505), .B(n20476), .S(n19606), .Z(n9840) );
  NAND3_X1 U12953 ( .A1(n9837), .A2(n9836), .A3(n20505), .ZN(n9839) );
  XNOR2_X1 U12954 ( .A(n9842), .B(n9841), .ZN(n10611) );
  XNOR2_X1 U12955 ( .A(n10613), .B(n9843), .ZN(n10010) );
  XNOR2_X1 U12956 ( .A(n10010), .B(n10611), .ZN(n9850) );
  INV_X1 U12957 ( .A(n9844), .ZN(n9845) );
  XNOR2_X1 U12958 ( .A(n9845), .B(n10094), .ZN(n9848) );
  XNOR2_X1 U12959 ( .A(n9846), .B(n19321), .ZN(n9847) );
  XNOR2_X1 U12960 ( .A(n9848), .B(n9847), .ZN(n9849) );
  INV_X1 U12961 ( .A(n11365), .ZN(n10676) );
  INV_X1 U12962 ( .A(n10382), .ZN(n9851) );
  XNOR2_X1 U12963 ( .A(n9851), .B(n10542), .ZN(n9852) );
  XNOR2_X1 U12964 ( .A(n9854), .B(n16424), .ZN(n9855) );
  XNOR2_X1 U12965 ( .A(n10598), .B(n10205), .ZN(n9858) );
  XNOR2_X1 U12966 ( .A(n10107), .B(n2424), .ZN(n9857) );
  XNOR2_X1 U12967 ( .A(n9857), .B(n9858), .ZN(n9859) );
  XNOR2_X1 U12968 ( .A(n10571), .B(n10163), .ZN(n10600) );
  INV_X1 U12969 ( .A(n9883), .ZN(n10852) );
  XNOR2_X1 U12970 ( .A(n10558), .B(n10436), .ZN(n9992) );
  XNOR2_X1 U12971 ( .A(n10498), .B(n9861), .ZN(n10158) );
  XNOR2_X1 U12973 ( .A(n9862), .B(n2087), .ZN(n9864) );
  XNOR2_X1 U12974 ( .A(n10087), .B(n10349), .ZN(n9863) );
  INV_X1 U12976 ( .A(n11234), .ZN(n10851) );
  NOR2_X1 U12977 ( .A1(n10852), .A2(n10851), .ZN(n9874) );
  XNOR2_X1 U12978 ( .A(n10229), .B(Key[60]), .ZN(n9867) );
  XNOR2_X1 U12979 ( .A(n9867), .B(n9868), .ZN(n9871) );
  XNOR2_X1 U12980 ( .A(n9977), .B(n9869), .ZN(n9870) );
  XNOR2_X1 U12981 ( .A(n9871), .B(n9870), .ZN(n9873) );
  XNOR2_X1 U12982 ( .A(n20115), .B(n10173), .ZN(n9872) );
  XNOR2_X1 U12983 ( .A(n9872), .B(n10473), .ZN(n10609) );
  XNOR2_X1 U12984 ( .A(n9873), .B(n10609), .ZN(n10675) );
  BUF_X2 U12985 ( .A(n10675), .Z(n11230) );
  INV_X1 U12986 ( .A(n10490), .ZN(n9876) );
  XNOR2_X1 U12987 ( .A(n9876), .B(n10150), .ZN(n10580) );
  XNOR2_X1 U12988 ( .A(n19945), .B(n10360), .ZN(n9877) );
  INV_X1 U12990 ( .A(n10578), .ZN(n10550) );
  XNOR2_X1 U12991 ( .A(n878), .B(n10550), .ZN(n10004) );
  XNOR2_X1 U12992 ( .A(n9879), .B(n17466), .ZN(n9880) );
  INV_X1 U12994 ( .A(n11231), .ZN(n10854) );
  INV_X1 U12995 ( .A(n12509), .ZN(n11834) );
  NAND2_X1 U12996 ( .A1(n11834), .A2(n12359), .ZN(n9885) );
  XNOR2_X1 U12997 ( .A(n13746), .B(n12696), .ZN(n13444) );
  XNOR2_X1 U12998 ( .A(n11801), .B(n13444), .ZN(n10634) );
  XNOR2_X1 U12999 ( .A(n10171), .B(n10262), .ZN(n9889) );
  XNOR2_X1 U13000 ( .A(n10231), .B(n2216), .ZN(n9888) );
  XNOR2_X1 U13001 ( .A(n9889), .B(n9888), .ZN(n9893) );
  XNOR2_X1 U13002 ( .A(n872), .B(n20484), .ZN(n10373) );
  INV_X1 U13003 ( .A(n10373), .ZN(n9891) );
  XNOR2_X1 U13004 ( .A(n9891), .B(n10475), .ZN(n9892) );
  INV_X1 U13006 ( .A(n9894), .ZN(n10222) );
  XNOR2_X1 U13007 ( .A(n10222), .B(n2420), .ZN(n9895) );
  XNOR2_X1 U13008 ( .A(n20228), .B(n9895), .ZN(n9900) );
  XNOR2_X1 U13009 ( .A(n20134), .B(n10320), .ZN(n10381) );
  XNOR2_X1 U13010 ( .A(n19839), .B(n10028), .ZN(n9898) );
  XNOR2_X1 U13011 ( .A(n10381), .B(n9898), .ZN(n9899) );
  XNOR2_X1 U13012 ( .A(n9900), .B(n9899), .ZN(n9919) );
  INV_X1 U13013 ( .A(n10359), .ZN(n9901) );
  XNOR2_X1 U13014 ( .A(n9901), .B(n9902), .ZN(n10410) );
  XNOR2_X1 U13015 ( .A(n19829), .B(n10410), .ZN(n9907) );
  XNOR2_X1 U13016 ( .A(n10151), .B(n10270), .ZN(n9905) );
  XNOR2_X1 U13017 ( .A(n10213), .B(n18006), .ZN(n9904) );
  XNOR2_X1 U13018 ( .A(n9905), .B(n9904), .ZN(n9906) );
  XNOR2_X1 U13019 ( .A(n10395), .B(n10501), .ZN(n9912) );
  XNOR2_X1 U13020 ( .A(n19990), .B(n645), .ZN(n9909) );
  XNOR2_X1 U13021 ( .A(n9910), .B(n9909), .ZN(n9911) );
  XNOR2_X1 U13022 ( .A(n9912), .B(n9911), .ZN(n11216) );
  XNOR2_X1 U13023 ( .A(n10186), .B(n19871), .ZN(n9914) );
  XNOR2_X1 U13024 ( .A(n9914), .B(n10508), .ZN(n9918) );
  XNOR2_X1 U13025 ( .A(n10298), .B(n10367), .ZN(n10403) );
  INV_X1 U13026 ( .A(n10403), .ZN(n9916) );
  XNOR2_X1 U13027 ( .A(n10247), .B(n18090), .ZN(n9915) );
  XNOR2_X1 U13028 ( .A(n9916), .B(n9915), .ZN(n9917) );
  XNOR2_X1 U13029 ( .A(n9918), .B(n9917), .ZN(n11475) );
  NAND2_X1 U13030 ( .A1(n9920), .A2(n11475), .ZN(n9921) );
  XNOR2_X1 U13031 ( .A(n10567), .B(n10204), .ZN(n9925) );
  XNOR2_X1 U13032 ( .A(n9923), .B(n9922), .ZN(n10515) );
  INV_X1 U13033 ( .A(n10515), .ZN(n9924) );
  XNOR2_X1 U13034 ( .A(n9925), .B(n9924), .ZN(n9929) );
  XNOR2_X1 U13035 ( .A(n9926), .B(n10332), .ZN(n10391) );
  XNOR2_X1 U13036 ( .A(n10054), .B(n2417), .ZN(n9927) );
  XNOR2_X1 U13037 ( .A(n10391), .B(n9927), .ZN(n9928) );
  NAND2_X1 U13038 ( .A1(n9930), .A2(n11079), .ZN(n12498) );
  INV_X1 U13039 ( .A(n10755), .ZN(n11522) );
  OAI21_X1 U13040 ( .B1(n11528), .B2(n11530), .A(n19999), .ZN(n9931) );
  XNOR2_X1 U13041 ( .A(n10422), .B(n9935), .ZN(n9936) );
  XNOR2_X1 U13042 ( .A(n9936), .B(n10342), .ZN(n9940) );
  XNOR2_X1 U13043 ( .A(n9937), .B(n9978), .ZN(n9938) );
  XNOR2_X1 U13044 ( .A(n10473), .B(n9938), .ZN(n9939) );
  XNOR2_X1 U13045 ( .A(n10043), .B(n19018), .ZN(n9942) );
  INV_X1 U13046 ( .A(n9991), .ZN(n9941) );
  XNOR2_X1 U13047 ( .A(n9942), .B(n9941), .ZN(n9943) );
  XNOR2_X1 U13048 ( .A(n10088), .B(n10498), .ZN(n10587) );
  XNOR2_X1 U13049 ( .A(n9943), .B(n10587), .ZN(n9945) );
  XNOR2_X1 U13050 ( .A(n9945), .B(n9944), .ZN(n10883) );
  INV_X1 U13051 ( .A(n10484), .ZN(n9946) );
  XNOR2_X1 U13052 ( .A(n10031), .B(n9986), .ZN(n9949) );
  XNOR2_X1 U13053 ( .A(n9947), .B(n17089), .ZN(n9948) );
  XNOR2_X1 U13054 ( .A(n9949), .B(n9948), .ZN(n9950) );
  XNOR2_X1 U13055 ( .A(n9952), .B(n10579), .ZN(n9955) );
  XNOR2_X1 U13056 ( .A(n19717), .B(n17535), .ZN(n9953) );
  XNOR2_X1 U13057 ( .A(n9953), .B(n10079), .ZN(n9954) );
  XNOR2_X1 U13058 ( .A(n9954), .B(n9955), .ZN(n9956) );
  XNOR2_X1 U13059 ( .A(n9957), .B(n20211), .ZN(n9959) );
  XNOR2_X1 U13060 ( .A(n10008), .B(n2233), .ZN(n9958) );
  XNOR2_X1 U13061 ( .A(n9958), .B(n9959), .ZN(n9962) );
  XNOR2_X1 U13062 ( .A(n9960), .B(n10404), .ZN(n9961) );
  XNOR2_X1 U13063 ( .A(n9962), .B(n9961), .ZN(n9964) );
  INV_X1 U13064 ( .A(n10371), .ZN(n9963) );
  NAND2_X1 U13065 ( .A1(n11182), .A2(n10882), .ZN(n9972) );
  XNOR2_X1 U13066 ( .A(n10514), .B(n10105), .ZN(n9966) );
  XNOR2_X1 U13067 ( .A(n10594), .B(n10388), .ZN(n9965) );
  XNOR2_X1 U13068 ( .A(n9965), .B(n9966), .ZN(n9970) );
  XNOR2_X1 U13069 ( .A(n9967), .B(n2305), .ZN(n9968) );
  XNOR2_X1 U13070 ( .A(n10334), .B(n9968), .ZN(n9969) );
  NAND2_X1 U13071 ( .A1(n11566), .A2(n11466), .ZN(n9971) );
  MUX2_X1 U13072 ( .A(n9972), .B(n9971), .S(n11568), .Z(n9973) );
  INV_X1 U13073 ( .A(n9974), .ZN(n9976) );
  XNOR2_X1 U13074 ( .A(n9976), .B(n9975), .ZN(n9982) );
  XNOR2_X1 U13075 ( .A(n9977), .B(n20115), .ZN(n9980) );
  XNOR2_X1 U13076 ( .A(n9978), .B(n2306), .ZN(n9979) );
  XNOR2_X1 U13077 ( .A(n9979), .B(n9980), .ZN(n9981) );
  XNOR2_X1 U13078 ( .A(n10542), .B(n9983), .ZN(n10618) );
  INV_X1 U13079 ( .A(n9984), .ZN(n9985) );
  XNOR2_X1 U13080 ( .A(n10618), .B(n9985), .ZN(n9990) );
  XNOR2_X1 U13081 ( .A(n10219), .B(n9986), .ZN(n9989) );
  XNOR2_X1 U13082 ( .A(n9987), .B(n16030), .ZN(n9988) );
  NAND2_X1 U13083 ( .A1(n11515), .A2(n10742), .ZN(n11575) );
  XNOR2_X1 U13084 ( .A(n10240), .B(n9991), .ZN(n9993) );
  XNOR2_X1 U13085 ( .A(n9992), .B(n9993), .ZN(n9997) );
  XNOR2_X1 U13086 ( .A(n9994), .B(n19205), .ZN(n9995) );
  INV_X1 U13087 ( .A(n9998), .ZN(n10001) );
  XNOR2_X1 U13088 ( .A(n9999), .B(n10079), .ZN(n10000) );
  XNOR2_X1 U13089 ( .A(n10001), .B(n10000), .ZN(n10006) );
  INV_X1 U13090 ( .A(n10002), .ZN(n10214) );
  XNOR2_X1 U13091 ( .A(n10214), .B(n2455), .ZN(n10003) );
  XNOR2_X1 U13092 ( .A(n10004), .B(n10003), .ZN(n10005) );
  XNOR2_X1 U13094 ( .A(n10254), .B(n10008), .ZN(n10009) );
  XNOR2_X1 U13095 ( .A(n10010), .B(n10009), .ZN(n10015) );
  INV_X1 U13096 ( .A(n10011), .ZN(n10013) );
  XNOR2_X1 U13097 ( .A(n10249), .B(n18726), .ZN(n10012) );
  XNOR2_X1 U13098 ( .A(n10013), .B(n10012), .ZN(n10014) );
  XNOR2_X1 U13101 ( .A(n10016), .B(n20176), .ZN(n10018) );
  XNOR2_X1 U13102 ( .A(n10018), .B(n10017), .ZN(n10022) );
  XNOR2_X1 U13103 ( .A(n10105), .B(n19806), .ZN(n10020) );
  XNOR2_X1 U13104 ( .A(n10571), .B(n1148), .ZN(n10019) );
  XNOR2_X1 U13105 ( .A(n10020), .B(n10019), .ZN(n10021) );
  XNOR2_X1 U13106 ( .A(n10022), .B(n10021), .ZN(n11510) );
  NOR2_X1 U13107 ( .A1(n11510), .A2(n11514), .ZN(n10740) );
  INV_X1 U13108 ( .A(n12498), .ZN(n12497) );
  XNOR2_X1 U13109 ( .A(n10404), .B(n19457), .ZN(n10024) );
  XNOR2_X1 U13110 ( .A(n10406), .B(n10024), .ZN(n10025) );
  XNOR2_X1 U13111 ( .A(n10026), .B(n10442), .ZN(n10370) );
  XNOR2_X1 U13112 ( .A(n10028), .B(n10382), .ZN(n10029) );
  XNOR2_X1 U13113 ( .A(n10220), .B(n10030), .ZN(n10033) );
  XNOR2_X1 U13114 ( .A(n10031), .B(n18308), .ZN(n10032) );
  XNOR2_X1 U13115 ( .A(n10033), .B(n10032), .ZN(n10034) );
  XNOR2_X1 U13116 ( .A(n10035), .B(n10034), .ZN(n10060) );
  INV_X1 U13117 ( .A(n10060), .ZN(n11482) );
  INV_X1 U13118 ( .A(n10036), .ZN(n10374) );
  XNOR2_X1 U13119 ( .A(n10037), .B(n10262), .ZN(n10038) );
  XNOR2_X1 U13120 ( .A(n10374), .B(n10038), .ZN(n10042) );
  XNOR2_X1 U13121 ( .A(n10174), .B(n456), .ZN(n10040) );
  XNOR2_X1 U13122 ( .A(n10340), .B(n10040), .ZN(n10041) );
  INV_X1 U13123 ( .A(n10043), .ZN(n10044) );
  XNOR2_X1 U13124 ( .A(n10044), .B(n10430), .ZN(n10047) );
  XNOR2_X1 U13125 ( .A(n10347), .B(n10047), .ZN(n10051) );
  XNOR2_X1 U13126 ( .A(n19990), .B(n17989), .ZN(n10049) );
  XNOR2_X1 U13127 ( .A(n10397), .B(n10049), .ZN(n10050) );
  XNOR2_X1 U13128 ( .A(n10051), .B(n10050), .ZN(n10745) );
  XNOR2_X1 U13129 ( .A(n10052), .B(n10388), .ZN(n10115) );
  INV_X1 U13130 ( .A(n10392), .ZN(n10053) );
  XNOR2_X1 U13131 ( .A(n10115), .B(n10053), .ZN(n10058) );
  XNOR2_X1 U13132 ( .A(n10114), .B(n10166), .ZN(n10458) );
  INV_X1 U13133 ( .A(n10458), .ZN(n10056) );
  XNOR2_X1 U13134 ( .A(n10054), .B(n632), .ZN(n10055) );
  XNOR2_X1 U13135 ( .A(n10056), .B(n10055), .ZN(n10057) );
  XNOR2_X1 U13136 ( .A(n10058), .B(n10057), .ZN(n10896) );
  NAND2_X1 U13137 ( .A1(n19897), .A2(n11480), .ZN(n10748) );
  NAND2_X1 U13138 ( .A1(n11073), .A2(n10748), .ZN(n10066) );
  INV_X1 U13139 ( .A(n10745), .ZN(n11481) );
  XNOR2_X1 U13140 ( .A(n10409), .B(n10356), .ZN(n10065) );
  XNOR2_X1 U13141 ( .A(n1057), .B(n10270), .ZN(n10063) );
  XNOR2_X1 U13142 ( .A(n9952), .B(n17787), .ZN(n10062) );
  XNOR2_X1 U13143 ( .A(n10063), .B(n10062), .ZN(n10064) );
  NAND2_X1 U13144 ( .A1(n11481), .A2(n10897), .ZN(n11479) );
  NAND2_X1 U13145 ( .A1(n10066), .A2(n11479), .ZN(n10067) );
  INV_X1 U13146 ( .A(n10761), .ZN(n10889) );
  INV_X1 U13147 ( .A(n11546), .ZN(n11547) );
  NAND2_X1 U13148 ( .A1(n11546), .A2(n11550), .ZN(n10069) );
  NAND3_X1 U13149 ( .A1(n1859), .A2(n12005), .A3(n12502), .ZN(n10070) );
  XNOR2_X1 U13150 ( .A(n19818), .B(n18284), .ZN(n10074) );
  XNOR2_X1 U13151 ( .A(n10072), .B(n10382), .ZN(n10073) );
  XNOR2_X1 U13152 ( .A(n10074), .B(n10073), .ZN(n10076) );
  XNOR2_X1 U13153 ( .A(n10318), .B(n10417), .ZN(n10075) );
  INV_X1 U13154 ( .A(n10112), .ZN(n11125) );
  INV_X1 U13155 ( .A(n19945), .ZN(n10078) );
  XNOR2_X1 U13156 ( .A(n10078), .B(n10579), .ZN(n10081) );
  INV_X1 U13157 ( .A(n10213), .ZN(n10080) );
  XNOR2_X1 U13158 ( .A(n10080), .B(n10079), .ZN(n10357) );
  XNOR2_X1 U13159 ( .A(n10357), .B(n10081), .ZN(n10084) );
  XNOR2_X1 U13160 ( .A(n10551), .B(n17170), .ZN(n10082) );
  XNOR2_X1 U13161 ( .A(n10462), .B(n10082), .ZN(n10083) );
  XNOR2_X1 U13162 ( .A(n10557), .B(n10087), .ZN(n10090) );
  XNOR2_X1 U13163 ( .A(n10088), .B(n18011), .ZN(n10089) );
  XNOR2_X1 U13164 ( .A(n10090), .B(n10089), .ZN(n10091) );
  MUX2_X1 U13165 ( .A(n11125), .B(n10814), .S(n1317), .Z(n10104) );
  XNOR2_X1 U13166 ( .A(n20210), .B(n1904), .ZN(n10093) );
  INV_X1 U13167 ( .A(n929), .ZN(n10092) );
  XNOR2_X1 U13168 ( .A(n10093), .B(n10092), .ZN(n10097) );
  XNOR2_X1 U13169 ( .A(n10094), .B(n10402), .ZN(n10095) );
  XNOR2_X1 U13170 ( .A(n10447), .B(n10095), .ZN(n10096) );
  INV_X1 U13171 ( .A(n11358), .ZN(n10103) );
  XNOR2_X1 U13173 ( .A(n20456), .B(n10099), .ZN(n10102) );
  XNOR2_X1 U13174 ( .A(n10526), .B(n649), .ZN(n10100) );
  XNOR2_X1 U13175 ( .A(n10343), .B(n10100), .ZN(n10101) );
  XNOR2_X1 U13176 ( .A(n10453), .B(n10106), .ZN(n10111) );
  XNOR2_X1 U13177 ( .A(n10204), .B(n10570), .ZN(n10109) );
  XNOR2_X1 U13178 ( .A(n10107), .B(n1869), .ZN(n10108) );
  XNOR2_X1 U13179 ( .A(n10109), .B(n10108), .ZN(n10110) );
  XNOR2_X1 U13180 ( .A(n10111), .B(n10110), .ZN(n11356) );
  INV_X1 U13181 ( .A(n11356), .ZN(n11127) );
  NAND2_X1 U13182 ( .A1(n11127), .A2(n10813), .ZN(n10113) );
  XNOR2_X1 U13183 ( .A(n10595), .B(n10114), .ZN(n10116) );
  XNOR2_X1 U13184 ( .A(n10116), .B(n10115), .ZN(n10120) );
  XNOR2_X1 U13185 ( .A(n10570), .B(n18768), .ZN(n10117) );
  XNOR2_X1 U13186 ( .A(n10118), .B(n10117), .ZN(n10119) );
  XNOR2_X1 U13187 ( .A(n10120), .B(n10119), .ZN(n11238) );
  INV_X1 U13188 ( .A(n11238), .ZN(n11355) );
  XNOR2_X1 U13189 ( .A(n10589), .B(n19436), .ZN(n10121) );
  XNOR2_X1 U13190 ( .A(n10396), .B(n10121), .ZN(n10124) );
  XNOR2_X1 U13191 ( .A(n10347), .B(n10122), .ZN(n10123) );
  XNOR2_X1 U13192 ( .A(n10123), .B(n10124), .ZN(n10779) );
  INV_X1 U13193 ( .A(n10779), .ZN(n11239) );
  XNOR2_X1 U13194 ( .A(n10126), .B(n10358), .ZN(n10128) );
  XNOR2_X1 U13195 ( .A(n10582), .B(n2413), .ZN(n10127) );
  XNOR2_X1 U13196 ( .A(n10128), .B(n10127), .ZN(n10129) );
  XNOR2_X1 U13197 ( .A(n10130), .B(n10129), .ZN(n11240) );
  INV_X1 U13198 ( .A(n10131), .ZN(n10133) );
  XNOR2_X1 U13199 ( .A(n10612), .B(n18988), .ZN(n10132) );
  XNOR2_X1 U13200 ( .A(n10133), .B(n10132), .ZN(n10136) );
  XNOR2_X1 U13201 ( .A(n10134), .B(n10370), .ZN(n10135) );
  INV_X1 U13202 ( .A(n11349), .ZN(n11055) );
  INV_X1 U13203 ( .A(n10604), .ZN(n10137) );
  XNOR2_X1 U13204 ( .A(n10137), .B(n2108), .ZN(n10139) );
  XNOR2_X1 U13205 ( .A(n10139), .B(n10138), .ZN(n10141) );
  XNOR2_X1 U13206 ( .A(n10376), .B(n10340), .ZN(n10140) );
  XNOR2_X1 U13207 ( .A(n10140), .B(n10141), .ZN(n11347) );
  INV_X1 U13208 ( .A(n11347), .ZN(n11350) );
  NAND2_X1 U13209 ( .A1(n11347), .A2(n10798), .ZN(n10142) );
  NAND2_X1 U13210 ( .A1(n11060), .A2(n10142), .ZN(n10148) );
  XNOR2_X1 U13211 ( .A(n10379), .B(n10319), .ZN(n10147) );
  XNOR2_X1 U13212 ( .A(n10286), .B(n9462), .ZN(n10145) );
  XNOR2_X1 U13213 ( .A(n10143), .B(n18439), .ZN(n10144) );
  XNOR2_X1 U13214 ( .A(n10145), .B(n10144), .ZN(n10146) );
  INV_X1 U13215 ( .A(n11057), .ZN(n11348) );
  MUX2_X2 U13216 ( .A(n10149), .B(n10148), .S(n11348), .Z(n12334) );
  XNOR2_X1 U13217 ( .A(n10151), .B(n10150), .ZN(n10153) );
  XNOR2_X1 U13218 ( .A(n19718), .B(n2082), .ZN(n10152) );
  XNOR2_X1 U13219 ( .A(n10153), .B(n10152), .ZN(n10156) );
  XNOR2_X1 U13220 ( .A(n1057), .B(n10271), .ZN(n10464) );
  XNOR2_X1 U13221 ( .A(n10548), .B(n10464), .ZN(n10155) );
  XNOR2_X1 U13222 ( .A(n260), .B(n10430), .ZN(n10159) );
  XNOR2_X1 U13223 ( .A(n10158), .B(n10159), .ZN(n10162) );
  XNOR2_X1 U13224 ( .A(n10431), .B(n19052), .ZN(n10160) );
  XNOR2_X1 U13225 ( .A(n10563), .B(n10160), .ZN(n10161) );
  INV_X1 U13226 ( .A(n11428), .ZN(n11425) );
  XNOR2_X1 U13227 ( .A(n10514), .B(n10163), .ZN(n10164) );
  XNOR2_X1 U13228 ( .A(n10165), .B(n10164), .ZN(n10170) );
  INV_X1 U13229 ( .A(n10568), .ZN(n10168) );
  XNOR2_X1 U13230 ( .A(n10166), .B(n2035), .ZN(n10167) );
  XNOR2_X1 U13231 ( .A(n10168), .B(n10167), .ZN(n10169) );
  AOI21_X1 U13232 ( .B1(n11105), .B2(n11425), .A(n11106), .ZN(n10193) );
  XNOR2_X1 U13233 ( .A(n10473), .B(n10171), .ZN(n10172) );
  XNOR2_X1 U13234 ( .A(n10524), .B(n10172), .ZN(n10177) );
  XNOR2_X1 U13235 ( .A(n10173), .B(n2369), .ZN(n10175) );
  XNOR2_X1 U13236 ( .A(n10264), .B(n10174), .ZN(n10427) );
  XNOR2_X1 U13237 ( .A(n10427), .B(n10175), .ZN(n10176) );
  XNOR2_X1 U13238 ( .A(n10177), .B(n10176), .ZN(n11104) );
  INV_X1 U13239 ( .A(n11104), .ZN(n11427) );
  XNOR2_X1 U13240 ( .A(n10289), .B(n10220), .ZN(n10415) );
  XNOR2_X1 U13241 ( .A(n10484), .B(n2445), .ZN(n10178) );
  XNOR2_X1 U13242 ( .A(n10415), .B(n10178), .ZN(n10184) );
  XNOR2_X1 U13243 ( .A(n19839), .B(n10180), .ZN(n10181) );
  XNOR2_X1 U13244 ( .A(n10182), .B(n10181), .ZN(n10183) );
  XNOR2_X1 U13245 ( .A(n10185), .B(n10186), .ZN(n10187) );
  XNOR2_X1 U13246 ( .A(n10187), .B(n10611), .ZN(n10190) );
  XNOR2_X1 U13247 ( .A(n10445), .B(n18203), .ZN(n10188) );
  XNOR2_X1 U13248 ( .A(n10535), .B(n10188), .ZN(n10189) );
  INV_X1 U13249 ( .A(n11106), .ZN(n11424) );
  NAND3_X1 U13250 ( .A1(n11425), .A2(n11430), .A3(n11424), .ZN(n10191) );
  NAND2_X1 U13251 ( .A1(n12334), .A2(n11990), .ZN(n12333) );
  OAI21_X1 U13252 ( .B1(n12338), .B2(n12334), .A(n12333), .ZN(n10317) );
  AOI21_X1 U13254 ( .B1(n11337), .B2(n11263), .A(n3669), .ZN(n10198) );
  NOR2_X1 U13255 ( .A1(n11267), .A2(n11265), .ZN(n10797) );
  NOR2_X1 U13256 ( .A1(n11339), .A2(n9830), .ZN(n10196) );
  INV_X1 U13257 ( .A(n11263), .ZN(n10195) );
  OAI21_X1 U13258 ( .B1(n10797), .B2(n10196), .A(n10195), .ZN(n10197) );
  INV_X1 U13259 ( .A(n11992), .ZN(n12337) );
  XNOR2_X1 U13260 ( .A(n19806), .B(n10200), .ZN(n10202) );
  XNOR2_X1 U13261 ( .A(n10201), .B(n10202), .ZN(n10209) );
  XNOR2_X1 U13262 ( .A(n10203), .B(n10204), .ZN(n10207) );
  XNOR2_X1 U13263 ( .A(n10205), .B(n20064), .ZN(n10206) );
  XNOR2_X1 U13264 ( .A(n10207), .B(n10206), .ZN(n10208) );
  XNOR2_X1 U13265 ( .A(n10209), .B(n10208), .ZN(n11460) );
  INV_X1 U13266 ( .A(n11460), .ZN(n11048) );
  XNOR2_X1 U13270 ( .A(n10213), .B(n10360), .ZN(n10216) );
  XNOR2_X1 U13271 ( .A(n10214), .B(n2055), .ZN(n10215) );
  XNOR2_X1 U13272 ( .A(n10216), .B(n10215), .ZN(n10217) );
  XNOR2_X1 U13274 ( .A(n10219), .B(n10220), .ZN(n10221) );
  XNOR2_X1 U13275 ( .A(n10618), .B(n10221), .ZN(n10227) );
  XNOR2_X1 U13276 ( .A(n10222), .B(n2446), .ZN(n10225) );
  INV_X1 U13277 ( .A(n10223), .ZN(n10224) );
  XNOR2_X1 U13278 ( .A(n10225), .B(n10224), .ZN(n10226) );
  XNOR2_X1 U13279 ( .A(n10226), .B(n10227), .ZN(n10259) );
  XNOR2_X1 U13280 ( .A(n10229), .B(n10421), .ZN(n10230) );
  XNOR2_X1 U13281 ( .A(n10603), .B(n10230), .ZN(n10235) );
  XNOR2_X1 U13282 ( .A(n10231), .B(n106), .ZN(n10232) );
  XNOR2_X1 U13283 ( .A(n10233), .B(n10232), .ZN(n10234) );
  XNOR2_X1 U13284 ( .A(n10235), .B(n10234), .ZN(n10808) );
  XNOR2_X1 U13285 ( .A(n10237), .B(n10236), .ZN(n10591) );
  INV_X1 U13286 ( .A(n10591), .ZN(n10239) );
  XNOR2_X1 U13287 ( .A(n10239), .B(n10238), .ZN(n10244) );
  XNOR2_X1 U13288 ( .A(n10240), .B(n10349), .ZN(n10241) );
  XNOR2_X1 U13289 ( .A(n10242), .B(n10241), .ZN(n10243) );
  INV_X1 U13290 ( .A(n11120), .ZN(n11881) );
  NAND2_X1 U13291 ( .A1(n11881), .A2(n11460), .ZN(n10245) );
  NAND3_X1 U13292 ( .A1(n10246), .A2(n10788), .A3(n10245), .ZN(n10260) );
  XNOR2_X1 U13293 ( .A(n10249), .B(n15479), .ZN(n10250) );
  XNOR2_X1 U13294 ( .A(n10251), .B(n10250), .ZN(n10256) );
  INV_X1 U13295 ( .A(n10252), .ZN(n10253) );
  XNOR2_X1 U13296 ( .A(n10254), .B(n10253), .ZN(n10255) );
  XNOR2_X1 U13297 ( .A(n10256), .B(n10255), .ZN(n10258) );
  XNOR2_X1 U13298 ( .A(n10258), .B(n10257), .ZN(n11884) );
  NAND2_X1 U13299 ( .A1(n10786), .A2(n10259), .ZN(n11050) );
  INV_X1 U13300 ( .A(n11884), .ZN(n11459) );
  INV_X1 U13301 ( .A(n12339), .ZN(n11974) );
  INV_X1 U13302 ( .A(n12338), .ZN(n10314) );
  XNOR2_X1 U13303 ( .A(n10261), .B(n10262), .ZN(n10263) );
  XNOR2_X1 U13304 ( .A(n10373), .B(n10263), .ZN(n10269) );
  XNOR2_X1 U13305 ( .A(n10604), .B(n10264), .ZN(n10267) );
  XNOR2_X1 U13306 ( .A(n10265), .B(n2122), .ZN(n10266) );
  XNOR2_X1 U13307 ( .A(n10267), .B(n10266), .ZN(n10268) );
  INV_X1 U13308 ( .A(n190), .ZN(n11254) );
  XNOR2_X1 U13309 ( .A(n10271), .B(n10270), .ZN(n10272) );
  XNOR2_X1 U13310 ( .A(n10410), .B(n10272), .ZN(n10278) );
  XNOR2_X1 U13311 ( .A(n10273), .B(n10582), .ZN(n10276) );
  XNOR2_X1 U13312 ( .A(n10274), .B(n2296), .ZN(n10275) );
  XNOR2_X1 U13313 ( .A(n10276), .B(n10275), .ZN(n10277) );
  XNOR2_X1 U13314 ( .A(n10395), .B(n10279), .ZN(n10285) );
  XNOR2_X1 U13315 ( .A(n10280), .B(n10431), .ZN(n10283) );
  XNOR2_X1 U13316 ( .A(n10281), .B(n2410), .ZN(n10282) );
  XNOR2_X1 U13317 ( .A(n10283), .B(n10282), .ZN(n10284) );
  XNOR2_X1 U13318 ( .A(n10285), .B(n10284), .ZN(n11321) );
  XNOR2_X1 U13319 ( .A(n10286), .B(n10320), .ZN(n10288) );
  XNOR2_X1 U13320 ( .A(n10287), .B(n10288), .ZN(n10293) );
  XNOR2_X1 U13321 ( .A(n10289), .B(n2395), .ZN(n10291) );
  XNOR2_X1 U13322 ( .A(n10290), .B(n10291), .ZN(n10292) );
  INV_X1 U13324 ( .A(n11257), .ZN(n11327) );
  INV_X1 U13325 ( .A(n2284), .ZN(n18664) );
  XNOR2_X1 U13326 ( .A(n19785), .B(n18664), .ZN(n10295) );
  XNOR2_X1 U13327 ( .A(n10296), .B(n10367), .ZN(n10297) );
  XNOR2_X1 U13328 ( .A(n10298), .B(n10445), .ZN(n10300) );
  XNOR2_X1 U13329 ( .A(n10300), .B(n19871), .ZN(n10301) );
  XNOR2_X1 U13330 ( .A(n10302), .B(n10301), .ZN(n11256) );
  INV_X1 U13331 ( .A(n11256), .ZN(n11322) );
  XNOR2_X1 U13332 ( .A(n10517), .B(n10391), .ZN(n10308) );
  XNOR2_X1 U13333 ( .A(n10303), .B(n2337), .ZN(n10306) );
  XNOR2_X1 U13334 ( .A(n10304), .B(n10456), .ZN(n10305) );
  XNOR2_X1 U13335 ( .A(n10306), .B(n10305), .ZN(n10307) );
  OAI21_X1 U13336 ( .B1(n10310), .B2(n11322), .A(n10309), .ZN(n10311) );
  NOR2_X1 U13337 ( .A1(n11992), .A2(n12335), .ZN(n10313) );
  XNOR2_X1 U13338 ( .A(n13588), .B(n13352), .ZN(n13289) );
  INV_X1 U13339 ( .A(n13289), .ZN(n10632) );
  XNOR2_X1 U13340 ( .A(n10318), .B(n10319), .ZN(n10324) );
  XNOR2_X1 U13341 ( .A(n10320), .B(n2381), .ZN(n10322) );
  XNOR2_X1 U13342 ( .A(n10321), .B(n10322), .ZN(n10323) );
  INV_X1 U13344 ( .A(n10328), .ZN(n10326) );
  INV_X1 U13345 ( .A(n18304), .ZN(n10325) );
  OAI21_X1 U13346 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10331) );
  NAND3_X1 U13347 ( .A1(n10329), .A2(n18304), .A3(n10328), .ZN(n10330) );
  NAND2_X1 U13348 ( .A1(n10331), .A2(n10330), .ZN(n10333) );
  XNOR2_X1 U13349 ( .A(n10333), .B(n20161), .ZN(n10336) );
  INV_X1 U13350 ( .A(n10334), .ZN(n10335) );
  XNOR2_X1 U13351 ( .A(n10336), .B(n10335), .ZN(n10338) );
  XNOR2_X1 U13352 ( .A(n10339), .B(n19216), .ZN(n10341) );
  XNOR2_X1 U13353 ( .A(n10341), .B(n10340), .ZN(n10345) );
  XNOR2_X1 U13354 ( .A(n10343), .B(n10342), .ZN(n10344) );
  XNOR2_X1 U13355 ( .A(n10345), .B(n10344), .ZN(n11087) );
  NAND2_X1 U13356 ( .A1(n11455), .A2(n11454), .ZN(n10346) );
  OAI21_X1 U13357 ( .B1(n11455), .B2(n1812), .A(n10346), .ZN(n10366) );
  XNOR2_X1 U13358 ( .A(n10348), .B(n10347), .ZN(n10355) );
  XNOR2_X1 U13359 ( .A(n10349), .B(n2392), .ZN(n10353) );
  XNOR2_X1 U13360 ( .A(n10351), .B(n10350), .ZN(n10352) );
  XNOR2_X1 U13361 ( .A(n10353), .B(n10352), .ZN(n10354) );
  NOR2_X1 U13362 ( .A1(n11452), .A2(n11455), .ZN(n10365) );
  XNOR2_X1 U13363 ( .A(n10357), .B(n10356), .ZN(n10364) );
  XNOR2_X1 U13364 ( .A(n928), .B(n18170), .ZN(n10362) );
  XNOR2_X1 U13365 ( .A(n10359), .B(n10360), .ZN(n10361) );
  XNOR2_X1 U13366 ( .A(n10362), .B(n10361), .ZN(n10363) );
  XNOR2_X1 U13367 ( .A(n10367), .B(n16366), .ZN(n10369) );
  BUF_X2 U13368 ( .A(n11088), .Z(n11455) );
  NAND2_X1 U13369 ( .A1(n11455), .A2(n11114), .ZN(n10372) );
  XNOR2_X1 U13370 ( .A(n10374), .B(n10373), .ZN(n10378) );
  XNOR2_X1 U13371 ( .A(n10528), .B(n19027), .ZN(n10375) );
  XNOR2_X1 U13372 ( .A(n10376), .B(n10375), .ZN(n10377) );
  INV_X1 U13373 ( .A(n10379), .ZN(n10380) );
  XNOR2_X1 U13374 ( .A(n10380), .B(n10381), .ZN(n10386) );
  XNOR2_X1 U13375 ( .A(n10482), .B(n10382), .ZN(n10384) );
  XNOR2_X1 U13376 ( .A(n10384), .B(n10383), .ZN(n10385) );
  XNOR2_X1 U13377 ( .A(n10387), .B(n10388), .ZN(n10390) );
  XNOR2_X1 U13378 ( .A(n10570), .B(n18055), .ZN(n10389) );
  XNOR2_X1 U13379 ( .A(n10390), .B(n10389), .ZN(n10394) );
  XNOR2_X1 U13380 ( .A(n10392), .B(n10391), .ZN(n10393) );
  XNOR2_X1 U13381 ( .A(n10394), .B(n10393), .ZN(n11132) );
  XNOR2_X1 U13382 ( .A(n10395), .B(n10396), .ZN(n10400) );
  XNOR2_X1 U13383 ( .A(n10561), .B(n18078), .ZN(n10398) );
  XNOR2_X1 U13384 ( .A(n10397), .B(n10398), .ZN(n10399) );
  XNOR2_X1 U13385 ( .A(n10400), .B(n10399), .ZN(n10724) );
  AOI22_X1 U13386 ( .A1(n11133), .A2(n11131), .B1(n19837), .B2(n10724), .ZN(
        n11054) );
  INV_X1 U13387 ( .A(n11131), .ZN(n11420) );
  NOR2_X1 U13388 ( .A1(n11133), .A2(n11420), .ZN(n10414) );
  XNOR2_X1 U13389 ( .A(n10401), .B(n10402), .ZN(n10534) );
  XNOR2_X1 U13390 ( .A(n10534), .B(n10403), .ZN(n10408) );
  XNOR2_X1 U13391 ( .A(n10404), .B(n16035), .ZN(n10405) );
  XNOR2_X1 U13392 ( .A(n10406), .B(n10405), .ZN(n10407) );
  XNOR2_X1 U13394 ( .A(n10409), .B(n10410), .ZN(n10411) );
  OAI21_X1 U13395 ( .B1(n11054), .B2(n10414), .A(n10413), .ZN(n11997) );
  INV_X1 U13396 ( .A(n11997), .ZN(n12515) );
  XNOR2_X1 U13397 ( .A(n10416), .B(n10415), .ZN(n10420) );
  XNOR2_X1 U13398 ( .A(n10417), .B(n10418), .ZN(n10419) );
  XNOR2_X1 U13399 ( .A(n10420), .B(n10419), .ZN(n10450) );
  XNOR2_X1 U13400 ( .A(n10422), .B(n10421), .ZN(n10424) );
  XNOR2_X1 U13401 ( .A(n10424), .B(n20456), .ZN(n10429) );
  XNOR2_X1 U13402 ( .A(n10425), .B(n16651), .ZN(n10426) );
  XNOR2_X1 U13403 ( .A(n10427), .B(n10426), .ZN(n10428) );
  INV_X1 U13404 ( .A(n10430), .ZN(n10432) );
  XNOR2_X1 U13405 ( .A(n10432), .B(n10431), .ZN(n10434) );
  XNOR2_X1 U13406 ( .A(n10434), .B(n10433), .ZN(n10440) );
  INV_X1 U13407 ( .A(n18830), .ZN(n10435) );
  XNOR2_X1 U13408 ( .A(n10436), .B(n10435), .ZN(n10437) );
  XOR2_X1 U13409 ( .A(n10438), .B(n10437), .Z(n10439) );
  XNOR2_X1 U13411 ( .A(n10441), .B(n10442), .ZN(n10443) );
  XNOR2_X1 U13412 ( .A(n10444), .B(n10443), .ZN(n10449) );
  XNOR2_X1 U13413 ( .A(n10445), .B(n18433), .ZN(n10446) );
  XNOR2_X1 U13414 ( .A(n10447), .B(n10446), .ZN(n10448) );
  XNOR2_X1 U13415 ( .A(n10449), .B(n10448), .ZN(n11446) );
  NOR2_X1 U13416 ( .A1(n11446), .A2(n11202), .ZN(n10452) );
  INV_X1 U13417 ( .A(n19920), .ZN(n10451) );
  INV_X1 U13418 ( .A(n10453), .ZN(n10455) );
  XNOR2_X1 U13419 ( .A(n10455), .B(n10454), .ZN(n10460) );
  XNOR2_X1 U13420 ( .A(n10456), .B(n2275), .ZN(n10457) );
  XNOR2_X1 U13421 ( .A(n10458), .B(n10457), .ZN(n10459) );
  NAND2_X1 U13422 ( .A1(n11202), .A2(n10845), .ZN(n10468) );
  XNOR2_X1 U13423 ( .A(n10461), .B(n18984), .ZN(n10463) );
  XNOR2_X1 U13424 ( .A(n10463), .B(n10462), .ZN(n10467) );
  XNOR2_X1 U13425 ( .A(n10464), .B(n10465), .ZN(n10466) );
  XNOR2_X1 U13426 ( .A(n10467), .B(n10466), .ZN(n10726) );
  INV_X1 U13427 ( .A(n11995), .ZN(n12325) );
  XNOR2_X1 U13428 ( .A(n10472), .B(n18691), .ZN(n10474) );
  XNOR2_X1 U13429 ( .A(n10474), .B(n10473), .ZN(n10476) );
  XNOR2_X1 U13430 ( .A(n10476), .B(n10475), .ZN(n10479) );
  INV_X1 U13431 ( .A(n10477), .ZN(n10478) );
  XNOR2_X1 U13432 ( .A(n10480), .B(n10481), .ZN(n10488) );
  XNOR2_X1 U13433 ( .A(n10482), .B(n10483), .ZN(n10486) );
  XNOR2_X1 U13434 ( .A(n10484), .B(n18070), .ZN(n10485) );
  XNOR2_X1 U13435 ( .A(n10486), .B(n10485), .ZN(n10487) );
  XNOR2_X1 U13436 ( .A(n10488), .B(n10487), .ZN(n10513) );
  INV_X1 U13437 ( .A(n10489), .ZN(n10496) );
  XNOR2_X1 U13438 ( .A(n10490), .B(n2310), .ZN(n10492) );
  XNOR2_X1 U13439 ( .A(n10492), .B(n10491), .ZN(n10493) );
  XNOR2_X1 U13440 ( .A(n10494), .B(n10493), .ZN(n10495) );
  XNOR2_X1 U13441 ( .A(n10497), .B(n19243), .ZN(n10500) );
  INV_X1 U13442 ( .A(n10498), .ZN(n10499) );
  XNOR2_X1 U13443 ( .A(n10500), .B(n10499), .ZN(n10502) );
  XNOR2_X1 U13444 ( .A(n10502), .B(n10501), .ZN(n10504) );
  XNOR2_X1 U13445 ( .A(n10504), .B(n10503), .ZN(n11115) );
  NOR2_X1 U13446 ( .A1(n11116), .A2(n11115), .ZN(n10505) );
  XNOR2_X1 U13447 ( .A(n10506), .B(n2454), .ZN(n10507) );
  XNOR2_X1 U13448 ( .A(n10509), .B(n10508), .ZN(n10512) );
  INV_X1 U13449 ( .A(n10510), .ZN(n10511) );
  AND2_X1 U13450 ( .A1(n11037), .A2(n11440), .ZN(n11117) );
  XNOR2_X1 U13451 ( .A(n10566), .B(n10514), .ZN(n10516) );
  XNOR2_X1 U13452 ( .A(n10515), .B(n10516), .ZN(n10521) );
  INV_X1 U13453 ( .A(n10517), .ZN(n10519) );
  XNOR2_X1 U13454 ( .A(n10572), .B(n20682), .ZN(n10518) );
  XNOR2_X1 U13455 ( .A(n10519), .B(n10518), .ZN(n10520) );
  OAI21_X1 U13457 ( .B1(n11117), .B2(n11035), .A(n11116), .ZN(n10522) );
  XNOR2_X1 U13459 ( .A(n10524), .B(n10525), .ZN(n10532) );
  XNOR2_X1 U13460 ( .A(n10527), .B(n10526), .ZN(n10530) );
  XNOR2_X1 U13461 ( .A(n10528), .B(n18809), .ZN(n10529) );
  XNOR2_X1 U13462 ( .A(n10530), .B(n10529), .ZN(n10531) );
  XNOR2_X2 U13463 ( .A(n10532), .B(n10531), .ZN(n11193) );
  XNOR2_X1 U13464 ( .A(n10534), .B(n10533), .ZN(n10539) );
  XNOR2_X1 U13465 ( .A(n10613), .B(n18887), .ZN(n10537) );
  INV_X1 U13466 ( .A(n10535), .ZN(n10536) );
  XNOR2_X1 U13467 ( .A(n10536), .B(n10537), .ZN(n10538) );
  XNOR2_X1 U13468 ( .A(n10540), .B(n10541), .ZN(n10547) );
  XNOR2_X1 U13469 ( .A(n865), .B(n311), .ZN(n10545) );
  INV_X1 U13470 ( .A(n10543), .ZN(n10544) );
  XNOR2_X1 U13471 ( .A(n10544), .B(n10545), .ZN(n10546) );
  NAND2_X1 U13472 ( .A1(n11186), .A2(n19983), .ZN(n10903) );
  XNOR2_X1 U13473 ( .A(n10548), .B(n10549), .ZN(n10556) );
  XNOR2_X1 U13474 ( .A(n10550), .B(n2032), .ZN(n10554) );
  XNOR2_X1 U13475 ( .A(n10552), .B(n10551), .ZN(n10553) );
  XNOR2_X1 U13476 ( .A(n10554), .B(n10553), .ZN(n10555) );
  XNOR2_X1 U13477 ( .A(n10557), .B(n10558), .ZN(n10560) );
  XNOR2_X1 U13478 ( .A(n10560), .B(n10559), .ZN(n10565) );
  XNOR2_X1 U13479 ( .A(n10561), .B(n19336), .ZN(n10562) );
  XNOR2_X1 U13480 ( .A(n10562), .B(n10563), .ZN(n10564) );
  XNOR2_X1 U13481 ( .A(n10564), .B(n10565), .ZN(n10575) );
  XNOR2_X1 U13482 ( .A(n10566), .B(n10567), .ZN(n10569) );
  XNOR2_X1 U13483 ( .A(n10571), .B(n10570), .ZN(n10574) );
  XNOR2_X1 U13484 ( .A(n10572), .B(n2376), .ZN(n10573) );
  OAI21_X1 U13485 ( .B1(n11500), .B2(n11499), .A(n11192), .ZN(n10577) );
  INV_X1 U13486 ( .A(n10575), .ZN(n11188) );
  NAND2_X1 U13487 ( .A1(n11188), .A2(n11192), .ZN(n11502) );
  INV_X1 U13488 ( .A(n11502), .ZN(n10576) );
  NAND2_X1 U13489 ( .A1(n11995), .A2(n11820), .ZN(n10627) );
  XNOR2_X1 U13490 ( .A(n10578), .B(n10579), .ZN(n10581) );
  XNOR2_X1 U13491 ( .A(n10581), .B(n10580), .ZN(n10586) );
  XNOR2_X1 U13492 ( .A(n10582), .B(n19180), .ZN(n10583) );
  XNOR2_X1 U13493 ( .A(n10584), .B(n10583), .ZN(n10585) );
  INV_X1 U13494 ( .A(n11491), .ZN(n11495) );
  XNOR2_X1 U13495 ( .A(n10588), .B(n10587), .ZN(n10593) );
  XNOR2_X1 U13496 ( .A(n10589), .B(n19140), .ZN(n10590) );
  XNOR2_X1 U13497 ( .A(n10591), .B(n10590), .ZN(n10592) );
  XNOR2_X1 U13498 ( .A(n10594), .B(n10595), .ZN(n10597) );
  XNOR2_X1 U13499 ( .A(n10596), .B(n10597), .ZN(n10602) );
  INV_X1 U13500 ( .A(Key[124]), .ZN(n18517) );
  XNOR2_X1 U13501 ( .A(n10598), .B(n18517), .ZN(n10599) );
  XNOR2_X1 U13502 ( .A(n10600), .B(n10599), .ZN(n10601) );
  INV_X1 U13504 ( .A(n10603), .ZN(n10608) );
  XNOR2_X1 U13505 ( .A(n10606), .B(n10605), .ZN(n10607) );
  XNOR2_X1 U13506 ( .A(n10608), .B(n10607), .ZN(n10610) );
  XNOR2_X1 U13507 ( .A(n961), .B(n10611), .ZN(n10617) );
  XNOR2_X1 U13508 ( .A(n10613), .B(n10612), .ZN(n10616) );
  XNOR2_X1 U13509 ( .A(n20210), .B(n2096), .ZN(n10615) );
  XNOR2_X1 U13510 ( .A(n10619), .B(n10618), .ZN(n10622) );
  NOR2_X1 U13511 ( .A1(n11494), .A2(n11493), .ZN(n10623) );
  INV_X1 U13513 ( .A(n10625), .ZN(n12326) );
  NAND2_X1 U13514 ( .A1(n12513), .A2(n12326), .ZN(n10626) );
  OAI22_X1 U13515 ( .A1(n20073), .A2(n10627), .B1(n10626), .B2(n13275), .ZN(
        n10629) );
  AOI21_X1 U13516 ( .B1(n13275), .B2(n10630), .A(n10629), .ZN(n12962) );
  INV_X1 U13517 ( .A(n12962), .ZN(n13590) );
  INV_X1 U13518 ( .A(n2100), .ZN(n15021) );
  XNOR2_X1 U13519 ( .A(n13590), .B(n15021), .ZN(n10631) );
  XNOR2_X1 U13520 ( .A(n10632), .B(n10631), .ZN(n10633) );
  XNOR2_X1 U13521 ( .A(n10633), .B(n10634), .ZN(n14775) );
  INV_X1 U13522 ( .A(n14775), .ZN(n14057) );
  AOI21_X1 U13523 ( .B1(n11528), .B2(n11521), .A(n10635), .ZN(n10636) );
  INV_X1 U13524 ( .A(n11528), .ZN(n10921) );
  MUX2_X1 U13525 ( .A(n10636), .B(n10924), .S(n10755), .Z(n10637) );
  NOR2_X1 U13526 ( .A1(n10638), .A2(n10640), .ZN(n10932) );
  NOR2_X1 U13527 ( .A1(n11168), .A2(n11539), .ZN(n10639) );
  OAI211_X1 U13528 ( .C1(n11534), .C2(n11170), .A(n11538), .B(n11168), .ZN(
        n10641) );
  OAI21_X1 U13529 ( .B1(n10737), .B2(n11169), .A(n10641), .ZN(n12422) );
  NAND2_X1 U13530 ( .A1(n12415), .A2(n12422), .ZN(n11312) );
  AOI22_X1 U13531 ( .A1(n1721), .A2(n20366), .B1(n10642), .B2(n10960), .ZN(
        n10644) );
  NAND2_X1 U13532 ( .A1(n11142), .A2(n10642), .ZN(n10957) );
  MUX2_X1 U13533 ( .A(n10960), .B(n10957), .S(n11145), .Z(n10643) );
  OAI21_X2 U13534 ( .B1(n10644), .B2(n10701), .A(n10643), .ZN(n12416) );
  NAND2_X1 U13537 ( .A1(n12416), .A2(n20352), .ZN(n11311) );
  NAND2_X1 U13538 ( .A1(n11161), .A2(n10649), .ZN(n10654) );
  NAND2_X1 U13539 ( .A1(n10650), .A2(n11159), .ZN(n10651) );
  MUX2_X1 U13540 ( .A(n10652), .B(n10651), .S(n10945), .Z(n10653) );
  INV_X1 U13542 ( .A(n11602), .ZN(n12419) );
  AOI21_X1 U13543 ( .B1(n11312), .B2(n11311), .A(n12419), .ZN(n10659) );
  AOI21_X1 U13546 ( .B1(n12083), .B2(n12415), .A(n20352), .ZN(n10658) );
  NAND2_X1 U13548 ( .A1(n11659), .A2(n11830), .ZN(n11954) );
  NAND2_X1 U13549 ( .A1(n11957), .A2(n11954), .ZN(n10660) );
  XNOR2_X1 U13550 ( .A(n13088), .B(n13192), .ZN(n11975) );
  AOI22_X1 U13551 ( .A1(n11254), .A2(n11253), .B1(n11256), .B2(n11255), .ZN(
        n10663) );
  NAND2_X1 U13552 ( .A1(n11256), .A2(n11257), .ZN(n10664) );
  MUX2_X1 U13553 ( .A(n11255), .B(n10664), .S(n191), .Z(n10665) );
  INV_X1 U13554 ( .A(n11395), .ZN(n11296) );
  NAND2_X1 U13555 ( .A1(n2724), .A2(n10667), .ZN(n10668) );
  INV_X1 U13556 ( .A(n10986), .ZN(n11398) );
  INV_X1 U13557 ( .A(n11397), .ZN(n11295) );
  MUX2_X1 U13558 ( .A(n10668), .B(n11398), .S(n11295), .Z(n10669) );
  NAND2_X1 U13559 ( .A1(n12099), .A2(n12435), .ZN(n10687) );
  MUX2_X1 U13560 ( .A(n11267), .B(n11265), .S(n11339), .Z(n10674) );
  NAND2_X1 U13561 ( .A1(n11263), .A2(n11265), .ZN(n10671) );
  NAND2_X1 U13562 ( .A1(n10673), .A2(n9830), .ZN(n10670) );
  MUX2_X1 U13563 ( .A(n10671), .B(n10670), .S(n11343), .Z(n10672) );
  INV_X1 U13564 ( .A(n10675), .ZN(n10818) );
  NOR2_X1 U13565 ( .A1(n10852), .A2(n11231), .ZN(n10678) );
  MUX2_X1 U13566 ( .A(n10679), .B(n10678), .S(n11366), .Z(n10682) );
  NAND2_X1 U13567 ( .A1(n10818), .A2(n11234), .ZN(n10680) );
  NOR2_X1 U13568 ( .A1(n12437), .A2(n12440), .ZN(n11065) );
  AOI21_X2 U13569 ( .B1(n10687), .B2(n10686), .A(n11065), .ZN(n13618) );
  MUX2_X1 U13570 ( .A(n11408), .B(n10688), .S(n19736), .Z(n10692) );
  NAND2_X1 U13571 ( .A1(n11000), .A2(n11278), .ZN(n11410) );
  INV_X1 U13572 ( .A(n11410), .ZN(n10690) );
  NOR2_X1 U13573 ( .A1(n11278), .A2(n11413), .ZN(n10689) );
  AOI22_X1 U13574 ( .A1(n10690), .A2(n11411), .B1(n10689), .B2(n11408), .ZN(
        n10691) );
  INV_X1 U13575 ( .A(n12631), .ZN(n12629) );
  MUX2_X1 U13576 ( .A(n10947), .B(n10693), .S(n19779), .Z(n10695) );
  NOR2_X1 U13577 ( .A1(n9559), .A2(n10694), .ZN(n10999) );
  NOR2_X1 U13578 ( .A1(n10980), .A2(n11294), .ZN(n10697) );
  NOR2_X1 U13579 ( .A1(n20235), .A2(n11290), .ZN(n10696) );
  NAND2_X1 U13581 ( .A1(n11292), .A2(n11403), .ZN(n10698) );
  AOI21_X1 U13582 ( .B1(n10698), .B2(n11293), .A(n11291), .ZN(n10699) );
  NOR2_X2 U13583 ( .A1(n10700), .A2(n10699), .ZN(n12634) );
  OAI22_X1 U13584 ( .A1(n11145), .A2(n1749), .B1(n20366), .B2(n10701), .ZN(
        n10703) );
  NAND3_X1 U13586 ( .A1(n11148), .A2(n11147), .A3(n11009), .ZN(n10704) );
  NAND2_X1 U13587 ( .A1(n11009), .A2(n10953), .ZN(n11152) );
  INV_X1 U13589 ( .A(n10709), .ZN(n11869) );
  OAI21_X1 U13590 ( .B1(n20601), .B2(n11866), .A(n11869), .ZN(n10710) );
  INV_X1 U13591 ( .A(n10711), .ZN(n10712) );
  INV_X1 U13592 ( .A(n11871), .ZN(n11388) );
  NAND2_X1 U13593 ( .A1(n10712), .A2(n11388), .ZN(n10713) );
  INV_X1 U13594 ( .A(n12634), .ZN(n10716) );
  XNOR2_X1 U13595 ( .A(n13415), .B(n11975), .ZN(n10795) );
  NAND2_X1 U13596 ( .A1(n10717), .A2(n11076), .ZN(n10718) );
  INV_X1 U13597 ( .A(n11191), .ZN(n11501) );
  NOR2_X1 U13598 ( .A1(n11500), .A2(n11501), .ZN(n10719) );
  NOR2_X1 U13600 ( .A1(n11193), .A2(n19983), .ZN(n10721) );
  NOR2_X1 U13601 ( .A1(n11192), .A2(n11188), .ZN(n10720) );
  AOI22_X1 U13602 ( .A1(n10721), .A2(n11186), .B1(n10720), .B2(n11193), .ZN(
        n10722) );
  INV_X1 U13603 ( .A(n12648), .ZN(n12645) );
  INV_X1 U13604 ( .A(n11132), .ZN(n11417) );
  INV_X1 U13605 ( .A(n11446), .ZN(n10847) );
  MUX2_X1 U13606 ( .A(n10847), .B(n11093), .S(n19920), .Z(n10728) );
  MUX2_X2 U13607 ( .A(n10728), .B(n10727), .S(n11094), .Z(n12684) );
  INV_X1 U13608 ( .A(n10730), .ZN(n11069) );
  NAND2_X1 U13609 ( .A1(n11069), .A2(n11489), .ZN(n10732) );
  NAND2_X1 U13610 ( .A1(n19505), .A2(n19719), .ZN(n10731) );
  INV_X1 U13611 ( .A(n11456), .ZN(n11091) );
  OAI21_X1 U13612 ( .B1(n10734), .B2(n11091), .A(n10733), .ZN(n10736) );
  AOI21_X1 U13613 ( .B1(n10734), .B2(n11114), .A(n11455), .ZN(n10735) );
  NOR2_X1 U13614 ( .A1(n10736), .A2(n10735), .ZN(n12430) );
  AND2_X2 U13615 ( .A1(n10739), .A2(n10738), .ZN(n12759) );
  INV_X1 U13616 ( .A(n12759), .ZN(n12410) );
  INV_X1 U13617 ( .A(n11514), .ZN(n10906) );
  INV_X1 U13618 ( .A(n11515), .ZN(n10935) );
  INV_X1 U13619 ( .A(n10740), .ZN(n10741) );
  OAI21_X1 U13620 ( .B1(n10906), .B2(n11513), .A(n10741), .ZN(n10743) );
  INV_X1 U13622 ( .A(n10896), .ZN(n11483) );
  AOI21_X1 U13623 ( .B1(n11487), .B2(n11483), .A(n20233), .ZN(n10750) );
  NAND2_X1 U13624 ( .A1(n10745), .A2(n20233), .ZN(n10747) );
  AOI21_X1 U13625 ( .B1(n10748), .B2(n10747), .A(n3500), .ZN(n10749) );
  NOR2_X1 U13626 ( .A1(n898), .A2(n11568), .ZN(n10754) );
  NAND2_X1 U13627 ( .A1(n10883), .A2(n11566), .ZN(n10753) );
  INV_X1 U13628 ( .A(n10883), .ZN(n11567) );
  NAND2_X1 U13629 ( .A1(n11567), .A2(n11466), .ZN(n10751) );
  AOI22_X1 U13631 ( .A1(n12410), .A2(n12754), .B1(n254), .B2(n12407), .ZN(
        n11315) );
  NAND2_X1 U13633 ( .A1(n10755), .A2(n11527), .ZN(n10757) );
  INV_X1 U13634 ( .A(n12754), .ZN(n10766) );
  NAND3_X1 U13635 ( .A1(n10889), .A2(n10760), .A3(n11546), .ZN(n10763) );
  INV_X1 U13636 ( .A(n12407), .ZN(n11313) );
  OAI21_X1 U13637 ( .B1(n12389), .B2(n11313), .A(n254), .ZN(n10765) );
  NAND2_X1 U13638 ( .A1(n10766), .A2(n10765), .ZN(n10767) );
  INV_X1 U13639 ( .A(n11430), .ZN(n10768) );
  NOR2_X1 U13640 ( .A1(n19830), .A2(n10768), .ZN(n10770) );
  MUX2_X1 U13641 ( .A(n10770), .B(n10769), .S(n11041), .Z(n10773) );
  INV_X1 U13642 ( .A(n11105), .ZN(n11429) );
  NAND2_X1 U13644 ( .A1(n11105), .A2(n19830), .ZN(n11109) );
  NOR2_X2 U13646 ( .A1(n10773), .A2(n10772), .ZN(n12639) );
  OAI21_X1 U13647 ( .B1(n10802), .B2(n10774), .A(n11257), .ZN(n10778) );
  INV_X1 U13648 ( .A(n11255), .ZN(n10775) );
  MUX2_X1 U13649 ( .A(n10776), .B(n10775), .S(n11253), .Z(n10777) );
  NAND2_X1 U13650 ( .A1(n10778), .A2(n10777), .ZN(n12453) );
  NAND2_X1 U13651 ( .A1(n11238), .A2(n10779), .ZN(n11236) );
  OAI211_X1 U13652 ( .C1(n11349), .C2(n11057), .A(n11239), .B(n10798), .ZN(
        n10780) );
  NAND2_X1 U13653 ( .A1(n11347), .A2(n11057), .ZN(n11237) );
  OAI211_X1 U13654 ( .C1(n11057), .C2(n11236), .A(n10780), .B(n11237), .ZN(
        n12449) );
  NAND2_X1 U13655 ( .A1(n12453), .A2(n12449), .ZN(n11946) );
  INV_X1 U13656 ( .A(n11115), .ZN(n11439) );
  NAND2_X1 U13657 ( .A1(n11439), .A2(n11035), .ZN(n10782) );
  NAND2_X1 U13658 ( .A1(n11034), .A2(n11440), .ZN(n10781) );
  NAND2_X1 U13659 ( .A1(n10782), .A2(n10781), .ZN(n10833) );
  OAI21_X1 U13660 ( .B1(n11438), .B2(n11115), .A(n11035), .ZN(n10784) );
  NAND2_X1 U13661 ( .A1(n12637), .A2(n12642), .ZN(n10792) );
  MUX2_X1 U13662 ( .A(n11886), .B(n11880), .S(n11120), .Z(n10789) );
  NAND2_X1 U13663 ( .A1(n12636), .A2(n12449), .ZN(n12089) );
  INV_X1 U13664 ( .A(n12089), .ZN(n10790) );
  INV_X1 U13665 ( .A(n12453), .ZN(n12450) );
  INV_X1 U13666 ( .A(n12642), .ZN(n12452) );
  OAI21_X1 U13667 ( .B1(n10790), .B2(n12450), .A(n12452), .ZN(n10791) );
  XNOR2_X1 U13669 ( .A(n13617), .B(n13336), .ZN(n13305) );
  XNOR2_X1 U13670 ( .A(n13305), .B(n10793), .ZN(n10794) );
  NOR2_X1 U13671 ( .A1(n11337), .A2(n11263), .ZN(n10796) );
  AND2_X1 U13672 ( .A1(n11355), .A2(n10798), .ZN(n10799) );
  AND2_X1 U13673 ( .A1(n11239), .A2(n11347), .ZN(n10800) );
  INV_X1 U13674 ( .A(n10800), .ZN(n10801) );
  NAND2_X1 U13675 ( .A1(n12212), .A2(n12208), .ZN(n11639) );
  NAND2_X1 U13676 ( .A1(n10805), .A2(n10804), .ZN(n10807) );
  AND2_X1 U13677 ( .A1(n11321), .A2(n11253), .ZN(n11324) );
  AOI21_X1 U13678 ( .B1(n11124), .B2(n10809), .A(n11459), .ZN(n10812) );
  AOI21_X1 U13679 ( .B1(n10810), .B2(n11048), .A(n11883), .ZN(n10811) );
  NOR2_X1 U13680 ( .A1(n20099), .A2(n11125), .ZN(n10816) );
  NOR2_X1 U13681 ( .A1(n11127), .A2(n10813), .ZN(n10815) );
  OAI22_X1 U13682 ( .A1(n10818), .A2(n1601), .B1(n11231), .B2(n11234), .ZN(
        n10820) );
  INV_X1 U13683 ( .A(n11235), .ZN(n10819) );
  NOR2_X1 U13684 ( .A1(n9883), .A2(n10854), .ZN(n11638) );
  INV_X1 U13685 ( .A(n11638), .ZN(n11808) );
  NOR2_X1 U13686 ( .A1(n11811), .A2(n10821), .ZN(n10822) );
  NAND2_X1 U13687 ( .A1(n913), .A2(n3051), .ZN(n11200) );
  NAND2_X1 U13688 ( .A1(n11199), .A2(n11200), .ZN(n10825) );
  OAI21_X1 U13689 ( .B1(n19719), .B2(n19913), .A(n913), .ZN(n10824) );
  INV_X1 U13690 ( .A(n12061), .ZN(n11637) );
  NAND3_X1 U13691 ( .A1(n11042), .A2(n11106), .A3(n11105), .ZN(n10828) );
  NOR2_X1 U13693 ( .A1(n1378), .A2(n11430), .ZN(n10826) );
  INV_X1 U13695 ( .A(n12202), .ZN(n12591) );
  NOR2_X1 U13696 ( .A1(n11637), .A2(n12591), .ZN(n10844) );
  INV_X1 U13699 ( .A(n12594), .ZN(n12590) );
  OAI211_X1 U13700 ( .C1(n11037), .C2(n11440), .A(n11115), .B(n11438), .ZN(
        n10835) );
  NAND2_X1 U13701 ( .A1(n11451), .A2(n11455), .ZN(n10843) );
  INV_X1 U13702 ( .A(n11088), .ZN(n10839) );
  NAND2_X1 U13703 ( .A1(n10839), .A2(n11452), .ZN(n10838) );
  OAI21_X1 U13704 ( .B1(n11451), .B2(n11452), .A(n10838), .ZN(n10841) );
  NAND2_X1 U13705 ( .A1(n10839), .A2(n11113), .ZN(n11112) );
  NAND2_X1 U13706 ( .A1(n11112), .A2(n11114), .ZN(n10840) );
  OAI21_X1 U13707 ( .B1(n10841), .B2(n11114), .A(n10840), .ZN(n10842) );
  AOI21_X1 U13708 ( .B1(n10845), .B2(n11445), .A(n11443), .ZN(n10846) );
  INV_X1 U13709 ( .A(n10845), .ZN(n11444) );
  XNOR2_X1 U13710 ( .A(n13577), .B(n10849), .ZN(n13357) );
  INV_X1 U13711 ( .A(n13357), .ZN(n10881) );
  INV_X1 U13712 ( .A(n11670), .ZN(n12185) );
  NOR2_X1 U13713 ( .A1(n11841), .A2(n20427), .ZN(n11844) );
  NAND2_X1 U13714 ( .A1(n11844), .A2(n11670), .ZN(n10850) );
  INV_X1 U13715 ( .A(n11369), .ZN(n10853) );
  NOR2_X1 U13716 ( .A1(n10854), .A2(n11234), .ZN(n10855) );
  NAND2_X1 U13718 ( .A1(n10986), .A2(n11397), .ZN(n10859) );
  AOI21_X1 U13719 ( .B1(n19756), .B2(n12057), .A(n874), .ZN(n10879) );
  INV_X1 U13720 ( .A(n19750), .ZN(n11867) );
  NAND2_X1 U13721 ( .A1(n20601), .A2(n11866), .ZN(n11305) );
  INV_X1 U13722 ( .A(n11305), .ZN(n10863) );
  NAND2_X1 U13724 ( .A1(n10868), .A2(n10867), .ZN(n12615) );
  NAND2_X1 U13725 ( .A1(n11380), .A2(n12103), .ZN(n10866) );
  NAND2_X1 U13726 ( .A1(n10864), .A2(n12101), .ZN(n10865) );
  MUX2_X1 U13727 ( .A(n10866), .B(n10865), .S(n11381), .Z(n11632) );
  NAND4_X1 U13728 ( .A1(n11632), .A2(n10868), .A3(n11633), .A4(n10867), .ZN(
        n10869) );
  OAI22_X1 U13729 ( .A1(n19756), .A2(n12053), .B1(n10869), .B2(n12240), .ZN(
        n10878) );
  OAI22_X1 U13730 ( .A1(n10978), .A2(n19506), .B1(n11402), .B2(n3588), .ZN(
        n10871) );
  OAI22_X1 U13731 ( .A1(n11293), .A2(n20235), .B1(n11403), .B2(n11291), .ZN(
        n10870) );
  INV_X1 U13732 ( .A(n11632), .ZN(n10875) );
  INV_X1 U13733 ( .A(n10873), .ZN(n10874) );
  NOR2_X1 U13734 ( .A1(n10875), .A2(n10874), .ZN(n10876) );
  XNOR2_X1 U13735 ( .A(n13827), .B(n19854), .ZN(n10880) );
  XNOR2_X1 U13736 ( .A(n10881), .B(n10880), .ZN(n10977) );
  INV_X1 U13737 ( .A(n10882), .ZN(n11469) );
  MUX2_X1 U13738 ( .A(n11568), .B(n10884), .S(n10883), .Z(n10888) );
  NAND2_X1 U13739 ( .A1(n11565), .A2(n11569), .ZN(n10887) );
  INV_X1 U13740 ( .A(n927), .ZN(n11467) );
  INV_X1 U13741 ( .A(n11466), .ZN(n11564) );
  NOR2_X1 U13742 ( .A1(n11467), .A2(n10885), .ZN(n10886) );
  OAI22_X1 U13744 ( .A1(n647), .A2(n10926), .B1(n10889), .B2(n11547), .ZN(
        n10890) );
  NAND2_X1 U13745 ( .A1(n11544), .A2(n647), .ZN(n10892) );
  INV_X1 U13746 ( .A(n11217), .ZN(n10895) );
  MUX2_X1 U13747 ( .A(n19897), .B(n10896), .S(n10060), .Z(n10900) );
  INV_X1 U13748 ( .A(n10898), .ZN(n10899) );
  AOI22_X1 U13749 ( .A1(n11193), .A2(n19983), .B1(n11188), .B2(n11500), .ZN(
        n10901) );
  NOR2_X1 U13750 ( .A1(n10901), .A2(n11186), .ZN(n10905) );
  AOI21_X1 U13751 ( .B1(n10903), .B2(n19998), .A(n11500), .ZN(n10904) );
  NOR2_X1 U13752 ( .A1(n10905), .A2(n10904), .ZN(n12601) );
  NAND2_X1 U13753 ( .A1(n12609), .A2(n12601), .ZN(n10911) );
  NAND3_X1 U13755 ( .A1(n20106), .A2(n20639), .A3(n11572), .ZN(n10910) );
  NAND3_X1 U13756 ( .A1(n11510), .A2(n19864), .A3(n10936), .ZN(n10909) );
  NAND3_X1 U13757 ( .A1(n10935), .A2(n11510), .A3(n10906), .ZN(n10907) );
  INV_X1 U13759 ( .A(n10913), .ZN(n11557) );
  MUX2_X1 U13760 ( .A(n11556), .B(n11557), .S(n10914), .Z(n10918) );
  INV_X1 U13761 ( .A(n11553), .ZN(n11163) );
  NAND2_X1 U13762 ( .A1(n11556), .A2(n11559), .ZN(n10915) );
  MUX2_X1 U13763 ( .A(n10916), .B(n10915), .S(n20479), .Z(n10917) );
  OAI21_X1 U13764 ( .B1(n10918), .B2(n19564), .A(n10917), .ZN(n12232) );
  NAND2_X1 U13765 ( .A1(n12230), .A2(n12232), .ZN(n12048) );
  MUX2_X1 U13766 ( .A(n11523), .B(n19999), .S(n2470), .Z(n10922) );
  NOR2_X1 U13767 ( .A1(n10922), .A2(n10921), .ZN(n12223) );
  INV_X1 U13768 ( .A(n12121), .ZN(n10944) );
  NAND2_X1 U13769 ( .A1(n258), .A2(n10926), .ZN(n10927) );
  NAND3_X1 U13770 ( .A1(n11548), .A2(n258), .A3(n11549), .ZN(n10929) );
  AND3_X2 U13771 ( .A1(n10931), .A2(n10930), .A3(n10929), .ZN(n12122) );
  INV_X1 U13772 ( .A(n12122), .ZN(n12226) );
  NAND2_X1 U13773 ( .A1(n10932), .A2(n11533), .ZN(n10933) );
  NOR2_X1 U13774 ( .A1(n20639), .A2(n10935), .ZN(n10940) );
  OAI21_X1 U13775 ( .B1(n11573), .B2(n19864), .A(n10936), .ZN(n10939) );
  NAND2_X1 U13776 ( .A1(n11573), .A2(n11513), .ZN(n10937) );
  INV_X1 U13778 ( .A(n12228), .ZN(n10941) );
  XNOR2_X1 U13780 ( .A(n13058), .B(n13580), .ZN(n12791) );
  NAND2_X1 U13781 ( .A1(n10946), .A2(n10693), .ZN(n10996) );
  OAI21_X1 U13782 ( .B1(n11284), .B2(n11283), .A(n10693), .ZN(n10948) );
  NAND2_X1 U13783 ( .A1(n10948), .A2(n10947), .ZN(n10949) );
  NAND2_X1 U13784 ( .A1(n12130), .A2(n12126), .ZN(n11760) );
  MUX2_X1 U13785 ( .A(n11010), .B(n20470), .S(n10951), .Z(n10955) );
  NAND2_X1 U13786 ( .A1(n3382), .A2(n10952), .ZN(n10954) );
  MUX2_X1 U13787 ( .A(n10955), .B(n10954), .S(n10953), .Z(n10956) );
  INV_X1 U13788 ( .A(n12127), .ZN(n11701) );
  INV_X1 U13789 ( .A(n10957), .ZN(n10959) );
  NAND2_X1 U13791 ( .A1(n11176), .A2(n11178), .ZN(n10965) );
  OAI211_X1 U13792 ( .C1(n19878), .C2(n11178), .A(n11174), .B(n3789), .ZN(
        n10964) );
  OAI211_X1 U13793 ( .C1(n10966), .C2(n11178), .A(n10965), .B(n10964), .ZN(
        n12128) );
  NOR2_X1 U13794 ( .A1(n11586), .A2(n12128), .ZN(n10967) );
  AND2_X1 U13795 ( .A1(n12126), .A2(n12128), .ZN(n10972) );
  AOI21_X1 U13796 ( .B1(n11163), .B2(n20479), .A(n11559), .ZN(n10971) );
  OAI22_X1 U13797 ( .A1(n19957), .A2(n19564), .B1(n10913), .B2(n11556), .ZN(
        n10970) );
  OAI211_X2 U13798 ( .C1(n11701), .C2(n11760), .A(n10974), .B(n10973), .ZN(
        n13020) );
  XNOR2_X1 U13799 ( .A(n13020), .B(n2164), .ZN(n10975) );
  XNOR2_X1 U13800 ( .A(n12791), .B(n10975), .ZN(n10976) );
  XNOR2_X1 U13801 ( .A(n10977), .B(n10976), .ZN(n13901) );
  NOR2_X1 U13802 ( .A1(n11292), .A2(n11294), .ZN(n10982) );
  NOR2_X1 U13803 ( .A1(n10980), .A2(n11290), .ZN(n10981) );
  MUX2_X1 U13804 ( .A(n10982), .B(n10981), .S(n11403), .Z(n10983) );
  NAND2_X1 U13805 ( .A1(n10985), .A2(n11297), .ZN(n10989) );
  OAI21_X1 U13806 ( .B1(n11394), .B2(n11397), .A(n10986), .ZN(n10987) );
  NAND2_X1 U13807 ( .A1(n10987), .A2(n11395), .ZN(n10988) );
  NAND2_X1 U13808 ( .A1(n11686), .A2(n11683), .ZN(n11018) );
  NOR2_X1 U13809 ( .A1(n11388), .A2(n10990), .ZN(n10992) );
  MUX2_X1 U13811 ( .A(n10992), .B(n10991), .S(n11869), .Z(n10994) );
  NOR2_X1 U13812 ( .A1(n11871), .A2(n11390), .ZN(n11385) );
  NAND2_X1 U13813 ( .A1(n11385), .A2(n11302), .ZN(n11874) );
  INV_X1 U13814 ( .A(n11874), .ZN(n10993) );
  NAND2_X1 U13815 ( .A1(n20462), .A2(n11922), .ZN(n11007) );
  NOR2_X1 U13816 ( .A1(n19851), .A2(n11278), .ZN(n11002) );
  NOR2_X1 U13817 ( .A1(n11277), .A2(n10688), .ZN(n11001) );
  OAI21_X1 U13818 ( .B1(n11002), .B2(n11001), .A(n937), .ZN(n11004) );
  NAND3_X1 U13819 ( .A1(n11408), .A2(n11278), .A3(n11413), .ZN(n11003) );
  NAND2_X1 U13820 ( .A1(n11007), .A2(n12579), .ZN(n11008) );
  AOI21_X1 U13821 ( .B1(n11009), .B2(n3382), .A(n11149), .ZN(n11015) );
  NOR2_X1 U13822 ( .A1(n11148), .A2(n11010), .ZN(n11012) );
  OAI21_X1 U13823 ( .B1(n11013), .B2(n11012), .A(n11011), .ZN(n11014) );
  OAI21_X1 U13824 ( .B1(n11016), .B2(n11015), .A(n11014), .ZN(n11863) );
  INV_X1 U13825 ( .A(n12502), .ZN(n11020) );
  NAND3_X1 U13826 ( .A1(n11020), .A2(n12004), .A3(n201), .ZN(n11022) );
  INV_X1 U13827 ( .A(n12499), .ZN(n11019) );
  OAI211_X1 U13828 ( .C1(n12497), .C2(n12500), .A(n11022), .B(n11021), .ZN(
        n11024) );
  NOR2_X1 U13829 ( .A1(n12345), .A2(n12500), .ZN(n11023) );
  NAND2_X1 U13830 ( .A1(n12419), .A2(n20351), .ZN(n11025) );
  OAI21_X1 U13831 ( .B1(n12419), .B2(n12084), .A(n11025), .ZN(n11028) );
  INV_X1 U13832 ( .A(n12416), .ZN(n12418) );
  INV_X1 U13833 ( .A(n12422), .ZN(n11603) );
  NOR2_X1 U13834 ( .A1(n11603), .A2(n12084), .ZN(n11026) );
  AOI22_X1 U13835 ( .A1(n11026), .A2(n12419), .B1(n12415), .B2(n12084), .ZN(
        n11027) );
  OAI21_X2 U13836 ( .B1(n11028), .B2(n12418), .A(n11027), .ZN(n13657) );
  XNOR2_X1 U13837 ( .A(n11029), .B(n13657), .ZN(n13076) );
  INV_X1 U13838 ( .A(n13076), .ZN(n11103) );
  INV_X1 U13839 ( .A(n12354), .ZN(n11031) );
  NAND3_X1 U13840 ( .A1(n12001), .A2(n12352), .A3(n11031), .ZN(n11033) );
  XNOR2_X1 U13841 ( .A(n13715), .B(n2344), .ZN(n11064) );
  NOR2_X1 U13842 ( .A1(n11034), .A2(n11439), .ZN(n11036) );
  INV_X1 U13843 ( .A(n11035), .ZN(n11119) );
  INV_X1 U13844 ( .A(n11037), .ZN(n11436) );
  NOR3_X1 U13845 ( .A1(n11435), .A2(n11440), .A3(n11436), .ZN(n11891) );
  INV_X1 U13846 ( .A(n11038), .ZN(n11040) );
  NAND2_X1 U13847 ( .A1(n1039), .A2(n1317), .ZN(n11039) );
  INV_X1 U13848 ( .A(n12261), .ZN(n12563) );
  NAND2_X1 U13849 ( .A1(n11428), .A2(n11105), .ZN(n11043) );
  MUX2_X1 U13850 ( .A(n11043), .B(n11042), .S(n11041), .Z(n11047) );
  NOR2_X1 U13851 ( .A1(n11428), .A2(n1378), .ZN(n11045) );
  NOR2_X1 U13852 ( .A1(n19830), .A2(n11105), .ZN(n11044) );
  AOI22_X1 U13853 ( .A1(n11045), .A2(n11427), .B1(n11044), .B2(n11106), .ZN(
        n11046) );
  NAND2_X1 U13854 ( .A1(n11047), .A2(n11046), .ZN(n11061) );
  OAI21_X1 U13855 ( .B1(n11129), .B2(n11051), .A(n19837), .ZN(n11052) );
  OAI21_X2 U13856 ( .B1(n11054), .B2(n19959), .A(n11053), .ZN(n12262) );
  OAI21_X1 U13857 ( .B1(n12563), .B2(n12016), .A(n12565), .ZN(n11063) );
  NOR2_X1 U13858 ( .A1(n11346), .A2(n11239), .ZN(n11056) );
  AOI22_X1 U13859 ( .A1(n11056), .A2(n11055), .B1(n11346), .B2(n11238), .ZN(
        n11059) );
  NAND3_X1 U13860 ( .A1(n11349), .A2(n11057), .A3(n11346), .ZN(n11058) );
  OAI211_X1 U13861 ( .C1(n11060), .C2(n11348), .A(n11059), .B(n11058), .ZN(
        n12264) );
  INV_X1 U13862 ( .A(n11061), .ZN(n12562) );
  XNOR2_X1 U13864 ( .A(n11064), .B(n13321), .ZN(n11101) );
  NAND2_X1 U13865 ( .A1(n11943), .A2(n12441), .ZN(n11066) );
  NOR2_X1 U13866 ( .A1(n11066), .A2(n11065), .ZN(n11068) );
  MUX2_X1 U13867 ( .A(n19505), .B(n19913), .S(n11495), .Z(n11071) );
  INV_X1 U13869 ( .A(n11198), .ZN(n11072) );
  AND2_X1 U13870 ( .A1(n11072), .A2(n20539), .ZN(n12252) );
  AOI21_X1 U13871 ( .B1(n10745), .B2(n11210), .A(n11483), .ZN(n11075) );
  NAND2_X1 U13872 ( .A1(n11073), .A2(n3500), .ZN(n11074) );
  NAND2_X1 U13874 ( .A1(n12250), .A2(n20153), .ZN(n12570) );
  INV_X1 U13875 ( .A(n12570), .ZN(n13144) );
  INV_X1 U13876 ( .A(n11076), .ZN(n11218) );
  NAND2_X1 U13877 ( .A1(n11218), .A2(n204), .ZN(n11077) );
  NAND2_X1 U13878 ( .A1(n11475), .A2(n11219), .ZN(n11078) );
  INV_X1 U13879 ( .A(n12253), .ZN(n13145) );
  NOR2_X1 U13880 ( .A1(n11501), .A2(n11193), .ZN(n11505) );
  NOR2_X1 U13881 ( .A1(n11193), .A2(n11500), .ZN(n11081) );
  INV_X1 U13882 ( .A(n11193), .ZN(n11187) );
  INV_X1 U13883 ( .A(n11186), .ZN(n11503) );
  MUX2_X1 U13884 ( .A(n11083), .B(n11082), .S(n11501), .Z(n11084) );
  NAND2_X1 U13886 ( .A1(n11112), .A2(n11458), .ZN(n11086) );
  INV_X1 U13887 ( .A(n11452), .ZN(n11089) );
  OAI22_X1 U13888 ( .A1(n11089), .A2(n11110), .B1(n11455), .B2(n11454), .ZN(
        n11090) );
  NOR2_X1 U13889 ( .A1(n13147), .A2(n12255), .ZN(n11092) );
  OAI21_X1 U13890 ( .B1(n13146), .B2(n13145), .A(n11092), .ZN(n11099) );
  NAND3_X1 U13891 ( .A1(n11209), .A2(n11201), .A3(n11094), .ZN(n11096) );
  NAND3_X1 U13892 ( .A1(n11445), .A2(n11202), .A3(n11444), .ZN(n11095) );
  NAND4_X1 U13893 ( .A1(n11097), .A2(n11448), .A3(n11096), .A4(n11095), .ZN(
        n12254) );
  INV_X1 U13894 ( .A(n12254), .ZN(n13141) );
  OAI21_X1 U13895 ( .B1(n13141), .B2(n12258), .A(n13147), .ZN(n11098) );
  XNOR2_X1 U13896 ( .A(n13319), .B(n13280), .ZN(n11100) );
  XNOR2_X1 U13897 ( .A(n11101), .B(n11100), .ZN(n11102) );
  INV_X1 U13898 ( .A(n14780), .ZN(n14077) );
  NOR2_X1 U13899 ( .A1(n14077), .A2(n20518), .ZN(n11319) );
  NOR2_X1 U13901 ( .A1(n11106), .A2(n11105), .ZN(n11107) );
  NAND2_X1 U13902 ( .A1(n11452), .A2(n11110), .ZN(n11111) );
  NAND2_X1 U13903 ( .A1(n12138), .A2(n12137), .ZN(n11139) );
  AND2_X1 U13904 ( .A1(n11120), .A2(n11880), .ZN(n11121) );
  OAI21_X1 U13905 ( .B1(n11121), .B2(n11883), .A(n85), .ZN(n11123) );
  NAND2_X1 U13906 ( .A1(n11121), .A2(n909), .ZN(n11122) );
  NAND3_X1 U13907 ( .A1(n12470), .A2(n11915), .A3(n12137), .ZN(n11138) );
  NAND2_X1 U13908 ( .A1(n20099), .A2(n11125), .ZN(n11126) );
  NAND3_X1 U13909 ( .A1(n205), .A2(n19837), .A3(n11131), .ZN(n11135) );
  NOR2_X1 U13910 ( .A1(n12463), .A2(n12386), .ZN(n11136) );
  NAND2_X1 U13911 ( .A1(n12470), .A2(n11136), .ZN(n11137) );
  INV_X1 U13912 ( .A(n12281), .ZN(n11167) );
  OAI21_X1 U13913 ( .B1(n11148), .B2(n11147), .A(n11149), .ZN(n11154) );
  NAND2_X1 U13914 ( .A1(n20470), .A2(n11149), .ZN(n11151) );
  NAND2_X1 U13916 ( .A1(n11557), .A2(n11559), .ZN(n11554) );
  OR2_X1 U13917 ( .A1(n11554), .A2(n20479), .ZN(n11165) );
  NAND2_X1 U13918 ( .A1(n19564), .A2(n10968), .ZN(n11555) );
  OAI211_X1 U13919 ( .C1(n11163), .C2(n20479), .A(n10913), .B(n11162), .ZN(
        n11164) );
  AND3_X1 U13920 ( .A1(n11555), .A2(n11165), .A3(n11164), .ZN(n12279) );
  NAND2_X1 U13921 ( .A1(n11717), .A2(n12279), .ZN(n12044) );
  INV_X1 U13922 ( .A(n12044), .ZN(n11166) );
  OAI21_X1 U13923 ( .B1(n11167), .B2(n12040), .A(n11166), .ZN(n11181) );
  NAND2_X1 U13924 ( .A1(n11171), .A2(n11532), .ZN(n12035) );
  INV_X1 U13925 ( .A(n12035), .ZN(n11172) );
  INV_X1 U13926 ( .A(n12279), .ZN(n12042) );
  AOI21_X1 U13927 ( .B1(n12282), .B2(n12042), .A(n12040), .ZN(n11180) );
  NOR2_X1 U13928 ( .A1(n11176), .A2(n11175), .ZN(n11179) );
  AND2_X1 U13929 ( .A1(n12040), .A2(n12041), .ZN(n11775) );
  XNOR2_X1 U13930 ( .A(n13330), .B(n13833), .ZN(n11229) );
  INV_X1 U13931 ( .A(n11182), .ZN(n11183) );
  OAI22_X1 U13932 ( .A1(n11183), .A2(n11564), .B1(n11566), .B2(n11469), .ZN(
        n11184) );
  NAND2_X1 U13933 ( .A1(n11184), .A2(n11567), .ZN(n11185) );
  NOR2_X1 U13935 ( .A1(n11500), .A2(n11188), .ZN(n11189) );
  MUX2_X1 U13937 ( .A(n11193), .B(n11192), .S(n11191), .Z(n11194) );
  AOI21_X1 U13938 ( .B1(n11446), .B2(n19920), .A(n11202), .ZN(n11207) );
  INV_X1 U13939 ( .A(n11203), .ZN(n11206) );
  INV_X1 U13940 ( .A(n11204), .ZN(n11205) );
  OAI21_X1 U13941 ( .B1(n11207), .B2(n11206), .A(n11205), .ZN(n11208) );
  NAND2_X1 U13942 ( .A1(n11708), .A2(n12394), .ZN(n12785) );
  INV_X1 U13943 ( .A(n12785), .ZN(n11225) );
  NAND2_X1 U13944 ( .A1(n3500), .A2(n11482), .ZN(n11213) );
  NAND2_X1 U13945 ( .A1(n11481), .A2(n11483), .ZN(n11212) );
  MUX2_X1 U13946 ( .A(n11213), .B(n11212), .S(n19897), .Z(n11214) );
  NAND2_X1 U13947 ( .A1(n11217), .A2(n11475), .ZN(n11221) );
  OAI211_X1 U13948 ( .C1(n11474), .C2(n11222), .A(n11221), .B(n11220), .ZN(
        n11930) );
  BUF_X2 U13949 ( .A(n11930), .Z(n12473) );
  NOR2_X1 U13950 ( .A1(n12478), .A2(n12473), .ZN(n11223) );
  INV_X1 U13951 ( .A(n12784), .ZN(n11224) );
  OAI21_X1 U13952 ( .B1(n11225), .B2(n11224), .A(n18355), .ZN(n11227) );
  NAND3_X1 U13953 ( .A1(n12785), .A2(n621), .A3(n12784), .ZN(n11226) );
  NAND2_X1 U13954 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  XNOR2_X1 U13955 ( .A(n11229), .B(n11228), .ZN(n11318) );
  NOR2_X1 U13956 ( .A1(n9883), .A2(n11231), .ZN(n11232) );
  NOR2_X1 U13957 ( .A1(n11235), .A2(n11234), .ZN(n11243) );
  NAND2_X1 U13958 ( .A1(n11237), .A2(n11236), .ZN(n11242) );
  OAI21_X1 U13959 ( .B1(n11239), .B2(n10798), .A(n11238), .ZN(n11241) );
  NOR2_X1 U13960 ( .A1(n12381), .A2(n20191), .ZN(n11270) );
  NOR2_X1 U13961 ( .A1(n20191), .A2(n11243), .ZN(n11251) );
  AOI21_X1 U13962 ( .B1(n11373), .B2(n11244), .A(n11376), .ZN(n11246) );
  NOR2_X1 U13963 ( .A1(n2861), .A2(n11330), .ZN(n11245) );
  MUX2_X1 U13964 ( .A(n11246), .B(n11245), .S(n11377), .Z(n11248) );
  INV_X1 U13965 ( .A(n11375), .ZN(n11247) );
  MUX2_X1 U13966 ( .A(n11381), .B(n11271), .S(n11380), .Z(n11250) );
  AOI22_X1 U13967 ( .A1(n11252), .A2(n11251), .B1(n12269), .B2(n20497), .ZN(
        n12271) );
  NAND2_X1 U13969 ( .A1(n11253), .A2(n11255), .ZN(n11258) );
  INV_X1 U13970 ( .A(n11258), .ZN(n11262) );
  OAI21_X1 U13971 ( .B1(n11321), .B2(n11255), .A(n11254), .ZN(n11261) );
  NAND2_X1 U13972 ( .A1(n191), .A2(n11256), .ZN(n11259) );
  MUX2_X1 U13973 ( .A(n11259), .B(n11258), .S(n11257), .Z(n11260) );
  NOR2_X1 U13974 ( .A1(n11267), .A2(n11263), .ZN(n11336) );
  OAI21_X1 U13975 ( .B1(n11343), .B2(n11264), .A(n11337), .ZN(n11268) );
  AND2_X1 U13976 ( .A1(n11339), .A2(n9830), .ZN(n11335) );
  OAI21_X1 U13977 ( .B1(n12369), .B2(n12373), .A(n12377), .ZN(n11269) );
  OAI21_X1 U13978 ( .B1(n11270), .B2(n12271), .A(n11269), .ZN(n13120) );
  NAND2_X1 U13979 ( .A1(n11276), .A2(n11410), .ZN(n11280) );
  OAI211_X1 U13980 ( .C1(n11411), .C2(n11278), .A(n11408), .B(n11277), .ZN(
        n11279) );
  OAI21_X1 U13982 ( .B1(n11284), .B2(n9559), .A(n11283), .ZN(n11285) );
  OAI21_X1 U13983 ( .B1(n11287), .B2(n11286), .A(n11285), .ZN(n11288) );
  MUX2_X1 U13984 ( .A(n11296), .B(n11399), .S(n11295), .Z(n11301) );
  NAND2_X1 U13985 ( .A1(n11297), .A2(n11399), .ZN(n11299) );
  NAND2_X1 U13986 ( .A1(n11394), .A2(n11398), .ZN(n11298) );
  MUX2_X1 U13987 ( .A(n11299), .B(n11298), .S(n11395), .Z(n11300) );
  INV_X1 U13988 ( .A(n12488), .ZN(n12812) );
  NAND2_X1 U13989 ( .A1(n11303), .A2(n11302), .ZN(n11309) );
  NAND3_X1 U13990 ( .A1(n11305), .A2(n11388), .A3(n11304), .ZN(n11308) );
  NAND3_X1 U13991 ( .A1(n20517), .A2(n11867), .A3(n20601), .ZN(n11307) );
  OAI211_X1 U13992 ( .C1(n12399), .C2(n12807), .A(n12812), .B(n12487), .ZN(
        n11310) );
  OAI211_X1 U13993 ( .C1(n12807), .C2(n11693), .A(n11911), .B(n11310), .ZN(
        n13431) );
  XNOR2_X1 U13994 ( .A(n13120), .B(n13431), .ZN(n13329) );
  INV_X1 U13995 ( .A(n13329), .ZN(n11316) );
  NOR2_X1 U13996 ( .A1(n12754), .A2(n12759), .ZN(n12757) );
  OAI21_X1 U13997 ( .B1(n11315), .B2(n12757), .A(n11314), .ZN(n13079) );
  XNOR2_X1 U13998 ( .A(n13031), .B(n13079), .ZN(n11965) );
  XNOR2_X1 U13999 ( .A(n11316), .B(n11965), .ZN(n11317) );
  AOI22_X1 U14002 ( .A1(n191), .A2(n11324), .B1(n11323), .B2(n11327), .ZN(
        n11326) );
  INV_X1 U14003 ( .A(n11709), .ZN(n12311) );
  OAI21_X1 U14004 ( .B1(n11331), .B2(n2611), .A(n2861), .ZN(n11334) );
  MUX2_X1 U14005 ( .A(n11330), .B(n11329), .S(n11332), .Z(n11333) );
  NAND2_X1 U14006 ( .A1(n12311), .A2(n20486), .ZN(n11363) );
  NAND2_X1 U14007 ( .A1(n11341), .A2(n11340), .ZN(n11342) );
  AOI21_X1 U14008 ( .B1(n11343), .B2(n11265), .A(n11342), .ZN(n11344) );
  MUX2_X1 U14009 ( .A(n11347), .B(n11348), .S(n11346), .Z(n11354) );
  NAND2_X1 U14011 ( .A1(n11355), .A2(n11239), .ZN(n11351) );
  MUX2_X1 U14012 ( .A(n11352), .B(n11351), .S(n11350), .Z(n11353) );
  NAND2_X1 U14013 ( .A1(n11358), .A2(n19949), .ZN(n11361) );
  NAND2_X1 U14014 ( .A1(n11367), .A2(n11366), .ZN(n11368) );
  MUX2_X1 U14015 ( .A(n12312), .B(n12148), .S(n19952), .Z(n11370) );
  NOR2_X1 U14016 ( .A1(n11370), .A2(n12311), .ZN(n11371) );
  INV_X1 U14017 ( .A(n13099), .ZN(n11416) );
  NAND2_X1 U14018 ( .A1(n202), .A2(n11377), .ZN(n11374) );
  NAND2_X1 U14019 ( .A1(n11377), .A2(n11376), .ZN(n11379) );
  AOI21_X1 U14020 ( .B1(n11379), .B2(n202), .A(n11378), .ZN(n12548) );
  NOR2_X1 U14022 ( .A1(n12542), .A2(n12543), .ZN(n12310) );
  INV_X1 U14023 ( .A(n11385), .ZN(n11386) );
  NAND2_X1 U14025 ( .A1(n11388), .A2(n11870), .ZN(n11392) );
  MUX2_X1 U14026 ( .A(n20517), .B(n11866), .S(n11389), .Z(n11391) );
  MUX2_X1 U14027 ( .A(n11399), .B(n11397), .S(n11394), .Z(n11396) );
  NAND3_X1 U14028 ( .A1(n11399), .A2(n11398), .A3(n11397), .ZN(n11400) );
  NOR2_X1 U14029 ( .A1(n10978), .A2(n11405), .ZN(n11407) );
  AOI22_X1 U14030 ( .A1(n12310), .A2(n2160), .B1(n11795), .B2(n12305), .ZN(
        n11415) );
  INV_X1 U14031 ( .A(n11411), .ZN(n11412) );
  AND2_X1 U14032 ( .A1(n11413), .A2(n937), .ZN(n12549) );
  NAND2_X1 U14033 ( .A1(n11415), .A2(n11414), .ZN(n13756) );
  XNOR2_X1 U14034 ( .A(n11416), .B(n13756), .ZN(n13347) );
  NAND2_X1 U14035 ( .A1(n11419), .A2(n1680), .ZN(n11422) );
  INV_X1 U14036 ( .A(n12524), .ZN(n12165) );
  AOI21_X1 U14037 ( .B1(n11425), .B2(n11424), .A(n19830), .ZN(n11434) );
  NOR2_X1 U14038 ( .A1(n11427), .A2(n1378), .ZN(n11433) );
  OAI211_X1 U14039 ( .C1(n19830), .C2(n11430), .A(n11429), .B(n11428), .ZN(
        n11432) );
  INV_X1 U14041 ( .A(n12167), .ZN(n12520) );
  MUX2_X1 U14042 ( .A(n11438), .B(n11436), .S(n11435), .Z(n11442) );
  NAND2_X1 U14043 ( .A1(n11445), .A2(n11444), .ZN(n11447) );
  NAND3_X1 U14044 ( .A1(n11456), .A2(n11455), .A3(n11454), .ZN(n11457) );
  MUX2_X1 U14045 ( .A(n11883), .B(n11880), .S(n11884), .Z(n11463) );
  INV_X1 U14046 ( .A(n12168), .ZN(n11464) );
  NAND2_X1 U14047 ( .A1(n898), .A2(n11469), .ZN(n11468) );
  NAND2_X1 U14048 ( .A1(n11467), .A2(n11466), .ZN(n11471) );
  MUX2_X1 U14049 ( .A(n11468), .B(n11471), .S(n11568), .Z(n11473) );
  NAND2_X1 U14050 ( .A1(n11471), .A2(n11470), .ZN(n11472) );
  OAI211_X1 U14051 ( .C1(n11481), .C2(n11480), .A(n11486), .B(n11479), .ZN(
        n11485) );
  NAND3_X1 U14052 ( .A1(n11483), .A2(n20233), .A3(n11482), .ZN(n11484) );
  OAI211_X2 U14053 ( .C1(n11486), .C2(n11487), .A(n11485), .B(n11484), .ZN(
        n12534) );
  NAND2_X1 U14054 ( .A1(n19719), .A2(n3051), .ZN(n11490) );
  NAND2_X1 U14055 ( .A1(n20539), .A2(n11493), .ZN(n11497) );
  NOR2_X1 U14056 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  NAND2_X1 U14057 ( .A1(n11500), .A2(n11499), .ZN(n11504) );
  MUX2_X1 U14058 ( .A(n11504), .B(n11502), .S(n11501), .Z(n11508) );
  NOR2_X1 U14059 ( .A1(n11504), .A2(n11503), .ZN(n11506) );
  NOR2_X1 U14060 ( .A1(n11506), .A2(n11505), .ZN(n11507) );
  NAND2_X1 U14061 ( .A1(n11508), .A2(n11507), .ZN(n12532) );
  MUX2_X1 U14062 ( .A(n12535), .B(n243), .S(n12534), .Z(n11519) );
  NAND2_X1 U14063 ( .A1(n11512), .A2(n20639), .ZN(n11518) );
  XNOR2_X1 U14065 ( .A(n13569), .B(n13347), .ZN(n11593) );
  NOR2_X1 U14066 ( .A1(n11528), .A2(n11521), .ZN(n11525) );
  NOR2_X1 U14067 ( .A1(n11522), .A2(n11527), .ZN(n11524) );
  NAND3_X1 U14068 ( .A1(n11528), .A2(n11527), .A3(n11526), .ZN(n11529) );
  OAI21_X1 U14069 ( .B1(n11531), .B2(n11530), .A(n11529), .ZN(n11742) );
  NOR2_X2 U14070 ( .A1(n11741), .A2(n11742), .ZN(n12299) );
  NAND2_X1 U14072 ( .A1(n731), .A2(n11538), .ZN(n11541) );
  MUX2_X1 U14074 ( .A(n11549), .B(n11548), .S(n11547), .Z(n11551) );
  AOI21_X1 U14076 ( .B1(n11555), .B2(n11554), .A(n11553), .ZN(n11562) );
  NAND2_X1 U14077 ( .A1(n11557), .A2(n11556), .ZN(n11560) );
  AOI21_X1 U14078 ( .B1(n11560), .B2(n11559), .A(n19564), .ZN(n11561) );
  INV_X1 U14079 ( .A(n11563), .ZN(n12304) );
  NOR2_X1 U14080 ( .A1(n12299), .A2(n11782), .ZN(n11739) );
  AOI21_X1 U14081 ( .B1(n11565), .B2(n11564), .A(n927), .ZN(n11744) );
  NAND2_X1 U14082 ( .A1(n11567), .A2(n927), .ZN(n11571) );
  NAND2_X1 U14083 ( .A1(n11569), .A2(n11568), .ZN(n11570) );
  AOI21_X1 U14084 ( .B1(n11571), .B2(n11570), .A(n898), .ZN(n11740) );
  AND2_X1 U14085 ( .A1(n12304), .A2(n12274), .ZN(n11578) );
  INV_X1 U14086 ( .A(n12033), .ZN(n11577) );
  INV_X1 U14087 ( .A(n13063), .ZN(n11585) );
  NAND2_X1 U14088 ( .A1(n12281), .A2(n12041), .ZN(n11581) );
  AND2_X1 U14089 ( .A1(n11580), .A2(n11581), .ZN(n11584) );
  OAI21_X1 U14090 ( .B1(n11582), .B2(n11776), .A(n12278), .ZN(n11583) );
  XNOR2_X1 U14091 ( .A(n11585), .B(n12863), .ZN(n11862) );
  INV_X1 U14092 ( .A(n12128), .ZN(n11642) );
  OAI21_X1 U14093 ( .B1(n882), .B2(n12126), .A(n12130), .ZN(n11588) );
  INV_X1 U14094 ( .A(n11586), .ZN(n11763) );
  NAND2_X1 U14095 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  XNOR2_X1 U14096 ( .A(n13425), .B(n1840), .ZN(n11591) );
  XNOR2_X1 U14097 ( .A(n11862), .B(n11591), .ZN(n11592) );
  NAND2_X1 U14098 ( .A1(n14216), .A2(n14781), .ZN(n14852) );
  INV_X1 U14099 ( .A(n14852), .ZN(n11594) );
  AND2_X1 U14100 ( .A1(n12408), .A2(n12389), .ZN(n12756) );
  NOR2_X1 U14101 ( .A1(n12409), .A2(n12759), .ZN(n11595) );
  NOR2_X1 U14102 ( .A1(n12389), .A2(n12407), .ZN(n12755) );
  XNOR2_X1 U14103 ( .A(n19792), .B(n19027), .ZN(n11609) );
  INV_X1 U14104 ( .A(n11951), .ZN(n11955) );
  INV_X1 U14105 ( .A(n11659), .ZN(n11600) );
  NAND3_X1 U14106 ( .A1(n11955), .A2(n1578), .A3(n11600), .ZN(n11601) );
  NOR2_X1 U14107 ( .A1(n11602), .A2(n20351), .ZN(n12082) );
  NAND2_X1 U14110 ( .A1(n11605), .A2(n12084), .ZN(n11606) );
  XNOR2_X1 U14111 ( .A(n13368), .B(n13277), .ZN(n13582) );
  XNOR2_X1 U14112 ( .A(n13582), .B(n11609), .ZN(n11626) );
  NAND2_X1 U14114 ( .A1(n12684), .A2(n12648), .ZN(n11610) );
  MUX2_X1 U14115 ( .A(n11611), .B(n11610), .S(n12686), .Z(n11612) );
  INV_X1 U14116 ( .A(n13707), .ZN(n13019) );
  INV_X1 U14117 ( .A(n12449), .ZN(n12635) );
  NAND2_X1 U14118 ( .A1(n11948), .A2(n12642), .ZN(n11617) );
  INV_X1 U14119 ( .A(n12455), .ZN(n12640) );
  NOR2_X1 U14120 ( .A1(n12640), .A2(n12635), .ZN(n11616) );
  NAND3_X1 U14121 ( .A1(n20458), .A2(n2256), .A3(n12450), .ZN(n11615) );
  NAND2_X1 U14122 ( .A1(n12637), .A2(n12452), .ZN(n11614) );
  XNOR2_X1 U14124 ( .A(n13019), .B(n13774), .ZN(n13233) );
  NOR2_X1 U14125 ( .A1(n12634), .A2(n11618), .ZN(n11620) );
  NAND2_X1 U14126 ( .A1(n11618), .A2(n12630), .ZN(n11619) );
  MUX2_X1 U14127 ( .A(n11942), .B(n12437), .S(n12440), .Z(n11624) );
  NOR2_X1 U14128 ( .A1(n12440), .A2(n11942), .ZN(n11623) );
  XNOR2_X1 U14129 ( .A(n13706), .B(n13776), .ZN(n13475) );
  XNOR2_X1 U14130 ( .A(n13233), .B(n13475), .ZN(n11625) );
  AOI21_X1 U14131 ( .B1(n12603), .B2(n12237), .A(n12072), .ZN(n11631) );
  INV_X1 U14132 ( .A(n11628), .ZN(n11629) );
  NAND2_X1 U14133 ( .A1(n12242), .A2(n12240), .ZN(n12054) );
  INV_X1 U14134 ( .A(n12054), .ZN(n11635) );
  INV_X1 U14135 ( .A(n12616), .ZN(n12059) );
  XNOR2_X1 U14136 ( .A(n12986), .B(n13734), .ZN(n11641) );
  INV_X1 U14137 ( .A(n12201), .ZN(n12593) );
  INV_X1 U14138 ( .A(n12200), .ZN(n12592) );
  OAI211_X1 U14139 ( .C1(n11637), .C2(n12593), .A(n193), .B(n12592), .ZN(
        n11636) );
  OAI211_X1 U14140 ( .C1(n11978), .C2(n11637), .A(n11636), .B(n11979), .ZN(
        n13029) );
  NOR2_X1 U14141 ( .A1(n12211), .A2(n19726), .ZN(n12214) );
  XNOR2_X1 U14142 ( .A(n13029), .B(n11640), .ZN(n13237) );
  XNOR2_X1 U14143 ( .A(n11641), .B(n13237), .ZN(n11655) );
  NAND2_X1 U14144 ( .A1(n12129), .A2(n12128), .ZN(n11702) );
  OR2_X1 U14145 ( .A1(n11702), .A2(n12126), .ZN(n11645) );
  NAND4_X1 U14146 ( .A1(n11703), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n12671) );
  INV_X1 U14147 ( .A(n12671), .ZN(n13391) );
  NAND2_X1 U14148 ( .A1(n12121), .A2(n12230), .ZN(n12049) );
  INV_X1 U14150 ( .A(n12232), .ZN(n11646) );
  OAI21_X1 U14151 ( .B1(n12049), .B2(n19694), .A(n11648), .ZN(n13484) );
  XNOR2_X1 U14152 ( .A(n13391), .B(n13484), .ZN(n13612) );
  NOR2_X1 U14153 ( .A1(n12180), .A2(n256), .ZN(n11652) );
  NAND2_X1 U14154 ( .A1(n11841), .A2(n20427), .ZN(n11651) );
  XNOR2_X1 U14155 ( .A(n13612), .B(n11653), .ZN(n11654) );
  XNOR2_X1 U14156 ( .A(n11654), .B(n11655), .ZN(n14806) );
  NOR2_X1 U14158 ( .A1(n11828), .A2(n11829), .ZN(n11657) );
  MUX2_X1 U14159 ( .A(n11659), .B(n11830), .S(n11829), .Z(n11660) );
  INV_X1 U14160 ( .A(n13134), .ZN(n12087) );
  XNOR2_X1 U14161 ( .A(n12087), .B(n13572), .ZN(n13464) );
  MUX2_X1 U14162 ( .A(n12008), .B(n12509), .S(n12506), .Z(n11663) );
  INV_X1 U14163 ( .A(n12359), .ZN(n11661) );
  NAND2_X1 U14165 ( .A1(n11992), .A2(n965), .ZN(n11664) );
  XNOR2_X1 U14166 ( .A(n12940), .B(n13651), .ZN(n13243) );
  NAND2_X1 U14167 ( .A1(n11841), .A2(n11670), .ZN(n11671) );
  MUX2_X1 U14168 ( .A(n12179), .B(n11673), .S(n12180), .Z(n11675) );
  MUX2_X1 U14169 ( .A(n12514), .B(n11997), .S(n11995), .Z(n11677) );
  XNOR2_X1 U14170 ( .A(n13397), .B(n13687), .ZN(n11681) );
  MUX2_X1 U14171 ( .A(n201), .B(n12499), .S(n12004), .Z(n11679) );
  XNOR2_X1 U14172 ( .A(n12979), .B(n19243), .ZN(n11680) );
  XNOR2_X1 U14173 ( .A(n11681), .B(n11680), .ZN(n11682) );
  INV_X1 U14174 ( .A(n14806), .ZN(n14811) );
  NAND2_X1 U14175 ( .A1(n11863), .A2(n11922), .ZN(n12578) );
  INV_X1 U14176 ( .A(n12578), .ZN(n11685) );
  NOR2_X1 U14177 ( .A1(n11926), .A2(n12577), .ZN(n11684) );
  NAND2_X1 U14179 ( .A1(n11686), .A2(n11922), .ZN(n11865) );
  INV_X1 U14180 ( .A(n11863), .ZN(n11923) );
  NAND2_X1 U14181 ( .A1(n11865), .A2(n11863), .ZN(n11687) );
  NAND2_X1 U14182 ( .A1(n11687), .A2(n11926), .ZN(n11688) );
  OAI21_X1 U14183 ( .B1(n12229), .B2(n12122), .A(n12228), .ZN(n11690) );
  NAND2_X1 U14184 ( .A1(n11690), .A2(n12121), .ZN(n11691) );
  XNOR2_X1 U14185 ( .A(n13622), .B(n13193), .ZN(n11698) );
  NAND2_X1 U14186 ( .A1(n11911), .A2(n11693), .ZN(n11696) );
  NAND2_X1 U14187 ( .A1(n12488), .A2(n12809), .ZN(n11694) );
  NAND2_X1 U14188 ( .A1(n11694), .A2(n12811), .ZN(n11695) );
  XNOR2_X1 U14189 ( .A(n13339), .B(n18433), .ZN(n11697) );
  XNOR2_X1 U14190 ( .A(n11698), .B(n11697), .ZN(n11716) );
  INV_X1 U14191 ( .A(n12386), .ZN(n12384) );
  NAND2_X1 U14192 ( .A1(n12384), .A2(n12137), .ZN(n12383) );
  INV_X1 U14193 ( .A(n12138), .ZN(n12468) );
  NOR2_X1 U14194 ( .A1(n12138), .A2(n857), .ZN(n11699) );
  OR3_X1 U14195 ( .A1(n12138), .A2(n12470), .A3(n11915), .ZN(n11700) );
  XNOR2_X1 U14198 ( .A(n13222), .B(n13623), .ZN(n11714) );
  NAND2_X1 U14199 ( .A1(n12478), .A2(n11930), .ZN(n11706) );
  NAND2_X1 U14200 ( .A1(n11706), .A2(n12142), .ZN(n11707) );
  INV_X1 U14201 ( .A(n12312), .ZN(n12154) );
  INV_X1 U14202 ( .A(n12152), .ZN(n11710) );
  AOI21_X1 U14203 ( .B1(n12153), .B2(n20186), .A(n11710), .ZN(n11713) );
  INV_X1 U14204 ( .A(n12148), .ZN(n12155) );
  OAI21_X1 U14205 ( .B1(n12148), .B2(n19952), .A(n11711), .ZN(n12315) );
  XNOR2_X1 U14206 ( .A(n13138), .B(n13048), .ZN(n13227) );
  INV_X1 U14207 ( .A(n13227), .ZN(n13727) );
  XNOR2_X1 U14208 ( .A(n13727), .B(n11714), .ZN(n11715) );
  NAND2_X1 U14210 ( .A1(n12041), .A2(n12279), .ZN(n11721) );
  OR2_X1 U14211 ( .A1(n11717), .A2(n12280), .ZN(n11777) );
  OAI21_X1 U14212 ( .B1(n12283), .B2(n11776), .A(n11777), .ZN(n11718) );
  NOR2_X1 U14213 ( .A1(n12281), .A2(n12040), .ZN(n11719) );
  NAND2_X1 U14214 ( .A1(n11719), .A2(n876), .ZN(n11720) );
  XNOR2_X1 U14215 ( .A(n13491), .B(n18170), .ZN(n11724) );
  NAND2_X1 U14216 ( .A1(n12634), .A2(n11618), .ZN(n11962) );
  NAND2_X1 U14217 ( .A1(n12630), .A2(n11722), .ZN(n11961) );
  NAND3_X1 U14218 ( .A1(n11961), .A2(n12632), .A3(n1371), .ZN(n11723) );
  XNOR2_X1 U14219 ( .A(n11724), .B(n13517), .ZN(n11729) );
  NOR2_X1 U14220 ( .A1(n12267), .A2(n12262), .ZN(n11725) );
  INV_X1 U14221 ( .A(n11726), .ZN(n11727) );
  XNOR2_X1 U14222 ( .A(n11729), .B(n13248), .ZN(n11756) );
  NAND2_X1 U14223 ( .A1(n12373), .A2(n20191), .ZN(n11855) );
  INV_X1 U14224 ( .A(n11855), .ZN(n11731) );
  INV_X1 U14225 ( .A(n11856), .ZN(n12371) );
  XNOR2_X1 U14226 ( .A(n13745), .B(n13642), .ZN(n11754) );
  INV_X1 U14227 ( .A(n13149), .ZN(n11734) );
  NAND2_X1 U14228 ( .A1(n244), .A2(n12254), .ZN(n11733) );
  NOR2_X1 U14229 ( .A1(n13146), .A2(n20153), .ZN(n11735) );
  NOR2_X1 U14230 ( .A1(n12029), .A2(n12304), .ZN(n11738) );
  INV_X1 U14231 ( .A(n12275), .ZN(n12272) );
  AOI22_X1 U14232 ( .A1(n11739), .A2(n12274), .B1(n11738), .B2(n12272), .ZN(
        n11752) );
  INV_X1 U14233 ( .A(n12299), .ZN(n12028) );
  INV_X1 U14234 ( .A(n11740), .ZN(n11749) );
  INV_X1 U14235 ( .A(n11741), .ZN(n11746) );
  INV_X1 U14236 ( .A(n11742), .ZN(n11743) );
  AND2_X1 U14237 ( .A1(n11744), .A2(n11743), .ZN(n11745) );
  NAND2_X1 U14238 ( .A1(n11746), .A2(n11745), .ZN(n11747) );
  OAI211_X1 U14239 ( .C1(n12028), .C2(n11749), .A(n11748), .B(n11747), .ZN(
        n11750) );
  NAND2_X1 U14240 ( .A1(n11750), .A2(n920), .ZN(n11751) );
  NAND2_X1 U14241 ( .A1(n11752), .A2(n11751), .ZN(n12846) );
  XNOR2_X1 U14242 ( .A(n13695), .B(n12846), .ZN(n11753) );
  XNOR2_X1 U14243 ( .A(n11754), .B(n11753), .ZN(n11755) );
  NOR2_X1 U14244 ( .A1(n14807), .A2(n14593), .ZN(n14809) );
  INV_X1 U14245 ( .A(n14593), .ZN(n14590) );
  INV_X1 U14247 ( .A(n12543), .ZN(n11757) );
  NAND2_X1 U14248 ( .A1(n11795), .A2(n12543), .ZN(n11758) );
  AOI21_X1 U14249 ( .B1(n11760), .B2(n11759), .A(n882), .ZN(n11767) );
  INV_X1 U14250 ( .A(n11761), .ZN(n11762) );
  NAND2_X1 U14251 ( .A1(n11763), .A2(n11762), .ZN(n11765) );
  NOR2_X1 U14252 ( .A1(n882), .A2(n12129), .ZN(n11764) );
  NOR2_X1 U14253 ( .A1(n11765), .A2(n11764), .ZN(n11766) );
  NOR2_X1 U14254 ( .A1(n11767), .A2(n11766), .ZN(n12077) );
  XNOR2_X1 U14255 ( .A(n13717), .B(n12077), .ZN(n13153) );
  INV_X1 U14256 ( .A(n13153), .ZN(n13499) );
  OAI21_X1 U14257 ( .B1(n11768), .B2(n12522), .A(n12525), .ZN(n11771) );
  NOR2_X1 U14258 ( .A1(n12528), .A2(n12288), .ZN(n12292) );
  NAND2_X1 U14259 ( .A1(n12165), .A2(n182), .ZN(n11770) );
  XNOR2_X1 U14260 ( .A(n19697), .B(n13255), .ZN(n13714) );
  NAND2_X1 U14261 ( .A1(n12311), .A2(n20186), .ZN(n11773) );
  NOR2_X1 U14263 ( .A1(n11777), .A2(n12281), .ZN(n11778) );
  NOR2_X1 U14264 ( .A1(n3801), .A2(n11778), .ZN(n11779) );
  XNOR2_X1 U14265 ( .A(n13601), .B(n13539), .ZN(n11787) );
  OAI211_X1 U14266 ( .C1(n12029), .C2(n11782), .A(n12028), .B(n11781), .ZN(
        n11785) );
  INV_X1 U14267 ( .A(n12029), .ZN(n12300) );
  OAI21_X1 U14268 ( .B1(n12300), .B2(n12298), .A(n12299), .ZN(n11784) );
  NOR2_X1 U14269 ( .A1(n12300), .A2(n11782), .ZN(n11783) );
  XNOR2_X1 U14270 ( .A(n13602), .B(n18284), .ZN(n11786) );
  XNOR2_X1 U14271 ( .A(n11787), .B(n11786), .ZN(n11788) );
  NOR2_X1 U14272 ( .A1(n907), .A2(n12167), .ZN(n11794) );
  INV_X1 U14273 ( .A(n11795), .ZN(n11800) );
  OAI211_X1 U14274 ( .C1(n11977), .C2(n250), .A(n11796), .B(n2160), .ZN(n11799) );
  XNOR2_X1 U14275 ( .A(n13126), .B(n13810), .ZN(n13641) );
  XNOR2_X1 U14276 ( .A(n13641), .B(n11801), .ZN(n11819) );
  INV_X1 U14277 ( .A(n12807), .ZN(n12490) );
  OAI21_X1 U14278 ( .B1(n12812), .B2(n12811), .A(n953), .ZN(n11802) );
  NAND2_X1 U14279 ( .A1(n12811), .A2(n12809), .ZN(n12397) );
  MUX2_X1 U14280 ( .A(n12490), .B(n11802), .S(n12397), .Z(n11803) );
  INV_X1 U14282 ( .A(n13519), .ZN(n11816) );
  NAND3_X1 U14283 ( .A1(n11810), .A2(n11809), .A3(n11808), .ZN(n11812) );
  INV_X1 U14284 ( .A(n12209), .ZN(n12213) );
  OAI21_X1 U14285 ( .B1(n11812), .B2(n11811), .A(n2428), .ZN(n11815) );
  NAND3_X1 U14286 ( .A1(n12209), .A2(n12206), .A3(n19726), .ZN(n11813) );
  OAI211_X2 U14287 ( .C1(n11815), .C2(n12065), .A(n11814), .B(n11813), .ZN(
        n13351) );
  XNOR2_X1 U14288 ( .A(n13351), .B(n11816), .ZN(n13447) );
  INV_X1 U14289 ( .A(n13447), .ZN(n13375) );
  XNOR2_X1 U14290 ( .A(n13375), .B(n11817), .ZN(n11818) );
  INV_X1 U14291 ( .A(n12513), .ZN(n11996) );
  NAND2_X1 U14292 ( .A1(n13275), .A2(n11820), .ZN(n11822) );
  NAND2_X1 U14293 ( .A1(n12514), .A2(n11995), .ZN(n11821) );
  OAI21_X1 U14294 ( .B1(n11996), .B2(n11995), .A(n11823), .ZN(n13404) );
  AOI21_X1 U14295 ( .B1(n12339), .B2(n11990), .A(n11992), .ZN(n11826) );
  NAND3_X1 U14296 ( .A1(n12338), .A2(n11974), .A3(n12335), .ZN(n11825) );
  OAI211_X1 U14297 ( .C1(n12338), .C2(n11826), .A(n11825), .B(n11824), .ZN(
        n13108) );
  XNOR2_X1 U14298 ( .A(n13404), .B(n13108), .ZN(n13440) );
  NOR2_X1 U14299 ( .A1(n11827), .A2(n11829), .ZN(n11833) );
  OAI21_X1 U14300 ( .B1(n11952), .B2(n11828), .A(n11951), .ZN(n11832) );
  NAND2_X1 U14301 ( .A1(n12509), .A2(n12009), .ZN(n11836) );
  NAND2_X1 U14302 ( .A1(n12008), .A2(n11836), .ZN(n11838) );
  NAND2_X1 U14303 ( .A1(n12507), .A2(n12508), .ZN(n11837) );
  NAND2_X1 U14304 ( .A1(n11838), .A2(n11837), .ZN(n11839) );
  NAND2_X1 U14305 ( .A1(n11840), .A2(n11839), .ZN(n13405) );
  XNOR2_X1 U14306 ( .A(n13843), .B(n13405), .ZN(n12993) );
  NAND2_X1 U14307 ( .A1(n252), .A2(n256), .ZN(n11842) );
  AOI21_X1 U14308 ( .B1(n11843), .B2(n11842), .A(n12181), .ZN(n11848) );
  INV_X1 U14309 ( .A(n11844), .ZN(n11846) );
  OAI21_X1 U14310 ( .B1(n11846), .B2(n252), .A(n11845), .ZN(n11847) );
  XNOR2_X1 U14311 ( .A(n13409), .B(n13711), .ZN(n11850) );
  XNOR2_X1 U14312 ( .A(n13715), .B(n18075), .ZN(n11849) );
  XNOR2_X1 U14313 ( .A(n11850), .B(n11849), .ZN(n11851) );
  AND2_X1 U14314 ( .A1(n12374), .A2(n20191), .ZN(n11853) );
  NAND2_X1 U14315 ( .A1(n12381), .A2(n11853), .ZN(n11854) );
  OAI21_X1 U14316 ( .B1(n12381), .B2(n11855), .A(n11854), .ZN(n11858) );
  NOR2_X1 U14317 ( .A1(n13147), .A2(n13141), .ZN(n12251) );
  INV_X1 U14318 ( .A(n12251), .ZN(n11860) );
  AOI21_X1 U14319 ( .B1(n13147), .B2(n12255), .A(n13145), .ZN(n11859) );
  NAND2_X1 U14320 ( .A1(n11860), .A2(n11859), .ZN(n11861) );
  NOR2_X1 U14321 ( .A1(n12258), .A2(n20153), .ZN(n12573) );
  XNOR2_X1 U14322 ( .A(n13064), .B(n12471), .ZN(n13428) );
  NAND2_X1 U14323 ( .A1(n20462), .A2(n11863), .ZN(n11864) );
  NAND2_X1 U14324 ( .A1(n11865), .A2(n11864), .ZN(n11878) );
  NAND3_X1 U14325 ( .A1(n20517), .A2(n11866), .A3(n20160), .ZN(n11873) );
  NAND2_X1 U14326 ( .A1(n11870), .A2(n11867), .ZN(n11868) );
  OAI211_X1 U14327 ( .C1(n20160), .C2(n11870), .A(n11869), .B(n11868), .ZN(
        n11872) );
  NAND3_X1 U14328 ( .A1(n11874), .A2(n11873), .A3(n11872), .ZN(n11875) );
  NAND2_X1 U14329 ( .A1(n11926), .A2(n11875), .ZN(n11876) );
  OAI21_X1 U14330 ( .B1(n20462), .B2(n11926), .A(n11876), .ZN(n11877) );
  XNOR2_X1 U14331 ( .A(n13848), .B(n345), .ZN(n11899) );
  INV_X1 U14332 ( .A(n11879), .ZN(n11890) );
  OAI21_X1 U14333 ( .B1(n11881), .B2(n11880), .A(n85), .ZN(n11889) );
  NOR2_X1 U14334 ( .A1(n11883), .A2(n85), .ZN(n11885) );
  AOI22_X1 U14335 ( .A1(n11887), .A2(n11886), .B1(n11885), .B2(n909), .ZN(
        n11888) );
  NOR3_X1 U14336 ( .A1(n11892), .A2(n11891), .A3(n12262), .ZN(n12568) );
  MUX2_X1 U14337 ( .A(n3401), .B(n12630), .S(n12631), .Z(n11897) );
  XNOR2_X1 U14338 ( .A(n13422), .B(n13686), .ZN(n11898) );
  XNOR2_X1 U14339 ( .A(n11899), .B(n11898), .ZN(n11900) );
  OAI21_X1 U14340 ( .B1(n12148), .B2(n20186), .A(n12313), .ZN(n11907) );
  NAND2_X1 U14341 ( .A1(n11709), .A2(n12312), .ZN(n11903) );
  AOI21_X1 U14343 ( .B1(n11905), .B2(n11710), .A(n11904), .ZN(n11906) );
  NOR2_X1 U14344 ( .A1(n12807), .A2(n12811), .ZN(n11909) );
  MUX2_X1 U14345 ( .A(n11910), .B(n11909), .S(n12487), .Z(n11914) );
  NOR2_X2 U14347 ( .A1(n11914), .A2(n11913), .ZN(n13230) );
  XNOR2_X1 U14348 ( .A(n12859), .B(n13230), .ZN(n13005) );
  INV_X1 U14349 ( .A(n13005), .ZN(n11929) );
  INV_X1 U14350 ( .A(n12470), .ZN(n12139) );
  NOR2_X1 U14351 ( .A1(n12139), .A2(n12463), .ZN(n11921) );
  OAI21_X1 U14352 ( .B1(n11915), .B2(n12137), .A(n12138), .ZN(n11920) );
  NAND4_X1 U14353 ( .A1(n12459), .A2(n12460), .A3(n12382), .A4(n11916), .ZN(
        n11917) );
  INV_X1 U14354 ( .A(n11918), .ZN(n11919) );
  INV_X1 U14355 ( .A(n11922), .ZN(n12574) );
  MUX2_X1 U14356 ( .A(n12577), .B(n20462), .S(n12574), .Z(n11927) );
  NAND3_X1 U14357 ( .A1(n20462), .A2(n12577), .A3(n11923), .ZN(n11925) );
  XNOR2_X1 U14358 ( .A(n20155), .B(n13453), .ZN(n11928) );
  XNOR2_X1 U14359 ( .A(n11929), .B(n11928), .ZN(n11936) );
  INV_X1 U14360 ( .A(n11930), .ZN(n12472) );
  NOR2_X1 U14361 ( .A1(n12142), .A2(n12473), .ZN(n11932) );
  XNOR2_X1 U14362 ( .A(n13058), .B(n13528), .ZN(n11934) );
  XNOR2_X1 U14363 ( .A(n13020), .B(n2341), .ZN(n11933) );
  XNOR2_X1 U14364 ( .A(n11934), .B(n11933), .ZN(n11935) );
  AOI22_X1 U14366 ( .A1(n14627), .A2(n14146), .B1(n14192), .B2(n19875), .ZN(
        n11989) );
  NOR2_X1 U14367 ( .A1(n12110), .A2(n11942), .ZN(n11937) );
  NAND2_X1 U14368 ( .A1(n11939), .A2(n12441), .ZN(n11940) );
  INV_X1 U14369 ( .A(n12093), .ZN(n11945) );
  XNOR2_X1 U14370 ( .A(n13390), .B(n12713), .ZN(n11950) );
  NAND2_X1 U14371 ( .A1(n20457), .A2(n12639), .ZN(n12088) );
  INV_X1 U14372 ( .A(n12088), .ZN(n11949) );
  OAI21_X1 U14373 ( .B1(n11949), .B2(n11948), .A(n11947), .ZN(n13121) );
  INV_X1 U14374 ( .A(n13121), .ZN(n13672) );
  XNOR2_X1 U14375 ( .A(n11950), .B(n13672), .ZN(n13436) );
  INV_X1 U14376 ( .A(n13436), .ZN(n11968) );
  NOR2_X1 U14377 ( .A1(n11952), .A2(n11951), .ZN(n11959) );
  NAND2_X1 U14378 ( .A1(n1578), .A2(n11953), .ZN(n11958) );
  XNOR2_X1 U14380 ( .A(n13736), .B(n2023), .ZN(n11964) );
  OAI211_X1 U14381 ( .C1(n11962), .C2(n12630), .A(n11961), .B(n11960), .ZN(
        n11963) );
  XNOR2_X1 U14382 ( .A(n11964), .B(n20222), .ZN(n11966) );
  XNOR2_X1 U14383 ( .A(n11966), .B(n11965), .ZN(n11967) );
  XNOR2_X2 U14384 ( .A(n11968), .B(n11967), .ZN(n14623) );
  OR2_X1 U14385 ( .A1(n12338), .A2(n3813), .ZN(n11973) );
  XNOR2_X1 U14386 ( .A(n13534), .B(n19887), .ZN(n13416) );
  XNOR2_X1 U14387 ( .A(n13416), .B(n11975), .ZN(n11987) );
  NOR2_X1 U14388 ( .A1(n250), .A2(n12305), .ZN(n11976) );
  OAI21_X1 U14389 ( .B1(n11977), .B2(n12305), .A(n12547), .ZN(n12307) );
  AOI21_X1 U14390 ( .B1(n12589), .B2(n12200), .A(n12202), .ZN(n11981) );
  XNOR2_X1 U14392 ( .A(n13103), .B(n13725), .ZN(n11985) );
  AND2_X1 U14393 ( .A1(n12616), .A2(n12615), .ZN(n12246) );
  OAI21_X1 U14394 ( .B1(n12246), .B2(n19784), .A(n12240), .ZN(n11982) );
  XNOR2_X1 U14395 ( .A(n20260), .B(n2307), .ZN(n11984) );
  XNOR2_X1 U14396 ( .A(n11985), .B(n11984), .ZN(n11986) );
  XNOR2_X1 U14397 ( .A(n11987), .B(n11986), .ZN(n14000) );
  OR2_X1 U14398 ( .A1(n12339), .A2(n11990), .ZN(n11991) );
  NAND3_X1 U14399 ( .A1(n11991), .A2(n12338), .A3(n12332), .ZN(n11994) );
  OAI21_X1 U14400 ( .B1(n13275), .B2(n12326), .A(n12322), .ZN(n12000) );
  NAND2_X1 U14401 ( .A1(n11996), .A2(n12326), .ZN(n11999) );
  NAND2_X1 U14404 ( .A1(n12352), .A2(n12349), .ZN(n12175) );
  OR2_X1 U14405 ( .A1(n12352), .A2(n12354), .ZN(n12003) );
  XNOR2_X1 U14406 ( .A(n13736), .B(n13795), .ZN(n12913) );
  OR2_X1 U14407 ( .A1(n12499), .A2(n12004), .ZN(n12346) );
  AOI21_X1 U14408 ( .B1(n12509), .B2(n12359), .A(n12009), .ZN(n12007) );
  AND2_X1 U14409 ( .A1(n12359), .A2(n12009), .ZN(n12364) );
  INV_X1 U14410 ( .A(n12508), .ZN(n12010) );
  XNOR2_X1 U14411 ( .A(n13673), .B(n2417), .ZN(n12013) );
  XNOR2_X1 U14412 ( .A(n12014), .B(n12013), .ZN(n12015) );
  INV_X1 U14413 ( .A(n14203), .ZN(n14206) );
  NAND2_X1 U14414 ( .A1(n13145), .A2(n12254), .ZN(n12017) );
  OAI21_X1 U14416 ( .B1(n12020), .B2(n12369), .A(n12381), .ZN(n12026) );
  NAND2_X1 U14417 ( .A1(n12373), .A2(n12369), .ZN(n12023) );
  NAND3_X1 U14418 ( .A1(n12376), .A2(n19504), .A3(n20191), .ZN(n12022) );
  OAI21_X1 U14419 ( .B1(n12381), .B2(n12023), .A(n12022), .ZN(n12024) );
  INV_X1 U14420 ( .A(n12024), .ZN(n12025) );
  INV_X1 U14421 ( .A(n13369), .ZN(n12027) );
  NOR2_X1 U14422 ( .A1(n12028), .A2(n12274), .ZN(n12031) );
  NOR2_X1 U14423 ( .A1(n12272), .A2(n12029), .ZN(n12030) );
  AND2_X1 U14424 ( .A1(n12304), .A2(n12273), .ZN(n12032) );
  NAND3_X1 U14425 ( .A1(n12037), .A2(n12036), .A3(n12035), .ZN(n12038) );
  OAI21_X1 U14426 ( .B1(n12039), .B2(n12038), .A(n12280), .ZN(n12046) );
  OAI21_X1 U14427 ( .B1(n12281), .B2(n876), .A(n12040), .ZN(n12045) );
  AOI21_X1 U14428 ( .B1(n12280), .B2(n12042), .A(n12041), .ZN(n12043) );
  AOI22_X2 U14429 ( .A1(n12046), .A2(n12045), .B1(n12044), .B2(n12043), .ZN(
        n13783) );
  XNOR2_X1 U14430 ( .A(n13018), .B(n13783), .ZN(n12559) );
  NAND2_X1 U14431 ( .A1(n12047), .A2(n12228), .ZN(n12120) );
  NAND3_X1 U14432 ( .A1(n12049), .A2(n12120), .A3(n12048), .ZN(n12052) );
  NAND2_X1 U14433 ( .A1(n12229), .A2(n1952), .ZN(n12051) );
  NOR3_X1 U14434 ( .A1(n1952), .A2(n12047), .A3(n12122), .ZN(n12050) );
  INV_X1 U14435 ( .A(n12615), .ZN(n12053) );
  NAND2_X1 U14436 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  NAND3_X1 U14437 ( .A1(n12057), .A2(n2053), .A3(n19756), .ZN(n12058) );
  XNOR2_X1 U14438 ( .A(n13658), .B(n13260), .ZN(n12920) );
  OAI21_X1 U14439 ( .B1(n12592), .B2(n12593), .A(n193), .ZN(n12063) );
  NOR2_X1 U14441 ( .A1(n12595), .A2(n20430), .ZN(n12062) );
  INV_X1 U14442 ( .A(n13027), .ZN(n12071) );
  INV_X1 U14443 ( .A(n12065), .ZN(n12069) );
  NOR2_X1 U14444 ( .A1(n2712), .A2(n19726), .ZN(n12066) );
  AND2_X1 U14445 ( .A1(n948), .A2(n12211), .ZN(n12189) );
  INV_X1 U14447 ( .A(n13710), .ZN(n12070) );
  XNOR2_X1 U14448 ( .A(n13206), .B(n12920), .ZN(n12081) );
  NOR2_X1 U14449 ( .A1(n19971), .A2(n12237), .ZN(n12075) );
  INV_X1 U14450 ( .A(n12601), .ZN(n12608) );
  INV_X1 U14451 ( .A(n12077), .ZN(n13772) );
  XNOR2_X1 U14452 ( .A(n13772), .B(n17686), .ZN(n12078) );
  XNOR2_X1 U14453 ( .A(n12079), .B(n12078), .ZN(n12080) );
  XNOR2_X1 U14454 ( .A(n12081), .B(n12080), .ZN(n13908) );
  INV_X1 U14455 ( .A(n13908), .ZN(n12196) );
  MUX2_X1 U14456 ( .A(n14206), .B(n14612), .S(n12196), .Z(n12199) );
  XNOR2_X1 U14457 ( .A(n12087), .B(n12906), .ZN(n13754) );
  NAND2_X1 U14458 ( .A1(n12642), .A2(n20458), .ZN(n12457) );
  NAND2_X1 U14459 ( .A1(n12457), .A2(n12088), .ZN(n12092) );
  NAND2_X1 U14460 ( .A1(n12642), .A2(n19861), .ZN(n12091) );
  AOI21_X1 U14461 ( .B1(n2256), .B2(n12453), .A(n20458), .ZN(n12090) );
  AOI22_X1 U14463 ( .A1(n12095), .A2(n12094), .B1(n12093), .B2(n12684), .ZN(
        n12098) );
  NOR2_X1 U14464 ( .A1(n12684), .A2(n12686), .ZN(n12096) );
  NAND2_X1 U14465 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  XNOR2_X1 U14466 ( .A(n13065), .B(n13462), .ZN(n13218) );
  XNOR2_X1 U14467 ( .A(n13754), .B(n13218), .ZN(n12117) );
  XNOR2_X1 U14468 ( .A(n940), .B(n13427), .ZN(n12115) );
  INV_X1 U14469 ( .A(n12099), .ZN(n12438) );
  INV_X1 U14470 ( .A(n12100), .ZN(n12102) );
  NOR2_X1 U14471 ( .A1(n12102), .A2(n12101), .ZN(n12106) );
  MUX2_X1 U14472 ( .A(n12106), .B(n12105), .S(n12104), .Z(n12108) );
  NOR2_X1 U14473 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  NAND3_X1 U14474 ( .A1(n1099), .A2(n12440), .A3(n12110), .ZN(n12111) );
  XNOR2_X1 U14475 ( .A(n13398), .B(n17989), .ZN(n12114) );
  XNOR2_X1 U14476 ( .A(n12115), .B(n12114), .ZN(n12116) );
  XNOR2_X1 U14477 ( .A(n12117), .B(n12116), .ZN(n14011) );
  INV_X1 U14478 ( .A(n13745), .ZN(n12118) );
  XNOR2_X1 U14479 ( .A(n12119), .B(n12118), .ZN(n12135) );
  INV_X1 U14480 ( .A(n12120), .ZN(n12125) );
  OAI21_X1 U14481 ( .B1(n12122), .B2(n12228), .A(n12121), .ZN(n12124) );
  NOR2_X1 U14483 ( .A1(n12129), .A2(n12128), .ZN(n12131) );
  XNOR2_X1 U14484 ( .A(n12697), .B(n13250), .ZN(n12614) );
  XNOR2_X1 U14485 ( .A(n12135), .B(n12614), .ZN(n12161) );
  AOI21_X1 U14486 ( .B1(n12382), .B2(n12463), .A(n12138), .ZN(n12136) );
  OAI21_X1 U14487 ( .B1(n12470), .B2(n12382), .A(n12136), .ZN(n12140) );
  AND2_X1 U14488 ( .A1(n857), .A2(n12137), .ZN(n12466) );
  NOR2_X1 U14489 ( .A1(n12137), .A2(n12386), .ZN(n12467) );
  NAND2_X1 U14490 ( .A1(n2550), .A2(n12479), .ZN(n12145) );
  INV_X1 U14491 ( .A(n12142), .ZN(n12474) );
  NAND2_X1 U14492 ( .A1(n12478), .A2(n12474), .ZN(n12143) );
  NAND3_X1 U14493 ( .A1(n12480), .A2(n12393), .A3(n12143), .ZN(n12144) );
  NOR2_X1 U14496 ( .A1(n12148), .A2(n12147), .ZN(n12151) );
  MUX2_X1 U14498 ( .A(n12154), .B(n12153), .S(n20486), .Z(n12156) );
  NOR2_X1 U14499 ( .A1(n12156), .A2(n12155), .ZN(n12157) );
  XNOR2_X1 U14501 ( .A(n12159), .B(n13643), .ZN(n13187) );
  INV_X1 U14502 ( .A(n13187), .ZN(n12160) );
  NAND2_X1 U14504 ( .A1(n19488), .A2(n14011), .ZN(n14614) );
  NAND2_X1 U14505 ( .A1(n3811), .A2(n12537), .ZN(n12164) );
  AND2_X1 U14506 ( .A1(n12162), .A2(n12532), .ZN(n12295) );
  OAI21_X1 U14507 ( .B1(n12165), .B2(n12520), .A(n907), .ZN(n12166) );
  NOR2_X1 U14508 ( .A1(n3256), .A2(n12166), .ZN(n12171) );
  NAND2_X1 U14509 ( .A1(n12168), .A2(n12167), .ZN(n12289) );
  INV_X1 U14510 ( .A(n12289), .ZN(n12169) );
  NAND2_X1 U14511 ( .A1(n12169), .A2(n182), .ZN(n12170) );
  XNOR2_X1 U14513 ( .A(n13721), .B(n12173), .ZN(n13191) );
  INV_X1 U14514 ( .A(n13191), .ZN(n12186) );
  AND2_X1 U14515 ( .A1(n11030), .A2(n19769), .ZN(n12177) );
  INV_X1 U14516 ( .A(n12175), .ZN(n12176) );
  AOI22_X1 U14517 ( .A1(n12355), .A2(n12177), .B1(n12176), .B2(n11030), .ZN(
        n12178) );
  AOI21_X1 U14518 ( .B1(n12180), .B2(n256), .A(n12179), .ZN(n12184) );
  INV_X1 U14519 ( .A(n12745), .ZN(n12889) );
  XNOR2_X1 U14520 ( .A(n13047), .B(n12889), .ZN(n12504) );
  XNOR2_X1 U14521 ( .A(n12186), .B(n12504), .ZN(n12195) );
  AOI21_X1 U14522 ( .B1(n12188), .B2(n12187), .A(n12212), .ZN(n12190) );
  XNOR2_X1 U14523 ( .A(n13383), .B(n13725), .ZN(n12193) );
  XNOR2_X1 U14524 ( .A(n13339), .B(n2384), .ZN(n12192) );
  XNOR2_X1 U14525 ( .A(n12193), .B(n12192), .ZN(n12194) );
  XNOR2_X2 U14526 ( .A(n12195), .B(n12194), .ZN(n14611) );
  INV_X1 U14527 ( .A(n14611), .ZN(n14208) );
  NAND3_X1 U14528 ( .A1(n14614), .A2(n14208), .A3(n19488), .ZN(n12198) );
  NAND3_X1 U14529 ( .A1(n14612), .A2(n12196), .A3(n14611), .ZN(n12197) );
  NOR2_X1 U14531 ( .A1(n15474), .A2(n15769), .ZN(n15245) );
  MUX2_X1 U14532 ( .A(n12200), .B(n20430), .S(n12595), .Z(n12205) );
  NAND3_X1 U14533 ( .A1(n12209), .A2(n2712), .A3(n12208), .ZN(n12217) );
  NAND3_X1 U14534 ( .A1(n12212), .A2(n12211), .A3(n12210), .ZN(n12216) );
  NAND2_X1 U14535 ( .A1(n12214), .A2(n12213), .ZN(n12215) );
  XNOR2_X1 U14536 ( .A(n13295), .B(n2087), .ZN(n12219) );
  NAND2_X1 U14537 ( .A1(n12225), .A2(n12224), .ZN(n12231) );
  NAND2_X1 U14538 ( .A1(n12231), .A2(n12047), .ZN(n12236) );
  NAND3_X1 U14539 ( .A1(n12230), .A2(n12229), .A3(n12228), .ZN(n12234) );
  XNOR2_X1 U14540 ( .A(n13425), .B(n19869), .ZN(n13852) );
  MUX2_X1 U14541 ( .A(n12600), .B(n12601), .S(n12609), .Z(n12238) );
  OAI21_X1 U14542 ( .B1(n12616), .B2(n19784), .A(n12242), .ZN(n12618) );
  NAND2_X1 U14543 ( .A1(n12241), .A2(n12243), .ZN(n12245) );
  OAI211_X1 U14544 ( .C1(n12618), .C2(n12246), .A(n12245), .B(n12244), .ZN(
        n13688) );
  XNOR2_X1 U14545 ( .A(n13688), .B(n13755), .ZN(n12247) );
  XNOR2_X1 U14546 ( .A(n13397), .B(n12247), .ZN(n12248) );
  OAI21_X1 U14547 ( .B1(n12251), .B2(n244), .A(n12250), .ZN(n12260) );
  AOI22_X1 U14548 ( .A1(n12255), .A2(n12254), .B1(n12253), .B2(n12252), .ZN(
        n12256) );
  OAI21_X1 U14549 ( .B1(n13145), .B2(n12257), .A(n12256), .ZN(n12569) );
  OAI21_X1 U14551 ( .B1(n12563), .B2(n12562), .A(n12264), .ZN(n12265) );
  NAND2_X1 U14552 ( .A1(n12265), .A2(n248), .ZN(n12266) );
  INV_X1 U14553 ( .A(n12373), .ZN(n12370) );
  AOI21_X1 U14554 ( .B1(n12374), .B2(n12269), .A(n19504), .ZN(n12270) );
  OAI22_X1 U14555 ( .A1(n12271), .A2(n12370), .B1(n12381), .B2(n12270), .ZN(
        n13724) );
  NAND2_X1 U14556 ( .A1(n12272), .A2(n12304), .ZN(n12302) );
  NAND2_X1 U14557 ( .A1(n12274), .A2(n12273), .ZN(n12303) );
  NAND2_X1 U14558 ( .A1(n12302), .A2(n12303), .ZN(n12276) );
  XNOR2_X1 U14559 ( .A(n19883), .B(n13724), .ZN(n12277) );
  XNOR2_X1 U14560 ( .A(n13303), .B(n12277), .ZN(n12287) );
  XNOR2_X1 U14561 ( .A(n13335), .B(n12284), .ZN(n13817) );
  INV_X1 U14564 ( .A(n12522), .ZN(n12291) );
  OAI21_X1 U14565 ( .B1(n12531), .B2(n20363), .A(n12293), .ZN(n12297) );
  NAND2_X1 U14566 ( .A1(n924), .A2(n20363), .ZN(n12296) );
  XNOR2_X1 U14567 ( .A(n19946), .B(n13791), .ZN(n12957) );
  OAI211_X1 U14568 ( .C1(n12300), .C2(n12304), .A(n12299), .B(n12298), .ZN(
        n12301) );
  OAI211_X1 U14569 ( .C1(n12304), .C2(n12303), .A(n12302), .B(n12301), .ZN(
        n13328) );
  NAND2_X1 U14570 ( .A1(n250), .A2(n12305), .ZN(n12309) );
  NAND2_X1 U14571 ( .A1(n12307), .A2(n12306), .ZN(n12308) );
  OAI21_X1 U14572 ( .B1(n12310), .B2(n12309), .A(n12308), .ZN(n13735) );
  XNOR2_X1 U14573 ( .A(n13735), .B(n13328), .ZN(n13551) );
  XNOR2_X1 U14574 ( .A(n13551), .B(n12957), .ZN(n12319) );
  XNOR2_X1 U14575 ( .A(n13309), .B(n13833), .ZN(n12317) );
  XNOR2_X1 U14576 ( .A(n13391), .B(n2203), .ZN(n12316) );
  XNOR2_X1 U14577 ( .A(n12317), .B(n12316), .ZN(n12318) );
  INV_X1 U14578 ( .A(n13275), .ZN(n12324) );
  NAND2_X1 U14579 ( .A1(n13270), .A2(n13275), .ZN(n12328) );
  XNOR2_X1 U14582 ( .A(n19796), .B(n18396), .ZN(n12331) );
  XNOR2_X1 U14583 ( .A(n13368), .B(n13827), .ZN(n12330) );
  XNOR2_X1 U14584 ( .A(n12330), .B(n12331), .ZN(n12368) );
  INV_X1 U14585 ( .A(n12334), .ZN(n12336) );
  NAND2_X1 U14586 ( .A1(n12340), .A2(n12339), .ZN(n12341) );
  NOR2_X1 U14588 ( .A1(n12354), .A2(n12349), .ZN(n12351) );
  INV_X1 U14590 ( .A(n12506), .ZN(n12361) );
  NAND2_X1 U14591 ( .A1(n12508), .A2(n12359), .ZN(n12360) );
  OAI22_X1 U14592 ( .A1(n916), .A2(n12361), .B1(n12507), .B2(n12360), .ZN(
        n12366) );
  NOR3_X1 U14593 ( .A1(n12506), .A2(n12364), .A3(n3798), .ZN(n12365) );
  XNOR2_X1 U14594 ( .A(n13826), .B(n13781), .ZN(n13527) );
  NAND2_X1 U14595 ( .A1(n12370), .A2(n12369), .ZN(n12380) );
  NAND2_X1 U14596 ( .A1(n12371), .A2(n12373), .ZN(n12379) );
  AND2_X1 U14597 ( .A1(n12386), .A2(n12463), .ZN(n12387) );
  INV_X1 U14598 ( .A(n12992), .ZN(n13768) );
  AOI21_X1 U14600 ( .B1(n12754), .B2(n12409), .A(n12759), .ZN(n12392) );
  NAND2_X1 U14601 ( .A1(n12389), .A2(n12407), .ZN(n12390) );
  XNOR2_X1 U14602 ( .A(n13544), .B(n13657), .ZN(n13846) );
  XNOR2_X1 U14603 ( .A(n13282), .B(n13846), .ZN(n12406) );
  NAND2_X1 U14604 ( .A1(n12472), .A2(n12478), .ZN(n12396) );
  NAND3_X1 U14605 ( .A1(n12479), .A2(n12473), .A3(n19833), .ZN(n12395) );
  XNOR2_X1 U14606 ( .A(n13601), .B(n13259), .ZN(n12404) );
  OAI21_X1 U14607 ( .B1(n953), .B2(n12399), .A(n12807), .ZN(n12402) );
  NAND2_X1 U14608 ( .A1(n12487), .A2(n12488), .ZN(n12398) );
  AND2_X1 U14609 ( .A1(n12398), .A2(n12397), .ZN(n12401) );
  NOR2_X1 U14610 ( .A1(n253), .A2(n12809), .ZN(n12400) );
  AOI21_X1 U14611 ( .B1(n12402), .B2(n12401), .A(n12400), .ZN(n13541) );
  INV_X1 U14612 ( .A(n13541), .ZN(n13716) );
  XNOR2_X1 U14613 ( .A(n13716), .B(n2263), .ZN(n12403) );
  XNOR2_X1 U14614 ( .A(n12404), .B(n12403), .ZN(n12405) );
  XNOR2_X1 U14615 ( .A(n12406), .B(n12405), .ZN(n13891) );
  NOR2_X1 U14616 ( .A1(n12412), .A2(n12759), .ZN(n12413) );
  NOR2_X2 U14617 ( .A1(n12414), .A2(n12413), .ZN(n13251) );
  OAI21_X1 U14618 ( .B1(n12417), .B2(n12416), .A(n12415), .ZN(n12426) );
  NAND2_X1 U14619 ( .A1(n12418), .A2(n20351), .ZN(n12420) );
  OR2_X1 U14620 ( .A1(n12420), .A2(n12419), .ZN(n12425) );
  NOR2_X1 U14621 ( .A1(n12422), .A2(n20352), .ZN(n12423) );
  NAND2_X1 U14622 ( .A1(n257), .A2(n12423), .ZN(n12424) );
  OAI211_X1 U14623 ( .C1(n12427), .C2(n12426), .A(n12425), .B(n12424), .ZN(
        n13168) );
  XNOR2_X1 U14624 ( .A(n12696), .B(n13168), .ZN(n13807) );
  NOR3_X1 U14625 ( .A1(n12684), .A2(n12645), .A3(n12686), .ZN(n12432) );
  AND3_X1 U14626 ( .A1(n12684), .A2(n12430), .A3(n12429), .ZN(n12431) );
  AOI21_X1 U14627 ( .B1(n12434), .B2(n12685), .A(n12433), .ZN(n12448) );
  INV_X1 U14628 ( .A(n12435), .ZN(n12436) );
  NAND2_X1 U14629 ( .A1(n12440), .A2(n12439), .ZN(n12445) );
  MUX2_X1 U14630 ( .A(n12445), .B(n12444), .S(n12443), .Z(n12446) );
  NAND2_X1 U14631 ( .A1(n12450), .A2(n12449), .ZN(n12451) );
  NAND2_X1 U14632 ( .A1(n19861), .A2(n12453), .ZN(n12641) );
  MUX2_X1 U14633 ( .A(n20457), .B(n12454), .S(n12641), .Z(n12456) );
  XNOR2_X1 U14634 ( .A(n12458), .B(n19689), .ZN(n13291) );
  NOR2_X1 U14635 ( .A1(n14850), .A2(n14851), .ZN(n15655) );
  INV_X1 U14636 ( .A(n15655), .ZN(n15658) );
  INV_X1 U14637 ( .A(n12459), .ZN(n12462) );
  NAND2_X1 U14638 ( .A1(n12460), .A2(n991), .ZN(n12461) );
  NOR2_X1 U14639 ( .A1(n12462), .A2(n12461), .ZN(n12464) );
  AOI22_X1 U14640 ( .A1(n12465), .A2(n12464), .B1(n12463), .B2(n12137), .ZN(
        n12469) );
  INV_X1 U14641 ( .A(n12471), .ZN(n13343) );
  XNOR2_X1 U14642 ( .A(n12863), .B(n13427), .ZN(n13035) );
  XNOR2_X1 U14643 ( .A(n12864), .B(n13035), .ZN(n12496) );
  NOR2_X1 U14644 ( .A1(n12480), .A2(n12472), .ZN(n12476) );
  NOR2_X1 U14645 ( .A1(n12474), .A2(n12473), .ZN(n12475) );
  INV_X1 U14647 ( .A(n12478), .ZN(n12483) );
  NAND2_X1 U14648 ( .A1(n12480), .A2(n12479), .ZN(n12482) );
  OAI22_X1 U14649 ( .A1(n12484), .A2(n12483), .B1(n12482), .B2(n19833), .ZN(
        n12485) );
  NOR2_X2 U14650 ( .A1(n12486), .A2(n12485), .ZN(n13512) );
  XNOR2_X1 U14651 ( .A(n13512), .B(n12906), .ZN(n12494) );
  NOR2_X1 U14652 ( .A1(n953), .A2(n12487), .ZN(n12491) );
  MUX2_X1 U14653 ( .A(n12811), .B(n12488), .S(n12809), .Z(n12489) );
  XNOR2_X1 U14654 ( .A(n13396), .B(n17999), .ZN(n12493) );
  XNOR2_X1 U14655 ( .A(n12494), .B(n12493), .ZN(n12495) );
  INV_X1 U14656 ( .A(n14789), .ZN(n14343) );
  OAI21_X1 U14657 ( .B1(n12500), .B2(n12499), .A(n12498), .ZN(n12501) );
  XNOR2_X1 U14658 ( .A(n19887), .B(n13468), .ZN(n13340) );
  XNOR2_X1 U14659 ( .A(n13340), .B(n12504), .ZN(n12519) );
  OR2_X1 U14660 ( .A1(n12509), .A2(n12508), .ZN(n12511) );
  XNOR2_X1 U14661 ( .A(n13192), .B(n18854), .ZN(n12516) );
  XNOR2_X1 U14662 ( .A(n12517), .B(n12516), .ZN(n12518) );
  XNOR2_X1 U14663 ( .A(n12519), .B(n12518), .ZN(n14792) );
  NOR2_X1 U14664 ( .A1(n12523), .A2(n12520), .ZN(n12521) );
  NOR2_X1 U14665 ( .A1(n12522), .A2(n12521), .ZN(n12529) );
  NOR3_X1 U14666 ( .A1(n12524), .A2(n907), .A3(n12523), .ZN(n12527) );
  AOI211_X4 U14667 ( .C1(n12529), .C2(n3256), .A(n12527), .B(n12526), .ZN(
        n13173) );
  XNOR2_X1 U14668 ( .A(n13173), .B(n13020), .ZN(n12541) );
  INV_X1 U14669 ( .A(n12530), .ZN(n12539) );
  OAI21_X1 U14670 ( .B1(n12531), .B2(n12532), .A(n12533), .ZN(n12538) );
  NOR2_X1 U14671 ( .A1(n12534), .A2(n12533), .ZN(n12536) );
  XNOR2_X1 U14672 ( .A(n12541), .B(n12540), .ZN(n12561) );
  NAND2_X1 U14673 ( .A1(n12543), .A2(n12542), .ZN(n12546) );
  AOI21_X1 U14674 ( .B1(n12547), .B2(n12546), .A(n12555), .ZN(n12558) );
  INV_X1 U14675 ( .A(n12548), .ZN(n12550) );
  NAND2_X1 U14676 ( .A1(n12550), .A2(n3615), .ZN(n12551) );
  NOR3_X1 U14677 ( .A1(n12553), .A2(n12552), .A3(n12551), .ZN(n12556) );
  MUX2_X1 U14678 ( .A(n12556), .B(n12555), .S(n12554), .Z(n12557) );
  INV_X1 U14679 ( .A(n13451), .ZN(n13359) );
  XNOR2_X1 U14680 ( .A(n13017), .B(n13359), .ZN(n13366) );
  XNOR2_X1 U14681 ( .A(n12559), .B(n13366), .ZN(n12560) );
  INV_X1 U14682 ( .A(n14790), .ZN(n13897) );
  NAND2_X1 U14683 ( .A1(n12563), .A2(n12562), .ZN(n12567) );
  OAI21_X1 U14684 ( .B1(n12568), .B2(n12567), .A(n12566), .ZN(n13834) );
  XNOR2_X1 U14685 ( .A(n13834), .B(n13390), .ZN(n12870) );
  AND2_X1 U14687 ( .A1(n20462), .A2(n12574), .ZN(n12582) );
  NAND2_X1 U14688 ( .A1(n12576), .A2(n12577), .ZN(n12581) );
  NAND2_X1 U14689 ( .A1(n12578), .A2(n12577), .ZN(n12580) );
  AOI22_X1 U14690 ( .A1(n12582), .A2(n12581), .B1(n12580), .B2(n12579), .ZN(
        n12715) );
  INV_X1 U14691 ( .A(n12715), .ZN(n13607) );
  XNOR2_X1 U14692 ( .A(n13479), .B(n13607), .ZN(n12583) );
  XNOR2_X1 U14693 ( .A(n12870), .B(n12583), .ZN(n12588) );
  XNOR2_X1 U14694 ( .A(n13795), .B(n18819), .ZN(n12586) );
  INV_X1 U14695 ( .A(n13031), .ZN(n12584) );
  XNOR2_X1 U14696 ( .A(n12584), .B(n13677), .ZN(n12585) );
  XNOR2_X1 U14697 ( .A(n12586), .B(n12585), .ZN(n12587) );
  AOI22_X1 U14699 ( .A1(n14343), .A2(n20141), .B1(n13897), .B2(n14787), .ZN(
        n12657) );
  INV_X1 U14700 ( .A(n12596), .ZN(n12599) );
  OAI21_X1 U14701 ( .B1(n12592), .B2(n12591), .A(n12590), .ZN(n12598) );
  OAI21_X1 U14702 ( .B1(n12599), .B2(n12598), .A(n12597), .ZN(n13376) );
  NAND2_X1 U14703 ( .A1(n12601), .A2(n12600), .ZN(n12605) );
  NAND2_X1 U14704 ( .A1(n12607), .A2(n12606), .ZN(n12612) );
  NAND3_X1 U14705 ( .A1(n12610), .A2(n12609), .A3(n12608), .ZN(n12611) );
  XNOR2_X1 U14706 ( .A(n13042), .B(n13351), .ZN(n12624) );
  MUX2_X1 U14707 ( .A(n12616), .B(n12615), .S(n19784), .Z(n12622) );
  OR2_X1 U14708 ( .A1(n12618), .A2(n19784), .ZN(n12621) );
  XNOR2_X1 U14709 ( .A(n20253), .B(n2368), .ZN(n12623) );
  XNOR2_X1 U14710 ( .A(n12624), .B(n12623), .ZN(n12625) );
  NAND2_X1 U14711 ( .A1(n12627), .A2(n14791), .ZN(n14344) );
  INV_X1 U14712 ( .A(n14344), .ZN(n12655) );
  NOR2_X1 U14713 ( .A1(n3403), .A2(n20184), .ZN(n12633) );
  XNOR2_X1 U14714 ( .A(n13405), .B(n13659), .ZN(n13437) );
  INV_X1 U14715 ( .A(n13437), .ZN(n12652) );
  NAND2_X1 U14718 ( .A1(n12645), .A2(n3649), .ZN(n12651) );
  NOR2_X1 U14719 ( .A1(n12648), .A2(n12647), .ZN(n12649) );
  NAND2_X1 U14720 ( .A1(n12684), .A2(n12649), .ZN(n12650) );
  XNOR2_X1 U14721 ( .A(n20489), .B(n13543), .ZN(n13844) );
  XNOR2_X1 U14722 ( .A(n13844), .B(n12652), .ZN(n12653) );
  XNOR2_X1 U14723 ( .A(n12653), .B(n12654), .ZN(n14103) );
  INV_X1 U14727 ( .A(n14849), .ZN(n15660) );
  NAND2_X1 U14729 ( .A1(n15659), .A2(n15655), .ZN(n12660) );
  NAND2_X1 U14730 ( .A1(n12660), .A2(n15660), .ZN(n12661) );
  XNOR2_X1 U14731 ( .A(n13397), .B(n13512), .ZN(n13097) );
  XNOR2_X1 U14732 ( .A(n13757), .B(n13427), .ZN(n12665) );
  XNOR2_X1 U14733 ( .A(n12665), .B(n13097), .ZN(n12668) );
  XNOR2_X1 U14734 ( .A(n13756), .B(n13295), .ZN(n13573) );
  XNOR2_X1 U14735 ( .A(n13063), .B(n2448), .ZN(n12666) );
  XNOR2_X1 U14736 ( .A(n13573), .B(n12666), .ZN(n12667) );
  XNOR2_X1 U14737 ( .A(n12668), .B(n12667), .ZN(n13940) );
  XNOR2_X1 U14738 ( .A(n13079), .B(n13791), .ZN(n12670) );
  XNOR2_X1 U14739 ( .A(n13677), .B(n2401), .ZN(n12669) );
  XNOR2_X1 U14740 ( .A(n12670), .B(n12669), .ZN(n12672) );
  XNOR2_X1 U14741 ( .A(n13479), .B(n12671), .ZN(n13550) );
  XNOR2_X1 U14742 ( .A(n13309), .B(n13431), .ZN(n13080) );
  XNOR2_X1 U14743 ( .A(n13468), .B(n13622), .ZN(n13536) );
  XNOR2_X1 U14744 ( .A(n13536), .B(n19899), .ZN(n12678) );
  XNOR2_X1 U14747 ( .A(n13088), .B(n13618), .ZN(n12675) );
  XNOR2_X1 U14748 ( .A(n12676), .B(n12675), .ZN(n12677) );
  MUX2_X1 U14749 ( .A(n2039), .B(n19939), .S(n14052), .Z(n12695) );
  INV_X1 U14750 ( .A(n19797), .ZN(n12679) );
  XNOR2_X1 U14751 ( .A(n13058), .B(n16242), .ZN(n12680) );
  XNOR2_X1 U14752 ( .A(n13070), .B(n13517), .ZN(n13374) );
  INV_X1 U14753 ( .A(n13746), .ZN(n12683) );
  XNOR2_X1 U14754 ( .A(n12683), .B(n13518), .ZN(n13353) );
  XNOR2_X1 U14755 ( .A(n13353), .B(n13374), .ZN(n12691) );
  XNOR2_X1 U14756 ( .A(n12697), .B(n13584), .ZN(n12689) );
  XNOR2_X1 U14757 ( .A(n13747), .B(n610), .ZN(n12688) );
  XNOR2_X1 U14758 ( .A(n12689), .B(n12688), .ZN(n12690) );
  XNOR2_X1 U14759 ( .A(n12691), .B(n12690), .ZN(n13939) );
  XNOR2_X1 U14760 ( .A(n13543), .B(n13767), .ZN(n13322) );
  XNOR2_X1 U14761 ( .A(n13282), .B(n13322), .ZN(n12694) );
  XNOR2_X1 U14762 ( .A(n13409), .B(n13601), .ZN(n13110) );
  XNOR2_X1 U14763 ( .A(n13659), .B(n18084), .ZN(n12692) );
  XNOR2_X1 U14764 ( .A(n13110), .B(n12692), .ZN(n12693) );
  XNOR2_X1 U14765 ( .A(n12694), .B(n12693), .ZN(n14355) );
  INV_X1 U14766 ( .A(n14355), .ZN(n14418) );
  XNOR2_X1 U14767 ( .A(n12697), .B(n12696), .ZN(n13640) );
  XNOR2_X1 U14768 ( .A(n13352), .B(n13585), .ZN(n13812) );
  XNOR2_X1 U14769 ( .A(n13812), .B(n13640), .ZN(n12701) );
  XNOR2_X1 U14770 ( .A(n13590), .B(n12846), .ZN(n12699) );
  XNOR2_X1 U14771 ( .A(n19892), .B(n16487), .ZN(n12698) );
  XNOR2_X1 U14772 ( .A(n12699), .B(n12698), .ZN(n12700) );
  XNOR2_X1 U14773 ( .A(n12701), .B(n12700), .ZN(n14469) );
  INV_X1 U14774 ( .A(n14469), .ZN(n14369) );
  XNOR2_X1 U14775 ( .A(n13085), .B(n13047), .ZN(n13633) );
  XNOR2_X1 U14776 ( .A(n13619), .B(n13336), .ZN(n13816) );
  XNOR2_X1 U14777 ( .A(n13816), .B(n13633), .ZN(n12706) );
  INV_X1 U14778 ( .A(n13534), .ZN(n12702) );
  XNOR2_X1 U14779 ( .A(n12702), .B(n13624), .ZN(n12704) );
  XNOR2_X1 U14780 ( .A(n13193), .B(n2356), .ZN(n12703) );
  XNOR2_X1 U14781 ( .A(n12704), .B(n12703), .ZN(n12705) );
  NOR2_X1 U14782 ( .A1(n14369), .A2(n14468), .ZN(n12727) );
  XNOR2_X1 U14783 ( .A(n13017), .B(n2306), .ZN(n12707) );
  XNOR2_X1 U14784 ( .A(n12707), .B(n19792), .ZN(n12708) );
  XNOR2_X1 U14785 ( .A(n12708), .B(n13357), .ZN(n12712) );
  XNOR2_X1 U14786 ( .A(n13528), .B(n12709), .ZN(n13057) );
  XNOR2_X1 U14791 ( .A(n12986), .B(n632), .ZN(n12714) );
  XNOR2_X1 U14792 ( .A(n13120), .B(n12715), .ZN(n13838) );
  XNOR2_X1 U14793 ( .A(n13404), .B(n13321), .ZN(n13542) );
  XNOR2_X1 U14794 ( .A(n13842), .B(n13542), .ZN(n12719) );
  XNOR2_X1 U14795 ( .A(n13657), .B(n13659), .ZN(n12717) );
  XNOR2_X1 U14796 ( .A(n19697), .B(n311), .ZN(n12716) );
  XNOR2_X1 U14797 ( .A(n12717), .B(n12716), .ZN(n12718) );
  XNOR2_X1 U14798 ( .A(n12719), .B(n12718), .ZN(n14462) );
  INV_X1 U14799 ( .A(n14468), .ZN(n12725) );
  XNOR2_X1 U14800 ( .A(n13344), .B(n13064), .ZN(n13510) );
  XNOR2_X1 U14801 ( .A(n13396), .B(n13099), .ZN(n13853) );
  INV_X1 U14802 ( .A(n13853), .ZN(n12720) );
  XNOR2_X1 U14803 ( .A(n12720), .B(n13510), .ZN(n12724) );
  XNOR2_X1 U14804 ( .A(n13427), .B(n12979), .ZN(n12722) );
  XNOR2_X1 U14805 ( .A(n13425), .B(n19018), .ZN(n12721) );
  XNOR2_X1 U14806 ( .A(n12722), .B(n12721), .ZN(n12723) );
  XNOR2_X1 U14807 ( .A(n12724), .B(n12723), .ZN(n13921) );
  XNOR2_X1 U14808 ( .A(n13484), .B(n13795), .ZN(n12729) );
  XNOR2_X1 U14809 ( .A(n12729), .B(n12728), .ZN(n12733) );
  XNOR2_X1 U14810 ( .A(n12986), .B(n20222), .ZN(n12731) );
  XNOR2_X1 U14811 ( .A(n13673), .B(n13121), .ZN(n12915) );
  INV_X1 U14812 ( .A(n12915), .ZN(n12730) );
  XNOR2_X1 U14813 ( .A(n12730), .B(n12731), .ZN(n12732) );
  XNOR2_X1 U14814 ( .A(n12732), .B(n12733), .ZN(n14826) );
  INV_X1 U14815 ( .A(n13440), .ZN(n12734) );
  XNOR2_X1 U14816 ( .A(n12734), .B(n12920), .ZN(n12739) );
  INV_X1 U14817 ( .A(n19697), .ZN(n12735) );
  INV_X1 U14818 ( .A(n13843), .ZN(n13258) );
  XNOR2_X1 U14819 ( .A(n13258), .B(n12735), .ZN(n12737) );
  XNOR2_X1 U14820 ( .A(n13602), .B(Key[63]), .ZN(n12736) );
  XNOR2_X1 U14821 ( .A(n12737), .B(n12736), .ZN(n12738) );
  XNOR2_X1 U14822 ( .A(n13572), .B(n12979), .ZN(n12741) );
  XNOR2_X1 U14825 ( .A(n20237), .B(n12741), .ZN(n12744) );
  XNOR2_X1 U14827 ( .A(n13064), .B(n19140), .ZN(n12742) );
  XNOR2_X1 U14828 ( .A(n13649), .B(n12742), .ZN(n12743) );
  INV_X1 U14829 ( .A(n12996), .ZN(n12746) );
  XNOR2_X1 U14830 ( .A(n13631), .B(n12746), .ZN(n12750) );
  XNOR2_X1 U14831 ( .A(n20482), .B(n13623), .ZN(n12748) );
  XNOR2_X1 U14832 ( .A(n13193), .B(n19457), .ZN(n12747) );
  XNOR2_X1 U14833 ( .A(n12748), .B(n12747), .ZN(n12749) );
  NOR2_X1 U14834 ( .A1(n14347), .A2(n2684), .ZN(n14833) );
  XNOR2_X1 U14835 ( .A(n13491), .B(n13643), .ZN(n12961) );
  XNOR2_X1 U14836 ( .A(n13641), .B(n12961), .ZN(n12753) );
  XNOR2_X1 U14837 ( .A(n12846), .B(n13250), .ZN(n13012) );
  XNOR2_X1 U14838 ( .A(n19892), .B(n18006), .ZN(n12751) );
  XNOR2_X1 U14839 ( .A(n13012), .B(n12751), .ZN(n12752) );
  XNOR2_X1 U14840 ( .A(n13453), .B(n13369), .ZN(n13668) );
  XNOR2_X1 U14841 ( .A(n13002), .B(n13277), .ZN(n12760) );
  XNOR2_X1 U14842 ( .A(n933), .B(n12760), .ZN(n12764) );
  XNOR2_X1 U14843 ( .A(n13230), .B(n13528), .ZN(n12762) );
  XNOR2_X1 U14844 ( .A(n13783), .B(n18809), .ZN(n12761) );
  XNOR2_X1 U14845 ( .A(n12762), .B(n12761), .ZN(n12763) );
  OAI21_X1 U14846 ( .B1(n14827), .B2(n14826), .A(n19985), .ZN(n12765) );
  NAND2_X1 U14847 ( .A1(n19496), .A2(n12765), .ZN(n12766) );
  MUX2_X1 U14848 ( .A(n15341), .B(n12768), .S(n12842), .Z(n12875) );
  XNOR2_X1 U14849 ( .A(n13248), .B(n12769), .ZN(n13744) );
  XNOR2_X1 U14850 ( .A(n13168), .B(n2423), .ZN(n12771) );
  XNOR2_X1 U14851 ( .A(n13490), .B(n12771), .ZN(n12773) );
  XNOR2_X1 U14852 ( .A(n13070), .B(n20123), .ZN(n12772) );
  XNOR2_X1 U14853 ( .A(n12773), .B(n12772), .ZN(n12774) );
  XNOR2_X1 U14854 ( .A(n12774), .B(n13744), .ZN(n12876) );
  INV_X1 U14855 ( .A(n12876), .ZN(n14094) );
  XNOR2_X1 U14856 ( .A(n13617), .B(n13088), .ZN(n12775) );
  XNOR2_X1 U14857 ( .A(n13761), .B(n12775), .ZN(n12779) );
  XNOR2_X1 U14858 ( .A(n13335), .B(n13048), .ZN(n12777) );
  XNOR2_X1 U14859 ( .A(n13339), .B(n19321), .ZN(n12776) );
  XOR2_X1 U14860 ( .A(n12777), .B(n12776), .Z(n12778) );
  XNOR2_X1 U14862 ( .A(n13293), .B(n13687), .ZN(n12905) );
  INV_X1 U14863 ( .A(n12905), .ZN(n12780) );
  XNOR2_X1 U14864 ( .A(n13134), .B(n19869), .ZN(n13348) );
  XNOR2_X1 U14865 ( .A(n12780), .B(n13348), .ZN(n12783) );
  XNOR2_X1 U14866 ( .A(n12940), .B(n13688), .ZN(n13753) );
  XNOR2_X1 U14867 ( .A(n13063), .B(n1386), .ZN(n12781) );
  XNOR2_X1 U14868 ( .A(n13753), .B(n12781), .ZN(n12782) );
  NAND2_X1 U14869 ( .A1(n19485), .A2(n13931), .ZN(n14093) );
  XNOR2_X1 U14870 ( .A(n13312), .B(n13079), .ZN(n12787) );
  XNOR2_X1 U14871 ( .A(n12787), .B(n12786), .ZN(n12790) );
  INV_X1 U14872 ( .A(n13551), .ZN(n12788) );
  XNOR2_X1 U14873 ( .A(n12788), .B(n13237), .ZN(n12789) );
  XNOR2_X1 U14874 ( .A(n13233), .B(n13527), .ZN(n12794) );
  XNOR2_X1 U14875 ( .A(n13776), .B(n17804), .ZN(n12792) );
  XNOR2_X1 U14876 ( .A(n12791), .B(n12792), .ZN(n12793) );
  XNOR2_X1 U14877 ( .A(n12794), .B(n12793), .ZN(n13930) );
  INV_X1 U14879 ( .A(n13930), .ZN(n14336) );
  XNOR2_X1 U14880 ( .A(n13255), .B(n13280), .ZN(n12921) );
  XNOR2_X1 U14881 ( .A(n13772), .B(n13544), .ZN(n13325) );
  XNOR2_X1 U14882 ( .A(n13325), .B(n12921), .ZN(n12799) );
  INV_X1 U14883 ( .A(n13409), .ZN(n12795) );
  XNOR2_X1 U14884 ( .A(n12795), .B(n13539), .ZN(n12797) );
  XNOR2_X1 U14885 ( .A(n13716), .B(n17733), .ZN(n12796) );
  XNOR2_X1 U14886 ( .A(n12797), .B(n12796), .ZN(n12798) );
  XNOR2_X1 U14887 ( .A(n12798), .B(n12799), .ZN(n12879) );
  INV_X1 U14888 ( .A(n12879), .ZN(n14092) );
  NAND2_X1 U14889 ( .A1(n14334), .A2(n14342), .ZN(n12801) );
  XNOR2_X1 U14891 ( .A(n13511), .B(n18011), .ZN(n12803) );
  XNOR2_X1 U14892 ( .A(n12803), .B(n13572), .ZN(n12804) );
  XNOR2_X1 U14893 ( .A(n13755), .B(n940), .ZN(n12938) );
  XNOR2_X1 U14894 ( .A(n12938), .B(n12804), .ZN(n12806) );
  XNOR2_X1 U14895 ( .A(n13651), .B(n13218), .ZN(n12805) );
  NAND2_X1 U14896 ( .A1(n12807), .A2(n12809), .ZN(n12808) );
  OAI211_X1 U14897 ( .C1(n3586), .C2(n12809), .A(n12811), .B(n12808), .ZN(
        n12810) );
  INV_X1 U14898 ( .A(n12810), .ZN(n12815) );
  AOI21_X1 U14899 ( .B1(n953), .B2(n12812), .A(n12811), .ZN(n12814) );
  XNOR2_X1 U14900 ( .A(n13251), .B(n13287), .ZN(n12965) );
  INV_X1 U14901 ( .A(n12965), .ZN(n12817) );
  INV_X1 U14902 ( .A(n13446), .ZN(n12816) );
  XNOR2_X1 U14903 ( .A(n12816), .B(n13642), .ZN(n13489) );
  INV_X1 U14904 ( .A(n13489), .ZN(n13694) );
  XNOR2_X1 U14905 ( .A(n12817), .B(n13694), .ZN(n12822) );
  INV_X1 U14906 ( .A(n13168), .ZN(n12818) );
  XNOR2_X1 U14907 ( .A(n13491), .B(n12818), .ZN(n12820) );
  XNOR2_X1 U14908 ( .A(n13644), .B(n2082), .ZN(n12819) );
  XNOR2_X1 U14909 ( .A(n12820), .B(n12819), .ZN(n12821) );
  XNOR2_X1 U14910 ( .A(n12822), .B(n12821), .ZN(n14087) );
  INV_X1 U14911 ( .A(n14087), .ZN(n14821) );
  XNOR2_X1 U14912 ( .A(n19883), .B(n13725), .ZN(n12823) );
  XNOR2_X1 U14913 ( .A(n13335), .B(n2454), .ZN(n12825) );
  INV_X1 U14914 ( .A(n13138), .ZN(n13635) );
  XNOR2_X1 U14915 ( .A(n13635), .B(n13623), .ZN(n12824) );
  NOR2_X1 U14916 ( .A1(n14821), .A2(n14818), .ZN(n14328) );
  XNOR2_X1 U14917 ( .A(n13778), .B(n13702), .ZN(n12950) );
  XNOR2_X1 U14918 ( .A(n12826), .B(n12950), .ZN(n12830) );
  XNOR2_X1 U14919 ( .A(n20440), .B(n13706), .ZN(n12828) );
  XNOR2_X1 U14920 ( .A(n13277), .B(n106), .ZN(n12827) );
  XNOR2_X1 U14921 ( .A(n12828), .B(n12827), .ZN(n12829) );
  XNOR2_X1 U14922 ( .A(n12831), .B(n19102), .ZN(n12832) );
  XNOR2_X1 U14923 ( .A(n12832), .B(n13717), .ZN(n12833) );
  XNOR2_X1 U14924 ( .A(n13206), .B(n12833), .ZN(n12835) );
  XNOR2_X1 U14925 ( .A(n12834), .B(n13711), .ZN(n12971) );
  XNOR2_X1 U14926 ( .A(n12835), .B(n12971), .ZN(n14325) );
  NOR2_X1 U14927 ( .A1(n14823), .A2(n14352), .ZN(n14330) );
  AOI21_X1 U14928 ( .B1(n19693), .B2(n14328), .A(n14330), .ZN(n12841) );
  INV_X1 U14929 ( .A(n14325), .ZN(n12932) );
  XNOR2_X1 U14931 ( .A(n12914), .B(n13734), .ZN(n13238) );
  XNOR2_X1 U14932 ( .A(n13199), .B(n13238), .ZN(n12838) );
  XNOR2_X1 U14933 ( .A(n13736), .B(n13484), .ZN(n13311) );
  XNOR2_X1 U14934 ( .A(n13328), .B(n18768), .ZN(n12836) );
  XNOR2_X1 U14935 ( .A(n13311), .B(n12836), .ZN(n12837) );
  XNOR2_X1 U14936 ( .A(n12838), .B(n12837), .ZN(n12931) );
  INV_X1 U14937 ( .A(n12931), .ZN(n14326) );
  NOR2_X1 U14938 ( .A1(n14352), .A2(n912), .ZN(n14817) );
  INV_X1 U14939 ( .A(n14817), .ZN(n12839) );
  OAI211_X1 U14940 ( .C1(n12932), .C2(n14326), .A(n14350), .B(n12839), .ZN(
        n12840) );
  INV_X1 U14941 ( .A(n12842), .ZN(n15468) );
  INV_X1 U14942 ( .A(n13351), .ZN(n12843) );
  XNOR2_X1 U14943 ( .A(n13251), .B(n12843), .ZN(n12845) );
  XNOR2_X1 U14944 ( .A(n13810), .B(n18984), .ZN(n12844) );
  XNOR2_X1 U14945 ( .A(n12845), .B(n12844), .ZN(n12848) );
  XNOR2_X1 U14946 ( .A(n13644), .B(n13376), .ZN(n13073) );
  XNOR2_X1 U14947 ( .A(n13042), .B(n12846), .ZN(n13693) );
  XNOR2_X1 U14948 ( .A(n13073), .B(n13693), .ZN(n12847) );
  INV_X1 U14949 ( .A(n14453), .ZN(n14179) );
  XNOR2_X1 U14950 ( .A(n20260), .B(n13136), .ZN(n13815) );
  XNOR2_X1 U14951 ( .A(n13193), .B(n13192), .ZN(n13722) );
  XNOR2_X1 U14952 ( .A(n13815), .B(n13722), .ZN(n12853) );
  INV_X1 U14953 ( .A(n12997), .ZN(n12849) );
  XNOR2_X1 U14954 ( .A(n12945), .B(n12849), .ZN(n12851) );
  XNOR2_X1 U14955 ( .A(n12851), .B(n12850), .ZN(n12852) );
  INV_X1 U14956 ( .A(n13715), .ZN(n12854) );
  XNOR2_X1 U14957 ( .A(n19697), .B(n12854), .ZN(n12856) );
  XNOR2_X1 U14958 ( .A(n13259), .B(n2446), .ZN(n12855) );
  XNOR2_X1 U14959 ( .A(n12856), .B(n12855), .ZN(n12857) );
  AOI21_X1 U14961 ( .B1(n14179), .B2(n1364), .A(n14451), .ZN(n12873) );
  XNOR2_X1 U14962 ( .A(n13173), .B(n13230), .ZN(n13823) );
  XNOR2_X1 U14963 ( .A(n12859), .B(n19216), .ZN(n12860) );
  XNOR2_X1 U14964 ( .A(n13823), .B(n12860), .ZN(n12862) );
  XNOR2_X1 U14965 ( .A(n12863), .B(n12979), .ZN(n13684) );
  XNOR2_X1 U14966 ( .A(n12864), .B(n13684), .ZN(n12867) );
  XNOR2_X1 U14967 ( .A(n13065), .B(n13848), .ZN(n13650) );
  XNOR2_X1 U14968 ( .A(n13755), .B(n18078), .ZN(n12865) );
  XNOR2_X1 U14969 ( .A(n13650), .B(n12865), .ZN(n12866) );
  INV_X1 U14970 ( .A(n14450), .ZN(n14454) );
  XNOR2_X1 U14971 ( .A(n12914), .B(n20682), .ZN(n12868) );
  XNOR2_X1 U14972 ( .A(n13733), .B(n12868), .ZN(n12872) );
  INV_X1 U14973 ( .A(n13081), .ZN(n12869) );
  XNOR2_X1 U14974 ( .A(n12869), .B(n20223), .ZN(n13676) );
  XNOR2_X1 U14975 ( .A(n13676), .B(n12870), .ZN(n12871) );
  INV_X1 U14976 ( .A(n15339), .ZN(n14896) );
  NAND2_X1 U14977 ( .A1(n14092), .A2(n14336), .ZN(n12877) );
  NAND2_X1 U14978 ( .A1(n12880), .A2(n13931), .ZN(n12881) );
  INV_X1 U14979 ( .A(n14052), .ZN(n14357) );
  MUX2_X1 U14980 ( .A(n14357), .B(n14419), .S(n19939), .Z(n12884) );
  NAND3_X1 U14981 ( .A1(n14357), .A2(n14355), .A3(n14419), .ZN(n12883) );
  NAND3_X1 U14982 ( .A1(n2039), .A2(n14359), .A3(n14422), .ZN(n12882) );
  MUX2_X1 U14985 ( .A(n14369), .B(n19531), .S(n3252), .Z(n12887) );
  MUX2_X1 U14986 ( .A(n14465), .B(n19819), .S(n19657), .Z(n12886) );
  INV_X1 U14987 ( .A(n12888), .ZN(n15165) );
  XNOR2_X1 U14988 ( .A(n12889), .B(n12945), .ZN(n13764) );
  XNOR2_X1 U14989 ( .A(n13764), .B(n13631), .ZN(n12893) );
  XNOR2_X1 U14990 ( .A(n13617), .B(n13725), .ZN(n12891) );
  XNOR2_X1 U14991 ( .A(n13048), .B(n1904), .ZN(n12890) );
  XNOR2_X1 U14992 ( .A(n12891), .B(n12890), .ZN(n12892) );
  XNOR2_X1 U14993 ( .A(n12893), .B(n12892), .ZN(n12910) );
  INV_X1 U14994 ( .A(n12910), .ZN(n14441) );
  XNOR2_X1 U14995 ( .A(n20123), .B(n13643), .ZN(n12895) );
  XNOR2_X1 U14996 ( .A(n12895), .B(n12894), .ZN(n12899) );
  XNOR2_X1 U14997 ( .A(n13250), .B(n2413), .ZN(n12897) );
  INV_X1 U14998 ( .A(n13251), .ZN(n12896) );
  XNOR2_X1 U14999 ( .A(n12898), .B(n12899), .ZN(n12911) );
  XNOR2_X1 U15000 ( .A(n13019), .B(n13580), .ZN(n12901) );
  XNOR2_X1 U15001 ( .A(n13783), .B(n2122), .ZN(n12900) );
  XNOR2_X1 U15002 ( .A(n12901), .B(n12900), .ZN(n12904) );
  INV_X1 U15003 ( .A(n12950), .ZN(n12902) );
  XNOR2_X1 U15004 ( .A(n13668), .B(n12902), .ZN(n12903) );
  XNOR2_X1 U15005 ( .A(n12905), .B(n12938), .ZN(n12909) );
  XNOR2_X1 U15006 ( .A(n12906), .B(n18863), .ZN(n12907) );
  XNOR2_X1 U15007 ( .A(n13649), .B(n12907), .ZN(n12908) );
  XNOR2_X1 U15008 ( .A(n13312), .B(n19734), .ZN(n12912) );
  XNOR2_X1 U15009 ( .A(n12912), .B(n12913), .ZN(n12918) );
  XNOR2_X1 U15010 ( .A(n12914), .B(n2424), .ZN(n12916) );
  XNOR2_X1 U15011 ( .A(n12915), .B(n12916), .ZN(n12917) );
  XNOR2_X1 U15012 ( .A(n12918), .B(n12917), .ZN(n14167) );
  INV_X1 U15013 ( .A(n14167), .ZN(n12919) );
  XNOR2_X1 U15014 ( .A(n12921), .B(n12920), .ZN(n12925) );
  XNOR2_X1 U15016 ( .A(n13259), .B(n2192), .ZN(n12922) );
  XNOR2_X1 U15017 ( .A(n12923), .B(n12922), .ZN(n12924) );
  XNOR2_X1 U15018 ( .A(n12925), .B(n12924), .ZN(n13918) );
  AOI22_X1 U15019 ( .A1(n14439), .A2(n12926), .B1(n3516), .B2(n20262), .ZN(
        n12927) );
  NAND2_X1 U15020 ( .A1(n15165), .A2(n15379), .ZN(n15375) );
  MUX2_X1 U15021 ( .A(n13559), .B(n1363), .S(n14455), .Z(n12930) );
  NAND2_X1 U15023 ( .A1(n231), .A2(n19513), .ZN(n15031) );
  NAND2_X1 U15024 ( .A1(n15375), .A2(n15031), .ZN(n12935) );
  AOI21_X1 U15025 ( .B1(n235), .B2(n12931), .A(n14352), .ZN(n12934) );
  AND2_X1 U15026 ( .A1(n12932), .A2(n12931), .ZN(n14085) );
  OAI21_X1 U15027 ( .B1(n14086), .B2(n14085), .A(n19821), .ZN(n12933) );
  XNOR2_X1 U15029 ( .A(n12937), .B(n13572), .ZN(n12939) );
  XNOR2_X1 U15030 ( .A(n12938), .B(n12939), .ZN(n12943) );
  XNOR2_X1 U15031 ( .A(n13398), .B(n12940), .ZN(n13215) );
  XNOR2_X1 U15032 ( .A(n13757), .B(n18146), .ZN(n12941) );
  XNOR2_X1 U15033 ( .A(n13215), .B(n12941), .ZN(n12942) );
  XNOR2_X1 U15034 ( .A(n13222), .B(n13762), .ZN(n12944) );
  XNOR2_X1 U15035 ( .A(n13725), .B(n13623), .ZN(n13302) );
  XNOR2_X1 U15036 ( .A(n13302), .B(n12944), .ZN(n12949) );
  XNOR2_X1 U15037 ( .A(n13624), .B(n19923), .ZN(n12947) );
  XNOR2_X1 U15038 ( .A(n19883), .B(n18065), .ZN(n12946) );
  XNOR2_X1 U15039 ( .A(n12947), .B(n12946), .ZN(n12948) );
  XNOR2_X1 U15040 ( .A(n12949), .B(n12948), .ZN(n12973) );
  INV_X1 U15041 ( .A(n12973), .ZN(n14509) );
  NOR2_X1 U15042 ( .A1(n20473), .A2(n14509), .ZN(n14636) );
  XNOR2_X1 U15043 ( .A(n13577), .B(n13774), .ZN(n13525) );
  XNOR2_X1 U15044 ( .A(n12950), .B(n13525), .ZN(n12954) );
  XNOR2_X1 U15045 ( .A(n13369), .B(n13277), .ZN(n12952) );
  XNOR2_X1 U15046 ( .A(n19796), .B(n2280), .ZN(n12951) );
  XNOR2_X1 U15047 ( .A(n12952), .B(n12951), .ZN(n12953) );
  XNOR2_X1 U15049 ( .A(n13792), .B(n12955), .ZN(n12956) );
  XNOR2_X1 U15050 ( .A(n12956), .B(n12957), .ZN(n12960) );
  XNOR2_X1 U15051 ( .A(n13673), .B(Key[94]), .ZN(n12958) );
  XNOR2_X1 U15052 ( .A(n13311), .B(n12958), .ZN(n12959) );
  XNOR2_X1 U15053 ( .A(n12960), .B(n12959), .ZN(n14642) );
  NOR2_X1 U15054 ( .A1(n14642), .A2(n14641), .ZN(n14031) );
  AOI22_X1 U15055 ( .A1(n14636), .A2(n19703), .B1(n14031), .B2(n14509), .ZN(
        n12976) );
  XNOR2_X1 U15056 ( .A(n12961), .B(n13248), .ZN(n12968) );
  XNOR2_X1 U15057 ( .A(n12964), .B(n13747), .ZN(n12966) );
  XNOR2_X1 U15058 ( .A(n12965), .B(n12966), .ZN(n12967) );
  XNOR2_X1 U15060 ( .A(n12992), .B(n19222), .ZN(n12969) );
  XNOR2_X1 U15061 ( .A(n12969), .B(n13321), .ZN(n12970) );
  XNOR2_X1 U15062 ( .A(n13658), .B(n13539), .ZN(n13207) );
  XNOR2_X1 U15064 ( .A(n12977), .B(n13687), .ZN(n12978) );
  XNOR2_X1 U15065 ( .A(n20442), .B(n12978), .ZN(n12983) );
  XNOR2_X1 U15066 ( .A(n12471), .B(n2123), .ZN(n12981) );
  XNOR2_X1 U15067 ( .A(n12979), .B(n13462), .ZN(n12980) );
  XNOR2_X1 U15068 ( .A(n12981), .B(n12980), .ZN(n12982) );
  XNOR2_X1 U15070 ( .A(n13791), .B(n20223), .ZN(n12985) );
  XNOR2_X1 U15071 ( .A(n13029), .B(n12984), .ZN(n13732) );
  XNOR2_X1 U15072 ( .A(n12985), .B(n13732), .ZN(n12990) );
  XNOR2_X1 U15073 ( .A(n13795), .B(n12986), .ZN(n12988) );
  XNOR2_X1 U15074 ( .A(n13390), .B(n347), .ZN(n12987) );
  XNOR2_X1 U15075 ( .A(n12987), .B(n12988), .ZN(n12989) );
  XNOR2_X1 U15076 ( .A(n12990), .B(n12989), .ZN(n14525) );
  NOR2_X1 U15077 ( .A1(n20443), .A2(n19831), .ZN(n13008) );
  XNOR2_X1 U15078 ( .A(n13260), .B(n17024), .ZN(n12991) );
  XNOR2_X1 U15079 ( .A(n13714), .B(n12991), .ZN(n12995) );
  XNOR2_X1 U15080 ( .A(n13710), .B(n12992), .ZN(n13497) );
  XNOR2_X1 U15081 ( .A(n12993), .B(n13497), .ZN(n12994) );
  XNOR2_X1 U15082 ( .A(n13721), .B(n13762), .ZN(n13470) );
  XNOR2_X1 U15083 ( .A(n13470), .B(n12996), .ZN(n13001) );
  XNOR2_X1 U15084 ( .A(n12999), .B(n12998), .ZN(n13000) );
  XNOR2_X1 U15086 ( .A(n13783), .B(n642), .ZN(n13004) );
  XNOR2_X1 U15087 ( .A(n13005), .B(n13004), .ZN(n13006) );
  XNOR2_X1 U15089 ( .A(n13695), .B(n13810), .ZN(n13011) );
  XNOR2_X1 U15090 ( .A(n13747), .B(n17466), .ZN(n13010) );
  XNOR2_X1 U15091 ( .A(n13011), .B(n13010), .ZN(n13015) );
  XNOR2_X1 U15092 ( .A(n13446), .B(n13351), .ZN(n13013) );
  XOR2_X1 U15093 ( .A(n13013), .B(n13012), .Z(n13014) );
  NAND3_X1 U15094 ( .A1(n14522), .A2(n14524), .A3(n20443), .ZN(n13016) );
  INV_X1 U15095 ( .A(n15684), .ZN(n15687) );
  NOR2_X1 U15096 ( .A1(n19978), .A2(n15687), .ZN(n13096) );
  INV_X1 U15097 ( .A(n19978), .ZN(n15779) );
  XNOR2_X1 U15098 ( .A(n13576), .B(n13114), .ZN(n13829) );
  XNOR2_X1 U15099 ( .A(n20199), .B(n13018), .ZN(n13666) );
  XNOR2_X1 U15100 ( .A(n13666), .B(n13829), .ZN(n13024) );
  XNOR2_X1 U15101 ( .A(n13019), .B(n13453), .ZN(n13022) );
  XNOR2_X1 U15102 ( .A(n13020), .B(n2369), .ZN(n13021) );
  XNOR2_X1 U15103 ( .A(n13022), .B(n13021), .ZN(n13023) );
  XNOR2_X1 U15105 ( .A(n13255), .B(n13659), .ZN(n13026) );
  XNOR2_X1 U15106 ( .A(n13715), .B(n2395), .ZN(n13025) );
  XNOR2_X1 U15107 ( .A(n13027), .B(n13108), .ZN(n13655) );
  XNOR2_X1 U15108 ( .A(n13842), .B(n13655), .ZN(n13028) );
  XNOR2_X1 U15109 ( .A(n19734), .B(n13677), .ZN(n13030) );
  XNOR2_X1 U15110 ( .A(n13030), .B(n13838), .ZN(n13034) );
  XNOR2_X1 U15111 ( .A(n13031), .B(n13081), .ZN(n13033) );
  XNOR2_X1 U15112 ( .A(n13121), .B(n1869), .ZN(n13032) );
  XNOR2_X1 U15113 ( .A(n19937), .B(n13687), .ZN(n13036) );
  XNOR2_X1 U15114 ( .A(n13036), .B(n13035), .ZN(n13039) );
  XNOR2_X1 U15115 ( .A(n13422), .B(n2317), .ZN(n13037) );
  XNOR2_X1 U15116 ( .A(n13853), .B(n13037), .ZN(n13038) );
  XNOR2_X2 U15117 ( .A(n13039), .B(n13038), .ZN(n14499) );
  INV_X1 U15118 ( .A(n14499), .ZN(n13040) );
  XNOR2_X1 U15119 ( .A(n13041), .B(n13126), .ZN(n13443) );
  XNOR2_X1 U15120 ( .A(n13443), .B(n13812), .ZN(n13046) );
  XNOR2_X1 U15121 ( .A(n13042), .B(n13695), .ZN(n13044) );
  XNOR2_X1 U15122 ( .A(n13644), .B(n2310), .ZN(n13043) );
  XNOR2_X1 U15123 ( .A(n13044), .B(n13043), .ZN(n13045) );
  XNOR2_X1 U15124 ( .A(n13046), .B(n13045), .ZN(n14305) );
  XNOR2_X1 U15126 ( .A(n13103), .B(n13047), .ZN(n13417) );
  XNOR2_X1 U15127 ( .A(n13816), .B(n13417), .ZN(n13052) );
  XNOR2_X1 U15128 ( .A(n13048), .B(n13192), .ZN(n13050) );
  XNOR2_X1 U15129 ( .A(n13050), .B(n13049), .ZN(n13051) );
  INV_X1 U15130 ( .A(n14497), .ZN(n14307) );
  XNOR2_X1 U15135 ( .A(n13579), .B(n13057), .ZN(n13062) );
  XNOR2_X1 U15136 ( .A(n13058), .B(n13173), .ZN(n13367) );
  XNOR2_X1 U15137 ( .A(n20199), .B(n2216), .ZN(n13060) );
  XNOR2_X1 U15138 ( .A(n13367), .B(n13060), .ZN(n13061) );
  XNOR2_X1 U15139 ( .A(n13400), .B(n13573), .ZN(n13069) );
  XNOR2_X1 U15141 ( .A(n19937), .B(n13425), .ZN(n13066) );
  XNOR2_X1 U15142 ( .A(n13067), .B(n13066), .ZN(n13068) );
  XNOR2_X2 U15143 ( .A(n13069), .B(n13068), .ZN(n14520) );
  XNOR2_X1 U15144 ( .A(n13070), .B(n13584), .ZN(n13072) );
  XNOR2_X1 U15145 ( .A(n19892), .B(n17787), .ZN(n13071) );
  XNOR2_X1 U15146 ( .A(n13072), .B(n13071), .ZN(n13075) );
  XNOR2_X1 U15147 ( .A(n13444), .B(n13073), .ZN(n13074) );
  XNOR2_X1 U15148 ( .A(n13074), .B(n13075), .ZN(n14321) );
  INV_X1 U15149 ( .A(n14321), .ZN(n14186) );
  XNOR2_X1 U15150 ( .A(n13404), .B(n2381), .ZN(n13077) );
  AOI22_X1 U15151 ( .A1(n15119), .A2(n14520), .B1(n14186), .B2(n14514), .ZN(
        n13094) );
  XNOR2_X1 U15152 ( .A(n13080), .B(n13389), .ZN(n13084) );
  XNOR2_X1 U15153 ( .A(n13081), .B(n13833), .ZN(n13082) );
  XNOR2_X1 U15155 ( .A(n13085), .B(n20482), .ZN(n13087) );
  XNOR2_X1 U15156 ( .A(n13087), .B(n13086), .ZN(n13091) );
  XNOR2_X1 U15157 ( .A(n13616), .B(n13618), .ZN(n13089) );
  XNOR2_X1 U15158 ( .A(n13382), .B(n13089), .ZN(n13090) );
  XNOR2_X1 U15159 ( .A(n13091), .B(n13090), .ZN(n13563) );
  INV_X1 U15160 ( .A(n13563), .ZN(n14516) );
  NAND2_X1 U15161 ( .A1(n14514), .A2(n14520), .ZN(n13092) );
  OAI21_X1 U15162 ( .B1(n14519), .B2(n14520), .A(n13092), .ZN(n13093) );
  INV_X1 U15163 ( .A(n15686), .ZN(n15685) );
  OAI21_X1 U15164 ( .B1(n13096), .B2(n13095), .A(n15685), .ZN(n13182) );
  XNOR2_X1 U15167 ( .A(n13422), .B(n2392), .ZN(n13100) );
  XNOR2_X1 U15168 ( .A(n13099), .B(n13688), .ZN(n13299) );
  XNOR2_X1 U15169 ( .A(n13100), .B(n13299), .ZN(n13101) );
  XNOR2_X1 U15170 ( .A(n13103), .B(n18887), .ZN(n13104) );
  XNOR2_X1 U15171 ( .A(n13536), .B(n13104), .ZN(n13107) );
  XNOR2_X1 U15172 ( .A(n13724), .B(n13336), .ZN(n13105) );
  XNOR2_X1 U15173 ( .A(n13382), .B(n13105), .ZN(n13106) );
  INV_X1 U15175 ( .A(n13981), .ZN(n14020) );
  XNOR2_X1 U15176 ( .A(n13319), .B(n13716), .ZN(n13284) );
  XNOR2_X1 U15177 ( .A(n13108), .B(n2445), .ZN(n13109) );
  XNOR2_X1 U15178 ( .A(n13284), .B(n13109), .ZN(n13113) );
  INV_X1 U15179 ( .A(n13110), .ZN(n13111) );
  XNOR2_X1 U15180 ( .A(n13844), .B(n13111), .ZN(n13112) );
  XNOR2_X1 U15181 ( .A(n13530), .B(n13367), .ZN(n13117) );
  XNOR2_X1 U15182 ( .A(n13453), .B(n16651), .ZN(n13115) );
  XNOR2_X1 U15183 ( .A(n13114), .B(n915), .ZN(n13267) );
  XNOR2_X1 U15184 ( .A(n13267), .B(n13115), .ZN(n13116) );
  XNOR2_X1 U15185 ( .A(n13117), .B(n13116), .ZN(n13118) );
  INV_X1 U15186 ( .A(n13118), .ZN(n14261) );
  INV_X1 U15187 ( .A(n13550), .ZN(n13119) );
  XNOR2_X1 U15188 ( .A(n13119), .B(n13389), .ZN(n13124) );
  XNOR2_X1 U15189 ( .A(n13121), .B(n18055), .ZN(n13122) );
  XNOR2_X1 U15190 ( .A(n13313), .B(n13122), .ZN(n13123) );
  XNOR2_X1 U15191 ( .A(n13124), .B(n13123), .ZN(n13980) );
  INV_X1 U15192 ( .A(n13980), .ZN(n14260) );
  NAND2_X1 U15193 ( .A1(n20424), .A2(n14260), .ZN(n13125) );
  OAI211_X1 U15194 ( .C1(n14262), .C2(n14020), .A(n14543), .B(n13125), .ZN(
        n13132) );
  XNOR2_X1 U15195 ( .A(n13126), .B(n13374), .ZN(n13131) );
  XNOR2_X1 U15196 ( .A(n13697), .B(n19180), .ZN(n13128) );
  INV_X1 U15197 ( .A(n13352), .ZN(n13127) );
  XNOR2_X1 U15198 ( .A(n13128), .B(n13127), .ZN(n13129) );
  XNOR2_X1 U15199 ( .A(n13808), .B(n13129), .ZN(n13130) );
  XNOR2_X1 U15200 ( .A(n13130), .B(n13131), .ZN(n14673) );
  INV_X1 U15201 ( .A(n14673), .ZN(n14266) );
  XNOR2_X1 U15202 ( .A(n13136), .B(n2382), .ZN(n13137) );
  INV_X1 U15204 ( .A(n13147), .ZN(n13142) );
  NOR2_X1 U15205 ( .A1(n13142), .A2(n13141), .ZN(n13143) );
  OAI21_X1 U15206 ( .B1(n13144), .B2(n13143), .A(n13146), .ZN(n13151) );
  NOR3_X1 U15207 ( .A1(n13147), .A2(n13146), .A3(n13145), .ZN(n13148) );
  NOR2_X1 U15208 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  NAND2_X1 U15209 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  XNOR2_X1 U15210 ( .A(n13152), .B(n13321), .ZN(n13595) );
  XNOR2_X1 U15211 ( .A(n13153), .B(n13595), .ZN(n13158) );
  XNOR2_X1 U15212 ( .A(n13154), .B(n19904), .ZN(n13156) );
  XNOR2_X1 U15213 ( .A(n13544), .B(n2420), .ZN(n13155) );
  XNOR2_X1 U15214 ( .A(n13156), .B(n13155), .ZN(n13157) );
  XNOR2_X1 U15215 ( .A(n13158), .B(n13157), .ZN(n14316) );
  INV_X1 U15216 ( .A(n13309), .ZN(n13608) );
  XNOR2_X1 U15217 ( .A(n13608), .B(n13834), .ZN(n13160) );
  XNOR2_X1 U15218 ( .A(n13328), .B(n2305), .ZN(n13159) );
  XNOR2_X1 U15219 ( .A(n13160), .B(n13159), .ZN(n13163) );
  XNOR2_X1 U15220 ( .A(n13161), .B(n13330), .ZN(n13610) );
  XNOR2_X1 U15221 ( .A(n13610), .B(n13486), .ZN(n13162) );
  NAND2_X1 U15222 ( .A1(n13166), .A2(n13165), .ZN(n14538) );
  XNOR2_X1 U15223 ( .A(n13376), .B(n19689), .ZN(n13167) );
  XNOR2_X1 U15224 ( .A(n13490), .B(n13167), .ZN(n13171) );
  XNOR2_X1 U15225 ( .A(n13642), .B(n2218), .ZN(n13169) );
  XNOR2_X1 U15226 ( .A(n13590), .B(n13168), .ZN(n13523) );
  XNOR2_X1 U15227 ( .A(n13169), .B(n13523), .ZN(n13170) );
  XNOR2_X1 U15228 ( .A(n13577), .B(n13266), .ZN(n13172) );
  XNOR2_X1 U15229 ( .A(n13475), .B(n13172), .ZN(n13177) );
  XNOR2_X1 U15230 ( .A(n13173), .B(n2442), .ZN(n13175) );
  XNOR2_X1 U15231 ( .A(n20440), .B(n13580), .ZN(n13174) );
  XNOR2_X1 U15232 ( .A(n13175), .B(n13174), .ZN(n13176) );
  OAI211_X1 U15233 ( .C1(n15687), .C2(n15683), .A(n13180), .B(n15686), .ZN(
        n13181) );
  XNOR2_X1 U15234 ( .A(n13183), .B(n17104), .ZN(n13184) );
  XNOR2_X1 U15235 ( .A(n20253), .B(n19158), .ZN(n13185) );
  XNOR2_X1 U15236 ( .A(n13186), .B(n13693), .ZN(n13188) );
  INV_X1 U15237 ( .A(n13619), .ZN(n13189) );
  XNOR2_X1 U15238 ( .A(n13222), .B(n13189), .ZN(n13190) );
  XNOR2_X1 U15239 ( .A(n13191), .B(n13190), .ZN(n13197) );
  XNOR2_X1 U15240 ( .A(n19923), .B(n13192), .ZN(n13195) );
  XNOR2_X1 U15241 ( .A(n13193), .B(n17993), .ZN(n13194) );
  XNOR2_X1 U15242 ( .A(n13195), .B(n13194), .ZN(n13196) );
  NOR2_X1 U15243 ( .A1(n14654), .A2(n20266), .ZN(n13221) );
  INV_X1 U15244 ( .A(n13673), .ZN(n13198) );
  XNOR2_X1 U15245 ( .A(n13198), .B(n13607), .ZN(n13388) );
  XNOR2_X1 U15246 ( .A(n13199), .B(n13388), .ZN(n13202) );
  XNOR2_X1 U15247 ( .A(n13792), .B(n2329), .ZN(n13200) );
  XNOR2_X1 U15248 ( .A(n13733), .B(n13200), .ZN(n13201) );
  XNOR2_X1 U15249 ( .A(n19697), .B(n2079), .ZN(n13205) );
  XNOR2_X1 U15250 ( .A(n13206), .B(n13207), .ZN(n13208) );
  INV_X1 U15251 ( .A(n13708), .ZN(n13212) );
  XNOR2_X1 U15252 ( .A(n13774), .B(n620), .ZN(n13210) );
  XNOR2_X1 U15253 ( .A(n13210), .B(n13576), .ZN(n13211) );
  XNOR2_X1 U15254 ( .A(n13212), .B(n13211), .ZN(n13214) );
  INV_X1 U15255 ( .A(n14022), .ZN(n14653) );
  INV_X1 U15256 ( .A(n13215), .ZN(n13216) );
  XNOR2_X1 U15257 ( .A(n13216), .B(n13684), .ZN(n13220) );
  XNOR2_X1 U15258 ( .A(n20469), .B(n17932), .ZN(n13217) );
  XNOR2_X1 U15259 ( .A(n13218), .B(n13217), .ZN(n13219) );
  INV_X1 U15260 ( .A(n13222), .ZN(n13223) );
  XNOR2_X1 U15261 ( .A(n13616), .B(n13223), .ZN(n13225) );
  INV_X1 U15262 ( .A(n13764), .ZN(n13224) );
  XNOR2_X1 U15263 ( .A(n13224), .B(n13225), .ZN(n13229) );
  XNOR2_X1 U15264 ( .A(n20260), .B(n2298), .ZN(n13226) );
  XOR2_X1 U15265 ( .A(n20226), .B(n13226), .Z(n13228) );
  XNOR2_X1 U15266 ( .A(n13231), .B(n13230), .ZN(n13665) );
  XNOR2_X1 U15267 ( .A(n13783), .B(n18779), .ZN(n13232) );
  XNOR2_X1 U15268 ( .A(n13665), .B(n13232), .ZN(n13236) );
  XNOR2_X1 U15270 ( .A(n13238), .B(n13237), .ZN(n13241) );
  XNOR2_X1 U15271 ( .A(n13309), .B(n20222), .ZN(n13239) );
  XNOR2_X1 U15272 ( .A(n13241), .B(n13240), .ZN(n14575) );
  MUX2_X1 U15273 ( .A(n14267), .B(n14574), .S(n14575), .Z(n13264) );
  XNOR2_X1 U15274 ( .A(n13295), .B(n2385), .ZN(n13242) );
  XNOR2_X1 U15275 ( .A(n20442), .B(n13243), .ZN(n13245) );
  INV_X1 U15276 ( .A(n14570), .ZN(n14738) );
  AND2_X1 U15277 ( .A1(n14571), .A2(n14738), .ZN(n14578) );
  XNOR2_X1 U15278 ( .A(n13642), .B(n13810), .ZN(n13247) );
  XNOR2_X1 U15279 ( .A(n13247), .B(n13248), .ZN(n13253) );
  XNOR2_X1 U15280 ( .A(n20123), .B(n17587), .ZN(n13249) );
  XNOR2_X1 U15281 ( .A(n13249), .B(n19689), .ZN(n13252) );
  XNOR2_X1 U15282 ( .A(n13251), .B(n13250), .ZN(n13750) );
  XNOR2_X1 U15283 ( .A(n13539), .B(n2375), .ZN(n13256) );
  XNOR2_X1 U15284 ( .A(n13257), .B(n13256), .ZN(n13262) );
  XNOR2_X1 U15285 ( .A(n13258), .B(n13717), .ZN(n13656) );
  XNOR2_X1 U15286 ( .A(n13260), .B(n13259), .ZN(n13769) );
  XNOR2_X1 U15287 ( .A(n13656), .B(n13769), .ZN(n13261) );
  XNOR2_X1 U15288 ( .A(n13702), .B(n456), .ZN(n13265) );
  XNOR2_X1 U15289 ( .A(n13266), .B(n13265), .ZN(n13268) );
  XNOR2_X1 U15290 ( .A(n13268), .B(n13267), .ZN(n13279) );
  INV_X1 U15291 ( .A(n13269), .ZN(n13273) );
  INV_X1 U15292 ( .A(n13270), .ZN(n13271) );
  NAND2_X1 U15293 ( .A1(n13271), .A2(n13275), .ZN(n13272) );
  XNOR2_X1 U15295 ( .A(n13276), .B(n13277), .ZN(n13278) );
  XNOR2_X1 U15296 ( .A(n13278), .B(n13580), .ZN(n13477) );
  INV_X1 U15297 ( .A(n13316), .ZN(n14704) );
  INV_X1 U15298 ( .A(n13280), .ZN(n13281) );
  XNOR2_X1 U15299 ( .A(n13281), .B(n13602), .ZN(n13501) );
  XNOR2_X1 U15300 ( .A(n13282), .B(n13501), .ZN(n13286) );
  XNOR2_X1 U15301 ( .A(n13711), .B(n17851), .ZN(n13283) );
  XNOR2_X1 U15302 ( .A(n13284), .B(n13283), .ZN(n13285) );
  NOR2_X1 U15303 ( .A1(n14704), .A2(n14563), .ZN(n13308) );
  XNOR2_X1 U15304 ( .A(n13491), .B(n17535), .ZN(n13288) );
  XNOR2_X1 U15305 ( .A(n13288), .B(n13287), .ZN(n13290) );
  XNOR2_X1 U15306 ( .A(n13290), .B(n13289), .ZN(n13292) );
  XNOR2_X1 U15307 ( .A(n13292), .B(n13291), .ZN(n14562) );
  INV_X1 U15308 ( .A(n14562), .ZN(n14706) );
  INV_X1 U15309 ( .A(n13293), .ZN(n13294) );
  XNOR2_X1 U15310 ( .A(n13757), .B(n13294), .ZN(n13463) );
  XNOR2_X1 U15311 ( .A(n13295), .B(n645), .ZN(n13297) );
  INV_X1 U15312 ( .A(n13686), .ZN(n13296) );
  XNOR2_X1 U15313 ( .A(n13297), .B(n13296), .ZN(n13298) );
  XNOR2_X1 U15315 ( .A(n13572), .B(n13299), .ZN(n13300) );
  NOR2_X1 U15316 ( .A1(n14706), .A2(n20498), .ZN(n13955) );
  XNOR2_X1 U15317 ( .A(n13303), .B(n13302), .ZN(n13307) );
  XNOR2_X1 U15318 ( .A(n13724), .B(n18726), .ZN(n13304) );
  XNOR2_X1 U15319 ( .A(n13305), .B(n13304), .ZN(n13306) );
  XNOR2_X2 U15320 ( .A(n13307), .B(n13306), .ZN(n14566) );
  XNOR2_X1 U15321 ( .A(n13309), .B(n2376), .ZN(n13310) );
  XNOR2_X1 U15322 ( .A(n13311), .B(n13310), .ZN(n13315) );
  XNOR2_X1 U15323 ( .A(n13483), .B(n13313), .ZN(n13314) );
  MUX2_X1 U15324 ( .A(n14275), .B(n14273), .S(n14566), .Z(n13317) );
  MUX2_X1 U15326 ( .A(n15673), .B(n234), .S(n15672), .Z(n13461) );
  INV_X1 U15327 ( .A(n13319), .ZN(n13320) );
  XNOR2_X1 U15328 ( .A(n13321), .B(n13320), .ZN(n13323) );
  XNOR2_X1 U15329 ( .A(n13323), .B(n13322), .ZN(n13327) );
  XNOR2_X1 U15330 ( .A(n13405), .B(n18439), .ZN(n13324) );
  XNOR2_X1 U15331 ( .A(n13325), .B(n13324), .ZN(n13326) );
  XNOR2_X1 U15332 ( .A(n13328), .B(n13479), .ZN(n13839) );
  XNOR2_X1 U15333 ( .A(n13839), .B(n13329), .ZN(n13334) );
  XNOR2_X1 U15334 ( .A(n13390), .B(n20064), .ZN(n13331) );
  XNOR2_X1 U15335 ( .A(n13331), .B(n13332), .ZN(n13333) );
  XNOR2_X1 U15336 ( .A(n13334), .B(n13333), .ZN(n14690) );
  NAND2_X1 U15338 ( .A1(n14385), .A2(n19895), .ZN(n14387) );
  INV_X1 U15339 ( .A(n16366), .ZN(n19296) );
  XNOR2_X1 U15340 ( .A(n13335), .B(n19296), .ZN(n13338) );
  XNOR2_X1 U15341 ( .A(n13624), .B(n13336), .ZN(n13337) );
  XNOR2_X1 U15342 ( .A(n13338), .B(n13337), .ZN(n13342) );
  XNOR2_X1 U15343 ( .A(n13339), .B(n13618), .ZN(n13760) );
  XNOR2_X1 U15344 ( .A(n13340), .B(n13760), .ZN(n13341) );
  NAND2_X1 U15345 ( .A1(n14387), .A2(n200), .ZN(n13365) );
  XNOR2_X1 U15346 ( .A(n13344), .B(n13343), .ZN(n13346) );
  INV_X1 U15347 ( .A(n13512), .ZN(n13849) );
  XNOR2_X1 U15348 ( .A(n13849), .B(n19052), .ZN(n13345) );
  XNOR2_X1 U15349 ( .A(n13347), .B(n13348), .ZN(n13349) );
  XNOR2_X1 U15350 ( .A(n13745), .B(n1969), .ZN(n13350) );
  XNOR2_X1 U15351 ( .A(n13350), .B(n13523), .ZN(n13356) );
  XNOR2_X1 U15352 ( .A(n13352), .B(n13351), .ZN(n13354) );
  XNOR2_X1 U15353 ( .A(n13354), .B(n13353), .ZN(n13355) );
  XNOR2_X1 U15354 ( .A(n13356), .B(n13355), .ZN(n14127) );
  INV_X1 U15355 ( .A(n14127), .ZN(n14695) );
  XNOR2_X1 U15356 ( .A(n13776), .B(n19854), .ZN(n13358) );
  XNOR2_X1 U15357 ( .A(n13357), .B(n13358), .ZN(n13363) );
  XNOR2_X1 U15358 ( .A(n13359), .B(n20440), .ZN(n13361) );
  XNOR2_X1 U15359 ( .A(n13361), .B(n13360), .ZN(n13362) );
  XNOR2_X1 U15360 ( .A(n13363), .B(n13362), .ZN(n13946) );
  NAND2_X1 U15364 ( .A1(n15221), .A2(n15667), .ZN(n15772) );
  XNOR2_X1 U15365 ( .A(n13367), .B(n13366), .ZN(n13373) );
  XNOR2_X1 U15366 ( .A(n13368), .B(n13369), .ZN(n13371) );
  XNOR2_X1 U15367 ( .A(n13528), .B(Key[60]), .ZN(n13370) );
  XNOR2_X1 U15368 ( .A(n13371), .B(n13370), .ZN(n13372) );
  XNOR2_X1 U15371 ( .A(n13375), .B(n13374), .ZN(n13380) );
  XNOR2_X1 U15372 ( .A(n13376), .B(n13643), .ZN(n13378) );
  XNOR2_X1 U15373 ( .A(n20253), .B(n18208), .ZN(n13377) );
  XNOR2_X1 U15374 ( .A(n13378), .B(n13377), .ZN(n13379) );
  XNOR2_X1 U15375 ( .A(n13380), .B(n13379), .ZN(n14727) );
  INV_X1 U15376 ( .A(n14727), .ZN(n14224) );
  XNOR2_X1 U15378 ( .A(n13382), .B(n19824), .ZN(n13387) );
  XNOR2_X1 U15379 ( .A(n13622), .B(n2284), .ZN(n13385) );
  XNOR2_X1 U15380 ( .A(n20170), .B(n19923), .ZN(n13384) );
  XOR2_X1 U15381 ( .A(n13384), .B(n13385), .Z(n13386) );
  XNOR2_X2 U15382 ( .A(n13387), .B(n13386), .ZN(n14729) );
  NAND2_X1 U15383 ( .A1(n14224), .A2(n14729), .ZN(n14227) );
  XNOR2_X1 U15384 ( .A(n13391), .B(n13390), .ZN(n13393) );
  INV_X1 U15386 ( .A(n14410), .ZN(n14730) );
  NOR2_X1 U15387 ( .A1(n20451), .A2(n14730), .ZN(n13403) );
  XNOR2_X1 U15388 ( .A(n13397), .B(n20469), .ZN(n13570) );
  XNOR2_X1 U15389 ( .A(n13398), .B(n18420), .ZN(n13399) );
  XNOR2_X1 U15390 ( .A(n13400), .B(n13399), .ZN(n13401) );
  INV_X1 U15391 ( .A(n14137), .ZN(n13953) );
  XNOR2_X1 U15392 ( .A(n13601), .B(n18997), .ZN(n13407) );
  XNOR2_X1 U15393 ( .A(n13404), .B(n13405), .ZN(n13406) );
  XNOR2_X1 U15394 ( .A(n13407), .B(n13406), .ZN(n13413) );
  XNOR2_X1 U15395 ( .A(n20489), .B(n13658), .ZN(n13411) );
  XNOR2_X1 U15396 ( .A(n13409), .B(n13596), .ZN(n13410) );
  XNOR2_X1 U15397 ( .A(n13411), .B(n13410), .ZN(n13412) );
  XNOR2_X1 U15398 ( .A(n13413), .B(n13412), .ZN(n14724) );
  XNOR2_X1 U15400 ( .A(n13415), .B(n13416), .ZN(n13421) );
  XNOR2_X1 U15401 ( .A(n19721), .B(n15479), .ZN(n13419) );
  INV_X1 U15402 ( .A(n13417), .ZN(n13418) );
  XNOR2_X1 U15403 ( .A(n13419), .B(n13418), .ZN(n13420) );
  XNOR2_X1 U15404 ( .A(n13422), .B(n2410), .ZN(n13424) );
  XNOR2_X1 U15405 ( .A(n13462), .B(n13756), .ZN(n13423) );
  XNOR2_X1 U15406 ( .A(n13424), .B(n13423), .ZN(n13430) );
  INV_X1 U15407 ( .A(n13425), .ZN(n13426) );
  XNOR2_X1 U15408 ( .A(n13426), .B(n13427), .ZN(n13652) );
  XNOR2_X1 U15409 ( .A(n13652), .B(n13428), .ZN(n13429) );
  XNOR2_X1 U15410 ( .A(n13430), .B(n13429), .ZN(n14553) );
  AND2_X1 U15411 ( .A1(n14553), .A2(n14679), .ZN(n14552) );
  INV_X1 U15412 ( .A(n14552), .ZN(n14682) );
  INV_X1 U15413 ( .A(n13431), .ZN(n13797) );
  XNOR2_X1 U15414 ( .A(n13434), .B(n13433), .ZN(n13435) );
  XNOR2_X1 U15415 ( .A(n13435), .B(n13436), .ZN(n14279) );
  INV_X1 U15416 ( .A(n14279), .ZN(n13976) );
  XNOR2_X1 U15417 ( .A(n13767), .B(n13657), .ZN(n13438) );
  XNOR2_X1 U15418 ( .A(n13438), .B(n13437), .ZN(n13442) );
  XNOR2_X1 U15419 ( .A(n13710), .B(n2208), .ZN(n13439) );
  XNOR2_X1 U15420 ( .A(n13440), .B(n13439), .ZN(n13441) );
  NAND2_X1 U15422 ( .A1(n13976), .A2(n14555), .ZN(n14680) );
  NAND2_X1 U15423 ( .A1(n14682), .A2(n14680), .ZN(n13459) );
  INV_X1 U15424 ( .A(n13443), .ZN(n13445) );
  XNOR2_X1 U15425 ( .A(n13444), .B(n13445), .ZN(n13450) );
  XNOR2_X1 U15426 ( .A(n13446), .B(n17170), .ZN(n13448) );
  XNOR2_X1 U15427 ( .A(n13448), .B(n13447), .ZN(n13449) );
  INV_X1 U15428 ( .A(n14554), .ZN(n14678) );
  XNOR2_X1 U15429 ( .A(n13451), .B(n2108), .ZN(n13452) );
  XNOR2_X1 U15430 ( .A(n13452), .B(n19854), .ZN(n13455) );
  XNOR2_X1 U15431 ( .A(n13703), .B(n13453), .ZN(n13454) );
  XOR2_X1 U15432 ( .A(n13455), .B(n13454), .Z(n13456) );
  XNOR2_X1 U15433 ( .A(n13456), .B(n13457), .ZN(n14556) );
  OAI21_X1 U15434 ( .B1(n14677), .B2(n14279), .A(n14555), .ZN(n13458) );
  INV_X1 U15435 ( .A(n14553), .ZN(n14550) );
  XNOR2_X1 U15437 ( .A(n13462), .B(n13651), .ZN(n13685) );
  XNOR2_X1 U15438 ( .A(n13463), .B(n13685), .ZN(n13467) );
  XNOR2_X1 U15439 ( .A(n13849), .B(n17095), .ZN(n13465) );
  XNOR2_X1 U15441 ( .A(n13623), .B(n484), .ZN(n13469) );
  INV_X1 U15442 ( .A(n13471), .ZN(n13472) );
  XNOR2_X1 U15443 ( .A(n13703), .B(n13474), .ZN(n13476) );
  XNOR2_X1 U15444 ( .A(n13475), .B(n13476), .ZN(n13478) );
  INV_X1 U15445 ( .A(n13479), .ZN(n13480) );
  XNOR2_X1 U15446 ( .A(n13480), .B(n13481), .ZN(n13482) );
  XNOR2_X1 U15447 ( .A(n13483), .B(n13482), .ZN(n13488) );
  XNOR2_X1 U15448 ( .A(n13484), .B(n404), .ZN(n13485) );
  XNOR2_X1 U15449 ( .A(n13486), .B(n13485), .ZN(n13487) );
  INV_X1 U15450 ( .A(n14426), .ZN(n14494) );
  NOR2_X1 U15451 ( .A1(n14494), .A2(n14424), .ZN(n14749) );
  XNOR2_X1 U15452 ( .A(n13490), .B(n13489), .ZN(n13496) );
  XNOR2_X1 U15453 ( .A(n13491), .B(n13747), .ZN(n13494) );
  INV_X1 U15454 ( .A(n13518), .ZN(n13492) );
  XNOR2_X1 U15455 ( .A(n13492), .B(n18848), .ZN(n13493) );
  XNOR2_X1 U15456 ( .A(n13494), .B(n13493), .ZN(n13495) );
  XNOR2_X1 U15457 ( .A(n13495), .B(n13496), .ZN(n14493) );
  INV_X1 U15458 ( .A(n14425), .ZN(n14427) );
  NOR2_X1 U15459 ( .A1(n14427), .A2(n19728), .ZN(n13504) );
  INV_X1 U15460 ( .A(n13497), .ZN(n13498) );
  XNOR2_X1 U15461 ( .A(n13499), .B(n13498), .ZN(n13503) );
  XNOR2_X1 U15462 ( .A(n13543), .B(n18177), .ZN(n13500) );
  XNOR2_X1 U15463 ( .A(n13501), .B(n13500), .ZN(n13502) );
  AOI22_X1 U15464 ( .A1(n14749), .A2(n1936), .B1(n13504), .B2(n14753), .ZN(
        n13505) );
  MUX2_X1 U15465 ( .A(n19742), .B(n14499), .S(n14305), .Z(n13509) );
  NOR2_X1 U15467 ( .A1(n15457), .A2(n19759), .ZN(n13561) );
  XNOR2_X1 U15468 ( .A(n13753), .B(n13510), .ZN(n13516) );
  XNOR2_X1 U15469 ( .A(n19869), .B(n18801), .ZN(n13513) );
  XNOR2_X1 U15470 ( .A(n13518), .B(n13517), .ZN(n13521) );
  XNOR2_X1 U15471 ( .A(n19892), .B(n2383), .ZN(n13520) );
  XNOR2_X1 U15472 ( .A(n13523), .B(n13522), .ZN(n13524) );
  XNOR2_X1 U15473 ( .A(n13524), .B(n13744), .ZN(n14434) );
  INV_X1 U15474 ( .A(n13525), .ZN(n13526) );
  XNOR2_X1 U15475 ( .A(n13526), .B(n13527), .ZN(n13532) );
  XNOR2_X1 U15476 ( .A(n13528), .B(n17637), .ZN(n13529) );
  XNOR2_X1 U15477 ( .A(n13530), .B(n13529), .ZN(n13531) );
  XNOR2_X1 U15478 ( .A(n13532), .B(n13531), .ZN(n14435) );
  XNOR2_X1 U15480 ( .A(n13533), .B(n13761), .ZN(n13538) );
  XNOR2_X1 U15481 ( .A(n20482), .B(n17791), .ZN(n13535) );
  XNOR2_X1 U15482 ( .A(n13536), .B(n13535), .ZN(n13537) );
  XNOR2_X1 U15483 ( .A(n13538), .B(n13537), .ZN(n14172) );
  OAI21_X1 U15484 ( .B1(n14487), .B2(n20263), .A(n14172), .ZN(n13555) );
  XNOR2_X1 U15487 ( .A(n13771), .B(n13542), .ZN(n13548) );
  XNOR2_X1 U15488 ( .A(n13601), .B(n16030), .ZN(n13546) );
  XNOR2_X1 U15489 ( .A(n13544), .B(n13543), .ZN(n13545) );
  XNOR2_X1 U15490 ( .A(n13545), .B(n13546), .ZN(n13547) );
  INV_X1 U15491 ( .A(n14172), .ZN(n14480) );
  XNOR2_X1 U15492 ( .A(n13792), .B(n2067), .ZN(n13549) );
  XNOR2_X1 U15493 ( .A(n13551), .B(n13550), .ZN(n13552) );
  XNOR2_X1 U15494 ( .A(n13552), .B(n13553), .ZN(n14171) );
  NAND2_X1 U15495 ( .A1(n14435), .A2(n14171), .ZN(n14302) );
  OAI21_X1 U15496 ( .B1(n3516), .B2(n14167), .A(n14442), .ZN(n13558) );
  NOR2_X1 U15497 ( .A1(n701), .A2(n13918), .ZN(n14440) );
  NAND3_X1 U15498 ( .A1(n3516), .A2(n20262), .A3(n14441), .ZN(n13556) );
  OAI21_X1 U15499 ( .B1(n14448), .B2(n14447), .A(n14451), .ZN(n13560) );
  INV_X1 U15502 ( .A(n15457), .ZN(n15460) );
  AOI21_X1 U15503 ( .B1(n15353), .B2(n13566), .A(n15460), .ZN(n13567) );
  NOR2_X2 U15504 ( .A1(n13568), .A2(n13567), .ZN(n16601) );
  INV_X1 U15505 ( .A(n13569), .ZN(n13571) );
  XNOR2_X1 U15506 ( .A(n13571), .B(n13570), .ZN(n13575) );
  XNOR2_X1 U15507 ( .A(n13572), .B(n19436), .ZN(n13574) );
  XNOR2_X1 U15508 ( .A(n13577), .B(n13576), .ZN(n13578) );
  XNOR2_X1 U15509 ( .A(n13579), .B(n13578), .ZN(n13583) );
  XNOR2_X1 U15510 ( .A(n13580), .B(n649), .ZN(n13581) );
  XNOR2_X1 U15511 ( .A(n13584), .B(n13517), .ZN(n13587) );
  XNOR2_X1 U15512 ( .A(n13746), .B(n13585), .ZN(n13586) );
  XNOR2_X1 U15513 ( .A(n13587), .B(n13586), .ZN(n13594) );
  XNOR2_X1 U15514 ( .A(n13491), .B(n2055), .ZN(n13592) );
  INV_X1 U15515 ( .A(n13588), .ZN(n13589) );
  XNOR2_X1 U15516 ( .A(n13590), .B(n13589), .ZN(n13591) );
  XNOR2_X1 U15517 ( .A(n13592), .B(n13591), .ZN(n13593) );
  NOR2_X1 U15519 ( .A1(n13994), .A2(n13996), .ZN(n13630) );
  INV_X1 U15521 ( .A(n13596), .ZN(n13597) );
  XNOR2_X1 U15522 ( .A(n13597), .B(n13767), .ZN(n13598) );
  XNOR2_X1 U15524 ( .A(n19904), .B(n13601), .ZN(n13604) );
  XNOR2_X1 U15525 ( .A(n13602), .B(n16424), .ZN(n13603) );
  XNOR2_X1 U15526 ( .A(n13604), .B(n13603), .ZN(n13605) );
  XNOR2_X1 U15527 ( .A(n13606), .B(n13605), .ZN(n14153) );
  INV_X1 U15528 ( .A(n14153), .ZN(n14594) );
  XNOR2_X1 U15529 ( .A(n13608), .B(n13607), .ZN(n13609) );
  XNOR2_X1 U15530 ( .A(n13610), .B(n13609), .ZN(n13614) );
  XNOR2_X1 U15531 ( .A(n13797), .B(n2337), .ZN(n13611) );
  XNOR2_X1 U15532 ( .A(n13612), .B(n13611), .ZN(n13613) );
  XNOR2_X1 U15533 ( .A(n13614), .B(n13613), .ZN(n14395) );
  AND2_X1 U15537 ( .A1(n13615), .A2(n14156), .ZN(n13629) );
  XNOR2_X1 U15538 ( .A(n13617), .B(n13616), .ZN(n13621) );
  XNOR2_X1 U15539 ( .A(n20170), .B(n13618), .ZN(n13620) );
  XNOR2_X1 U15540 ( .A(n13621), .B(n13620), .ZN(n13628) );
  XNOR2_X1 U15541 ( .A(n13622), .B(n18203), .ZN(n13626) );
  XNOR2_X1 U15542 ( .A(n13624), .B(n13623), .ZN(n13625) );
  XNOR2_X1 U15543 ( .A(n13626), .B(n13625), .ZN(n13627) );
  INV_X1 U15545 ( .A(n13631), .ZN(n13632) );
  XNOR2_X1 U15547 ( .A(n20260), .B(n13635), .ZN(n13637) );
  XNOR2_X1 U15548 ( .A(n13637), .B(n13636), .ZN(n13638) );
  INV_X1 U15549 ( .A(n14388), .ZN(n14715) );
  XNOR2_X1 U15550 ( .A(n13641), .B(n13640), .ZN(n13648) );
  XNOR2_X1 U15551 ( .A(n13643), .B(n13642), .ZN(n13646) );
  XNOR2_X1 U15552 ( .A(n13644), .B(n2394), .ZN(n13645) );
  XNOR2_X1 U15553 ( .A(n13646), .B(n13645), .ZN(n13647) );
  XNOR2_X1 U15554 ( .A(n13648), .B(n13647), .ZN(n14716) );
  NAND2_X1 U15555 ( .A1(n14715), .A2(n14716), .ZN(n14389) );
  XNOR2_X1 U15556 ( .A(n13651), .B(n17060), .ZN(n13653) );
  XNOR2_X1 U15557 ( .A(n13652), .B(n13653), .ZN(n13654) );
  XNOR2_X1 U15558 ( .A(n13656), .B(n13655), .ZN(n13663) );
  XNOR2_X1 U15559 ( .A(n13658), .B(n13657), .ZN(n13661) );
  XNOR2_X1 U15560 ( .A(n13659), .B(n17365), .ZN(n13660) );
  XNOR2_X1 U15561 ( .A(n13661), .B(n13660), .ZN(n13662) );
  NAND2_X1 U15563 ( .A1(n20213), .A2(n19843), .ZN(n13664) );
  OAI21_X1 U15564 ( .B1(n14389), .B2(n19843), .A(n13664), .ZN(n13683) );
  XNOR2_X1 U15565 ( .A(n13666), .B(n13665), .ZN(n13670) );
  XNOR2_X1 U15566 ( .A(n13827), .B(n2221), .ZN(n13667) );
  XNOR2_X1 U15567 ( .A(n13668), .B(n13667), .ZN(n13669) );
  NAND2_X1 U15568 ( .A1(n14716), .A2(n14717), .ZN(n13682) );
  XNOR2_X1 U15569 ( .A(n13833), .B(n13672), .ZN(n13675) );
  XNOR2_X1 U15570 ( .A(n13673), .B(n1996), .ZN(n13674) );
  XNOR2_X1 U15571 ( .A(n13675), .B(n13674), .ZN(n13681) );
  INV_X1 U15572 ( .A(n13676), .ZN(n13679) );
  XNOR2_X1 U15573 ( .A(n13734), .B(n13677), .ZN(n13678) );
  XNOR2_X1 U15574 ( .A(n13679), .B(n13678), .ZN(n13680) );
  INV_X1 U15575 ( .A(n14718), .ZN(n13963) );
  XNOR2_X1 U15577 ( .A(n13684), .B(n13685), .ZN(n13692) );
  XNOR2_X1 U15578 ( .A(n13686), .B(n13687), .ZN(n13690) );
  XNOR2_X1 U15579 ( .A(n13688), .B(n18366), .ZN(n13689) );
  XNOR2_X1 U15580 ( .A(n13690), .B(n13689), .ZN(n13691) );
  INV_X1 U15581 ( .A(n14378), .ZN(n14232) );
  XNOR2_X1 U15582 ( .A(n13694), .B(n13693), .ZN(n13701) );
  XNOR2_X1 U15585 ( .A(n13699), .B(n13698), .ZN(n13700) );
  XNOR2_X1 U15586 ( .A(n13701), .B(n13700), .ZN(n14700) );
  NOR2_X1 U15587 ( .A1(n14232), .A2(n14700), .ZN(n13731) );
  XNOR2_X1 U15588 ( .A(n20155), .B(n13703), .ZN(n13704) );
  INV_X1 U15589 ( .A(n915), .ZN(n13705) );
  XNOR2_X1 U15590 ( .A(n13707), .B(n13706), .ZN(n13709) );
  XNOR2_X1 U15591 ( .A(n13710), .B(n18308), .ZN(n13712) );
  XNOR2_X1 U15592 ( .A(n13712), .B(n13711), .ZN(n13713) );
  XNOR2_X1 U15593 ( .A(n13714), .B(n13713), .ZN(n13720) );
  XNOR2_X1 U15594 ( .A(n13716), .B(n13715), .ZN(n13718) );
  XNOR2_X1 U15595 ( .A(n13718), .B(n13717), .ZN(n13719) );
  NOR2_X1 U15596 ( .A1(n14120), .A2(n14228), .ZN(n13730) );
  XNOR2_X1 U15597 ( .A(n19721), .B(n2248), .ZN(n13723) );
  XNOR2_X1 U15598 ( .A(n13722), .B(n13723), .ZN(n13729) );
  XNOR2_X1 U15599 ( .A(n13724), .B(n13725), .ZN(n13726) );
  XNOR2_X1 U15600 ( .A(n13727), .B(n13726), .ZN(n13728) );
  XNOR2_X1 U15602 ( .A(n13733), .B(n13732), .ZN(n13740) );
  XNOR2_X1 U15603 ( .A(n13735), .B(n13734), .ZN(n13738) );
  INV_X1 U15604 ( .A(n1148), .ZN(n18587) );
  XNOR2_X1 U15605 ( .A(n13736), .B(n18587), .ZN(n13737) );
  XNOR2_X1 U15606 ( .A(n13738), .B(n13737), .ZN(n13739) );
  MUX2_X1 U15607 ( .A(n2769), .B(n14230), .S(n240), .Z(n13741) );
  NOR2_X1 U15608 ( .A1(n13741), .A2(n20204), .ZN(n13742) );
  NAND2_X1 U15609 ( .A1(n15228), .A2(n15677), .ZN(n15229) );
  OAI21_X1 U15610 ( .B1(n2005), .B2(n15679), .A(n15229), .ZN(n13806) );
  INV_X1 U15611 ( .A(n13744), .ZN(n13752) );
  XNOR2_X1 U15612 ( .A(n13746), .B(n13745), .ZN(n13749) );
  XNOR2_X1 U15613 ( .A(n13747), .B(n2032), .ZN(n13748) );
  XNOR2_X1 U15614 ( .A(n13751), .B(n13752), .ZN(n14406) );
  INV_X1 U15615 ( .A(n14406), .ZN(n14149) );
  XNOR2_X1 U15616 ( .A(n13755), .B(n18830), .ZN(n13759) );
  XNOR2_X1 U15617 ( .A(n13757), .B(n13756), .ZN(n13758) );
  XNOR2_X1 U15618 ( .A(n13761), .B(n13760), .ZN(n13766) );
  XNOR2_X1 U15619 ( .A(n13762), .B(n18090), .ZN(n13763) );
  XNOR2_X1 U15620 ( .A(n13764), .B(n13763), .ZN(n13765) );
  INV_X1 U15622 ( .A(n19907), .ZN(n14405) );
  NOR2_X1 U15623 ( .A1(n14148), .A2(n14405), .ZN(n13789) );
  XNOR2_X1 U15624 ( .A(n13768), .B(n13767), .ZN(n13770) );
  XNOR2_X1 U15625 ( .A(n13772), .B(n18070), .ZN(n13773) );
  INV_X1 U15626 ( .A(n13774), .ZN(n13775) );
  XNOR2_X1 U15627 ( .A(n13776), .B(n13775), .ZN(n13780) );
  XNOR2_X1 U15628 ( .A(n13778), .B(n19854), .ZN(n13779) );
  XNOR2_X1 U15629 ( .A(n13780), .B(n13779), .ZN(n13787) );
  XNOR2_X1 U15630 ( .A(n19797), .B(n915), .ZN(n13785) );
  XNOR2_X1 U15631 ( .A(n13783), .B(n2349), .ZN(n13784) );
  XNOR2_X1 U15632 ( .A(n13785), .B(n13784), .ZN(n13786) );
  XNOR2_X1 U15633 ( .A(n13787), .B(n13786), .ZN(n14112) );
  INV_X1 U15634 ( .A(n14112), .ZN(n14238) );
  NOR2_X1 U15635 ( .A1(n14236), .A2(n14238), .ZN(n13788) );
  AOI22_X1 U15636 ( .A1(n14149), .A2(n13789), .B1(n14405), .B2(n13788), .ZN(
        n13804) );
  XNOR2_X1 U15637 ( .A(n13790), .B(n13791), .ZN(n13794) );
  XNOR2_X1 U15638 ( .A(n13794), .B(n13793), .ZN(n13801) );
  XNOR2_X1 U15639 ( .A(n19946), .B(n13795), .ZN(n13799) );
  XNOR2_X1 U15640 ( .A(n13797), .B(n18304), .ZN(n13798) );
  XNOR2_X1 U15641 ( .A(n13799), .B(n13798), .ZN(n13800) );
  INV_X1 U15642 ( .A(n14239), .ZN(n14403) );
  MUX2_X1 U15643 ( .A(n19908), .B(n14238), .S(n14403), .Z(n13802) );
  NAND2_X1 U15644 ( .A1(n15682), .A2(n15442), .ZN(n13805) );
  NAND2_X1 U15645 ( .A1(n13806), .A2(n13805), .ZN(n13863) );
  INV_X1 U15646 ( .A(n13807), .ZN(n13809) );
  XNOR2_X1 U15647 ( .A(n13809), .B(n13808), .ZN(n13814) );
  XNOR2_X1 U15648 ( .A(n13810), .B(n19410), .ZN(n13811) );
  XNOR2_X1 U15649 ( .A(n13812), .B(n13811), .ZN(n13813) );
  XNOR2_X1 U15650 ( .A(n13816), .B(n13815), .ZN(n13822) );
  INV_X1 U15651 ( .A(n13817), .ZN(n13820) );
  XNOR2_X1 U15652 ( .A(n13818), .B(n18338), .ZN(n13819) );
  XNOR2_X1 U15653 ( .A(n13820), .B(n13819), .ZN(n13821) );
  INV_X1 U15654 ( .A(n13823), .ZN(n13825) );
  XNOR2_X1 U15655 ( .A(n13825), .B(n13824), .ZN(n13832) );
  INV_X1 U15656 ( .A(n13826), .ZN(n13828) );
  XNOR2_X1 U15657 ( .A(n13827), .B(n13828), .ZN(n13830) );
  XNOR2_X1 U15658 ( .A(n13830), .B(n13829), .ZN(n13831) );
  XNOR2_X2 U15659 ( .A(n13832), .B(n13831), .ZN(n14599) );
  XNOR2_X1 U15660 ( .A(n13834), .B(n13833), .ZN(n13837) );
  XNOR2_X1 U15661 ( .A(n20223), .B(n1911), .ZN(n13836) );
  XNOR2_X1 U15662 ( .A(n13837), .B(n13836), .ZN(n13841) );
  XNOR2_X1 U15663 ( .A(n13839), .B(n13838), .ZN(n13840) );
  XNOR2_X1 U15664 ( .A(n13840), .B(n13841), .ZN(n14249) );
  INV_X1 U15665 ( .A(n13844), .ZN(n13845) );
  XNOR2_X1 U15666 ( .A(n13845), .B(n13846), .ZN(n13847) );
  XNOR2_X1 U15667 ( .A(n13849), .B(n18278), .ZN(n13850) );
  XNOR2_X1 U15668 ( .A(n13853), .B(n13852), .ZN(n13854) );
  INV_X1 U15670 ( .A(n15312), .ZN(n13861) );
  INV_X1 U15671 ( .A(n13856), .ZN(n13857) );
  OAI21_X1 U15672 ( .B1(n13857), .B2(n14146), .A(n19875), .ZN(n13858) );
  INV_X1 U15673 ( .A(n15676), .ZN(n13859) );
  OAI21_X1 U15674 ( .B1(n13859), .B2(n15442), .A(n15679), .ZN(n13860) );
  XOR2_X1 U15675 ( .A(n16601), .B(n17288), .Z(n13864) );
  INV_X1 U15676 ( .A(n17223), .ZN(n16634) );
  MUX2_X1 U15677 ( .A(n15120), .B(n14520), .S(n14516), .Z(n13867) );
  NAND2_X1 U15678 ( .A1(n14186), .A2(n14520), .ZN(n13866) );
  NAND2_X1 U15679 ( .A1(n14499), .A2(n14497), .ZN(n14306) );
  NOR2_X1 U15680 ( .A1(n19742), .A2(n13868), .ZN(n13871) );
  NAND2_X1 U15681 ( .A1(n14305), .A2(n14307), .ZN(n13870) );
  MUX2_X1 U15682 ( .A(n19634), .B(n19831), .S(n14648), .Z(n13875) );
  AOI21_X1 U15683 ( .B1(n20380), .B2(n14651), .A(n237), .ZN(n13874) );
  NAND2_X1 U15684 ( .A1(n14648), .A2(n14524), .ZN(n13873) );
  INV_X1 U15685 ( .A(n14042), .ZN(n13887) );
  NOR2_X1 U15686 ( .A1(n15500), .A2(n19512), .ZN(n15160) );
  INV_X1 U15687 ( .A(n15500), .ZN(n15497) );
  INV_X1 U15688 ( .A(n14753), .ZN(n13880) );
  NAND2_X1 U15689 ( .A1(n14427), .A2(n19727), .ZN(n14750) );
  OAI21_X1 U15690 ( .B1(n14494), .B2(n19727), .A(n14750), .ZN(n13879) );
  NAND3_X1 U15691 ( .A1(n14494), .A2(n14424), .A3(n1936), .ZN(n13876) );
  OAI21_X1 U15692 ( .B1(n13877), .B2(n3156), .A(n13876), .ZN(n13878) );
  INV_X1 U15693 ( .A(n15195), .ZN(n14041) );
  NOR2_X1 U15694 ( .A1(n14482), .A2(n14435), .ZN(n13882) );
  MUX2_X1 U15695 ( .A(n13882), .B(n13881), .S(n14480), .Z(n13885) );
  INV_X1 U15696 ( .A(n14171), .ZN(n14483) );
  NOR3_X1 U15697 ( .A1(n14431), .A2(n13883), .A3(n14487), .ZN(n13884) );
  NOR2_X2 U15698 ( .A1(n13885), .A2(n13884), .ZN(n15501) );
  OAI211_X1 U15699 ( .C1(n15497), .C2(n14041), .A(n15501), .B(n15192), .ZN(
        n13886) );
  XNOR2_X1 U15700 ( .A(n16587), .B(n17686), .ZN(n13945) );
  NOR2_X1 U15701 ( .A1(n14813), .A2(n14807), .ZN(n13888) );
  NAND2_X1 U15702 ( .A1(n14199), .A2(n14810), .ZN(n14141) );
  MUX2_X1 U15703 ( .A(n14811), .B(n19781), .S(n14199), .Z(n13889) );
  NOR2_X1 U15704 ( .A1(n13889), .A2(n14812), .ZN(n13890) );
  NOR2_X1 U15705 ( .A1(n20500), .A2(n14800), .ZN(n13896) );
  NAND2_X1 U15706 ( .A1(n13893), .A2(n3497), .ZN(n13895) );
  INV_X1 U15707 ( .A(n14787), .ZN(n14346) );
  NOR2_X1 U15708 ( .A1(n14791), .A2(n12627), .ZN(n13900) );
  NOR2_X1 U15709 ( .A1(n14346), .A2(n12627), .ZN(n14100) );
  NAND2_X1 U15710 ( .A1(n14100), .A2(n14788), .ZN(n13899) );
  NAND2_X1 U15711 ( .A1(n14789), .A2(n12627), .ZN(n13898) );
  OAI211_X1 U15712 ( .C1(n14102), .C2(n13900), .A(n13899), .B(n13898), .ZN(
        n15861) );
  INV_X1 U15713 ( .A(n15861), .ZN(n15327) );
  INV_X1 U15714 ( .A(n13901), .ZN(n14076) );
  NOR2_X1 U15715 ( .A1(n877), .A2(n14076), .ZN(n13904) );
  NAND2_X1 U15716 ( .A1(n14077), .A2(n14782), .ZN(n13903) );
  NAND2_X1 U15718 ( .A1(n20408), .A2(n14076), .ZN(n13902) );
  INV_X1 U15719 ( .A(n14779), .ZN(n14216) );
  NOR2_X1 U15720 ( .A1(n13905), .A2(n14216), .ZN(n13906) );
  AOI21_X1 U15721 ( .B1(n14612), .B2(n14206), .A(n13908), .ZN(n13911) );
  INV_X1 U15722 ( .A(n14011), .ZN(n13907) );
  INV_X1 U15723 ( .A(n13909), .ZN(n14142) );
  OAI21_X1 U15724 ( .B1(n14207), .B2(n14142), .A(n19488), .ZN(n13910) );
  NOR2_X1 U15725 ( .A1(n15866), .A2(n15863), .ZN(n13912) );
  INV_X1 U15727 ( .A(n14827), .ZN(n14073) );
  MUX2_X1 U15728 ( .A(n13914), .B(n13913), .S(n14073), .Z(n13915) );
  NOR2_X1 U15729 ( .A1(n15720), .A2(n15861), .ZN(n15721) );
  NOR2_X1 U15732 ( .A1(n13918), .A2(n14441), .ZN(n13919) );
  NOR2_X1 U15733 ( .A1(n13921), .A2(n14465), .ZN(n13923) );
  NOR2_X1 U15734 ( .A1(n14462), .A2(n14468), .ZN(n13922) );
  MUX2_X1 U15735 ( .A(n13923), .B(n13922), .S(n19657), .Z(n13926) );
  NAND2_X1 U15736 ( .A1(n13921), .A2(n14468), .ZN(n14363) );
  NAND2_X1 U15737 ( .A1(n1363), .A2(n14449), .ZN(n13928) );
  NAND2_X1 U15738 ( .A1(n14450), .A2(n14449), .ZN(n14182) );
  NAND3_X1 U15739 ( .A1(n14448), .A2(n14455), .A3(n14451), .ZN(n13929) );
  OAI21_X1 U15740 ( .B1(n14182), .B2(n14453), .A(n13929), .ZN(n14755) );
  OAI21_X1 U15741 ( .B1(n13930), .B2(n14335), .A(n14092), .ZN(n13932) );
  NOR2_X1 U15742 ( .A1(n14424), .A2(n1936), .ZN(n13936) );
  OAI211_X1 U15743 ( .C1(n14424), .C2(n14493), .A(n19728), .B(n14753), .ZN(
        n13935) );
  NOR3_X1 U15744 ( .A1(n15187), .A2(n15505), .A3(n13933), .ZN(n13943) );
  NOR2_X1 U15745 ( .A1(n13939), .A2(n14359), .ZN(n13941) );
  NOR2_X1 U15746 ( .A1(n14054), .A2(n14357), .ZN(n14757) );
  NAND3_X1 U15747 ( .A1(n15187), .A2(n15188), .A3(n15507), .ZN(n13942) );
  XNOR2_X1 U15748 ( .A(n16931), .B(n19659), .ZN(n13944) );
  XNOR2_X1 U15749 ( .A(n13945), .B(n13944), .ZN(n14018) );
  INV_X1 U15750 ( .A(n13946), .ZN(n14691) );
  MUX2_X1 U15751 ( .A(n14385), .B(n19895), .S(n14691), .Z(n13948) );
  NAND2_X1 U15752 ( .A1(n14693), .A2(n14688), .ZN(n13947) );
  INV_X1 U15753 ( .A(n14021), .ZN(n14289) );
  INV_X1 U15754 ( .A(n15153), .ZN(n16012) );
  NOR2_X1 U15755 ( .A1(n14223), .A2(n14729), .ZN(n13952) );
  NOR2_X1 U15756 ( .A1(n14273), .A2(n14275), .ZN(n13954) );
  OAI21_X1 U15757 ( .B1(n13955), .B2(n13954), .A(n2282), .ZN(n13958) );
  NAND3_X1 U15758 ( .A1(n14705), .A2(n14563), .A3(n14566), .ZN(n13956) );
  INV_X1 U15760 ( .A(n15705), .ZN(n13961) );
  NAND3_X1 U15761 ( .A1(n14736), .A2(n14571), .A3(n14269), .ZN(n13960) );
  NAND3_X1 U15762 ( .A1(n14740), .A2(n20157), .A3(n14570), .ZN(n13959) );
  INV_X1 U15763 ( .A(n20119), .ZN(n15152) );
  MUX2_X1 U15764 ( .A(n13963), .B(n20213), .S(n3057), .Z(n13965) );
  NAND2_X1 U15765 ( .A1(n19843), .A2(n14715), .ZN(n13964) );
  NAND3_X1 U15766 ( .A1(n13965), .A2(n14389), .A3(n13964), .ZN(n13967) );
  NAND2_X1 U15767 ( .A1(n14716), .A2(n19862), .ZN(n13966) );
  AND2_X2 U15768 ( .A1(n13967), .A2(n13966), .ZN(n16009) );
  INV_X1 U15769 ( .A(n16009), .ZN(n13968) );
  INV_X1 U15770 ( .A(n17281), .ZN(n13992) );
  NOR2_X1 U15771 ( .A1(n14651), .A2(n14522), .ZN(n13971) );
  NAND2_X1 U15773 ( .A1(n14677), .A2(n13976), .ZN(n13979) );
  INV_X1 U15774 ( .A(n14679), .ZN(n14557) );
  AOI21_X1 U15775 ( .B1(n14554), .B2(n14553), .A(n14557), .ZN(n13977) );
  INV_X1 U15777 ( .A(n14281), .ZN(n14284) );
  NAND3_X1 U15779 ( .A1(n15870), .A2(n20178), .A3(n13989), .ZN(n13991) );
  INV_X1 U15780 ( .A(n14032), .ZN(n14640) );
  INV_X1 U15782 ( .A(n14642), .ZN(n13983) );
  NOR2_X1 U15783 ( .A1(n20473), .A2(n13983), .ZN(n13984) );
  MUX2_X1 U15784 ( .A(n13985), .B(n13984), .S(n19703), .Z(n13988) );
  INV_X1 U15785 ( .A(n14512), .ZN(n14034) );
  OAI22_X1 U15786 ( .A1(n14508), .A2(n14034), .B1(n13986), .B2(n14642), .ZN(
        n13987) );
  NOR2_X2 U15787 ( .A1(n13988), .A2(n13987), .ZN(n15875) );
  INV_X1 U15788 ( .A(n15875), .ZN(n15148) );
  NOR2_X1 U15789 ( .A1(n15876), .A2(n15709), .ZN(n15303) );
  XNOR2_X1 U15790 ( .A(n13992), .B(n16566), .ZN(n16713) );
  NAND2_X1 U15791 ( .A1(n15028), .A2(n15380), .ZN(n14874) );
  INV_X1 U15792 ( .A(n14874), .ZN(n15170) );
  NOR2_X1 U15793 ( .A1(n19513), .A2(n231), .ZN(n14872) );
  OAI21_X1 U15794 ( .B1(n15167), .B2(n15380), .A(n14872), .ZN(n13993) );
  MUX2_X1 U15796 ( .A(n19709), .B(n13994), .S(n14395), .Z(n13999) );
  NOR2_X1 U15797 ( .A1(n14594), .A2(n14396), .ZN(n13997) );
  MUX2_X1 U15798 ( .A(n13997), .B(n13996), .S(n19731), .Z(n13998) );
  AOI22_X1 U15799 ( .A1(n954), .A2(n14624), .B1(n15314), .B2(n14623), .ZN(
        n14004) );
  NOR2_X1 U15800 ( .A1(n14627), .A2(n14624), .ZN(n14003) );
  NAND3_X1 U15801 ( .A1(n14001), .A2(n14620), .A3(n14146), .ZN(n14002) );
  INV_X1 U15803 ( .A(n15695), .ZN(n15138) );
  NAND2_X1 U15804 ( .A1(n15701), .A2(n15138), .ZN(n14016) );
  NAND2_X1 U15805 ( .A1(n14381), .A2(n20204), .ZN(n14005) );
  OAI21_X1 U15806 ( .B1(n14120), .B2(n14229), .A(n20480), .ZN(n14006) );
  NAND2_X1 U15808 ( .A1(n14238), .A2(n19908), .ZN(n14240) );
  OAI21_X1 U15809 ( .B1(n14238), .B2(n14148), .A(n14240), .ZN(n14007) );
  NOR2_X1 U15810 ( .A1(n20005), .A2(n15698), .ZN(n14015) );
  MUX2_X1 U15811 ( .A(n14203), .B(n13908), .S(n3225), .Z(n14014) );
  XNOR2_X1 U15814 ( .A(n17275), .B(n16926), .ZN(n16523) );
  XNOR2_X1 U15815 ( .A(n16523), .B(n19903), .ZN(n14017) );
  XNOR2_X1 U15816 ( .A(n14017), .B(n14018), .ZN(n16633) );
  AOI21_X1 U15819 ( .B1(n14654), .B2(n241), .A(n14288), .ZN(n14025) );
  OAI211_X1 U15820 ( .C1(n14268), .C2(n14267), .A(n14269), .B(n1819), .ZN(
        n14027) );
  NAND2_X1 U15821 ( .A1(n14578), .A2(n14268), .ZN(n15487) );
  OAI21_X1 U15822 ( .B1(n15756), .B2(n15754), .A(n15758), .ZN(n14040) );
  MUX2_X1 U15823 ( .A(n14677), .B(n14554), .S(n14550), .Z(n14030) );
  INV_X1 U15824 ( .A(n14555), .ZN(n14028) );
  MUX2_X1 U15825 ( .A(n14279), .B(n14028), .S(n14677), .Z(n14029) );
  OAI21_X1 U15826 ( .B1(n14032), .B2(n14031), .A(n20473), .ZN(n14033) );
  NAND2_X1 U15827 ( .A1(n15491), .A2(n15760), .ZN(n14039) );
  NOR2_X1 U15828 ( .A1(n14667), .A2(n14662), .ZN(n14035) );
  NAND3_X1 U15829 ( .A1(n14663), .A2(n14316), .A3(n14664), .ZN(n14036) );
  AND3_X1 U15830 ( .A1(n14038), .A2(n14037), .A3(n14036), .ZN(n15490) );
  NOR2_X1 U15831 ( .A1(n15501), .A2(n15192), .ZN(n14930) );
  OAI21_X1 U15832 ( .B1(n14930), .B2(n15496), .A(n19813), .ZN(n14044) );
  NAND2_X1 U15833 ( .A1(n14042), .A2(n14041), .ZN(n14043) );
  NAND2_X1 U15834 ( .A1(n14044), .A2(n14043), .ZN(n16821) );
  XNOR2_X1 U15835 ( .A(n16821), .B(n16743), .ZN(n16396) );
  NOR2_X1 U15836 ( .A1(n14347), .A2(n14827), .ZN(n14045) );
  INV_X1 U15838 ( .A(n14049), .ZN(n14051) );
  AOI22_X2 U15839 ( .A1(n14341), .A2(n14051), .B1(n14093), .B2(n14050), .ZN(
        n15844) );
  NOR2_X1 U15840 ( .A1(n15845), .A2(n15844), .ZN(n14056) );
  NOR2_X1 U15841 ( .A1(n14419), .A2(n14357), .ZN(n14053) );
  OAI21_X1 U15843 ( .B1(n14056), .B2(n15266), .A(n15636), .ZN(n14068) );
  NAND2_X1 U15844 ( .A1(n20454), .A2(n14778), .ZN(n14058) );
  AOI21_X1 U15845 ( .B1(n14852), .B2(n14058), .A(n14057), .ZN(n14061) );
  NAND2_X1 U15846 ( .A1(n14076), .A2(n14778), .ZN(n14059) );
  AOI21_X1 U15847 ( .B1(n20454), .B2(n14059), .A(n14216), .ZN(n14060) );
  NOR2_X2 U15848 ( .A1(n14061), .A2(n14060), .ZN(n15846) );
  INV_X1 U15849 ( .A(n14788), .ZN(n14066) );
  MUX2_X1 U15850 ( .A(n14789), .B(n2412), .S(n14790), .Z(n14065) );
  NAND2_X1 U15852 ( .A1(n14791), .A2(n14792), .ZN(n14062) );
  MUX2_X1 U15853 ( .A(n14063), .B(n14062), .S(n14789), .Z(n14064) );
  NAND3_X1 U15854 ( .A1(n15847), .A2(n2146), .A3(n868), .ZN(n14067) );
  NOR2_X1 U15855 ( .A1(n15187), .A2(n15505), .ZN(n14069) );
  NOR2_X1 U15856 ( .A1(n15187), .A2(n1614), .ZN(n14070) );
  XNOR2_X1 U15858 ( .A(n16593), .B(n864), .ZN(n16185) );
  MUX2_X1 U15859 ( .A(n14073), .B(n14828), .S(n19496), .Z(n14075) );
  MUX2_X1 U15860 ( .A(n19859), .B(n19984), .S(n14827), .Z(n14074) );
  NAND2_X1 U15861 ( .A1(n14077), .A2(n14778), .ZN(n14078) );
  NOR2_X1 U15862 ( .A1(n14057), .A2(n20518), .ZN(n14079) );
  NAND2_X1 U15863 ( .A1(n14079), .A2(n14216), .ZN(n14080) );
  OAI21_X1 U15864 ( .B1(n14796), .B2(n14584), .A(n14799), .ZN(n14082) );
  INV_X1 U15865 ( .A(n15515), .ZN(n15745) );
  INV_X1 U15866 ( .A(n14085), .ZN(n14091) );
  INV_X1 U15867 ( .A(n14086), .ZN(n14089) );
  OAI211_X1 U15868 ( .C1(n19821), .C2(n14818), .A(n912), .B(n14326), .ZN(
        n14088) );
  AOI21_X1 U15869 ( .B1(n19485), .B2(n12876), .A(n14092), .ZN(n14098) );
  INV_X1 U15870 ( .A(n14093), .ZN(n14096) );
  NOR2_X1 U15871 ( .A1(n14336), .A2(n14335), .ZN(n14095) );
  NAND3_X1 U15873 ( .A1(n15521), .A2(n15516), .A3(n15741), .ZN(n14099) );
  OAI21_X1 U15874 ( .B1(n15748), .B2(n14982), .A(n14099), .ZN(n14108) );
  INV_X1 U15875 ( .A(n14100), .ZN(n14101) );
  NAND2_X1 U15876 ( .A1(n15746), .A2(n15516), .ZN(n15740) );
  INV_X1 U15877 ( .A(n15748), .ZN(n15181) );
  AOI21_X1 U15878 ( .B1(n15740), .B2(n15741), .A(n15181), .ZN(n14107) );
  MUX2_X1 U15879 ( .A(n14717), .B(n14718), .S(n3057), .Z(n14110) );
  MUX2_X1 U15880 ( .A(n14716), .B(n3057), .S(n13671), .Z(n14109) );
  NAND2_X1 U15882 ( .A1(n14239), .A2(n15423), .ZN(n14113) );
  MUX2_X1 U15883 ( .A(n14113), .B(n14240), .S(n14149), .Z(n14118) );
  INV_X1 U15884 ( .A(n14242), .ZN(n14116) );
  NOR2_X1 U15885 ( .A1(n14114), .A2(n15423), .ZN(n14115) );
  AOI21_X1 U15886 ( .B1(n14116), .B2(n19907), .A(n14115), .ZN(n14117) );
  NAND2_X1 U15887 ( .A1(n14232), .A2(n14381), .ZN(n14699) );
  OAI211_X1 U15888 ( .C1(n19503), .C2(n14381), .A(n14703), .B(n14229), .ZN(
        n14121) );
  NAND2_X1 U15889 ( .A1(n16126), .A2(n15608), .ZN(n14131) );
  NAND2_X1 U15890 ( .A1(n14691), .A2(n14385), .ZN(n14126) );
  INV_X1 U15891 ( .A(n14126), .ZN(n14124) );
  NAND2_X1 U15892 ( .A1(n14124), .A2(n19921), .ZN(n14130) );
  INV_X1 U15893 ( .A(n14385), .ZN(n14689) );
  NAND2_X1 U15894 ( .A1(n14689), .A2(n19895), .ZN(n14125) );
  NAND3_X1 U15895 ( .A1(n14693), .A2(n20466), .A3(n200), .ZN(n14128) );
  NAND3_X1 U15896 ( .A1(n14726), .A2(n14134), .A3(n14133), .ZN(n14136) );
  NAND3_X1 U15897 ( .A1(n20376), .A2(n14728), .A3(n14724), .ZN(n14135) );
  NAND2_X1 U15898 ( .A1(n15608), .A2(n16129), .ZN(n15734) );
  AOI21_X1 U15899 ( .B1(n16126), .B2(n15734), .A(n3431), .ZN(n14138) );
  OAI21_X1 U15900 ( .B1(n19488), .B2(n14611), .A(n14143), .ZN(n14145) );
  INV_X1 U15901 ( .A(n14207), .ZN(n14144) );
  AND2_X1 U15902 ( .A1(n19875), .A2(n14624), .ZN(n15320) );
  NAND2_X1 U15903 ( .A1(n15320), .A2(n14623), .ZN(n14147) );
  NAND2_X1 U15904 ( .A1(n14148), .A2(n19907), .ZN(n14400) );
  NAND3_X1 U15905 ( .A1(n14237), .A2(n14239), .A3(n14238), .ZN(n14151) );
  INV_X1 U15906 ( .A(n3822), .ZN(n15562) );
  NAND2_X1 U15907 ( .A1(n14598), .A2(n14395), .ZN(n14155) );
  MUX2_X1 U15908 ( .A(n14250), .B(n14599), .S(n1262), .Z(n14157) );
  NAND2_X1 U15909 ( .A1(n14157), .A2(n20377), .ZN(n14158) );
  INV_X1 U15910 ( .A(n15509), .ZN(n15560) );
  NOR2_X1 U15911 ( .A1(n15560), .A2(n15558), .ZN(n14160) );
  INV_X1 U15912 ( .A(n15510), .ZN(n15212) );
  INV_X1 U15913 ( .A(n15558), .ZN(n15513) );
  AOI22_X1 U15914 ( .A1(n14159), .A2(n14160), .B1(n15212), .B2(n15513), .ZN(
        n14161) );
  OAI21_X1 U15915 ( .B1(n20435), .B2(n15559), .A(n14161), .ZN(n16936) );
  INV_X1 U15916 ( .A(n2032), .ZN(n18294) );
  XNOR2_X1 U15917 ( .A(n16936), .B(n18294), .ZN(n14162) );
  XNOR2_X1 U15918 ( .A(n14163), .B(n14162), .ZN(n14164) );
  AOI21_X1 U15919 ( .B1(n16634), .B2(n20271), .A(n16170), .ZN(n14848) );
  MUX2_X1 U15920 ( .A(n19727), .B(n1936), .S(n20453), .Z(n14166) );
  NOR2_X1 U15921 ( .A1(n19728), .A2(n14490), .ZN(n14165) );
  NOR2_X1 U15922 ( .A1(n14434), .A2(n14480), .ZN(n14174) );
  AND2_X1 U15923 ( .A1(n14482), .A2(n14171), .ZN(n14303) );
  NAND2_X1 U15924 ( .A1(n14303), .A2(n14172), .ZN(n14173) );
  INV_X1 U15925 ( .A(n15309), .ZN(n14886) );
  AND2_X1 U15926 ( .A1(n15396), .A2(n14177), .ZN(n14190) );
  NOR2_X1 U15927 ( .A1(n14448), .A2(n14180), .ZN(n14178) );
  MUX2_X1 U15928 ( .A(n14179), .B(n14178), .S(n1364), .Z(n14183) );
  MUX2_X1 U15929 ( .A(n14448), .B(n14447), .S(n14180), .Z(n14181) );
  OAI21_X1 U15931 ( .B1(n14519), .B2(n14514), .A(n15119), .ZN(n14184) );
  OAI21_X1 U15932 ( .B1(n15311), .B2(n14188), .A(n14187), .ZN(n14189) );
  AOI21_X2 U15933 ( .B1(n14190), .B2(n15311), .A(n14189), .ZN(n17338) );
  AOI21_X1 U15934 ( .B1(n19875), .B2(n14620), .A(n15313), .ZN(n14191) );
  OAI21_X1 U15935 ( .B1(n14192), .B2(n19875), .A(n14191), .ZN(n14194) );
  NAND3_X1 U15936 ( .A1(n14192), .A2(n15313), .A3(n14623), .ZN(n14193) );
  INV_X1 U15937 ( .A(n14196), .ZN(n14198) );
  NOR2_X1 U15938 ( .A1(n14813), .A2(n14810), .ZN(n14197) );
  AOI22_X1 U15939 ( .A1(n14599), .A2(n20513), .B1(n14601), .B2(n20181), .ZN(
        n14201) );
  NAND2_X1 U15940 ( .A1(n19488), .A2(n14611), .ZN(n14204) );
  MUX2_X1 U15941 ( .A(n14204), .B(n14609), .S(n13907), .Z(n14210) );
  NAND2_X1 U15942 ( .A1(n19906), .A2(n13908), .ZN(n14608) );
  INV_X1 U15943 ( .A(n14608), .ZN(n14209) );
  OAI211_X1 U15944 ( .C1(n20500), .C2(n3497), .A(n14796), .B(n1938), .ZN(
        n14212) );
  NOR2_X1 U15945 ( .A1(n15070), .A2(n15618), .ZN(n15408) );
  INV_X1 U15946 ( .A(n15618), .ZN(n14214) );
  MUX2_X1 U15948 ( .A(n14216), .B(n14782), .S(n14775), .Z(n14219) );
  NAND3_X1 U15949 ( .A1(n14057), .A2(n14782), .A3(n14778), .ZN(n14218) );
  INV_X1 U15950 ( .A(n15405), .ZN(n15544) );
  INV_X1 U15951 ( .A(n15070), .ZN(n15620) );
  INV_X1 U15952 ( .A(n15071), .ZN(n15406) );
  NAND3_X1 U15953 ( .A1(n15544), .A2(n15620), .A3(n15406), .ZN(n14220) );
  OAI211_X1 U15954 ( .C1(n15619), .C2(n15616), .A(n14221), .B(n14220), .ZN(
        n16954) );
  XNOR2_X1 U15955 ( .A(n16954), .B(n17338), .ZN(n16584) );
  OAI21_X1 U15956 ( .B1(n20376), .B2(n14730), .A(n236), .ZN(n14222) );
  NAND2_X1 U15957 ( .A1(n14222), .A2(n14731), .ZN(n14226) );
  NAND2_X1 U15959 ( .A1(n14594), .A2(n2924), .ZN(n14233) );
  MUX2_X1 U15960 ( .A(n14234), .B(n14233), .S(n19761), .Z(n14235) );
  INV_X1 U15961 ( .A(n15430), .ZN(n15919) );
  OAI21_X1 U15962 ( .B1(n14242), .B2(n19908), .A(n14241), .ZN(n15426) );
  MUX2_X1 U15963 ( .A(n14718), .B(n3057), .S(n14717), .Z(n14247) );
  NAND2_X1 U15964 ( .A1(n3057), .A2(n14717), .ZN(n14244) );
  MUX2_X1 U15965 ( .A(n14245), .B(n14244), .S(n14715), .Z(n14246) );
  NAND2_X1 U15966 ( .A1(n15921), .A2(n15422), .ZN(n15920) );
  INV_X1 U15967 ( .A(n15422), .ZN(n15420) );
  NAND2_X1 U15968 ( .A1(n14248), .A2(n14599), .ZN(n14255) );
  INV_X1 U15969 ( .A(n14601), .ZN(n14251) );
  NAND3_X1 U15970 ( .A1(n20513), .A2(n14251), .A3(n19918), .ZN(n14253) );
  NAND2_X1 U15971 ( .A1(n14599), .A2(n20181), .ZN(n14252) );
  OAI21_X1 U15973 ( .B1(n15421), .B2(n15920), .A(n14257), .ZN(n14258) );
  NAND2_X1 U15974 ( .A1(n14674), .A2(n19652), .ZN(n14264) );
  INV_X1 U15975 ( .A(n14575), .ZN(n14569) );
  NAND2_X1 U15976 ( .A1(n14569), .A2(n14269), .ZN(n14737) );
  NAND3_X1 U15977 ( .A1(n14270), .A2(n14571), .A3(n14737), .ZN(n14271) );
  NAND2_X1 U15978 ( .A1(n14705), .A2(n14275), .ZN(n14274) );
  AOI21_X1 U15979 ( .B1(n14274), .B2(n14273), .A(n14566), .ZN(n14278) );
  NAND2_X1 U15980 ( .A1(n919), .A2(n14276), .ZN(n14277) );
  AND2_X1 U15981 ( .A1(n15400), .A2(n15536), .ZN(n14296) );
  MUX2_X1 U15983 ( .A(n14283), .B(n14282), .S(n14550), .Z(n14909) );
  NAND2_X1 U15984 ( .A1(n14284), .A2(n20120), .ZN(n14908) );
  NOR2_X1 U15985 ( .A1(n20471), .A2(n14656), .ZN(n14287) );
  INV_X1 U15986 ( .A(n14288), .ZN(n14660) );
  OAI21_X1 U15987 ( .B1(n14289), .B2(n20266), .A(n14547), .ZN(n14290) );
  NOR2_X1 U15988 ( .A1(n14660), .A2(n14290), .ZN(n14291) );
  NAND3_X1 U15989 ( .A1(n14688), .A2(n19895), .A3(n14695), .ZN(n14295) );
  AND2_X1 U15990 ( .A1(n19921), .A2(n14127), .ZN(n14384) );
  OAI21_X1 U15991 ( .B1(n14384), .B2(n14385), .A(n14691), .ZN(n14294) );
  OAI211_X1 U15992 ( .C1(n14696), .C2(n20466), .A(n14295), .B(n14294), .ZN(
        n15401) );
  INV_X1 U15993 ( .A(n15401), .ZN(n15538) );
  NAND3_X1 U15994 ( .A1(n15898), .A2(n15402), .A3(n15538), .ZN(n14298) );
  NAND2_X1 U15995 ( .A1(n19722), .A2(n14296), .ZN(n14297) );
  XNOR2_X1 U15996 ( .A(n16755), .B(n16836), .ZN(n17267) );
  XNOR2_X1 U15997 ( .A(n16584), .B(n17267), .ZN(n14376) );
  NOR2_X1 U15998 ( .A1(n14512), .A2(n14509), .ZN(n14639) );
  NAND2_X1 U15999 ( .A1(n14642), .A2(n14641), .ZN(n14299) );
  NOR2_X1 U16000 ( .A1(n14639), .A2(n14299), .ZN(n14300) );
  NOR2_X1 U16001 ( .A1(n14309), .A2(n14308), .ZN(n14312) );
  MUX2_X1 U16002 ( .A(n14648), .B(n14651), .S(n20443), .Z(n14311) );
  OAI21_X1 U16005 ( .B1(n14314), .B2(n14667), .A(n14313), .ZN(n14318) );
  AOI21_X1 U16006 ( .B1(n14316), .B2(n14315), .A(n14662), .ZN(n14317) );
  INV_X1 U16007 ( .A(n14903), .ZN(n15410) );
  MUX2_X1 U16008 ( .A(n14520), .B(n15121), .S(n15119), .Z(n14323) );
  NAND2_X1 U16009 ( .A1(n15120), .A2(n14520), .ZN(n14319) );
  OAI22_X1 U16010 ( .A1(n14321), .A2(n14320), .B1(n14319), .B2(n14514), .ZN(
        n14322) );
  XNOR2_X1 U16011 ( .A(n16373), .B(n18278), .ZN(n14374) );
  MUX2_X1 U16012 ( .A(n15469), .B(n15336), .S(n15465), .Z(n14324) );
  NAND2_X1 U16013 ( .A1(n14324), .A2(n15337), .ZN(n14333) );
  MUX2_X1 U16015 ( .A(n14329), .B(n14328), .S(n19693), .Z(n14331) );
  INV_X1 U16016 ( .A(n15470), .ZN(n15343) );
  NOR2_X1 U16017 ( .A1(n19583), .A2(n15339), .ZN(n14332) );
  NAND2_X1 U16018 ( .A1(n14336), .A2(n14335), .ZN(n14337) );
  NAND2_X1 U16019 ( .A1(n14338), .A2(n14342), .ZN(n14340) );
  MUX2_X1 U16020 ( .A(n14788), .B(n14344), .S(n14789), .Z(n14345) );
  MUX2_X1 U16021 ( .A(n3223), .B(n19496), .S(n14827), .Z(n14349) );
  NOR2_X1 U16022 ( .A1(n19859), .A2(n19986), .ZN(n14348) );
  NOR2_X1 U16023 ( .A1(n235), .A2(n14818), .ZN(n14351) );
  AOI22_X1 U16024 ( .A1(n14353), .A2(n20330), .B1(n14352), .B2(n14351), .ZN(
        n14354) );
  OAI21_X1 U16025 ( .B1(n2039), .B2(n14357), .A(n14356), .ZN(n14423) );
  INV_X1 U16026 ( .A(n14423), .ZN(n14362) );
  INV_X1 U16027 ( .A(n14358), .ZN(n14361) );
  OAI211_X1 U16028 ( .C1(n14422), .C2(n14359), .A(n14419), .B(n19939), .ZN(
        n14360) );
  OAI21_X2 U16029 ( .B1(n14362), .B2(n14361), .A(n14360), .ZN(n15907) );
  INV_X1 U16030 ( .A(n14363), .ZN(n14365) );
  NAND2_X1 U16032 ( .A1(n19531), .A2(n14462), .ZN(n14466) );
  NAND3_X1 U16033 ( .A1(n19531), .A2(n14468), .A3(n14369), .ZN(n14367) );
  AND2_X1 U16034 ( .A1(n14466), .A2(n14367), .ZN(n14368) );
  NOR2_X1 U16035 ( .A1(n15909), .A2(n15905), .ZN(n15077) );
  XNOR2_X1 U16036 ( .A(n16300), .B(n16406), .ZN(n14373) );
  XNOR2_X1 U16037 ( .A(n14374), .B(n14373), .ZN(n14375) );
  NAND2_X1 U16038 ( .A1(n17511), .A2(n20271), .ZN(n17509) );
  INV_X1 U16039 ( .A(n17509), .ZN(n16172) );
  INV_X1 U16040 ( .A(n15843), .ZN(n15267) );
  NOR2_X1 U16041 ( .A1(n15636), .A2(n15267), .ZN(n14377) );
  MUX2_X1 U16042 ( .A(n14700), .B(n14703), .S(n20204), .Z(n14383) );
  NAND2_X1 U16043 ( .A1(n14380), .A2(n14379), .ZN(n14382) );
  INV_X1 U16044 ( .A(n15838), .ZN(n15100) );
  NAND2_X1 U16045 ( .A1(n14693), .A2(n14384), .ZN(n14386) );
  NAND2_X1 U16046 ( .A1(n19862), .A2(n14723), .ZN(n14392) );
  MUX2_X1 U16047 ( .A(n19862), .B(n14723), .S(n14718), .Z(n14390) );
  MUX2_X1 U16048 ( .A(n14390), .B(n14389), .S(n19843), .Z(n14391) );
  OAI21_X1 U16049 ( .B1(n2926), .B2(n14394), .A(n19731), .ZN(n14399) );
  NAND2_X1 U16050 ( .A1(n14403), .A2(n15423), .ZN(n14404) );
  AOI21_X1 U16051 ( .B1(n14406), .B2(n14405), .A(n14404), .ZN(n14407) );
  NOR2_X1 U16052 ( .A1(n15627), .A2(n15628), .ZN(n14415) );
  NOR2_X1 U16053 ( .A1(n14408), .A2(n14729), .ZN(n14409) );
  NAND2_X1 U16054 ( .A1(n14409), .A2(n14726), .ZN(n15002) );
  NAND2_X1 U16055 ( .A1(n14410), .A2(n14724), .ZN(n14411) );
  NAND2_X1 U16056 ( .A1(n14731), .A2(n14411), .ZN(n14413) );
  MUX2_X1 U16057 ( .A(n14728), .B(n14413), .S(n14412), .Z(n15003) );
  AOI21_X1 U16058 ( .B1(n15002), .B2(n15003), .A(n15625), .ZN(n14414) );
  MUX2_X1 U16059 ( .A(n14415), .B(n14414), .S(n15838), .Z(n14416) );
  AOI21_X1 U16060 ( .B1(n14417), .B2(n15627), .A(n14416), .ZN(n17261) );
  XNOR2_X1 U16061 ( .A(n17261), .B(n17438), .ZN(n16514) );
  OAI21_X1 U16062 ( .B1(n19939), .B2(n14419), .A(n14418), .ZN(n14421) );
  NAND2_X1 U16063 ( .A1(n14424), .A2(n3156), .ZN(n14430) );
  NOR2_X1 U16064 ( .A1(n14426), .A2(n14425), .ZN(n14492) );
  INV_X1 U16065 ( .A(n14492), .ZN(n14429) );
  NAND2_X1 U16066 ( .A1(n14433), .A2(n14480), .ZN(n14438) );
  INV_X1 U16067 ( .A(n14434), .ZN(n14436) );
  NOR2_X1 U16068 ( .A1(n14436), .A2(n14435), .ZN(n14437) );
  INV_X1 U16069 ( .A(n15297), .ZN(n14446) );
  MUX2_X1 U16070 ( .A(n14442), .B(n12919), .S(n14441), .Z(n14444) );
  NOR2_X1 U16071 ( .A1(n14444), .A2(n14443), .ZN(n14445) );
  AOI21_X1 U16072 ( .B1(n15296), .B2(n14446), .A(n15294), .ZN(n14460) );
  NOR2_X1 U16073 ( .A1(n14452), .A2(n14451), .ZN(n14457) );
  NOR2_X1 U16074 ( .A1(n14454), .A2(n14453), .ZN(n14456) );
  MUX2_X1 U16075 ( .A(n14457), .B(n14456), .S(n1364), .Z(n14458) );
  MUX2_X1 U16076 ( .A(n15111), .B(n14460), .S(n14770), .Z(n14473) );
  NAND2_X1 U16077 ( .A1(n15294), .A2(n14461), .ZN(n15293) );
  INV_X1 U16078 ( .A(n19819), .ZN(n14464) );
  AOI21_X1 U16079 ( .B1(n14465), .B2(n14464), .A(n3252), .ZN(n14467) );
  MUX2_X1 U16080 ( .A(n14468), .B(n14467), .S(n14466), .Z(n14471) );
  NOR3_X1 U16081 ( .A1(n3299), .A2(n14469), .A3(n14468), .ZN(n14470) );
  NOR2_X1 U16083 ( .A1(n15293), .A2(n15110), .ZN(n14472) );
  NOR2_X2 U16084 ( .A1(n14473), .A2(n14472), .ZN(n16607) );
  NAND2_X1 U16086 ( .A1(n15909), .A2(n15905), .ZN(n14475) );
  NAND2_X1 U16087 ( .A1(n15008), .A2(n15907), .ZN(n14474) );
  NAND3_X1 U16088 ( .A1(n14475), .A2(n2578), .A3(n14474), .ZN(n14478) );
  INV_X1 U16089 ( .A(n14475), .ZN(n14476) );
  NAND2_X1 U16090 ( .A1(n14476), .A2(n15906), .ZN(n14477) );
  OAI211_X1 U16091 ( .C1(n2578), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        n16293) );
  XNOR2_X1 U16092 ( .A(n16607), .B(n16293), .ZN(n16175) );
  XNOR2_X1 U16093 ( .A(n16514), .B(n16175), .ZN(n14634) );
  NAND2_X1 U16094 ( .A1(n14482), .A2(n14480), .ZN(n14489) );
  INV_X1 U16097 ( .A(n15132), .ZN(n14838) );
  NOR2_X1 U16098 ( .A1(n14747), .A2(n14490), .ZN(n14491) );
  OR2_X2 U16099 ( .A1(n14496), .A2(n14495), .ZN(n15282) );
  MUX2_X1 U16100 ( .A(n14499), .B(n14498), .S(n14497), .Z(n14505) );
  NOR2_X1 U16104 ( .A1(n15282), .A2(n15284), .ZN(n15286) );
  INV_X1 U16105 ( .A(n15286), .ZN(n14534) );
  NAND2_X1 U16106 ( .A1(n13983), .A2(n14641), .ZN(n14507) );
  AOI22_X1 U16107 ( .A1(n14635), .A2(n14512), .B1(n19703), .B2(n14640), .ZN(
        n14511) );
  INV_X1 U16108 ( .A(n15130), .ZN(n14529) );
  INV_X1 U16109 ( .A(n14514), .ZN(n14515) );
  NOR2_X1 U16111 ( .A1(n951), .A2(n14522), .ZN(n14523) );
  NAND3_X1 U16112 ( .A1(n14525), .A2(n14648), .A3(n14524), .ZN(n14526) );
  NAND2_X1 U16113 ( .A1(n14652), .A2(n14526), .ZN(n14527) );
  NAND2_X1 U16114 ( .A1(n14529), .A2(n15127), .ZN(n14530) );
  NAND2_X1 U16115 ( .A1(n15281), .A2(n14530), .ZN(n14531) );
  NAND2_X1 U16116 ( .A1(n14531), .A2(n19848), .ZN(n14533) );
  NAND3_X1 U16117 ( .A1(n15282), .A2(n15018), .A3(n20474), .ZN(n14532) );
  NAND2_X1 U16118 ( .A1(n14673), .A2(n14539), .ZN(n14546) );
  NAND2_X1 U16119 ( .A1(n20424), .A2(n19652), .ZN(n14675) );
  NAND2_X1 U16120 ( .A1(n14544), .A2(n13981), .ZN(n14545) );
  INV_X1 U16121 ( .A(n15645), .ZN(n15831) );
  INV_X1 U16124 ( .A(n15256), .ZN(n15643) );
  MUX2_X1 U16125 ( .A(n14552), .B(n14551), .S(n14279), .Z(n14561) );
  NOR2_X1 U16126 ( .A1(n14554), .A2(n14553), .ZN(n14559) );
  NOR2_X1 U16127 ( .A1(n14556), .A2(n14555), .ZN(n14558) );
  MUX2_X1 U16128 ( .A(n14559), .B(n14558), .S(n14557), .Z(n14560) );
  INV_X1 U16129 ( .A(n15644), .ZN(n15829) );
  MUX2_X1 U16130 ( .A(n20498), .B(n14705), .S(n14562), .Z(n14567) );
  MUX2_X1 U16131 ( .A(n14564), .B(n14563), .S(n14704), .Z(n14565) );
  OAI21_X1 U16132 ( .B1(n14567), .B2(n14566), .A(n14565), .ZN(n15096) );
  NAND2_X1 U16133 ( .A1(n15829), .A2(n19891), .ZN(n15649) );
  NAND2_X1 U16135 ( .A1(n14569), .A2(n14736), .ZN(n14573) );
  NAND2_X1 U16136 ( .A1(n14571), .A2(n14570), .ZN(n14572) );
  AND2_X1 U16138 ( .A1(n15096), .A2(n15644), .ZN(n15259) );
  INV_X1 U16139 ( .A(n15259), .ZN(n14580) );
  AOI21_X1 U16140 ( .B1(n14581), .B2(n14580), .A(n15256), .ZN(n14582) );
  XNOR2_X1 U16141 ( .A(n16750), .B(n19704), .ZN(n16392) );
  NOR2_X1 U16142 ( .A1(n14796), .A2(n1351), .ZN(n14585) );
  AOI22_X1 U16143 ( .A1(n14585), .A2(n3439), .B1(n1351), .B2(n14799), .ZN(
        n14586) );
  NAND2_X1 U16144 ( .A1(n14587), .A2(n14199), .ZN(n14592) );
  INV_X1 U16145 ( .A(n14807), .ZN(n14589) );
  NOR2_X1 U16146 ( .A1(n15270), .A2(n15601), .ZN(n14618) );
  NAND3_X1 U16147 ( .A1(n20377), .A2(n2682), .A3(n14601), .ZN(n14607) );
  INV_X1 U16148 ( .A(n14603), .ZN(n14604) );
  NAND3_X1 U16149 ( .A1(n20513), .A2(n1262), .A3(n14604), .ZN(n14606) );
  INV_X1 U16150 ( .A(n15274), .ZN(n15114) );
  NOR2_X1 U16151 ( .A1(n15275), .A2(n15114), .ZN(n14617) );
  AOI21_X1 U16152 ( .B1(n14612), .B2(n13907), .A(n14611), .ZN(n14613) );
  NAND2_X1 U16153 ( .A1(n14614), .A2(n14613), .ZN(n14615) );
  NAND3_X1 U16156 ( .A1(n954), .A2(n19875), .A3(n14623), .ZN(n14622) );
  NAND3_X1 U16157 ( .A1(n15314), .A2(n14620), .A3(n15313), .ZN(n14621) );
  OAI211_X1 U16159 ( .C1(n954), .C2(n14627), .A(n14625), .B(n14624), .ZN(
        n14628) );
  NAND2_X1 U16160 ( .A1(n15276), .A2(n15271), .ZN(n14629) );
  INV_X1 U16161 ( .A(n15270), .ZN(n15009) );
  AOI21_X1 U16162 ( .B1(n15277), .B2(n14629), .A(n15009), .ZN(n14630) );
  NOR2_X2 U16163 ( .A1(n14631), .A2(n14630), .ZN(n16914) );
  INV_X1 U16164 ( .A(n649), .ZN(n19152) );
  XNOR2_X1 U16165 ( .A(n16914), .B(n19152), .ZN(n14632) );
  XNOR2_X1 U16166 ( .A(n16392), .B(n14632), .ZN(n14633) );
  OR2_X1 U16167 ( .A1(n14636), .A2(n14635), .ZN(n14646) );
  NOR2_X1 U16168 ( .A1(n14640), .A2(n14637), .ZN(n14638) );
  NOR2_X1 U16169 ( .A1(n14639), .A2(n14638), .ZN(n14645) );
  MUX2_X1 U16170 ( .A(n14642), .B(n14641), .S(n14640), .Z(n14643) );
  OAI22_X1 U16171 ( .A1(n14651), .A2(n951), .B1(n14648), .B2(n20380), .ZN(
        n14649) );
  AND2_X1 U16172 ( .A1(n15573), .A2(n15577), .ZN(n15793) );
  NOR2_X1 U16173 ( .A1(n14653), .A2(n14656), .ZN(n14655) );
  NAND3_X1 U16174 ( .A1(n14655), .A2(n14654), .A3(n14659), .ZN(n14661) );
  OAI21_X1 U16175 ( .B1(n20266), .B2(n14656), .A(n20471), .ZN(n14658) );
  NOR2_X1 U16176 ( .A1(n15793), .A2(n15574), .ZN(n14687) );
  NOR2_X1 U16177 ( .A1(n14663), .A2(n14662), .ZN(n14665) );
  INV_X1 U16178 ( .A(n15573), .ZN(n15791) );
  NOR2_X1 U16179 ( .A1(n15791), .A2(n15577), .ZN(n14685) );
  OR2_X1 U16180 ( .A1(n14680), .A2(n20120), .ZN(n14681) );
  NAND3_X1 U16181 ( .A1(n14683), .A2(n14682), .A3(n14681), .ZN(n15365) );
  INV_X1 U16182 ( .A(n15365), .ZN(n15572) );
  NOR2_X1 U16183 ( .A1(n15577), .A2(n15572), .ZN(n14684) );
  AOI22_X1 U16184 ( .A1(n15796), .A2(n14685), .B1(n14684), .B2(n860), .ZN(
        n14686) );
  NAND3_X1 U16186 ( .A1(n14689), .A2(n14688), .A3(n200), .ZN(n14694) );
  NAND2_X1 U16187 ( .A1(n14120), .A2(n2769), .ZN(n14698) );
  NAND2_X1 U16188 ( .A1(n14699), .A2(n14698), .ZN(n14701) );
  NAND2_X1 U16189 ( .A1(n14701), .A2(n14700), .ZN(n14702) );
  OAI21_X1 U16190 ( .B1(n14273), .B2(n14704), .A(n919), .ZN(n14713) );
  NOR2_X1 U16191 ( .A1(n14705), .A2(n2282), .ZN(n14712) );
  NAND2_X1 U16192 ( .A1(n14708), .A2(n20498), .ZN(n14711) );
  NAND2_X1 U16193 ( .A1(n14273), .A2(n14709), .ZN(n14710) );
  OAI211_X1 U16194 ( .C1(n14713), .C2(n14712), .A(n14711), .B(n14710), .ZN(
        n15801) );
  INV_X1 U16195 ( .A(n15801), .ZN(n15042) );
  OAI21_X1 U16196 ( .B1(n14716), .B2(n14715), .A(n19862), .ZN(n14720) );
  MUX2_X1 U16197 ( .A(n14720), .B(n14719), .S(n14718), .Z(n14721) );
  MUX2_X1 U16198 ( .A(n14731), .B(n14730), .S(n14729), .Z(n14733) );
  NOR2_X1 U16199 ( .A1(n14733), .A2(n20376), .ZN(n14734) );
  NAND2_X1 U16200 ( .A1(n14737), .A2(n14736), .ZN(n14739) );
  INV_X1 U16202 ( .A(n15802), .ZN(n14742) );
  AND2_X1 U16204 ( .A1(n15801), .A2(n15803), .ZN(n15564) );
  INV_X1 U16205 ( .A(n15567), .ZN(n15804) );
  AOI22_X1 U16206 ( .A1(n15564), .A2(n942), .B1(n15804), .B2(n15801), .ZN(
        n14744) );
  XNOR2_X1 U16207 ( .A(n17294), .B(n16853), .ZN(n16365) );
  NOR2_X1 U16208 ( .A1(n14747), .A2(n19727), .ZN(n14748) );
  NOR2_X1 U16209 ( .A1(n14749), .A2(n14748), .ZN(n14751) );
  MUX2_X1 U16210 ( .A(n14751), .B(n14750), .S(n1936), .Z(n14752) );
  NAND2_X1 U16211 ( .A1(n15189), .A2(n14935), .ZN(n14764) );
  INV_X1 U16212 ( .A(n14754), .ZN(n14761) );
  INV_X1 U16213 ( .A(n14755), .ZN(n14760) );
  INV_X1 U16214 ( .A(n14756), .ZN(n14759) );
  INV_X1 U16215 ( .A(n14757), .ZN(n14758) );
  NAND4_X1 U16216 ( .A1(n14761), .A2(n14760), .A3(n14759), .A4(n14758), .ZN(
        n14762) );
  AOI22_X1 U16217 ( .A1(n15504), .A2(n15506), .B1(n2288), .B2(n14762), .ZN(
        n14763) );
  AOI22_X2 U16218 ( .A1(n14763), .A2(n14764), .B1(n15506), .B2(n15822), .ZN(
        n16945) );
  INV_X1 U16219 ( .A(n15559), .ZN(n14966) );
  OAI21_X1 U16220 ( .B1(n15511), .B2(n15510), .A(n14159), .ZN(n14766) );
  OAI211_X1 U16221 ( .C1(n14966), .C2(n14964), .A(n14766), .B(n14765), .ZN(
        n17300) );
  INV_X1 U16222 ( .A(n17300), .ZN(n14767) );
  XNOR2_X1 U16223 ( .A(n16945), .B(n14767), .ZN(n16527) );
  XNOR2_X1 U16224 ( .A(n16365), .B(n16527), .ZN(n14844) );
  NOR2_X1 U16225 ( .A1(n15110), .A2(n15295), .ZN(n14769) );
  AOI21_X1 U16226 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n14774) );
  NAND2_X1 U16227 ( .A1(n15295), .A2(n15111), .ZN(n14772) );
  NOR2_X1 U16228 ( .A1(n15110), .A2(n14772), .ZN(n14773) );
  NAND3_X1 U16229 ( .A1(n877), .A2(n20518), .A3(n14775), .ZN(n14776) );
  OAI21_X1 U16230 ( .B1(n14852), .B2(n20408), .A(n14776), .ZN(n14786) );
  NOR2_X1 U16231 ( .A1(n877), .A2(n14778), .ZN(n14784) );
  NOR2_X1 U16232 ( .A1(n14781), .A2(n20454), .ZN(n14783) );
  MUX2_X1 U16233 ( .A(n14784), .B(n14783), .S(n14782), .Z(n14785) );
  MUX2_X1 U16234 ( .A(n14103), .B(n14787), .S(n14790), .Z(n14794) );
  MUX2_X1 U16235 ( .A(n14791), .B(n14790), .S(n14789), .Z(n14793) );
  NAND2_X1 U16236 ( .A1(n14796), .A2(n13891), .ZN(n14798) );
  AOI21_X1 U16237 ( .B1(n14798), .B2(n14797), .A(n14800), .ZN(n14805) );
  NAND3_X1 U16238 ( .A1(n1351), .A2(n3497), .A3(n14799), .ZN(n14803) );
  NAND2_X1 U16239 ( .A1(n14803), .A2(n14802), .ZN(n14804) );
  MUX2_X1 U16240 ( .A(n15582), .B(n3534), .S(n15812), .Z(n14836) );
  NOR2_X1 U16241 ( .A1(n14807), .A2(n14806), .ZN(n14808) );
  AOI22_X1 U16242 ( .A1(n14812), .A2(n14809), .B1(n14808), .B2(n14199), .ZN(
        n14816) );
  OAI21_X1 U16243 ( .B1(n239), .B2(n14814), .A(n14813), .ZN(n14815) );
  NAND2_X1 U16245 ( .A1(n14820), .A2(n12931), .ZN(n14822) );
  INV_X1 U16247 ( .A(n15583), .ZN(n15814) );
  NOR2_X1 U16248 ( .A1(n15814), .A2(n15582), .ZN(n15354) );
  OAI211_X1 U16250 ( .C1(n14828), .C2(n3223), .A(n14827), .B(n14826), .ZN(
        n14832) );
  NOR2_X1 U16251 ( .A1(n15354), .A2(n14834), .ZN(n14835) );
  XNOR2_X1 U16252 ( .A(n16964), .B(n17295), .ZN(n14842) );
  NAND2_X1 U16253 ( .A1(n15132), .A2(n15282), .ZN(n14837) );
  MUX2_X1 U16254 ( .A(n15017), .B(n20474), .S(n15018), .Z(n14839) );
  XNOR2_X1 U16255 ( .A(n16614), .B(n18988), .ZN(n14841) );
  XNOR2_X1 U16256 ( .A(n14842), .B(n14841), .ZN(n14843) );
  XNOR2_X1 U16257 ( .A(n14844), .B(n14843), .ZN(n17225) );
  INV_X1 U16258 ( .A(n17225), .ZN(n14845) );
  NAND2_X1 U16259 ( .A1(n14845), .A2(n19700), .ZN(n14846) );
  INV_X1 U16261 ( .A(n15769), .ZN(n15475) );
  INV_X1 U16262 ( .A(n14850), .ZN(n14854) );
  INV_X1 U16263 ( .A(n14851), .ZN(n14853) );
  NAND3_X1 U16264 ( .A1(n14854), .A2(n14853), .A3(n14852), .ZN(n14855) );
  NOR2_X1 U16265 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  NOR2_X2 U16266 ( .A1(n14859), .A2(n14858), .ZN(n16981) );
  INV_X1 U16267 ( .A(n15349), .ZN(n15348) );
  NOR2_X1 U16268 ( .A1(n20173), .A2(n15348), .ZN(n14861) );
  XNOR2_X1 U16270 ( .A(n16981), .B(n19927), .ZN(n16506) );
  INV_X1 U16271 ( .A(n15673), .ZN(n15775) );
  NAND2_X1 U16273 ( .A1(n15672), .A2(n15665), .ZN(n14864) );
  NAND2_X1 U16274 ( .A1(n13414), .A2(n20151), .ZN(n14863) );
  MUX2_X1 U16275 ( .A(n14864), .B(n14863), .S(n234), .Z(n14865) );
  INV_X1 U16276 ( .A(n14866), .ZN(n15783) );
  NAND3_X1 U16279 ( .A1(n15685), .A2(n15683), .A3(n15684), .ZN(n14869) );
  NAND3_X1 U16280 ( .A1(n15686), .A2(n19977), .A3(n20362), .ZN(n14868) );
  XNOR2_X1 U16281 ( .A(n17339), .B(n1054), .ZN(n17036) );
  XNOR2_X1 U16282 ( .A(n16506), .B(n17036), .ZN(n14885) );
  NOR2_X1 U16283 ( .A1(n15380), .A2(n15166), .ZN(n14871) );
  NOR2_X1 U16284 ( .A1(n14872), .A2(n14871), .ZN(n14873) );
  NOR3_X1 U16285 ( .A1(n15380), .A2(n15379), .A3(n20103), .ZN(n14876) );
  NOR2_X1 U16286 ( .A1(n15682), .A2(n15445), .ZN(n14880) );
  NOR3_X1 U16287 ( .A1(n15676), .A2(n15679), .A3(n15442), .ZN(n14879) );
  NOR2_X1 U16288 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  XNOR2_X1 U16289 ( .A(n897), .B(n17340), .ZN(n14883) );
  XNOR2_X1 U16290 ( .A(n16300), .B(n19140), .ZN(n14882) );
  XNOR2_X1 U16291 ( .A(n14883), .B(n14882), .ZN(n14884) );
  NOR2_X1 U16293 ( .A1(n15311), .A2(n15395), .ZN(n14889) );
  NAND2_X1 U16294 ( .A1(n15059), .A2(n15308), .ZN(n14990) );
  OAI21_X1 U16295 ( .B1(n14886), .B2(n15308), .A(n14990), .ZN(n14887) );
  NOR2_X1 U16296 ( .A1(n15546), .A2(n15619), .ZN(n14890) );
  NAND2_X1 U16297 ( .A1(n14890), .A2(n15406), .ZN(n14894) );
  NOR2_X1 U16298 ( .A1(n15405), .A2(n15618), .ZN(n14891) );
  OAI21_X1 U16299 ( .B1(n15073), .B2(n14891), .A(n15546), .ZN(n14893) );
  NAND3_X1 U16300 ( .A1(n14894), .A2(n14893), .A3(n14892), .ZN(n16999) );
  INV_X1 U16301 ( .A(n16999), .ZN(n16510) );
  XNOR2_X1 U16302 ( .A(n16999), .B(n14895), .ZN(n15953) );
  NAND2_X1 U16303 ( .A1(n15465), .A2(n14896), .ZN(n14897) );
  NAND2_X1 U16304 ( .A1(n15082), .A2(n3817), .ZN(n14898) );
  INV_X1 U16305 ( .A(n19467), .ZN(n14901) );
  INV_X1 U16306 ( .A(n14902), .ZN(n15550) );
  NAND2_X1 U16307 ( .A1(n15550), .A2(n14903), .ZN(n14904) );
  AND3_X1 U16308 ( .A1(n14905), .A2(n14978), .A3(n14904), .ZN(n14906) );
  NOR2_X2 U16309 ( .A1(n14907), .A2(n14906), .ZN(n17260) );
  INV_X1 U16310 ( .A(n15400), .ZN(n15537) );
  OAI21_X1 U16311 ( .B1(n15401), .B2(n15536), .A(n15537), .ZN(n14913) );
  NAND2_X1 U16314 ( .A1(n14909), .A2(n14908), .ZN(n15892) );
  XNOR2_X1 U16317 ( .A(n17378), .B(n17260), .ZN(n14914) );
  INV_X1 U16319 ( .A(n15859), .ZN(n14918) );
  INV_X1 U16320 ( .A(n15720), .ZN(n15862) );
  OAI21_X1 U16321 ( .B1(n15866), .B2(n15862), .A(n15863), .ZN(n14917) );
  MUX2_X1 U16322 ( .A(n15864), .B(n15861), .S(n15720), .Z(n14916) );
  XNOR2_X1 U16323 ( .A(n16420), .B(n17104), .ZN(n14928) );
  NOR2_X1 U16324 ( .A1(n15875), .A2(n15714), .ZN(n15713) );
  INV_X1 U16325 ( .A(n15870), .ZN(n15150) );
  MUX2_X1 U16326 ( .A(n15874), .B(n15876), .S(n20178), .Z(n14920) );
  NOR2_X1 U16327 ( .A1(n14920), .A2(n15148), .ZN(n14921) );
  NOR2_X2 U16328 ( .A1(n14922), .A2(n14921), .ZN(n17012) );
  INV_X1 U16329 ( .A(n15335), .ZN(n14923) );
  NAND2_X1 U16330 ( .A1(n16009), .A2(n19739), .ZN(n15880) );
  NAND3_X1 U16331 ( .A1(n14923), .A2(n16015), .A3(n15880), .ZN(n14926) );
  INV_X1 U16332 ( .A(n14924), .ZN(n14925) );
  NAND2_X1 U16333 ( .A1(n15885), .A2(n14925), .ZN(n16017) );
  XNOR2_X1 U16334 ( .A(n17012), .B(n14927), .ZN(n16418) );
  XNOR2_X1 U16335 ( .A(n14928), .B(n16418), .ZN(n14943) );
  INV_X1 U16337 ( .A(n15496), .ZN(n15191) );
  AND2_X1 U16338 ( .A1(n15501), .A2(n15191), .ZN(n14929) );
  OAI21_X1 U16339 ( .B1(n14930), .B2(n14929), .A(n15497), .ZN(n14933) );
  INV_X1 U16340 ( .A(n15501), .ZN(n14931) );
  NAND3_X1 U16341 ( .A1(n14931), .A2(n19512), .A3(n15500), .ZN(n14932) );
  MUX2_X1 U16342 ( .A(n15505), .B(n15503), .S(n15188), .Z(n14936) );
  XNOR2_X1 U16343 ( .A(n16602), .B(n16045), .ZN(n16232) );
  NOR2_X1 U16344 ( .A1(n20133), .A2(n15696), .ZN(n14940) );
  NOR2_X1 U16345 ( .A1(n20145), .A2(n15702), .ZN(n14939) );
  XNOR2_X1 U16346 ( .A(n19836), .B(n18768), .ZN(n14941) );
  XNOR2_X1 U16347 ( .A(n16232), .B(n14941), .ZN(n14942) );
  MUX2_X1 U16349 ( .A(n17210), .B(n20135), .S(n20092), .Z(n15027) );
  NAND2_X1 U16352 ( .A1(n15297), .A2(n14461), .ZN(n14945) );
  MUX2_X1 U16353 ( .A(n14946), .B(n14945), .S(n15296), .Z(n14947) );
  XNOR2_X1 U16354 ( .A(n16329), .B(n17733), .ZN(n14957) );
  INV_X1 U16355 ( .A(n15574), .ZN(n15794) );
  NAND2_X1 U16356 ( .A1(n859), .A2(n15572), .ZN(n14949) );
  NOR2_X1 U16357 ( .A1(n15577), .A2(n15573), .ZN(n14948) );
  NOR2_X1 U16358 ( .A1(n14949), .A2(n14948), .ZN(n14950) );
  NOR2_X2 U16359 ( .A1(n14951), .A2(n14950), .ZN(n17280) );
  INV_X1 U16360 ( .A(n17280), .ZN(n14956) );
  INV_X1 U16361 ( .A(n14952), .ZN(n15371) );
  AOI22_X1 U16362 ( .A1(n20183), .A2(n15371), .B1(n15370), .B2(n15566), .ZN(
        n15043) );
  NAND2_X1 U16363 ( .A1(n15803), .A2(n15042), .ZN(n14953) );
  NAND2_X1 U16364 ( .A1(n15808), .A2(n14953), .ZN(n14955) );
  XNOR2_X1 U16367 ( .A(n17026), .B(n14957), .ZN(n14971) );
  NOR2_X1 U16368 ( .A1(n15132), .A2(n15282), .ZN(n15287) );
  INV_X1 U16369 ( .A(n15018), .ZN(n15285) );
  NAND2_X1 U16370 ( .A1(n15285), .A2(n15127), .ZN(n14961) );
  INV_X1 U16371 ( .A(n15282), .ZN(n14959) );
  NAND2_X1 U16372 ( .A1(n15130), .A2(n15017), .ZN(n14958) );
  INV_X1 U16374 ( .A(n16927), .ZN(n14963) );
  NOR2_X1 U16375 ( .A1(n15814), .A2(n233), .ZN(n14962) );
  XNOR2_X1 U16376 ( .A(n14963), .B(n16969), .ZN(n16522) );
  NOR2_X1 U16377 ( .A1(n14159), .A2(n15509), .ZN(n14965) );
  OAI21_X1 U16378 ( .B1(n14966), .B2(n15562), .A(n14965), .ZN(n14967) );
  XNOR2_X1 U16379 ( .A(n16974), .B(n17366), .ZN(n16288) );
  XNOR2_X1 U16380 ( .A(n19849), .B(n16288), .ZN(n14970) );
  NAND2_X1 U16382 ( .A1(n15756), .A2(n15588), .ZN(n15992) );
  INV_X1 U16383 ( .A(n15992), .ZN(n14974) );
  OAI21_X1 U16384 ( .B1(n15755), .B2(n15588), .A(n15760), .ZN(n15989) );
  NOR2_X1 U16385 ( .A1(n15756), .A2(n15758), .ZN(n15991) );
  INV_X1 U16386 ( .A(n15991), .ZN(n14972) );
  NAND3_X1 U16387 ( .A1(n14972), .A2(n15992), .A3(n15587), .ZN(n14973) );
  OAI21_X1 U16388 ( .B1(n14974), .B2(n15989), .A(n14973), .ZN(n16078) );
  XNOR2_X1 U16391 ( .A(n16078), .B(n17327), .ZN(n17019) );
  NAND2_X1 U16392 ( .A1(n15409), .A2(n15549), .ZN(n14981) );
  OR2_X1 U16393 ( .A1(n15549), .A2(n15553), .ZN(n14980) );
  NOR2_X1 U16394 ( .A1(n15181), .A2(n19502), .ZN(n15522) );
  INV_X1 U16395 ( .A(n14982), .ZN(n14983) );
  AND2_X1 U16396 ( .A1(n15746), .A2(n15741), .ZN(n15180) );
  INV_X1 U16397 ( .A(n15516), .ZN(n15178) );
  NOR2_X1 U16398 ( .A1(n15178), .A2(n15182), .ZN(n14984) );
  INV_X1 U16399 ( .A(n15746), .ZN(n15742) );
  XNOR2_X1 U16400 ( .A(n16961), .B(n16944), .ZN(n16528) );
  XNOR2_X1 U16401 ( .A(n17019), .B(n16528), .ZN(n14995) );
  INV_X1 U16402 ( .A(n15277), .ZN(n14986) );
  NAND2_X1 U16403 ( .A1(n19662), .A2(n15395), .ZN(n14992) );
  INV_X1 U16405 ( .A(n2356), .ZN(n19264) );
  XNOR2_X1 U16406 ( .A(n16227), .B(n19264), .ZN(n14993) );
  XNOR2_X1 U16407 ( .A(n16284), .B(n14993), .ZN(n14994) );
  NAND2_X1 U16411 ( .A1(n15003), .A2(n15002), .ZN(n15840) );
  AND2_X1 U16412 ( .A1(n15628), .A2(n15627), .ZN(n15837) );
  NAND2_X1 U16413 ( .A1(n15837), .A2(n15840), .ZN(n15006) );
  OAI21_X1 U16414 ( .B1(n1288), .B2(n15839), .A(n15627), .ZN(n15004) );
  NAND2_X1 U16415 ( .A1(n15004), .A2(n15100), .ZN(n15005) );
  OAI211_X1 U16416 ( .C1(n15626), .C2(n15100), .A(n15006), .B(n15005), .ZN(
        n17360) );
  XNOR2_X1 U16417 ( .A(n16706), .B(n17360), .ZN(n16276) );
  INV_X1 U16418 ( .A(n15601), .ZN(n15112) );
  OAI21_X1 U16420 ( .B1(n15112), .B2(n15009), .A(n15113), .ZN(n15605) );
  NAND2_X1 U16421 ( .A1(n15601), .A2(n15600), .ZN(n15010) );
  AOI21_X1 U16422 ( .B1(n15270), .B2(n15010), .A(n20112), .ZN(n15011) );
  XNOR2_X1 U16424 ( .A(n15935), .B(n16236), .ZN(n15012) );
  XNOR2_X1 U16425 ( .A(n16276), .B(n15012), .ZN(n15025) );
  NAND2_X1 U16426 ( .A1(n15296), .A2(n15297), .ZN(n15013) );
  AOI21_X1 U16427 ( .B1(n15108), .B2(n15013), .A(n15110), .ZN(n15016) );
  NAND2_X1 U16428 ( .A1(n15296), .A2(n15295), .ZN(n15014) );
  AOI21_X1 U16429 ( .B1(n15297), .B2(n15014), .A(n15294), .ZN(n15015) );
  NOR2_X2 U16430 ( .A1(n15016), .A2(n15015), .ZN(n16938) );
  NAND2_X1 U16431 ( .A1(n15018), .A2(n15017), .ZN(n15283) );
  NAND2_X1 U16432 ( .A1(n15283), .A2(n20474), .ZN(n15019) );
  AOI22_X2 U16433 ( .A1(n15020), .A2(n15132), .B1(n15019), .B2(n19848), .ZN(
        n17253) );
  XNOR2_X1 U16434 ( .A(n16938), .B(n17253), .ZN(n15023) );
  XNOR2_X1 U16435 ( .A(n864), .B(n15021), .ZN(n15022) );
  XNOR2_X1 U16436 ( .A(n15023), .B(n15022), .ZN(n15024) );
  XNOR2_X1 U16437 ( .A(n15025), .B(n15024), .ZN(n16251) );
  INV_X1 U16438 ( .A(n15380), .ZN(n15164) );
  NOR2_X1 U16439 ( .A1(n15164), .A2(n15028), .ZN(n15029) );
  AOI21_X2 U16440 ( .B1(n15033), .B2(n15167), .A(n15032), .ZN(n16554) );
  XNOR2_X1 U16441 ( .A(n16554), .B(n16429), .ZN(n15038) );
  NAND2_X1 U16442 ( .A1(n15583), .A2(n3315), .ZN(n15034) );
  OAI21_X1 U16443 ( .B1(n15582), .B2(n15581), .A(n15583), .ZN(n15036) );
  XNOR2_X1 U16444 ( .A(n17358), .B(n19158), .ZN(n15037) );
  XNOR2_X1 U16445 ( .A(n15038), .B(n15037), .ZN(n15055) );
  OAI21_X1 U16446 ( .B1(n20449), .B2(n15138), .A(n20133), .ZN(n15040) );
  AOI21_X1 U16447 ( .B1(n15567), .B2(n15566), .A(n942), .ZN(n15041) );
  OAI22_X1 U16448 ( .A1(n15043), .A2(n15042), .B1(n20182), .B2(n15041), .ZN(
        n16707) );
  NOR2_X1 U16449 ( .A1(n15796), .A2(n15791), .ZN(n15044) );
  OAI21_X1 U16450 ( .B1(n15045), .B2(n15044), .A(n15577), .ZN(n15048) );
  OAI21_X1 U16451 ( .B1(n860), .B2(n15572), .A(n15574), .ZN(n15046) );
  NAND2_X1 U16452 ( .A1(n15046), .A2(n15796), .ZN(n15047) );
  NAND2_X1 U16453 ( .A1(n15048), .A2(n15047), .ZN(n16741) );
  INV_X1 U16454 ( .A(n15350), .ZN(n15050) );
  INV_X1 U16455 ( .A(n15459), .ZN(n15049) );
  AOI22_X1 U16456 ( .A1(n15050), .A2(n20173), .B1(n15348), .B2(n15049), .ZN(
        n15053) );
  NAND2_X1 U16457 ( .A1(n15459), .A2(n15350), .ZN(n15456) );
  OAI211_X1 U16458 ( .C1(n19759), .C2(n15350), .A(n15456), .B(n15353), .ZN(
        n15051) );
  XNOR2_X1 U16459 ( .A(n16741), .B(n16873), .ZN(n16355) );
  XNOR2_X1 U16460 ( .A(n16355), .B(n16822), .ZN(n15054) );
  XNOR2_X1 U16461 ( .A(n15054), .B(n15055), .ZN(n15220) );
  MUX2_X1 U16462 ( .A(n15553), .B(n15056), .S(n15551), .Z(n15058) );
  MUX2_X1 U16463 ( .A(n14903), .B(n20147), .S(n15549), .Z(n15057) );
  AOI22_X1 U16464 ( .A1(n15311), .A2(n15061), .B1(n15395), .B2(n15060), .ZN(
        n15063) );
  XNOR2_X1 U16466 ( .A(n16269), .B(n16690), .ZN(n15075) );
  NOR2_X1 U16468 ( .A1(n15402), .A2(n19838), .ZN(n15065) );
  NAND2_X1 U16469 ( .A1(n15065), .A2(n20006), .ZN(n15068) );
  NAND2_X1 U16470 ( .A1(n15066), .A2(n15898), .ZN(n15067) );
  AND3_X2 U16471 ( .A1(n15069), .A2(n15068), .A3(n15067), .ZN(n16770) );
  AND2_X1 U16472 ( .A1(n15070), .A2(n15618), .ZN(n15545) );
  NOR2_X1 U16473 ( .A1(n15546), .A2(n15071), .ZN(n15072) );
  XNOR2_X1 U16474 ( .A(n16770), .B(n17098), .ZN(n15074) );
  XNOR2_X1 U16475 ( .A(n15075), .B(n15074), .ZN(n15090) );
  INV_X1 U16477 ( .A(n15909), .ZN(n15915) );
  NOR2_X1 U16478 ( .A1(n15915), .A2(n15907), .ZN(n15076) );
  NAND3_X1 U16479 ( .A1(n15007), .A2(n15078), .A3(n15915), .ZN(n15079) );
  XNOR2_X1 U16480 ( .A(n16600), .B(n17411), .ZN(n15088) );
  NAND2_X1 U16481 ( .A1(n15081), .A2(n15430), .ZN(n15532) );
  NAND2_X1 U16482 ( .A1(n15082), .A2(n19676), .ZN(n15085) );
  NOR2_X1 U16483 ( .A1(n15921), .A2(n15422), .ZN(n15431) );
  XNOR2_X1 U16484 ( .A(n15087), .B(n15088), .ZN(n15089) );
  XNOR2_X2 U16485 ( .A(n15090), .B(n15089), .ZN(n17243) );
  MUX2_X1 U16486 ( .A(n15092), .B(n15091), .S(n15846), .Z(n15094) );
  MUX2_X1 U16487 ( .A(n15846), .B(n15845), .S(n15844), .Z(n15093) );
  XNOR2_X1 U16488 ( .A(n17035), .B(n16406), .ZN(n15106) );
  NOR2_X1 U16489 ( .A1(n15643), .A2(n15644), .ZN(n15095) );
  NOR2_X1 U16490 ( .A1(n19891), .A2(n15829), .ZN(n15097) );
  MUX2_X1 U16491 ( .A(n15258), .B(n15097), .S(n14997), .Z(n15098) );
  NOR2_X1 U16492 ( .A1(n15838), .A2(n15840), .ZN(n15105) );
  OAI21_X1 U16493 ( .B1(n15100), .B2(n15628), .A(n15625), .ZN(n15104) );
  NAND3_X1 U16494 ( .A1(n1288), .A2(n15836), .A3(n2472), .ZN(n15103) );
  NOR2_X1 U16495 ( .A1(n1288), .A2(n15628), .ZN(n15101) );
  XNOR2_X1 U16497 ( .A(n16835), .B(n15106), .ZN(n15137) );
  INV_X1 U16498 ( .A(n15296), .ZN(n15109) );
  NOR2_X1 U16500 ( .A1(n15275), .A2(n15270), .ZN(n15116) );
  NOR2_X1 U16501 ( .A1(n15601), .A2(n15276), .ZN(n15115) );
  MUX2_X1 U16502 ( .A(n15116), .B(n15115), .S(n15600), .Z(n15117) );
  XNOR2_X1 U16503 ( .A(n17269), .B(n17111), .ZN(n16546) );
  NAND3_X1 U16504 ( .A1(n15120), .A2(n15119), .A3(n20272), .ZN(n15124) );
  NAND4_X1 U16505 ( .A1(n15126), .A2(n15125), .A3(n15124), .A4(n15123), .ZN(
        n15128) );
  INV_X1 U16506 ( .A(n15129), .ZN(n15133) );
  NOR2_X1 U16507 ( .A1(n15282), .A2(n20474), .ZN(n15131) );
  INV_X1 U16508 ( .A(n645), .ZN(n15134) );
  XNOR2_X1 U16509 ( .A(n16893), .B(n15134), .ZN(n15135) );
  XNOR2_X1 U16510 ( .A(n16546), .B(n15135), .ZN(n15136) );
  XNOR2_X1 U16511 ( .A(n16945), .B(n2248), .ZN(n15145) );
  INV_X1 U16512 ( .A(n20449), .ZN(n15139) );
  NOR2_X1 U16513 ( .A1(n15139), .A2(n15138), .ZN(n15140) );
  NOR2_X1 U16514 ( .A1(n15701), .A2(n15696), .ZN(n15384) );
  MUX2_X1 U16515 ( .A(n15140), .B(n15384), .S(n15698), .Z(n15144) );
  OR2_X1 U16516 ( .A1(n15701), .A2(n15386), .ZN(n15142) );
  AOI22_X1 U16517 ( .A1(n15142), .A2(n15141), .B1(n15701), .B2(n15698), .ZN(
        n15143) );
  XNOR2_X1 U16519 ( .A(n19720), .B(n15145), .ZN(n15158) );
  NOR2_X1 U16520 ( .A1(n15712), .A2(n20178), .ZN(n15147) );
  NOR2_X1 U16522 ( .A1(n15147), .A2(n15146), .ZN(n15151) );
  NAND2_X1 U16524 ( .A1(n15152), .A2(n16015), .ZN(n15156) );
  OAI21_X1 U16525 ( .B1(n192), .B2(n20119), .A(n19739), .ZN(n15154) );
  OAI21_X2 U16526 ( .B1(n15156), .B2(n16016), .A(n15155), .ZN(n16854) );
  INV_X1 U16527 ( .A(n16854), .ZN(n15157) );
  XNOR2_X1 U16528 ( .A(n15157), .B(n16900), .ZN(n16342) );
  XNOR2_X1 U16529 ( .A(n16342), .B(n15158), .ZN(n15176) );
  OR2_X1 U16530 ( .A1(n15500), .A2(n15195), .ZN(n15162) );
  NOR2_X1 U16531 ( .A1(n15501), .A2(n15496), .ZN(n15190) );
  INV_X1 U16532 ( .A(n15190), .ZN(n15161) );
  INV_X1 U16533 ( .A(n15192), .ZN(n15499) );
  AND2_X1 U16534 ( .A1(n15501), .A2(n15499), .ZN(n15159) );
  OAI211_X1 U16535 ( .C1(n15378), .C2(n20467), .A(n15163), .B(n19513), .ZN(
        n15169) );
  OAI21_X1 U16536 ( .B1(n15167), .B2(n15166), .A(n15165), .ZN(n15168) );
  XNOR2_X1 U16537 ( .A(n17299), .B(n16615), .ZN(n15175) );
  INV_X1 U16538 ( .A(n15864), .ZN(n15329) );
  AOI21_X2 U16539 ( .B1(n15173), .B2(n15172), .A(n15171), .ZN(n17116) );
  INV_X1 U16540 ( .A(n17116), .ZN(n15174) );
  XNOR2_X1 U16541 ( .A(n15175), .B(n15174), .ZN(n15998) );
  INV_X1 U16542 ( .A(n20354), .ZN(n17484) );
  NAND2_X1 U16543 ( .A1(n15177), .A2(n17484), .ZN(n15254) );
  NOR2_X1 U16544 ( .A1(n15178), .A2(n15741), .ZN(n15179) );
  NAND2_X1 U16545 ( .A1(n15521), .A2(n19502), .ZN(n15184) );
  NAND3_X1 U16546 ( .A1(n15182), .A2(n15741), .A3(n15745), .ZN(n15183) );
  OAI21_X1 U16547 ( .B1(n15748), .B2(n15184), .A(n15183), .ZN(n15185) );
  XNOR2_X1 U16548 ( .A(n16608), .B(n17438), .ZN(n15199) );
  NAND2_X1 U16549 ( .A1(n15190), .A2(n15500), .ZN(n15198) );
  AOI21_X1 U16550 ( .B1(n19813), .B2(n15192), .A(n15191), .ZN(n15193) );
  AOI21_X1 U16551 ( .B1(n19512), .B2(n15501), .A(n15193), .ZN(n15197) );
  NOR2_X1 U16552 ( .A1(n15195), .A2(n19813), .ZN(n15196) );
  XNOR2_X1 U16553 ( .A(n16562), .B(n16746), .ZN(n15887) );
  XNOR2_X1 U16554 ( .A(n15199), .B(n15887), .ZN(n15219) );
  MUX2_X1 U16555 ( .A(n15495), .B(n16128), .S(n16129), .Z(n15203) );
  NOR2_X1 U16556 ( .A1(n16126), .A2(n15608), .ZN(n15200) );
  INV_X1 U16557 ( .A(n15758), .ZN(n15204) );
  OAI21_X1 U16558 ( .B1(n15758), .B2(n15754), .A(n15755), .ZN(n15207) );
  NAND2_X1 U16559 ( .A1(n15208), .A2(n15760), .ZN(n15206) );
  NAND3_X1 U16561 ( .A1(n15491), .A2(n2247), .A3(n15588), .ZN(n15205) );
  XNOR2_X1 U16562 ( .A(n16844), .B(n16747), .ZN(n15217) );
  NOR2_X1 U16563 ( .A1(n15559), .A2(n15513), .ZN(n15209) );
  NAND2_X1 U16564 ( .A1(n15212), .A2(n15560), .ZN(n15213) );
  AOI21_X1 U16565 ( .B1(n15211), .B2(n15213), .A(n15558), .ZN(n15214) );
  INV_X1 U16567 ( .A(n18779), .ZN(n18784) );
  XNOR2_X1 U16568 ( .A(n20477), .B(n18784), .ZN(n15216) );
  XNOR2_X1 U16569 ( .A(n15216), .B(n15217), .ZN(n15218) );
  INV_X1 U16570 ( .A(n15220), .ZN(n17483) );
  NAND2_X1 U16571 ( .A1(n17245), .A2(n17483), .ZN(n15252) );
  OR2_X1 U16572 ( .A1(n19884), .A2(n15221), .ZN(n15222) );
  AOI22_X1 U16573 ( .A1(n15438), .A2(n15222), .B1(n20151), .B2(n15770), .ZN(
        n15224) );
  NOR2_X1 U16574 ( .A1(n15222), .A2(n15673), .ZN(n15223) );
  OR2_X2 U16575 ( .A1(n15224), .A2(n15223), .ZN(n16760) );
  XNOR2_X1 U16576 ( .A(n16760), .B(n18997), .ZN(n15225) );
  INV_X1 U16577 ( .A(n15226), .ZN(n15227) );
  NAND2_X1 U16578 ( .A1(n15686), .A2(n15777), .ZN(n15451) );
  NOR2_X1 U16579 ( .A1(n15682), .A2(n15228), .ZN(n15449) );
  NAND3_X1 U16581 ( .A1(n15229), .A2(n15446), .A3(n1494), .ZN(n15230) );
  XNOR2_X1 U16582 ( .A(n16330), .B(n16861), .ZN(n16887) );
  INV_X1 U16584 ( .A(n15234), .ZN(n15236) );
  NAND2_X1 U16585 ( .A1(n15465), .A2(n15339), .ZN(n15338) );
  NAND2_X1 U16586 ( .A1(n15338), .A2(n15468), .ZN(n15233) );
  OAI21_X1 U16587 ( .B1(n15234), .B2(n15467), .A(n15233), .ZN(n15235) );
  OAI21_X1 U16588 ( .B1(n15470), .B2(n15236), .A(n15235), .ZN(n17367) );
  NAND2_X1 U16589 ( .A1(n15459), .A2(n15237), .ZN(n15238) );
  NAND2_X1 U16590 ( .A1(n15239), .A2(n15238), .ZN(n15242) );
  NOR2_X1 U16591 ( .A1(n19759), .A2(n1458), .ZN(n15240) );
  AOI22_X1 U16592 ( .A1(n15240), .A2(n15458), .B1(n1458), .B2(n15350), .ZN(
        n15241) );
  XNOR2_X1 U16593 ( .A(n17279), .B(n17367), .ZN(n15249) );
  INV_X1 U16594 ( .A(n15244), .ZN(n15248) );
  INV_X1 U16595 ( .A(n15245), .ZN(n15246) );
  XNOR2_X1 U16599 ( .A(n15250), .B(n15968), .ZN(n17480) );
  NOR2_X1 U16602 ( .A1(n18425), .A2(n18427), .ZN(n15255) );
  AOI21_X1 U16603 ( .B1(n19702), .B2(n18425), .A(n15255), .ZN(n15530) );
  MUX2_X1 U16604 ( .A(n15259), .B(n15258), .S(n14997), .Z(n15260) );
  AOI21_X2 U16605 ( .B1(n15261), .B2(n15829), .A(n15260), .ZN(n17099) );
  NOR2_X1 U16606 ( .A1(n15838), .A2(n15625), .ZN(n15265) );
  NAND2_X1 U16607 ( .A1(n15265), .A2(n15840), .ZN(n15263) );
  NAND3_X1 U16608 ( .A1(n1288), .A2(n15627), .A3(n15625), .ZN(n15262) );
  XNOR2_X1 U16609 ( .A(n17099), .B(n16987), .ZN(n16905) );
  MUX2_X1 U16610 ( .A(n15844), .B(n15266), .S(n15845), .Z(n15269) );
  MUX2_X1 U16611 ( .A(n15845), .B(n15267), .S(n15636), .Z(n15268) );
  XNOR2_X1 U16612 ( .A(n16905), .B(n16691), .ZN(n16577) );
  OAI211_X1 U16613 ( .C1(n20112), .C2(n15275), .A(n15272), .B(n15271), .ZN(
        n15280) );
  NOR2_X1 U16614 ( .A1(n15275), .A2(n15274), .ZN(n15599) );
  NAND2_X1 U16615 ( .A1(n15599), .A2(n15276), .ZN(n15279) );
  INV_X1 U16616 ( .A(Key[94]), .ZN(n19007) );
  INV_X1 U16617 ( .A(n15281), .ZN(n15290) );
  NAND2_X1 U16618 ( .A1(n15283), .A2(n15282), .ZN(n15289) );
  OAI22_X1 U16619 ( .A1(n15287), .A2(n15286), .B1(n15285), .B2(n19848), .ZN(
        n15288) );
  XNOR2_X1 U16621 ( .A(n15291), .B(n17102), .ZN(n15300) );
  NAND2_X1 U16622 ( .A1(n15293), .A2(n15292), .ZN(n15299) );
  NAND2_X1 U16623 ( .A1(n15294), .A2(n15295), .ZN(n15298) );
  XNOR2_X1 U16624 ( .A(n16600), .B(n16095), .ZN(n16384) );
  XNOR2_X1 U16625 ( .A(n15300), .B(n16384), .ZN(n15301) );
  XNOR2_X1 U16626 ( .A(n16577), .B(n15301), .ZN(n16166) );
  OAI21_X1 U16627 ( .B1(n15875), .B2(n198), .A(n15874), .ZN(n15304) );
  NAND2_X1 U16628 ( .A1(n20094), .A2(n15304), .ZN(n15305) );
  NAND2_X1 U16629 ( .A1(n15309), .A2(n15308), .ZN(n15394) );
  AND2_X1 U16630 ( .A1(n15312), .A2(n15676), .ZN(n15325) );
  NOR2_X1 U16631 ( .A1(n15314), .A2(n15313), .ZN(n15322) );
  INV_X1 U16632 ( .A(n15315), .ZN(n15318) );
  INV_X1 U16633 ( .A(n15316), .ZN(n15317) );
  NAND2_X1 U16634 ( .A1(n15318), .A2(n15317), .ZN(n15319) );
  MUX2_X1 U16635 ( .A(n15320), .B(n15319), .S(n2731), .Z(n15321) );
  INV_X1 U16636 ( .A(n15677), .ZN(n15447) );
  OAI211_X1 U16637 ( .C1(n15322), .C2(n15321), .A(n15447), .B(n15443), .ZN(
        n15323) );
  XNOR2_X1 U16638 ( .A(n20167), .B(n17358), .ZN(n15326) );
  XNOR2_X1 U16639 ( .A(n17141), .B(n15326), .ZN(n15347) );
  OAI21_X1 U16641 ( .B1(n15329), .B2(n15328), .A(n15866), .ZN(n15330) );
  AND2_X1 U16643 ( .A1(n901), .A2(n20119), .ZN(n15334) );
  XNOR2_X1 U16644 ( .A(n15979), .B(n19807), .ZN(n15345) );
  NAND2_X1 U16646 ( .A1(n15340), .A2(n15339), .ZN(n15342) );
  XNOR2_X1 U16647 ( .A(n19889), .B(n17787), .ZN(n15344) );
  XNOR2_X1 U16648 ( .A(n15345), .B(n15344), .ZN(n15346) );
  NAND2_X1 U16649 ( .A1(n20173), .A2(n15348), .ZN(n15462) );
  OAI21_X1 U16650 ( .B1(n15458), .B2(n15350), .A(n19759), .ZN(n15351) );
  XNOR2_X1 U16651 ( .A(n19954), .B(n16608), .ZN(n15362) );
  NAND2_X1 U16652 ( .A1(n15354), .A2(n233), .ZN(n15356) );
  NAND3_X1 U16653 ( .A1(n15815), .A2(n15582), .A3(n15583), .ZN(n15355) );
  NAND2_X1 U16654 ( .A1(n15356), .A2(n15355), .ZN(n15360) );
  NOR2_X1 U16655 ( .A1(n233), .A2(n15812), .ZN(n15358) );
  NOR2_X1 U16656 ( .A1(n3315), .A2(n15583), .ZN(n15357) );
  XNOR2_X1 U16657 ( .A(n16359), .B(n2369), .ZN(n15361) );
  XNOR2_X1 U16658 ( .A(n15362), .B(n15361), .ZN(n15393) );
  OAI21_X1 U16659 ( .B1(n860), .B2(n15573), .A(n15574), .ZN(n15363) );
  INV_X1 U16660 ( .A(n15363), .ZN(n15369) );
  NAND2_X1 U16661 ( .A1(n15364), .A2(n859), .ZN(n15368) );
  MUX2_X1 U16662 ( .A(n15566), .B(n15567), .S(n15370), .Z(n15374) );
  INV_X1 U16664 ( .A(n15565), .ZN(n15372) );
  XNOR2_X1 U16665 ( .A(n17127), .B(n16996), .ZN(n16882) );
  INV_X1 U16666 ( .A(n15375), .ZN(n15377) );
  NOR2_X1 U16667 ( .A1(n15379), .A2(n231), .ZN(n15376) );
  NOR2_X1 U16668 ( .A1(n15377), .A2(n15376), .ZN(n15383) );
  NAND2_X1 U16669 ( .A1(n15384), .A2(n20133), .ZN(n15391) );
  NAND2_X1 U16670 ( .A1(n15386), .A2(n15695), .ZN(n15387) );
  NAND3_X1 U16671 ( .A1(n15701), .A2(n15702), .A3(n15387), .ZN(n15390) );
  NAND3_X1 U16672 ( .A1(n15385), .A2(n15696), .A3(n15698), .ZN(n15389) );
  NAND3_X1 U16673 ( .A1(n15387), .A2(n15702), .A3(n15386), .ZN(n15388) );
  NAND4_X1 U16674 ( .A1(n15391), .A2(n15390), .A3(n15389), .A4(n15388), .ZN(
        n17442) );
  XNOR2_X1 U16675 ( .A(n17442), .B(n16840), .ZN(n16102) );
  XNOR2_X1 U16676 ( .A(n16882), .B(n16102), .ZN(n15392) );
  XNOR2_X1 U16677 ( .A(n15392), .B(n15393), .ZN(n16165) );
  NAND3_X1 U16678 ( .A1(n17505), .A2(n17501), .A3(n16165), .ZN(n16443) );
  OAI22_X1 U16679 ( .A1(n15397), .A2(n15396), .B1(n15395), .B2(n15394), .ZN(
        n15398) );
  XNOR2_X1 U16680 ( .A(n16761), .B(n17367), .ZN(n16380) );
  OAI211_X1 U16682 ( .C1(n20006), .C2(n15892), .A(n15402), .B(n15536), .ZN(
        n15404) );
  XNOR2_X1 U16683 ( .A(n17135), .B(n16380), .ZN(n15436) );
  XNOR2_X1 U16684 ( .A(n17133), .B(n2420), .ZN(n15434) );
  OR2_X1 U16685 ( .A1(n15417), .A2(n15416), .ZN(n15418) );
  OAI21_X2 U16686 ( .B1(n15912), .B2(n15419), .A(n15418), .ZN(n17276) );
  OAI21_X1 U16688 ( .B1(n15426), .B2(n15423), .A(n15422), .ZN(n15429) );
  INV_X1 U16689 ( .A(n15424), .ZN(n15425) );
  NOR2_X1 U16690 ( .A1(n15426), .A2(n15425), .ZN(n15428) );
  NAND2_X1 U16691 ( .A1(n15430), .A2(n15531), .ZN(n15427) );
  INV_X1 U16693 ( .A(n15431), .ZN(n15432) );
  AOI22_X2 U16694 ( .A1(n15917), .A2(n15534), .B1(n15433), .B2(n15432), .ZN(
        n16971) );
  XNOR2_X1 U16695 ( .A(n17276), .B(n16971), .ZN(n16567) );
  XNOR2_X1 U16696 ( .A(n15434), .B(n16567), .ZN(n15435) );
  XNOR2_X1 U16697 ( .A(n15436), .B(n15435), .ZN(n15485) );
  NOR2_X1 U16698 ( .A1(n15665), .A2(n19884), .ZN(n15437) );
  OAI21_X1 U16699 ( .B1(n15438), .B2(n15437), .A(n15673), .ZN(n15441) );
  AND2_X1 U16700 ( .A1(n19884), .A2(n15666), .ZN(n15439) );
  NAND2_X1 U16701 ( .A1(n15441), .A2(n15440), .ZN(n16134) );
  NAND2_X1 U16703 ( .A1(n15446), .A2(n15443), .ZN(n15444) );
  NAND2_X1 U16704 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  XNOR2_X1 U16705 ( .A(n16134), .B(n20481), .ZN(n16898) );
  NAND2_X1 U16706 ( .A1(n15783), .A2(n15684), .ZN(n15450) );
  OAI211_X1 U16710 ( .C1(n15459), .C2(n20173), .A(n15456), .B(n1458), .ZN(
        n15463) );
  NAND3_X1 U16711 ( .A1(n15460), .A2(n15459), .A3(n15458), .ZN(n15461) );
  AND3_X1 U16712 ( .A1(n15463), .A2(n15462), .A3(n15461), .ZN(n16367) );
  XNOR2_X1 U16713 ( .A(n16963), .B(n16367), .ZN(n15633) );
  XNOR2_X1 U16714 ( .A(n16898), .B(n15633), .ZN(n15483) );
  NOR2_X1 U16715 ( .A1(n15470), .A2(n15468), .ZN(n15471) );
  XNOR2_X1 U16716 ( .A(n16615), .B(n17298), .ZN(n15481) );
  NOR2_X1 U16717 ( .A1(n15766), .A2(n15769), .ZN(n15473) );
  AND2_X1 U16719 ( .A1(n12658), .A2(n15657), .ZN(n15654) );
  INV_X1 U16720 ( .A(n15654), .ZN(n15477) );
  NAND3_X1 U16721 ( .A1(n15475), .A2(n15658), .A3(n15653), .ZN(n15476) );
  XNOR2_X1 U16722 ( .A(n17401), .B(n17909), .ZN(n15480) );
  XNOR2_X1 U16723 ( .A(n15481), .B(n15480), .ZN(n15482) );
  XNOR2_X1 U16724 ( .A(n15483), .B(n15482), .ZN(n17498) );
  AOI21_X1 U16728 ( .B1(n1683), .B2(n2247), .A(n15755), .ZN(n15493) );
  NAND3_X1 U16729 ( .A1(n15488), .A2(n15757), .A3(n15487), .ZN(n15489) );
  NOR2_X1 U16730 ( .A1(n15759), .A2(n15489), .ZN(n15492) );
  NOR2_X1 U16731 ( .A1(n15491), .A2(n15490), .ZN(n15761) );
  NOR2_X1 U16732 ( .A1(n16126), .A2(n16128), .ZN(n15494) );
  NAND2_X1 U16733 ( .A1(n1019), .A2(n15503), .ZN(n15821) );
  NAND2_X1 U16734 ( .A1(n15506), .A2(n15505), .ZN(n15824) );
  OR2_X1 U16735 ( .A1(n15824), .A2(n13933), .ZN(n15508) );
  XNOR2_X1 U16736 ( .A(n16892), .B(n15726), .ZN(n15526) );
  NAND2_X1 U16737 ( .A1(n15511), .A2(n15513), .ZN(n15512) );
  XNOR2_X1 U16738 ( .A(n17035), .B(n19909), .ZN(n15524) );
  NOR2_X1 U16739 ( .A1(n15746), .A2(n15516), .ZN(n15595) );
  INV_X1 U16740 ( .A(n15741), .ZN(n15517) );
  NAND3_X1 U16741 ( .A1(n15517), .A2(n15742), .A3(n19502), .ZN(n15518) );
  XNOR2_X1 U16744 ( .A(n16335), .B(n2123), .ZN(n15523) );
  XNOR2_X1 U16745 ( .A(n15524), .B(n15523), .ZN(n15525) );
  OAI21_X1 U16747 ( .B1(n20168), .B2(n19815), .A(n19898), .ZN(n15527) );
  NAND2_X1 U16748 ( .A1(n15527), .A2(n16480), .ZN(n15528) );
  NAND2_X1 U16749 ( .A1(n15530), .A2(n15529), .ZN(n15930) );
  XNOR2_X1 U16750 ( .A(n17002), .B(n16236), .ZN(n15543) );
  OAI21_X1 U16752 ( .B1(n15539), .B2(n15538), .A(n15537), .ZN(n15542) );
  XNOR2_X1 U16753 ( .A(n17355), .B(n16181), .ZN(n17419) );
  XNOR2_X1 U16754 ( .A(n17419), .B(n15543), .ZN(n15557) );
  NOR2_X1 U16755 ( .A1(n15545), .A2(n15544), .ZN(n15548) );
  AOI21_X1 U16756 ( .B1(n15550), .B2(n15549), .A(n14903), .ZN(n15552) );
  XNOR2_X1 U16757 ( .A(n17359), .B(n16872), .ZN(n15555) );
  XNOR2_X1 U16758 ( .A(n19889), .B(n18984), .ZN(n15554) );
  XNOR2_X1 U16759 ( .A(n15555), .B(n15554), .ZN(n15556) );
  INV_X1 U16760 ( .A(n16666), .ZN(n17221) );
  INV_X1 U16762 ( .A(n15566), .ZN(n15800) );
  NAND3_X1 U16763 ( .A1(n15800), .A2(n15567), .A3(n15371), .ZN(n15568) );
  XNOR2_X1 U16765 ( .A(n17014), .B(n16788), .ZN(n15571) );
  AND2_X1 U16767 ( .A1(n15572), .A2(n15573), .ZN(n15576) );
  NAND2_X1 U16768 ( .A1(n15574), .A2(n15573), .ZN(n15575) );
  MUX2_X1 U16769 ( .A(n15576), .B(n15575), .S(n860), .Z(n15578) );
  XNOR2_X1 U16770 ( .A(n16095), .B(n19713), .ZN(n15579) );
  MUX2_X1 U16772 ( .A(n15582), .B(n15812), .S(n15815), .Z(n15585) );
  MUX2_X2 U16773 ( .A(n15585), .B(n15584), .S(n233), .Z(n17406) );
  XNOR2_X1 U16774 ( .A(n15586), .B(n16132), .ZN(n16639) );
  INV_X1 U16775 ( .A(n16641), .ZN(n15731) );
  INV_X1 U16776 ( .A(n16639), .ZN(n19385) );
  XNOR2_X1 U16777 ( .A(n16761), .B(n2381), .ZN(n15592) );
  MUX2_X1 U16779 ( .A(n15589), .B(n15755), .S(n15760), .Z(n15590) );
  XNOR2_X1 U16780 ( .A(n15592), .B(n16928), .ZN(n15598) );
  NAND2_X1 U16781 ( .A1(n3821), .A2(n15741), .ZN(n15597) );
  NAND2_X1 U16782 ( .A1(n15744), .A2(n15595), .ZN(n15596) );
  XNOR2_X1 U16784 ( .A(n16886), .B(n17133), .ZN(n16146) );
  XNOR2_X1 U16785 ( .A(n15598), .B(n16146), .ZN(n15613) );
  INV_X1 U16786 ( .A(n15599), .ZN(n15603) );
  NOR2_X1 U16787 ( .A1(n15601), .A2(n15600), .ZN(n15602) );
  NOR2_X1 U16788 ( .A1(n15608), .A2(n16129), .ZN(n15610) );
  NOR2_X1 U16789 ( .A1(n3427), .A2(n16128), .ZN(n15609) );
  AOI22_X1 U16790 ( .A1(n15733), .A2(n15610), .B1(n15609), .B2(n16126), .ZN(
        n15611) );
  XNOR2_X1 U16791 ( .A(n16970), .B(n16932), .ZN(n17431) );
  XNOR2_X1 U16792 ( .A(n17431), .B(n16329), .ZN(n15612) );
  OAI22_X1 U16793 ( .A1(n15616), .A2(n20138), .B1(n15620), .B2(n15614), .ZN(
        n15624) );
  INV_X1 U16794 ( .A(n15617), .ZN(n15622) );
  NAND3_X1 U16795 ( .A1(n15620), .A2(n15619), .A3(n15618), .ZN(n15621) );
  NAND2_X1 U16796 ( .A1(n15622), .A2(n15621), .ZN(n15623) );
  INV_X1 U16797 ( .A(n15840), .ZN(n15629) );
  NAND2_X1 U16798 ( .A1(n15629), .A2(n15625), .ZN(n15632) );
  NAND3_X1 U16799 ( .A1(n15629), .A2(n1288), .A3(n15628), .ZN(n15630) );
  OAI211_X1 U16800 ( .C1(n15838), .C2(n15632), .A(n15631), .B(n15630), .ZN(
        n16947) );
  XNOR2_X1 U16801 ( .A(n16947), .B(n16960), .ZN(n17399) );
  XNOR2_X1 U16802 ( .A(n17399), .B(n15633), .ZN(n15652) );
  NOR2_X1 U16804 ( .A1(n15844), .A2(n868), .ZN(n15634) );
  NAND2_X1 U16805 ( .A1(n15845), .A2(n15634), .ZN(n15638) );
  NOR2_X1 U16806 ( .A1(n15846), .A2(n868), .ZN(n15635) );
  XNOR2_X1 U16808 ( .A(n16227), .B(n16412), .ZN(n16902) );
  NAND3_X1 U16809 ( .A1(n15643), .A2(n15645), .A3(n15642), .ZN(n15648) );
  NAND3_X1 U16810 ( .A1(n15645), .A2(n15644), .A3(n19931), .ZN(n15647) );
  XNOR2_X1 U16811 ( .A(n17330), .B(n18478), .ZN(n15650) );
  XNOR2_X1 U16812 ( .A(n16902), .B(n15650), .ZN(n15651) );
  XNOR2_X1 U16813 ( .A(n15651), .B(n15652), .ZN(n19382) );
  INV_X1 U16814 ( .A(n19382), .ZN(n17218) );
  XNOR2_X1 U16815 ( .A(n16240), .B(n16840), .ZN(n15675) );
  NAND2_X1 U16816 ( .A1(n15654), .A2(n15653), .ZN(n15663) );
  NAND3_X1 U16817 ( .A1(n15659), .A2(n15658), .A3(n15657), .ZN(n15662) );
  NAND3_X1 U16818 ( .A1(n15768), .A2(n15769), .A3(n15660), .ZN(n15661) );
  INV_X1 U16819 ( .A(n19879), .ZN(n15773) );
  NAND3_X1 U16820 ( .A1(n15773), .A2(n15665), .A3(n13414), .ZN(n15669) );
  NAND2_X1 U16821 ( .A1(n19879), .A2(n20151), .ZN(n15674) );
  XNOR2_X1 U16822 ( .A(n16295), .B(n955), .ZN(n17440) );
  XNOR2_X1 U16823 ( .A(n15675), .B(n17440), .ZN(n15694) );
  NOR2_X1 U16824 ( .A1(n15679), .A2(n15677), .ZN(n15681) );
  INV_X1 U16825 ( .A(n15678), .ZN(n15680) );
  INV_X1 U16826 ( .A(n2122), .ZN(n18598) );
  XNOR2_X1 U16827 ( .A(n17444), .B(n18598), .ZN(n15692) );
  NAND2_X1 U16828 ( .A1(n19977), .A2(n15683), .ZN(n15785) );
  NAND3_X1 U16829 ( .A1(n19978), .A2(n15782), .A3(n15684), .ZN(n15690) );
  XNOR2_X1 U16830 ( .A(n16292), .B(n19798), .ZN(n16513) );
  XNOR2_X1 U16831 ( .A(n15692), .B(n16513), .ZN(n15693) );
  XNOR2_X1 U16832 ( .A(n15694), .B(n15693), .ZN(n19386) );
  MUX2_X1 U16833 ( .A(n15701), .B(n15696), .S(n15695), .Z(n15703) );
  AND2_X1 U16834 ( .A1(n15702), .A2(n15698), .ZN(n15700) );
  OAI21_X1 U16835 ( .B1(n15885), .B2(n15705), .A(n15704), .ZN(n15707) );
  INV_X1 U16836 ( .A(n15957), .ZN(n15708) );
  XNOR2_X1 U16837 ( .A(n17335), .B(n15708), .ZN(n17424) );
  INV_X1 U16838 ( .A(n15874), .ZN(n15871) );
  NAND3_X1 U16839 ( .A1(n15871), .A2(n20178), .A3(n15875), .ZN(n15710) );
  OAI21_X1 U16840 ( .B1(n15712), .B2(n15711), .A(n15710), .ZN(n15718) );
  INV_X1 U16841 ( .A(n15713), .ZN(n15716) );
  XNOR2_X1 U16842 ( .A(n16027), .B(n17095), .ZN(n15719) );
  XNOR2_X1 U16843 ( .A(n17424), .B(n15719), .ZN(n15728) );
  OAI21_X1 U16844 ( .B1(n15864), .B2(n15720), .A(n15863), .ZN(n15724) );
  NOR3_X1 U16845 ( .A1(n15866), .A2(n15722), .A3(n15721), .ZN(n15723) );
  XNOR2_X1 U16846 ( .A(n20102), .B(n16336), .ZN(n16891) );
  XNOR2_X1 U16847 ( .A(n16891), .B(n15726), .ZN(n15727) );
  XNOR2_X1 U16848 ( .A(n15727), .B(n15728), .ZN(n16665) );
  OAI211_X1 U16849 ( .C1(n19386), .C2(n16666), .A(n19383), .B(n1897), .ZN(
        n15729) );
  INV_X1 U16850 ( .A(n15729), .ZN(n15730) );
  NOR2_X1 U16851 ( .A1(n20003), .A2(n18412), .ZN(n18424) );
  OAI211_X1 U16852 ( .C1(n15495), .C2(n15737), .A(n15736), .B(n15735), .ZN(
        n16097) );
  XNOR2_X1 U16853 ( .A(n15739), .B(n16097), .ZN(n15753) );
  INV_X1 U16854 ( .A(n15740), .ZN(n15752) );
  NAND2_X1 U16855 ( .A1(n15742), .A2(n15741), .ZN(n15743) );
  NAND2_X1 U16856 ( .A1(n15743), .A2(n15745), .ZN(n15751) );
  NOR3_X1 U16857 ( .A1(n15748), .A2(n15182), .A3(n15745), .ZN(n15747) );
  AOI21_X1 U16858 ( .B1(n15749), .B2(n15748), .A(n15747), .ZN(n15750) );
  OAI21_X1 U16859 ( .B1(n15752), .B2(n15751), .A(n15750), .ZN(n16188) );
  XNOR2_X1 U16860 ( .A(n15753), .B(n16188), .ZN(n17101) );
  XNOR2_X1 U16861 ( .A(n16269), .B(n16095), .ZN(n16772) );
  XNOR2_X1 U16862 ( .A(n17101), .B(n16772), .ZN(n15764) );
  XNOR2_X1 U16863 ( .A(n17410), .B(n457), .ZN(n15762) );
  XNOR2_X1 U16864 ( .A(n15762), .B(n19820), .ZN(n15763) );
  XNOR2_X1 U16866 ( .A(n16742), .B(n16873), .ZN(n16071) );
  NAND2_X1 U16867 ( .A1(n15771), .A2(n15770), .ZN(n15776) );
  NAND2_X1 U16868 ( .A1(n15778), .A2(n19977), .ZN(n15787) );
  NAND3_X1 U16869 ( .A1(n15783), .A2(n15782), .A3(n20362), .ZN(n15784) );
  XNOR2_X1 U16871 ( .A(n16278), .B(n16939), .ZN(n17003) );
  XNOR2_X1 U16872 ( .A(n17003), .B(n16071), .ZN(n15790) );
  INV_X1 U16873 ( .A(n2347), .ZN(n19259) );
  XNOR2_X1 U16874 ( .A(n16554), .B(n19259), .ZN(n15788) );
  XNOR2_X1 U16875 ( .A(n19889), .B(n17416), .ZN(n16107) );
  XNOR2_X1 U16876 ( .A(n16107), .B(n15788), .ZN(n15789) );
  INV_X1 U16877 ( .A(n16540), .ZN(n19353) );
  NOR2_X1 U16878 ( .A1(n19354), .A2(n19353), .ZN(n16674) );
  MUX2_X1 U16879 ( .A(n860), .B(n1520), .S(n15365), .Z(n15797) );
  OAI21_X1 U16880 ( .B1(n15800), .B2(n15371), .A(n20182), .ZN(n15807) );
  NAND3_X1 U16882 ( .A1(n15804), .A2(n942), .A3(n15803), .ZN(n15805) );
  XNOR2_X1 U16883 ( .A(n17269), .B(n19674), .ZN(n15809) );
  XNOR2_X1 U16884 ( .A(n15810), .B(n15809), .ZN(n15827) );
  NAND2_X1 U16885 ( .A1(n15814), .A2(n15813), .ZN(n15817) );
  XNOR2_X1 U16886 ( .A(n17110), .B(n16893), .ZN(n16054) );
  AND2_X1 U16887 ( .A1(n15821), .A2(n15820), .ZN(n15826) );
  NAND2_X1 U16888 ( .A1(n15822), .A2(n1758), .ZN(n15823) );
  MUX2_X1 U16889 ( .A(n15824), .B(n15823), .S(n13933), .Z(n15825) );
  NAND2_X1 U16890 ( .A1(n15826), .A2(n15825), .ZN(n16081) );
  XNOR2_X1 U16891 ( .A(n16054), .B(n16081), .ZN(n16758) );
  NOR2_X1 U16892 ( .A1(n15829), .A2(n15828), .ZN(n15830) );
  OAI21_X1 U16893 ( .B1(n15642), .B2(n15831), .A(n15830), .ZN(n15834) );
  NAND2_X1 U16894 ( .A1(n15832), .A2(n15257), .ZN(n15833) );
  INV_X1 U16895 ( .A(n16975), .ZN(n15842) );
  XNOR2_X1 U16896 ( .A(n15842), .B(n16973), .ZN(n16214) );
  NAND2_X1 U16898 ( .A1(n15845), .A2(n15844), .ZN(n15850) );
  NAND3_X1 U16899 ( .A1(n15847), .A2(n15846), .A3(n2146), .ZN(n15849) );
  XNOR2_X1 U16901 ( .A(n16761), .B(n15852), .ZN(n16089) );
  XNOR2_X1 U16902 ( .A(n17279), .B(n2079), .ZN(n15853) );
  XNOR2_X1 U16903 ( .A(n15853), .B(n16089), .ZN(n15854) );
  XNOR2_X1 U16904 ( .A(n15854), .B(n15855), .ZN(n16672) );
  AND2_X1 U16905 ( .A1(n16672), .A2(n19349), .ZN(n15856) );
  OR2_X1 U16906 ( .A1(n16674), .A2(n15856), .ZN(n15929) );
  NAND2_X1 U16907 ( .A1(n15859), .A2(n15858), .ZN(n15869) );
  NOR2_X1 U16908 ( .A1(n15863), .A2(n15862), .ZN(n15865) );
  INV_X1 U16910 ( .A(n2442), .ZN(n18924) );
  XNOR2_X1 U16911 ( .A(n17124), .B(n18924), .ZN(n15886) );
  NOR2_X1 U16912 ( .A1(n15875), .A2(n15871), .ZN(n15872) );
  NOR2_X2 U16913 ( .A1(n15878), .A2(n15877), .ZN(n17439) );
  NAND2_X1 U16914 ( .A1(n16012), .A2(n20119), .ZN(n15884) );
  OAI21_X1 U16915 ( .B1(n16009), .B2(n901), .A(n15880), .ZN(n15881) );
  NAND2_X1 U16916 ( .A1(n15881), .A2(n3473), .ZN(n15883) );
  NAND3_X1 U16917 ( .A1(n16009), .A2(n16010), .A3(n16015), .ZN(n15882) );
  OAI211_X1 U16918 ( .C1(n15885), .C2(n15884), .A(n15883), .B(n15882), .ZN(
        n17128) );
  XNOR2_X1 U16919 ( .A(n17128), .B(n17439), .ZN(n16998) );
  XNOR2_X1 U16920 ( .A(n15886), .B(n16998), .ZN(n15889) );
  XNOR2_X1 U16921 ( .A(n16102), .B(n15887), .ZN(n15888) );
  NAND2_X1 U16922 ( .A1(n19352), .A2(n19348), .ZN(n15927) );
  INV_X1 U16923 ( .A(n15892), .ZN(n15895) );
  OAI22_X1 U16925 ( .A1(n15891), .A2(n15890), .B1(n15895), .B2(n19722), .ZN(
        n15902) );
  NAND2_X1 U16926 ( .A1(n19722), .A2(n15892), .ZN(n15899) );
  OAI21_X1 U16927 ( .B1(n15899), .B2(n15898), .A(n15897), .ZN(n15900) );
  INV_X1 U16928 ( .A(n15900), .ZN(n15901) );
  XNOR2_X1 U16929 ( .A(n16900), .B(n16283), .ZN(n15904) );
  XNOR2_X1 U16930 ( .A(n20104), .B(n18726), .ZN(n15903) );
  XNOR2_X1 U16931 ( .A(n15904), .B(n15903), .ZN(n15926) );
  AOI21_X1 U16932 ( .B1(n2723), .B2(n15906), .A(n15905), .ZN(n15914) );
  INV_X1 U16933 ( .A(n15907), .ZN(n15908) );
  NOR2_X1 U16934 ( .A1(n15909), .A2(n15908), .ZN(n15911) );
  OAI21_X1 U16935 ( .B1(n15912), .B2(n15911), .A(n15910), .ZN(n15913) );
  XNOR2_X1 U16936 ( .A(n16225), .B(n16367), .ZN(n16851) );
  AND2_X1 U16937 ( .A1(n15917), .A2(n15916), .ZN(n15924) );
  MUX2_X1 U16938 ( .A(n15920), .B(n15919), .S(n19752), .Z(n15923) );
  XNOR2_X1 U16939 ( .A(n16224), .B(n17401), .ZN(n17120) );
  XNOR2_X1 U16940 ( .A(n16851), .B(n17120), .ZN(n15925) );
  XNOR2_X1 U16941 ( .A(n15925), .B(n15926), .ZN(n19347) );
  INV_X1 U16942 ( .A(n19347), .ZN(n19351) );
  AOI21_X1 U16943 ( .B1(n15927), .B2(n19351), .A(n19349), .ZN(n15928) );
  NOR2_X1 U16944 ( .A1(n18400), .A2(n18423), .ZN(n18414) );
  XNOR2_X1 U16946 ( .A(n16181), .B(n20450), .ZN(n15934) );
  INV_X1 U16947 ( .A(n17466), .ZN(n15932) );
  XNOR2_X1 U16948 ( .A(n864), .B(n15932), .ZN(n15933) );
  XNOR2_X1 U16949 ( .A(n15934), .B(n15933), .ZN(n15938) );
  XNOR2_X1 U16950 ( .A(n15936), .B(n15935), .ZN(n16534) );
  XNOR2_X1 U16951 ( .A(n16938), .B(n16278), .ZN(n17418) );
  XNOR2_X1 U16952 ( .A(n17418), .B(n16534), .ZN(n15937) );
  XNOR2_X1 U16954 ( .A(n16932), .B(n17275), .ZN(n17028) );
  XNOR2_X1 U16955 ( .A(n16522), .B(n17028), .ZN(n15942) );
  XNOR2_X1 U16956 ( .A(n16974), .B(n16568), .ZN(n15940) );
  XNOR2_X1 U16957 ( .A(n16975), .B(n2208), .ZN(n15939) );
  XNOR2_X1 U16958 ( .A(n15940), .B(n15939), .ZN(n15941) );
  XNOR2_X1 U16960 ( .A(n16964), .B(n16283), .ZN(n15943) );
  XNOR2_X1 U16961 ( .A(n16528), .B(n15943), .ZN(n15946) );
  XNOR2_X1 U16962 ( .A(n16947), .B(n19929), .ZN(n17020) );
  XNOR2_X1 U16963 ( .A(n16134), .B(n2298), .ZN(n15944) );
  XNOR2_X1 U16964 ( .A(n17020), .B(n15944), .ZN(n15945) );
  XNOR2_X1 U16965 ( .A(n15946), .B(n15945), .ZN(n17080) );
  NAND2_X1 U16966 ( .A1(n17823), .A2(n17080), .ZN(n17828) );
  XNOR2_X1 U16967 ( .A(n17099), .B(n19783), .ZN(n15948) );
  XNOR2_X1 U16968 ( .A(n17288), .B(n18055), .ZN(n15947) );
  XNOR2_X1 U16969 ( .A(n15948), .B(n15947), .ZN(n15950) );
  XNOR2_X1 U16970 ( .A(n16602), .B(n17014), .ZN(n17409) );
  XNOR2_X1 U16971 ( .A(n17104), .B(n17410), .ZN(n16990) );
  XNOR2_X1 U16972 ( .A(n17409), .B(n16990), .ZN(n15949) );
  NOR2_X1 U16973 ( .A1(n17825), .A2(n17172), .ZN(n16777) );
  AOI21_X1 U16974 ( .B1(n20239), .B2(n17828), .A(n16777), .ZN(n15965) );
  XNOR2_X1 U16975 ( .A(n15951), .B(n17439), .ZN(n15952) );
  XNOR2_X1 U16976 ( .A(n947), .B(n955), .ZN(n17046) );
  XNOR2_X1 U16977 ( .A(n17046), .B(n15952), .ZN(n15954) );
  XNOR2_X1 U16978 ( .A(n15953), .B(n15954), .ZN(n16262) );
  INV_X1 U16979 ( .A(n17823), .ZN(n15962) );
  XNOR2_X1 U16980 ( .A(n16981), .B(n17109), .ZN(n15956) );
  XNOR2_X1 U16981 ( .A(n17425), .B(n16300), .ZN(n15955) );
  XNOR2_X1 U16982 ( .A(n15956), .B(n15955), .ZN(n15961) );
  XNOR2_X1 U16983 ( .A(n16836), .B(n17426), .ZN(n15959) );
  XNOR2_X1 U16984 ( .A(n902), .B(n19205), .ZN(n15958) );
  XNOR2_X1 U16985 ( .A(n15959), .B(n15958), .ZN(n15960) );
  XNOR2_X1 U16986 ( .A(n15961), .B(n15960), .ZN(n16263) );
  NAND2_X1 U16987 ( .A1(n15962), .A2(n17079), .ZN(n15963) );
  AOI21_X1 U16988 ( .B1(n16262), .B2(n20239), .A(n15963), .ZN(n15964) );
  XNOR2_X1 U16989 ( .A(n17280), .B(n19102), .ZN(n15966) );
  XNOR2_X1 U16990 ( .A(n15966), .B(n16971), .ZN(n15967) );
  XNOR2_X1 U16991 ( .A(n20098), .B(n16928), .ZN(n16521) );
  XNOR2_X1 U16992 ( .A(n15967), .B(n16521), .ZN(n15969) );
  XNOR2_X1 U16994 ( .A(n17291), .B(n19713), .ZN(n16518) );
  XNOR2_X1 U16995 ( .A(n15970), .B(n16690), .ZN(n16574) );
  XNOR2_X1 U16996 ( .A(n16574), .B(n16518), .ZN(n15974) );
  XNOR2_X1 U16997 ( .A(n17012), .B(n16987), .ZN(n15972) );
  XNOR2_X1 U16998 ( .A(n16600), .B(n2275), .ZN(n15971) );
  XNOR2_X1 U16999 ( .A(n15972), .B(n15971), .ZN(n15973) );
  NOR2_X1 U17001 ( .A1(n20275), .A2(n20507), .ZN(n16003) );
  INV_X1 U17002 ( .A(n20507), .ZN(n17074) );
  XNOR2_X1 U17003 ( .A(n17379), .B(n2164), .ZN(n15975) );
  XNOR2_X1 U17004 ( .A(n15975), .B(n16996), .ZN(n15976) );
  XNOR2_X1 U17005 ( .A(n16750), .B(n16562), .ZN(n17259) );
  XNOR2_X1 U17006 ( .A(n17259), .B(n15976), .ZN(n15978) );
  XNOR2_X1 U17007 ( .A(n20478), .B(n17260), .ZN(n17048) );
  XNOR2_X1 U17008 ( .A(n17048), .B(n16608), .ZN(n15977) );
  XNOR2_X1 U17009 ( .A(n16554), .B(n16743), .ZN(n17250) );
  XNOR2_X1 U17010 ( .A(n17358), .B(n17253), .ZN(n17040) );
  XNOR2_X1 U17011 ( .A(n17250), .B(n17040), .ZN(n15983) );
  INV_X1 U17012 ( .A(n2296), .ZN(n15980) );
  XNOR2_X1 U17013 ( .A(n17359), .B(n15980), .ZN(n15981) );
  XNOR2_X1 U17014 ( .A(n16553), .B(n15981), .ZN(n15982) );
  OAI21_X1 U17015 ( .B1(n17074), .B2(n20514), .A(n17872), .ZN(n16002) );
  XNOR2_X1 U17018 ( .A(n20372), .B(n16546), .ZN(n15988) );
  XNOR2_X1 U17019 ( .A(n16027), .B(n16980), .ZN(n15986) );
  XNOR2_X1 U17020 ( .A(n16755), .B(n17999), .ZN(n15985) );
  XNOR2_X1 U17021 ( .A(n15986), .B(n15985), .ZN(n15987) );
  NAND2_X1 U17022 ( .A1(n16003), .A2(n17676), .ZN(n16001) );
  INV_X1 U17023 ( .A(n17872), .ZN(n17868) );
  OAI21_X1 U17024 ( .B1(n15991), .B2(n15990), .A(n15989), .ZN(n15993) );
  NAND2_X1 U17025 ( .A1(n15993), .A2(n15992), .ZN(n17293) );
  XNOR2_X1 U17026 ( .A(n15994), .B(n2222), .ZN(n15995) );
  XNOR2_X1 U17027 ( .A(n15995), .B(n17293), .ZN(n15997) );
  XNOR2_X1 U17028 ( .A(n17294), .B(n16965), .ZN(n15996) );
  XNOR2_X1 U17029 ( .A(n15997), .B(n15996), .ZN(n15999) );
  XNOR2_X1 U17030 ( .A(n15998), .B(n15999), .ZN(n17867) );
  INV_X1 U17031 ( .A(n17867), .ZN(n17078) );
  OAI211_X1 U17033 ( .C1(n16003), .C2(n16002), .A(n16001), .B(n16000), .ZN(
        n16155) );
  XNOR2_X1 U17034 ( .A(n17378), .B(n17439), .ZN(n16294) );
  XNOR2_X1 U17035 ( .A(n19799), .B(n19216), .ZN(n16004) );
  XNOR2_X1 U17036 ( .A(n16607), .B(n16004), .ZN(n16005) );
  XNOR2_X1 U17037 ( .A(n16294), .B(n16005), .ZN(n16007) );
  XNOR2_X1 U17038 ( .A(n16844), .B(n16914), .ZN(n16390) );
  XNOR2_X1 U17039 ( .A(n16390), .B(n17438), .ZN(n16006) );
  XNOR2_X1 U17040 ( .A(n16007), .B(n16006), .ZN(n17898) );
  NAND3_X1 U17041 ( .A1(n16009), .A2(n19739), .A3(n16015), .ZN(n16014) );
  OAI21_X1 U17042 ( .B1(n16012), .B2(n901), .A(n16010), .ZN(n16013) );
  OAI211_X1 U17043 ( .C1(n16016), .C2(n16015), .A(n16014), .B(n16013), .ZN(
        n16018) );
  XNOR2_X1 U17044 ( .A(n16601), .B(n17347), .ZN(n16021) );
  INV_X1 U17045 ( .A(n404), .ZN(n16019) );
  XNOR2_X1 U17046 ( .A(n16021), .B(n16020), .ZN(n16024) );
  XNOR2_X1 U17047 ( .A(n17410), .B(n17348), .ZN(n16022) );
  XNOR2_X1 U17048 ( .A(n19860), .B(n16022), .ZN(n16023) );
  XNOR2_X1 U17049 ( .A(n16023), .B(n16024), .ZN(n16025) );
  NAND2_X1 U17050 ( .A1(n17898), .A2(n16025), .ZN(n17895) );
  INV_X1 U17051 ( .A(n16025), .ZN(n17069) );
  XNOR2_X1 U17052 ( .A(n17339), .B(n17426), .ZN(n16303) );
  XNOR2_X1 U17053 ( .A(n16695), .B(n18863), .ZN(n16026) );
  XNOR2_X1 U17054 ( .A(n16303), .B(n16026), .ZN(n16029) );
  XNOR2_X1 U17055 ( .A(n16406), .B(n20192), .ZN(n16953) );
  XNOR2_X1 U17056 ( .A(n20269), .B(n16584), .ZN(n16028) );
  NAND2_X1 U17059 ( .A1(n17895), .A2(n16783), .ZN(n16043) );
  XNOR2_X1 U17060 ( .A(n16928), .B(n16587), .ZN(n16200) );
  XNOR2_X1 U17061 ( .A(n16200), .B(n16711), .ZN(n17371) );
  INV_X1 U17062 ( .A(n16030), .ZN(n19422) );
  XNOR2_X1 U17063 ( .A(n16975), .B(n19422), .ZN(n16031) );
  XNOR2_X1 U17064 ( .A(n16031), .B(n16926), .ZN(n16032) );
  XNOR2_X1 U17065 ( .A(n16931), .B(n16861), .ZN(n16588) );
  XNOR2_X1 U17066 ( .A(n16032), .B(n16588), .ZN(n16033) );
  XNOR2_X1 U17067 ( .A(n17295), .B(n19720), .ZN(n16619) );
  XNOR2_X1 U17068 ( .A(n16945), .B(n16283), .ZN(n16034) );
  XNOR2_X1 U17069 ( .A(n16619), .B(n16034), .ZN(n16038) );
  XNOR2_X1 U17070 ( .A(n16614), .B(n17330), .ZN(n16196) );
  XNOR2_X1 U17071 ( .A(n20126), .B(n304), .ZN(n16036) );
  XNOR2_X1 U17072 ( .A(n16196), .B(n16036), .ZN(n16037) );
  XNOR2_X1 U17073 ( .A(n16038), .B(n16037), .ZN(n17892) );
  MUX2_X1 U17074 ( .A(n19910), .B(n17892), .S(n17896), .Z(n16042) );
  XNOR2_X1 U17075 ( .A(n16278), .B(n16487), .ZN(n16039) );
  XNOR2_X1 U17076 ( .A(n17357), .B(n16039), .ZN(n16041) );
  XNOR2_X1 U17077 ( .A(n17359), .B(n16429), .ZN(n16937) );
  XNOR2_X1 U17078 ( .A(n16936), .B(n16707), .ZN(n16596) );
  XNOR2_X1 U17079 ( .A(n19863), .B(n16596), .ZN(n16040) );
  XNOR2_X1 U17080 ( .A(n16769), .B(n16906), .ZN(n16049) );
  XNOR2_X1 U17081 ( .A(n17099), .B(n17014), .ZN(n16047) );
  XNOR2_X1 U17082 ( .A(n16047), .B(n16046), .ZN(n16048) );
  INV_X1 U17084 ( .A(n17666), .ZN(n17668) );
  NOR2_X1 U17085 ( .A1(n16052), .A2(n16051), .ZN(n16053) );
  XNOR2_X1 U17086 ( .A(n17424), .B(n16053), .ZN(n16056) );
  XNOR2_X1 U17087 ( .A(n17109), .B(n16336), .ZN(n16140) );
  XNOR2_X1 U17088 ( .A(n16054), .B(n16140), .ZN(n16055) );
  XNOR2_X1 U17089 ( .A(n19882), .B(n955), .ZN(n16058) );
  XNOR2_X1 U17090 ( .A(n19705), .B(n620), .ZN(n16057) );
  XNOR2_X1 U17091 ( .A(n16058), .B(n16057), .ZN(n16061) );
  INV_X1 U17092 ( .A(n17444), .ZN(n16059) );
  XNOR2_X1 U17093 ( .A(n17124), .B(n16059), .ZN(n16749) );
  XNOR2_X1 U17094 ( .A(n16746), .B(n16240), .ZN(n16878) );
  XNOR2_X1 U17095 ( .A(n16749), .B(n16878), .ZN(n16060) );
  XNOR2_X1 U17096 ( .A(n17399), .B(n17119), .ZN(n16065) );
  XNOR2_X1 U17097 ( .A(n16227), .B(n16900), .ZN(n16063) );
  XNOR2_X1 U17098 ( .A(n16853), .B(n294), .ZN(n16062) );
  XNOR2_X1 U17099 ( .A(n16063), .B(n16062), .ZN(n16064) );
  OAI22_X1 U17100 ( .A1(n17668), .A2(n17876), .B1(n17879), .B2(n19832), .ZN(
        n16070) );
  XNOR2_X1 U17101 ( .A(n16329), .B(n16566), .ZN(n16066) );
  XNOR2_X1 U17102 ( .A(n17431), .B(n16066), .ZN(n16069) );
  INV_X1 U17103 ( .A(n18439), .ZN(n18443) );
  XNOR2_X1 U17104 ( .A(n16568), .B(n18443), .ZN(n16067) );
  NAND2_X1 U17106 ( .A1(n16070), .A2(n17881), .ZN(n16076) );
  XNOR2_X1 U17107 ( .A(n16071), .B(n16871), .ZN(n16074) );
  XNOR2_X1 U17108 ( .A(n16821), .B(n17170), .ZN(n16072) );
  XNOR2_X1 U17109 ( .A(n20219), .B(n16072), .ZN(n16073) );
  NOR2_X1 U17110 ( .A1(n17666), .A2(n17878), .ZN(n17882) );
  AOI22_X1 U17112 ( .A1(n17882), .A2(n20217), .B1(n19930), .B2(n19832), .ZN(
        n16075) );
  XNOR2_X1 U17114 ( .A(n16853), .B(n17298), .ZN(n16719) );
  XNOR2_X1 U17115 ( .A(n16367), .B(n18433), .ZN(n16077) );
  XNOR2_X1 U17116 ( .A(n16719), .B(n16077), .ZN(n16080) );
  XNOR2_X1 U17117 ( .A(n16078), .B(n16854), .ZN(n16617) );
  XNOR2_X1 U17118 ( .A(n16617), .B(n17120), .ZN(n16079) );
  XNOR2_X1 U17119 ( .A(n16080), .B(n16079), .ZN(n17886) );
  INV_X1 U17120 ( .A(n16982), .ZN(n16219) );
  XNOR2_X1 U17121 ( .A(n16219), .B(n19909), .ZN(n17107) );
  XNOR2_X1 U17122 ( .A(n17107), .B(n16083), .ZN(n16087) );
  INV_X1 U17123 ( .A(n16373), .ZN(n16084) );
  XNOR2_X1 U17124 ( .A(n17270), .B(n19436), .ZN(n16085) );
  XNOR2_X1 U17125 ( .A(n16696), .B(n16085), .ZN(n16086) );
  XNOR2_X1 U17126 ( .A(n17280), .B(n18075), .ZN(n16088) );
  XNOR2_X1 U17127 ( .A(n16089), .B(n16088), .ZN(n16093) );
  XNOR2_X1 U17128 ( .A(n16973), .B(n16760), .ZN(n16090) );
  XNOR2_X1 U17129 ( .A(n16090), .B(n16091), .ZN(n16092) );
  NOR2_X1 U17130 ( .A1(n17886), .A2(n20185), .ZN(n16101) );
  XNOR2_X1 U17131 ( .A(n16094), .B(n16770), .ZN(n16096) );
  XNOR2_X1 U17132 ( .A(n16096), .B(n16828), .ZN(n16100) );
  XNOR2_X1 U17133 ( .A(n16097), .B(n17012), .ZN(n16098) );
  XNOR2_X1 U17134 ( .A(n16098), .B(n16691), .ZN(n16099) );
  XNOR2_X1 U17135 ( .A(n19900), .B(n17128), .ZN(n16117) );
  XNOR2_X1 U17136 ( .A(n16117), .B(n16102), .ZN(n16105) );
  XNOR2_X1 U17137 ( .A(n16359), .B(n19705), .ZN(n16702) );
  XNOR2_X1 U17138 ( .A(n17260), .B(n2349), .ZN(n16103) );
  XNOR2_X1 U17139 ( .A(n16702), .B(n16103), .ZN(n16104) );
  XNOR2_X1 U17140 ( .A(n16104), .B(n16105), .ZN(n16261) );
  XNOR2_X1 U17141 ( .A(n16821), .B(n17252), .ZN(n16705) );
  XNOR2_X1 U17142 ( .A(n16939), .B(n16741), .ZN(n16122) );
  XNOR2_X1 U17143 ( .A(n16705), .B(n16122), .ZN(n16109) );
  INV_X1 U17144 ( .A(n2151), .ZN(n18880) );
  XNOR2_X1 U17145 ( .A(n17253), .B(n18880), .ZN(n16106) );
  XNOR2_X1 U17146 ( .A(n16107), .B(n16106), .ZN(n16108) );
  NOR2_X1 U17147 ( .A1(n16261), .A2(n17890), .ZN(n16110) );
  NAND2_X1 U17148 ( .A1(n16110), .A2(n17891), .ZN(n16111) );
  OAI21_X1 U17149 ( .B1(n17600), .B2(n3825), .A(n16111), .ZN(n16114) );
  INV_X1 U17150 ( .A(n17600), .ZN(n16112) );
  INV_X1 U17151 ( .A(n17890), .ZN(n17663) );
  NOR2_X1 U17152 ( .A1(n16112), .A2(n17663), .ZN(n16113) );
  INV_X1 U17154 ( .A(n19170), .ZN(n18324) );
  NAND3_X1 U17155 ( .A1(n16115), .A2(n18324), .A3(n20394), .ZN(n16164) );
  XNOR2_X1 U17156 ( .A(n16292), .B(n17127), .ZN(n16116) );
  XNOR2_X1 U17157 ( .A(n16116), .B(n16240), .ZN(n16118) );
  XNOR2_X1 U17158 ( .A(n16118), .B(n16117), .ZN(n16121) );
  XNOR2_X1 U17160 ( .A(n16880), .B(n16119), .ZN(n16120) );
  XNOR2_X1 U17161 ( .A(n17002), .B(n17535), .ZN(n16123) );
  XNOR2_X1 U17162 ( .A(n16122), .B(n16123), .ZN(n16125) );
  XNOR2_X1 U17163 ( .A(n17360), .B(n16872), .ZN(n16182) );
  XNOR2_X1 U17164 ( .A(n16871), .B(n16182), .ZN(n16124) );
  NAND2_X1 U17165 ( .A1(n20264), .A2(n17840), .ZN(n16139) );
  XNOR2_X1 U17166 ( .A(n17349), .B(n1996), .ZN(n16130) );
  INV_X1 U17167 ( .A(n16126), .ZN(n16127) );
  XNOR2_X1 U17168 ( .A(n17099), .B(n16770), .ZN(n16131) );
  NAND2_X1 U17169 ( .A1(n16139), .A2(n17063), .ZN(n17201) );
  INV_X1 U17170 ( .A(n17840), .ZN(n16153) );
  XNOR2_X1 U17171 ( .A(n16224), .B(n17328), .ZN(n16946) );
  XNOR2_X1 U17172 ( .A(n16902), .B(n16946), .ZN(n16138) );
  XNOR2_X1 U17173 ( .A(n16963), .B(n16134), .ZN(n16136) );
  XNOR2_X1 U17174 ( .A(n16854), .B(n18203), .ZN(n16135) );
  XNOR2_X1 U17175 ( .A(n16136), .B(n16135), .ZN(n16137) );
  NAND2_X1 U17176 ( .A1(n16139), .A2(n16731), .ZN(n16152) );
  XNOR2_X1 U17177 ( .A(n17340), .B(n16407), .ZN(n16301) );
  XNOR2_X1 U17178 ( .A(n16301), .B(n16140), .ZN(n16144) );
  XNOR2_X1 U17179 ( .A(n19674), .B(n18420), .ZN(n16141) );
  XNOR2_X1 U17180 ( .A(n16142), .B(n16141), .ZN(n16143) );
  INV_X1 U17182 ( .A(n16973), .ZN(n16929) );
  XNOR2_X1 U17183 ( .A(n16145), .B(n16929), .ZN(n16147) );
  XNOR2_X1 U17184 ( .A(n16147), .B(n16146), .ZN(n16150) );
  XNOR2_X1 U17185 ( .A(n16568), .B(n16760), .ZN(n16148) );
  XNOR2_X1 U17186 ( .A(n16329), .B(n16148), .ZN(n16149) );
  NAND2_X1 U17187 ( .A1(n3826), .A2(n20423), .ZN(n16151) );
  NAND2_X1 U17188 ( .A1(n18157), .A2(n16155), .ZN(n18156) );
  NAND2_X1 U17189 ( .A1(n16154), .A2(n993), .ZN(n16163) );
  INV_X1 U17190 ( .A(n16155), .ZN(n18317) );
  NOR2_X1 U17191 ( .A1(n18317), .A2(n20460), .ZN(n16159) );
  INV_X1 U17195 ( .A(n16159), .ZN(n16160) );
  NAND4_X1 U17196 ( .A1(n18156), .A2(n16160), .A3(n2368), .A4(n19170), .ZN(
        n16161) );
  NAND4_X1 U17197 ( .A1(n16164), .A2(n16163), .A3(n20384), .A4(n16161), .ZN(
        Ciphertext[144]) );
  INV_X1 U17199 ( .A(n17501), .ZN(n16794) );
  NAND3_X1 U17201 ( .A1(n16794), .A2(n19815), .A3(n19924), .ZN(n16168) );
  NAND2_X1 U17202 ( .A1(n16794), .A2(n15485), .ZN(n16167) );
  NOR2_X1 U17205 ( .A1(n16634), .A2(n3573), .ZN(n16174) );
  OAI21_X1 U17206 ( .B1(n17508), .B2(n17507), .A(n16172), .ZN(n16173) );
  OAI21_X2 U17207 ( .B1(n16632), .B2(n16174), .A(n16173), .ZN(n18498) );
  XNOR2_X1 U17208 ( .A(n16880), .B(n17124), .ZN(n16176) );
  XNOR2_X1 U17209 ( .A(n16176), .B(n16175), .ZN(n16180) );
  XNOR2_X1 U17210 ( .A(n955), .B(n17377), .ZN(n16178) );
  XNOR2_X1 U17211 ( .A(n19799), .B(n19027), .ZN(n16177) );
  XNOR2_X1 U17212 ( .A(n16178), .B(n16177), .ZN(n16179) );
  XNOR2_X1 U17213 ( .A(n16180), .B(n16179), .ZN(n17565) );
  INV_X1 U17214 ( .A(n17565), .ZN(n17562) );
  XNOR2_X1 U17215 ( .A(n16742), .B(n16181), .ZN(n16183) );
  XNOR2_X1 U17216 ( .A(n16183), .B(n16182), .ZN(n16187) );
  XNOR2_X1 U17217 ( .A(n17359), .B(n2455), .ZN(n16184) );
  XNOR2_X1 U17218 ( .A(n16185), .B(n16184), .ZN(n16186) );
  XNOR2_X1 U17219 ( .A(n16187), .B(n16186), .ZN(n16320) );
  INV_X1 U17220 ( .A(n16320), .ZN(n18535) );
  XNOR2_X1 U17221 ( .A(n17104), .B(n17406), .ZN(n16190) );
  XNOR2_X1 U17222 ( .A(n16188), .B(n17348), .ZN(n16189) );
  XNOR2_X1 U17223 ( .A(n16190), .B(n16189), .ZN(n16194) );
  XNOR2_X1 U17224 ( .A(n16601), .B(n17014), .ZN(n16192) );
  XNOR2_X1 U17225 ( .A(n19836), .B(n621), .ZN(n16191) );
  XNOR2_X1 U17226 ( .A(n16191), .B(n16192), .ZN(n16193) );
  XNOR2_X1 U17227 ( .A(n16194), .B(n16193), .ZN(n16321) );
  INV_X1 U17228 ( .A(n16321), .ZN(n16790) );
  XNOR2_X1 U17229 ( .A(n16225), .B(n16412), .ZN(n16195) );
  XNOR2_X1 U17230 ( .A(n16284), .B(n16195), .ZN(n16199) );
  XNOR2_X1 U17231 ( .A(n16947), .B(n2454), .ZN(n16197) );
  XNOR2_X1 U17232 ( .A(n16197), .B(n16196), .ZN(n16198) );
  XNOR2_X1 U17233 ( .A(n16199), .B(n16198), .ZN(n17470) );
  XNOR2_X1 U17234 ( .A(n16200), .B(n16288), .ZN(n16204) );
  XNOR2_X1 U17235 ( .A(n16886), .B(n880), .ZN(n16202) );
  XNOR2_X1 U17236 ( .A(n16932), .B(n17089), .ZN(n16201) );
  XNOR2_X1 U17237 ( .A(n16202), .B(n16201), .ZN(n16203) );
  OAI22_X1 U17238 ( .A1(n18535), .A2(n16790), .B1(n17470), .B2(n18534), .ZN(
        n17163) );
  XNOR2_X1 U17240 ( .A(n902), .B(n17338), .ZN(n17034) );
  XNOR2_X1 U17241 ( .A(n16301), .B(n17034), .ZN(n16208) );
  XNOR2_X1 U17242 ( .A(n20192), .B(n911), .ZN(n16206) );
  XNOR2_X1 U17243 ( .A(n16300), .B(n2087), .ZN(n16205) );
  XNOR2_X1 U17244 ( .A(n16206), .B(n16205), .ZN(n16207) );
  INV_X1 U17245 ( .A(n17470), .ZN(n16209) );
  OAI21_X1 U17246 ( .B1(n17564), .B2(n20432), .A(n16209), .ZN(n16210) );
  NOR2_X1 U17247 ( .A1(n18500), .A2(n18485), .ZN(n17912) );
  XNOR2_X1 U17248 ( .A(n16927), .B(n2192), .ZN(n16213) );
  XNOR2_X1 U17249 ( .A(n16213), .B(n17276), .ZN(n16215) );
  XNOR2_X1 U17250 ( .A(n16215), .B(n16214), .ZN(n16218) );
  XNOR2_X1 U17251 ( .A(n16970), .B(n879), .ZN(n16216) );
  XNOR2_X1 U17252 ( .A(n16329), .B(n16216), .ZN(n16217) );
  XNOR2_X1 U17253 ( .A(n17335), .B(n17426), .ZN(n16979) );
  XNOR2_X1 U17254 ( .A(n16219), .B(n19928), .ZN(n16952) );
  XNOR2_X1 U17255 ( .A(n16979), .B(n16952), .ZN(n16223) );
  XNOR2_X1 U17256 ( .A(n16335), .B(n19018), .ZN(n16221) );
  XNOR2_X1 U17257 ( .A(n911), .B(n897), .ZN(n16220) );
  XNOR2_X1 U17258 ( .A(n16221), .B(n16220), .ZN(n16222) );
  XNOR2_X1 U17259 ( .A(n16224), .B(n16283), .ZN(n16962) );
  XNOR2_X1 U17260 ( .A(n16225), .B(n16960), .ZN(n16226) );
  XNOR2_X1 U17261 ( .A(n16962), .B(n16226), .ZN(n16230) );
  XNOR2_X1 U17262 ( .A(n17298), .B(n16227), .ZN(n16341) );
  XNOR2_X1 U17263 ( .A(n16944), .B(n17791), .ZN(n16228) );
  XNOR2_X1 U17264 ( .A(n16341), .B(n16228), .ZN(n16229) );
  XNOR2_X1 U17266 ( .A(n16988), .B(n16691), .ZN(n16231) );
  XNOR2_X1 U17267 ( .A(n16769), .B(n16231), .ZN(n16235) );
  INV_X1 U17268 ( .A(n20682), .ZN(n18631) );
  XNOR2_X1 U17269 ( .A(n17410), .B(n18631), .ZN(n16233) );
  XNOR2_X1 U17270 ( .A(n16233), .B(n16232), .ZN(n16234) );
  XNOR2_X1 U17271 ( .A(n16742), .B(n16939), .ZN(n17142) );
  XNOR2_X1 U17272 ( .A(n17252), .B(n16236), .ZN(n16353) );
  XNOR2_X1 U17273 ( .A(n17142), .B(n16353), .ZN(n16239) );
  INV_X1 U17274 ( .A(n2423), .ZN(n18506) );
  XNOR2_X1 U17275 ( .A(n17355), .B(n18506), .ZN(n16237) );
  XNOR2_X1 U17276 ( .A(n17418), .B(n16237), .ZN(n16238) );
  XNOR2_X1 U17277 ( .A(n16238), .B(n16239), .ZN(n16447) );
  INV_X1 U17278 ( .A(n16447), .ZN(n17495) );
  XNOR2_X1 U17279 ( .A(n17443), .B(n16240), .ZN(n16241) );
  XNOR2_X1 U17280 ( .A(n16749), .B(n16241), .ZN(n16245) );
  INV_X1 U17281 ( .A(n16242), .ZN(n19280) );
  XNOR2_X1 U17282 ( .A(n19743), .B(n19280), .ZN(n16243) );
  XNOR2_X1 U17283 ( .A(n16998), .B(n16243), .ZN(n16244) );
  XNOR2_X1 U17284 ( .A(n16245), .B(n16244), .ZN(n17491) );
  AND2_X1 U17285 ( .A1(n17495), .A2(n17491), .ZN(n16802) );
  NAND2_X1 U17286 ( .A1(n16802), .A2(n16801), .ZN(n16246) );
  OAI21_X1 U17287 ( .B1(n16247), .B2(n16801), .A(n16246), .ZN(n16249) );
  NAND2_X1 U17288 ( .A1(n16447), .A2(n17493), .ZN(n16800) );
  NOR2_X1 U17289 ( .A1(n16800), .A2(n17488), .ZN(n16248) );
  NAND2_X1 U17291 ( .A1(n17912), .A2(n19729), .ZN(n16257) );
  INV_X1 U17293 ( .A(n20135), .ZN(n17213) );
  NAND2_X1 U17294 ( .A1(n16465), .A2(n17211), .ZN(n16254) );
  NAND2_X1 U17295 ( .A1(n16465), .A2(n20135), .ZN(n16253) );
  INV_X1 U17296 ( .A(n17210), .ZN(n16658) );
  NAND3_X1 U17297 ( .A1(n16254), .A2(n16253), .A3(n16658), .ZN(n16255) );
  INV_X1 U17298 ( .A(n18495), .ZN(n18496) );
  NAND3_X1 U17299 ( .A1(n18496), .A2(n893), .A3(n19816), .ZN(n16256) );
  INV_X1 U17300 ( .A(n2023), .ZN(n16258) );
  XNOR2_X1 U17301 ( .A(n16259), .B(n16258), .ZN(Ciphertext[27]) );
  NAND2_X1 U17302 ( .A1(n17891), .A2(n20185), .ZN(n16260) );
  INV_X1 U17303 ( .A(n16261), .ZN(n17602) );
  OAI21_X1 U17305 ( .B1(n16262), .B2(n20239), .A(n17822), .ZN(n16264) );
  INV_X1 U17306 ( .A(n16263), .ZN(n17824) );
  NAND3_X1 U17307 ( .A1(n16262), .A2(n17079), .A3(n17823), .ZN(n16265) );
  INV_X1 U17308 ( .A(n19209), .ZN(n19202) );
  INV_X1 U17309 ( .A(n17898), .ZN(n17182) );
  AND2_X1 U17310 ( .A1(n17896), .A2(n17181), .ZN(n16266) );
  OAI21_X1 U17311 ( .B1(n17182), .B2(n19707), .A(n16266), .ZN(n16268) );
  NOR2_X1 U17312 ( .A1(n17892), .A2(n19910), .ZN(n17183) );
  INV_X1 U17313 ( .A(n16781), .ZN(n17897) );
  NAND2_X1 U17314 ( .A1(n17183), .A2(n17897), .ZN(n16267) );
  XNOR2_X1 U17315 ( .A(n16269), .B(n17104), .ZN(n16271) );
  XNOR2_X1 U17316 ( .A(n17406), .B(n17410), .ZN(n16270) );
  XNOR2_X1 U17317 ( .A(n16270), .B(n16271), .ZN(n16275) );
  XNOR2_X1 U17318 ( .A(n16992), .B(n17347), .ZN(n16273) );
  XNOR2_X1 U17319 ( .A(n19836), .B(n347), .ZN(n16272) );
  XNOR2_X1 U17320 ( .A(n16272), .B(n16273), .ZN(n16274) );
  XNOR2_X2 U17321 ( .A(n16275), .B(n16274), .ZN(n19402) );
  XNOR2_X1 U17322 ( .A(n17002), .B(n16872), .ZN(n16277) );
  XNOR2_X1 U17323 ( .A(n16276), .B(n16277), .ZN(n16282) );
  XNOR2_X1 U17324 ( .A(n864), .B(n16278), .ZN(n16280) );
  XNOR2_X1 U17325 ( .A(n16873), .B(n2383), .ZN(n16279) );
  XNOR2_X1 U17326 ( .A(n16280), .B(n16279), .ZN(n16281) );
  XNOR2_X1 U17327 ( .A(n16282), .B(n16281), .ZN(n17650) );
  XNOR2_X1 U17328 ( .A(n16412), .B(n16283), .ZN(n17400) );
  XNOR2_X1 U17329 ( .A(n16963), .B(n18887), .ZN(n16285) );
  XNOR2_X1 U17330 ( .A(n16975), .B(n16886), .ZN(n17435) );
  XNOR2_X1 U17331 ( .A(n16330), .B(n19222), .ZN(n16286) );
  XNOR2_X1 U17332 ( .A(n17435), .B(n16286), .ZN(n16290) );
  XNOR2_X1 U17333 ( .A(n17133), .B(n16711), .ZN(n16287) );
  XNOR2_X1 U17334 ( .A(n16288), .B(n16287), .ZN(n16289) );
  XNOR2_X1 U17335 ( .A(n16289), .B(n16290), .ZN(n17853) );
  NAND2_X1 U17336 ( .A1(n16306), .A2(n17853), .ZN(n16291) );
  XNOR2_X1 U17337 ( .A(n16293), .B(n19954), .ZN(n17125) );
  XNOR2_X1 U17338 ( .A(n16294), .B(n17125), .ZN(n16299) );
  XNOR2_X1 U17340 ( .A(n16297), .B(n16296), .ZN(n16298) );
  INV_X1 U17342 ( .A(n17853), .ZN(n17606) );
  XNOR2_X1 U17343 ( .A(n16507), .B(n16300), .ZN(n17108) );
  XNOR2_X1 U17344 ( .A(n17108), .B(n16301), .ZN(n16305) );
  XNOR2_X1 U17345 ( .A(n16893), .B(n2317), .ZN(n16302) );
  XNOR2_X1 U17346 ( .A(n16303), .B(n16302), .ZN(n16304) );
  XNOR2_X2 U17347 ( .A(n16305), .B(n16304), .ZN(n19404) );
  OAI21_X1 U17348 ( .B1(n17606), .B2(n19404), .A(n16306), .ZN(n16307) );
  MUX2_X1 U17349 ( .A(n3345), .B(n19930), .S(n17876), .Z(n16312) );
  NOR2_X1 U17350 ( .A1(n3345), .A2(n17879), .ZN(n16310) );
  NOR2_X1 U17351 ( .A1(n17881), .A2(n16308), .ZN(n16309) );
  MUX2_X1 U17352 ( .A(n16310), .B(n16309), .S(n19930), .Z(n16311) );
  AOI21_X2 U17353 ( .B1(n16308), .B2(n16312), .A(n16311), .ZN(n19210) );
  MUX2_X1 U17355 ( .A(n19973), .B(n20507), .S(n17868), .Z(n16317) );
  NAND2_X1 U17356 ( .A1(n20506), .A2(n17873), .ZN(n16315) );
  MUX2_X1 U17357 ( .A(n19190), .B(n19210), .S(n19842), .Z(n16318) );
  NAND2_X1 U17358 ( .A1(n16318), .A2(n19189), .ZN(n16319) );
  AND2_X1 U17359 ( .A1(n17564), .A2(n17470), .ZN(n16789) );
  INV_X1 U17360 ( .A(n18534), .ZN(n17468) );
  OAI21_X1 U17361 ( .B1(n17468), .B2(n17564), .A(n17471), .ZN(n16325) );
  NOR2_X1 U17362 ( .A1(n18539), .A2(n17471), .ZN(n16323) );
  NOR2_X1 U17363 ( .A1(n17564), .A2(n17471), .ZN(n16322) );
  AOI22_X1 U17364 ( .A1(n16323), .A2(n17565), .B1(n18539), .B2(n16322), .ZN(
        n16324) );
  OAI21_X2 U17365 ( .B1(n16325), .B2(n16789), .A(n16324), .ZN(n18568) );
  INV_X1 U17366 ( .A(n18568), .ZN(n16446) );
  INV_X1 U17367 ( .A(n17276), .ZN(n16326) );
  XNOR2_X1 U17368 ( .A(n19894), .B(n16326), .ZN(n16328) );
  XNOR2_X1 U17369 ( .A(n16931), .B(n2395), .ZN(n16327) );
  XNOR2_X1 U17370 ( .A(n16328), .B(n16327), .ZN(n16333) );
  XNOR2_X1 U17371 ( .A(n16329), .B(n16971), .ZN(n16885) );
  XNOR2_X1 U17372 ( .A(n16330), .B(n16760), .ZN(n16331) );
  INV_X1 U17373 ( .A(n16954), .ZN(n16334) );
  XNOR2_X1 U17374 ( .A(n16334), .B(n16335), .ZN(n17268) );
  XNOR2_X1 U17375 ( .A(n17268), .B(n16756), .ZN(n16340) );
  XNOR2_X1 U17376 ( .A(n17111), .B(n897), .ZN(n16338) );
  XNOR2_X1 U17377 ( .A(n16893), .B(n18801), .ZN(n16337) );
  XNOR2_X1 U17378 ( .A(n16338), .B(n16337), .ZN(n16339) );
  NOR2_X1 U17379 ( .A1(n20488), .A2(n18114), .ZN(n18116) );
  XNOR2_X1 U17380 ( .A(n16342), .B(n16341), .ZN(n16346) );
  XNOR2_X1 U17381 ( .A(n17116), .B(n17295), .ZN(n16344) );
  XNOR2_X1 U17382 ( .A(n16965), .B(n18065), .ZN(n16343) );
  XNOR2_X1 U17383 ( .A(n16344), .B(n16343), .ZN(n16345) );
  XNOR2_X1 U17384 ( .A(n16346), .B(n16345), .ZN(n17458) );
  INV_X1 U17385 ( .A(n16347), .ZN(n16599) );
  XNOR2_X1 U17386 ( .A(n16599), .B(n16691), .ZN(n16348) );
  XNOR2_X1 U17387 ( .A(n16348), .B(n16906), .ZN(n16352) );
  XNOR2_X1 U17388 ( .A(n16770), .B(n16987), .ZN(n16350) );
  XNOR2_X1 U17389 ( .A(n17098), .B(n18517), .ZN(n16349) );
  XNOR2_X1 U17390 ( .A(n16350), .B(n16349), .ZN(n16351) );
  OAI21_X1 U17391 ( .B1(n18116), .B2(n17559), .A(n18111), .ZN(n16364) );
  XNOR2_X1 U17393 ( .A(n16553), .B(n16353), .ZN(n16357) );
  XNOR2_X1 U17394 ( .A(n16936), .B(n2413), .ZN(n16354) );
  XNOR2_X1 U17395 ( .A(n16355), .B(n16354), .ZN(n16356) );
  NOR2_X1 U17397 ( .A1(n20488), .A2(n17458), .ZN(n16363) );
  XNOR2_X1 U17398 ( .A(n20477), .B(n16747), .ZN(n16847) );
  XNOR2_X1 U17399 ( .A(n19743), .B(n16914), .ZN(n17258) );
  XNOR2_X1 U17400 ( .A(n17258), .B(n16847), .ZN(n16362) );
  XNOR2_X1 U17401 ( .A(n16996), .B(n875), .ZN(n16360) );
  XNOR2_X1 U17402 ( .A(n16878), .B(n16360), .ZN(n16361) );
  INV_X1 U17403 ( .A(n18556), .ZN(n18199) );
  XNOR2_X1 U17404 ( .A(n16365), .B(n16619), .ZN(n16371) );
  XNOR2_X1 U17405 ( .A(n16615), .B(n16961), .ZN(n16369) );
  XNOR2_X1 U17406 ( .A(n16367), .B(n16366), .ZN(n16368) );
  XNOR2_X1 U17407 ( .A(n16369), .B(n16368), .ZN(n16370) );
  XNOR2_X1 U17408 ( .A(n16371), .B(n16370), .ZN(n17954) );
  XNOR2_X1 U17411 ( .A(n16373), .B(n16374), .ZN(n16834) );
  XNOR2_X1 U17412 ( .A(n17337), .B(n16834), .ZN(n16378) );
  XNOR2_X1 U17413 ( .A(n16954), .B(n16695), .ZN(n16376) );
  XNOR2_X1 U17414 ( .A(n16755), .B(n2410), .ZN(n16375) );
  XNOR2_X1 U17415 ( .A(n16376), .B(n16375), .ZN(n16377) );
  XNOR2_X1 U17416 ( .A(n16378), .B(n16377), .ZN(n17957) );
  OR2_X1 U17417 ( .A1(n17954), .A2(n17957), .ZN(n17552) );
  INV_X1 U17418 ( .A(n17552), .ZN(n16389) );
  XNOR2_X1 U17419 ( .A(n16969), .B(n2375), .ZN(n16379) );
  XNOR2_X1 U17420 ( .A(n16380), .B(n16379), .ZN(n16382) );
  XNOR2_X1 U17421 ( .A(n16588), .B(n16713), .ZN(n16381) );
  XNOR2_X1 U17422 ( .A(n16381), .B(n16382), .ZN(n16805) );
  AND2_X1 U17423 ( .A1(n18105), .A2(n17954), .ZN(n16388) );
  XNOR2_X1 U17425 ( .A(n16385), .B(n16384), .ZN(n16387) );
  XNOR2_X1 U17426 ( .A(n16386), .B(n17291), .ZN(n16693) );
  OAI21_X1 U17427 ( .B1(n16389), .B2(n16388), .A(n18103), .ZN(n16405) );
  INV_X1 U17428 ( .A(n18103), .ZN(n16404) );
  XNOR2_X1 U17429 ( .A(n16510), .B(n16608), .ZN(n16391) );
  XNOR2_X1 U17430 ( .A(n16391), .B(n16390), .ZN(n16395) );
  XNOR2_X1 U17434 ( .A(n16596), .B(n16396), .ZN(n16400) );
  XNOR2_X1 U17435 ( .A(n15935), .B(n17358), .ZN(n16398) );
  XNOR2_X1 U17436 ( .A(n19889), .B(n295), .ZN(n16397) );
  XNOR2_X1 U17437 ( .A(n16398), .B(n16397), .ZN(n16399) );
  XNOR2_X1 U17438 ( .A(n16399), .B(n16400), .ZN(n17955) );
  NOR2_X1 U17440 ( .A1(n17956), .A2(n18107), .ZN(n16403) );
  AND2_X1 U17441 ( .A1(n18107), .A2(n17957), .ZN(n16402) );
  INV_X1 U17442 ( .A(n17954), .ZN(n16401) );
  NAND2_X1 U17443 ( .A1(n18199), .A2(n18559), .ZN(n18201) );
  NAND2_X1 U17444 ( .A1(n18199), .A2(n18568), .ZN(n16453) );
  XNOR2_X1 U17445 ( .A(n20102), .B(n16406), .ZN(n17423) );
  XNOR2_X1 U17446 ( .A(n17423), .B(n17036), .ZN(n16411) );
  XNOR2_X1 U17447 ( .A(n16981), .B(n17269), .ZN(n16409) );
  XNOR2_X1 U17448 ( .A(n16836), .B(n18366), .ZN(n16408) );
  XNOR2_X1 U17449 ( .A(n16409), .B(n16408), .ZN(n16410) );
  INV_X1 U17450 ( .A(n18097), .ZN(n18094) );
  XNOR2_X1 U17451 ( .A(n17019), .B(n16527), .ZN(n16416) );
  XNOR2_X1 U17452 ( .A(n20104), .B(n16961), .ZN(n16414) );
  XNOR2_X1 U17453 ( .A(n16412), .B(n2307), .ZN(n16413) );
  XNOR2_X1 U17454 ( .A(n16414), .B(n16413), .ZN(n16415) );
  XNOR2_X1 U17455 ( .A(n16416), .B(n16415), .ZN(n18096) );
  XNOR2_X1 U17456 ( .A(n17406), .B(n18304), .ZN(n16417) );
  XNOR2_X1 U17457 ( .A(n16417), .B(n19820), .ZN(n16419) );
  XNOR2_X1 U17458 ( .A(n17288), .B(n17411), .ZN(n16421) );
  XNOR2_X1 U17459 ( .A(n16421), .B(n16420), .ZN(n16519) );
  XNOR2_X1 U17461 ( .A(n16969), .B(n16926), .ZN(n16423) );
  XNOR2_X1 U17462 ( .A(n17026), .B(n16423), .ZN(n16428) );
  XNOR2_X1 U17463 ( .A(n17275), .B(n16886), .ZN(n16426) );
  XNOR2_X1 U17464 ( .A(n17279), .B(n16424), .ZN(n16425) );
  XOR2_X1 U17465 ( .A(n16426), .B(n16425), .Z(n16427) );
  NOR2_X1 U17466 ( .A1(n18093), .A2(n20109), .ZN(n16434) );
  XNOR2_X1 U17467 ( .A(n16429), .B(n16872), .ZN(n17420) );
  XNOR2_X1 U17468 ( .A(n16534), .B(n17420), .ZN(n16433) );
  XNOR2_X1 U17469 ( .A(n16554), .B(n16706), .ZN(n16431) );
  XNOR2_X1 U17470 ( .A(n17253), .B(n18208), .ZN(n16430) );
  XNOR2_X1 U17471 ( .A(n16431), .B(n16430), .ZN(n16432) );
  XNOR2_X1 U17472 ( .A(n16510), .B(n16562), .ZN(n16435) );
  XNOR2_X1 U17473 ( .A(n16514), .B(n16435), .ZN(n16439) );
  XNOR2_X1 U17474 ( .A(n16880), .B(n17260), .ZN(n16437) );
  XNOR2_X1 U17475 ( .A(n17378), .B(n2221), .ZN(n16436) );
  XNOR2_X1 U17476 ( .A(n16437), .B(n16436), .ZN(n16438) );
  XNOR2_X1 U17477 ( .A(n16439), .B(n16438), .ZN(n18101) );
  AND2_X1 U17478 ( .A1(n18101), .A2(n160), .ZN(n18099) );
  MUX2_X1 U17479 ( .A(n17164), .B(n18099), .S(n19774), .Z(n16440) );
  NOR2_X1 U17481 ( .A1(n19815), .A2(n19898), .ZN(n16444) );
  NAND2_X1 U17482 ( .A1(n19815), .A2(n16165), .ZN(n16445) );
  NAND2_X1 U17483 ( .A1(n18565), .A2(n18556), .ZN(n16452) );
  OR2_X1 U17484 ( .A1(n18567), .A2(n18199), .ZN(n17997) );
  NAND2_X1 U17485 ( .A1(n17495), .A2(n17493), .ZN(n16449) );
  OAI21_X1 U17486 ( .B1(n17491), .B2(n17155), .A(n17488), .ZN(n16448) );
  MUX2_X1 U17487 ( .A(n16449), .B(n16448), .S(n17489), .Z(n16451) );
  INV_X1 U17489 ( .A(n2208), .ZN(n16454) );
  NAND4_X1 U17490 ( .A1(n16453), .A2(n19775), .A3(n16454), .A4(n16452), .ZN(
        n16457) );
  NAND2_X1 U17491 ( .A1(n18568), .A2(n16454), .ZN(n16455) );
  OR2_X1 U17492 ( .A1(n18201), .A2(n16455), .ZN(n16456) );
  OAI211_X1 U17493 ( .C1(n16459), .C2(n2208), .A(n16457), .B(n16456), .ZN(
        n16458) );
  AOI21_X1 U17494 ( .B1(n16460), .B2(n16459), .A(n16458), .ZN(Ciphertext[44])
         );
  NAND2_X1 U17495 ( .A1(n17243), .A2(n17245), .ZN(n16462) );
  NOR2_X1 U17496 ( .A1(n17243), .A2(n17483), .ZN(n17482) );
  MUX2_X1 U17497 ( .A(n17482), .B(n16463), .S(n17480), .Z(n16464) );
  NAND2_X1 U17499 ( .A1(n16660), .A2(n17208), .ZN(n16466) );
  INV_X1 U17501 ( .A(n17511), .ZN(n17512) );
  MUX2_X1 U17502 ( .A(n17512), .B(n17508), .S(n19956), .Z(n16469) );
  INV_X1 U17503 ( .A(n20271), .ZN(n17224) );
  MUX2_X1 U17504 ( .A(n17224), .B(n17510), .S(n19700), .Z(n16468) );
  INV_X1 U17505 ( .A(n17493), .ZN(n17154) );
  NOR2_X1 U17506 ( .A1(n17154), .A2(n17489), .ZN(n16470) );
  OAI21_X1 U17507 ( .B1(n16470), .B2(n17490), .A(n17491), .ZN(n16473) );
  OAI21_X1 U17508 ( .B1(n17488), .B2(n17489), .A(n17493), .ZN(n16471) );
  INV_X1 U17509 ( .A(n19814), .ZN(n17502) );
  NAND3_X1 U17510 ( .A1(n16794), .A2(n19898), .A3(n17502), .ZN(n16478) );
  OAI21_X1 U17511 ( .B1(n19815), .B2(n19924), .A(n17505), .ZN(n16477) );
  NAND2_X1 U17512 ( .A1(n15485), .A2(n19924), .ZN(n16476) );
  NAND3_X1 U17513 ( .A1(n16478), .A2(n16477), .A3(n16476), .ZN(n16479) );
  AOI21_X1 U17515 ( .B1(n16666), .B2(n19386), .A(n19382), .ZN(n16483) );
  NOR2_X1 U17516 ( .A1(n20463), .A2(n16665), .ZN(n16481) );
  OAI21_X1 U17517 ( .B1(n16641), .B2(n16481), .A(n17220), .ZN(n16482) );
  INV_X1 U17518 ( .A(n20232), .ZN(n16484) );
  AOI22_X1 U17519 ( .A1(n18469), .A2(n18464), .B1(n20148), .B2(n16484), .ZN(
        n16485) );
  NAND2_X1 U17520 ( .A1(n16486), .A2(n16485), .ZN(n16489) );
  INV_X1 U17521 ( .A(n16487), .ZN(n16488) );
  XNOR2_X1 U17522 ( .A(n16489), .B(n16488), .ZN(Ciphertext[18]) );
  OAI21_X1 U17523 ( .B1(n16491), .B2(n18406), .A(n16490), .ZN(n16493) );
  NOR2_X1 U17524 ( .A1(n18425), .A2(n15529), .ZN(n18409) );
  INV_X1 U17525 ( .A(n18427), .ZN(n18407) );
  XNOR2_X1 U17526 ( .A(n16494), .B(n2035), .ZN(Ciphertext[15]) );
  NAND2_X1 U17528 ( .A1(n19402), .A2(n19401), .ZN(n16495) );
  NAND2_X1 U17529 ( .A1(n16497), .A2(n16495), .ZN(n16496) );
  INV_X1 U17530 ( .A(n16497), .ZN(n16499) );
  NOR2_X1 U17531 ( .A1(n19401), .A2(n19403), .ZN(n16498) );
  NAND2_X1 U17532 ( .A1(n16499), .A2(n16498), .ZN(n16500) );
  AND2_X2 U17533 ( .A1(n16501), .A2(n16500), .ZN(n19329) );
  NOR2_X1 U17535 ( .A1(n20217), .A2(n19930), .ZN(n16505) );
  MUX2_X1 U17536 ( .A(n16308), .B(n17881), .S(n17876), .Z(n16503) );
  INV_X1 U17537 ( .A(n16503), .ZN(n16504) );
  OAI21_X1 U17538 ( .B1(n20162), .B2(n16505), .A(n16504), .ZN(n17539) );
  NAND2_X1 U17539 ( .A1(n17539), .A2(n17610), .ZN(n19333) );
  NOR2_X1 U17540 ( .A1(n19749), .A2(n19333), .ZN(n16581) );
  XNOR2_X1 U17541 ( .A(n20269), .B(n16506), .ZN(n16509) );
  INV_X1 U17542 ( .A(n2448), .ZN(n18473) );
  XNOR2_X1 U17543 ( .A(n16507), .B(n18473), .ZN(n16508) );
  INV_X1 U17544 ( .A(n19363), .ZN(n17863) );
  XNOR2_X1 U17545 ( .A(n16510), .B(n17443), .ZN(n16512) );
  XNOR2_X1 U17546 ( .A(n16750), .B(n17804), .ZN(n16511) );
  XNOR2_X1 U17547 ( .A(n16512), .B(n16511), .ZN(n16516) );
  XNOR2_X1 U17548 ( .A(n16514), .B(n16513), .ZN(n16515) );
  XNOR2_X1 U17549 ( .A(n16515), .B(n16516), .ZN(n16679) );
  INV_X1 U17550 ( .A(n16679), .ZN(n19361) );
  XNOR2_X1 U17551 ( .A(n16992), .B(n632), .ZN(n16517) );
  MUX2_X1 U17552 ( .A(n17863), .B(n19361), .S(n17861), .Z(n16539) );
  XNOR2_X1 U17553 ( .A(n19849), .B(n16521), .ZN(n16526) );
  XNOR2_X1 U17554 ( .A(n17133), .B(n2446), .ZN(n16524) );
  XNOR2_X1 U17555 ( .A(n16523), .B(n16524), .ZN(n16525) );
  NOR2_X1 U17556 ( .A1(n19362), .A2(n19938), .ZN(n17591) );
  XNOR2_X1 U17557 ( .A(n16528), .B(n16527), .ZN(n16532) );
  XNOR2_X1 U17558 ( .A(n17294), .B(n16963), .ZN(n16530) );
  XNOR2_X1 U17559 ( .A(n17330), .B(n484), .ZN(n16529) );
  XNOR2_X1 U17560 ( .A(n16530), .B(n16529), .ZN(n16531) );
  XNOR2_X1 U17561 ( .A(n16532), .B(n16531), .ZN(n17672) );
  AND2_X1 U17562 ( .A1(n19363), .A2(n17672), .ZN(n17592) );
  NOR2_X1 U17563 ( .A1(n17591), .A2(n17592), .ZN(n16538) );
  XNOR2_X1 U17564 ( .A(n16938), .B(n2082), .ZN(n16533) );
  XNOR2_X1 U17565 ( .A(n16937), .B(n16533), .ZN(n16537) );
  XNOR2_X1 U17566 ( .A(n20267), .B(n17002), .ZN(n16535) );
  XNOR2_X1 U17567 ( .A(n16535), .B(n16534), .ZN(n16536) );
  MUX2_X2 U17569 ( .A(n16539), .B(n16538), .S(n19360), .Z(n19340) );
  INV_X1 U17570 ( .A(n19340), .ZN(n16544) );
  NOR2_X1 U17572 ( .A1(n16636), .A2(n19351), .ZN(n16543) );
  NAND2_X1 U17573 ( .A1(n16672), .A2(n19347), .ZN(n17231) );
  NAND2_X1 U17574 ( .A1(n17234), .A2(n17231), .ZN(n16541) );
  XNOR2_X1 U17577 ( .A(n17338), .B(n17060), .ZN(n16545) );
  XNOR2_X1 U17578 ( .A(n16696), .B(n16545), .ZN(n16548) );
  XNOR2_X1 U17579 ( .A(n16892), .B(n16546), .ZN(n16547) );
  XNOR2_X1 U17580 ( .A(n16548), .B(n16547), .ZN(n16642) );
  XNOR2_X1 U17581 ( .A(n16719), .B(n16898), .ZN(n16552) );
  XNOR2_X1 U17582 ( .A(n20104), .B(n17116), .ZN(n16550) );
  XNOR2_X1 U17583 ( .A(n16614), .B(n18338), .ZN(n16549) );
  XNOR2_X1 U17584 ( .A(n16550), .B(n16549), .ZN(n16551) );
  XNOR2_X2 U17585 ( .A(n16552), .B(n16551), .ZN(n19372) );
  XNOR2_X1 U17586 ( .A(n16705), .B(n16553), .ZN(n16559) );
  XNOR2_X1 U17587 ( .A(n16554), .B(n20450), .ZN(n16557) );
  XNOR2_X1 U17588 ( .A(n16593), .B(n302), .ZN(n16556) );
  XNOR2_X1 U17589 ( .A(n16557), .B(n16556), .ZN(n16558) );
  INV_X1 U17590 ( .A(n19371), .ZN(n19375) );
  OAI21_X1 U17591 ( .B1(n20436), .B2(n19372), .A(n19375), .ZN(n16657) );
  INV_X1 U17592 ( .A(Key[60]), .ZN(n16560) );
  XNOR2_X1 U17593 ( .A(n20478), .B(n16560), .ZN(n16561) );
  XNOR2_X1 U17594 ( .A(n16702), .B(n16561), .ZN(n16565) );
  XNOR2_X1 U17595 ( .A(n16562), .B(n16607), .ZN(n16563) );
  XNOR2_X1 U17596 ( .A(n16563), .B(n16882), .ZN(n16564) );
  XNOR2_X1 U17597 ( .A(n16565), .B(n16564), .ZN(n19374) );
  NAND2_X1 U17598 ( .A1(n19374), .A2(n19666), .ZN(n16579) );
  XNOR2_X1 U17599 ( .A(n19894), .B(n16566), .ZN(n16859) );
  XNOR2_X1 U17600 ( .A(n16859), .B(n16567), .ZN(n16572) );
  XNOR2_X1 U17601 ( .A(n16587), .B(n16568), .ZN(n16570) );
  XNOR2_X1 U17602 ( .A(n17279), .B(n18070), .ZN(n16569) );
  XNOR2_X1 U17603 ( .A(n16570), .B(n16569), .ZN(n16571) );
  XNOR2_X1 U17604 ( .A(n16572), .B(n16571), .ZN(n19370) );
  XNOR2_X1 U17606 ( .A(n16601), .B(n16573), .ZN(n16575) );
  XNOR2_X1 U17607 ( .A(n16574), .B(n16575), .ZN(n16576) );
  OAI21_X1 U17608 ( .B1(n16581), .B2(n19315), .A(n19338), .ZN(n16623) );
  XNOR2_X1 U17609 ( .A(n16835), .B(n20494), .ZN(n16586) );
  XNOR2_X1 U17610 ( .A(n19927), .B(n19243), .ZN(n16583) );
  XNOR2_X1 U17611 ( .A(n16584), .B(n16583), .ZN(n16585) );
  XNOR2_X1 U17612 ( .A(n17367), .B(n16587), .ZN(n17029) );
  XNOR2_X1 U17613 ( .A(n17029), .B(n16588), .ZN(n16592) );
  XNOR2_X1 U17614 ( .A(n17280), .B(n16760), .ZN(n16590) );
  XNOR2_X1 U17615 ( .A(n16927), .B(n2344), .ZN(n16589) );
  XNOR2_X1 U17616 ( .A(n16590), .B(n16589), .ZN(n16591) );
  XNOR2_X1 U17617 ( .A(n16592), .B(n16591), .ZN(n17656) );
  XNOR2_X1 U17618 ( .A(n16938), .B(n18716), .ZN(n16595) );
  XNOR2_X1 U17619 ( .A(n16593), .B(n16741), .ZN(n16594) );
  XNOR2_X1 U17620 ( .A(n16595), .B(n16594), .ZN(n16598) );
  XNOR2_X1 U17621 ( .A(n17040), .B(n16596), .ZN(n16597) );
  XNOR2_X1 U17622 ( .A(n16599), .B(n17012), .ZN(n17286) );
  XNOR2_X1 U17623 ( .A(n17286), .B(n16829), .ZN(n16605) );
  XNOR2_X1 U17624 ( .A(n16600), .B(n16601), .ZN(n17345) );
  XNOR2_X1 U17625 ( .A(n16602), .B(n2203), .ZN(n16603) );
  XNOR2_X1 U17626 ( .A(n17345), .B(n16603), .ZN(n16604) );
  XNOR2_X1 U17627 ( .A(n16605), .B(n16604), .ZN(n19388) );
  AOI21_X1 U17628 ( .B1(n17656), .B2(n20172), .A(n19388), .ZN(n16606) );
  NAND2_X1 U17629 ( .A1(n16683), .A2(n16606), .ZN(n17537) );
  XNOR2_X1 U17630 ( .A(n16608), .B(n16607), .ZN(n17376) );
  XNOR2_X1 U17631 ( .A(n19900), .B(n16914), .ZN(n16609) );
  XNOR2_X1 U17632 ( .A(n17376), .B(n16609), .ZN(n16613) );
  XNOR2_X1 U17633 ( .A(n16844), .B(n17443), .ZN(n16611) );
  XNOR2_X1 U17634 ( .A(n17260), .B(n20593), .ZN(n16610) );
  XNOR2_X1 U17635 ( .A(n16611), .B(n16610), .ZN(n16612) );
  XNOR2_X1 U17636 ( .A(n16613), .B(n16612), .ZN(n17654) );
  XNOR2_X1 U17637 ( .A(n16615), .B(n16614), .ZN(n17325) );
  XNOR2_X1 U17638 ( .A(n16944), .B(n19457), .ZN(n16616) );
  XNOR2_X1 U17639 ( .A(n17325), .B(n16616), .ZN(n16621) );
  INV_X1 U17640 ( .A(n16617), .ZN(n16618) );
  XNOR2_X1 U17641 ( .A(n16618), .B(n16619), .ZN(n16620) );
  XNOR2_X1 U17642 ( .A(n16620), .B(n16621), .ZN(n19390) );
  INV_X1 U17644 ( .A(n19396), .ZN(n19391) );
  NAND3_X1 U17645 ( .A1(n19511), .A2(n19391), .A3(n20172), .ZN(n17536) );
  AND2_X1 U17646 ( .A1(n19329), .A2(n18311), .ZN(n17542) );
  OAI21_X1 U17647 ( .B1(n17542), .B2(n19333), .A(n19340), .ZN(n16622) );
  NAND2_X1 U17648 ( .A1(n16623), .A2(n16622), .ZN(n16625) );
  INV_X1 U17649 ( .A(n106), .ZN(n16624) );
  XNOR2_X1 U17650 ( .A(n16625), .B(n16624), .ZN(Ciphertext[179]) );
  MUX2_X1 U17651 ( .A(n16629), .B(n20092), .S(n17210), .Z(n16628) );
  NOR2_X1 U17652 ( .A1(n19975), .A2(n17208), .ZN(n16627) );
  NOR3_X1 U17653 ( .A1(n20092), .A2(n16629), .A3(n20135), .ZN(n16630) );
  INV_X1 U17654 ( .A(n17508), .ZN(n17513) );
  NOR2_X1 U17655 ( .A1(n16632), .A2(n17513), .ZN(n18340) );
  NOR2_X1 U17656 ( .A1(n18340), .A2(n18342), .ZN(n18287) );
  NOR2_X1 U17657 ( .A1(n18365), .A2(n18362), .ZN(n18286) );
  NOR2_X1 U17660 ( .A1(n19382), .A2(n16666), .ZN(n16640) );
  AOI22_X1 U17661 ( .A1(n16641), .A2(n19386), .B1(n16640), .B2(n1897), .ZN(
        n18341) );
  INV_X1 U17663 ( .A(n18290), .ZN(n18292) );
  INV_X1 U17664 ( .A(n19374), .ZN(n17240) );
  NAND2_X1 U17665 ( .A1(n17240), .A2(n19666), .ZN(n16654) );
  INV_X1 U17666 ( .A(n16642), .ZN(n19373) );
  NAND3_X1 U17668 ( .A1(n16654), .A2(n19373), .A3(n19647), .ZN(n17906) );
  MUX2_X1 U17669 ( .A(n17656), .B(n19390), .S(n19396), .Z(n16643) );
  INV_X1 U17670 ( .A(n16643), .ZN(n16647) );
  OAI21_X1 U17671 ( .B1(n19388), .B2(n17654), .A(n20004), .ZN(n16646) );
  INV_X1 U17672 ( .A(n17654), .ZN(n16644) );
  NOR2_X1 U17673 ( .A1(n16644), .A2(n19396), .ZN(n16645) );
  AOI21_X2 U17674 ( .B1(n16647), .B2(n16646), .A(n16645), .ZN(n18359) );
  OAI211_X1 U17675 ( .C1(n18292), .C2(n18358), .A(n18357), .B(n18359), .ZN(
        n16648) );
  OAI21_X1 U17676 ( .B1(n18286), .B2(n18357), .A(n16648), .ZN(n16650) );
  INV_X1 U17677 ( .A(n18358), .ZN(n18348) );
  NAND2_X1 U17678 ( .A1(n18348), .A2(n18359), .ZN(n17907) );
  NAND2_X1 U17679 ( .A1(n16650), .A2(n16649), .ZN(n16653) );
  INV_X1 U17680 ( .A(n16651), .ZN(n16652) );
  XNOR2_X1 U17681 ( .A(n16653), .B(n16652), .ZN(Ciphertext[5]) );
  AND2_X1 U17682 ( .A1(n19370), .A2(n16642), .ZN(n17596) );
  NAND2_X1 U17683 ( .A1(n19373), .A2(n19666), .ZN(n16655) );
  MUX2_X1 U17684 ( .A(n16655), .B(n16654), .S(n19733), .Z(n16656) );
  NAND2_X1 U17685 ( .A1(n16658), .A2(n17208), .ZN(n16659) );
  NAND2_X1 U17687 ( .A1(n16661), .A2(n20092), .ZN(n16664) );
  NAND2_X1 U17688 ( .A1(n16662), .A2(n17213), .ZN(n16663) );
  NOR2_X1 U17689 ( .A1(n19385), .A2(n17220), .ZN(n16667) );
  AND2_X1 U17690 ( .A1(n16665), .A2(n19382), .ZN(n16668) );
  MUX2_X1 U17691 ( .A(n16667), .B(n16668), .S(n3389), .Z(n16671) );
  OAI21_X1 U17692 ( .B1(n20463), .B2(n19382), .A(n19385), .ZN(n16669) );
  NOR2_X1 U17693 ( .A1(n16669), .A2(n16668), .ZN(n16670) );
  NOR2_X2 U17694 ( .A1(n16671), .A2(n16670), .ZN(n19459) );
  MUX2_X1 U17695 ( .A(n19349), .B(n19353), .S(n16672), .Z(n16677) );
  INV_X1 U17696 ( .A(n20240), .ZN(n16676) );
  NAND3_X1 U17697 ( .A1(n19349), .A2(n19353), .A3(n19351), .ZN(n16675) );
  INV_X1 U17698 ( .A(n18067), .ZN(n19462) );
  NAND2_X1 U17699 ( .A1(n19361), .A2(n19360), .ZN(n17595) );
  NAND2_X1 U17700 ( .A1(n17595), .A2(n20242), .ZN(n16681) );
  NAND2_X1 U17701 ( .A1(n17861), .A2(n19360), .ZN(n19365) );
  NAND2_X1 U17702 ( .A1(n20212), .A2(n19938), .ZN(n16678) );
  NAND2_X1 U17703 ( .A1(n19365), .A2(n16678), .ZN(n16680) );
  NAND3_X1 U17704 ( .A1(n19462), .A2(n19460), .A3(n19453), .ZN(n16682) );
  INV_X1 U17705 ( .A(n16683), .ZN(n16687) );
  INV_X1 U17706 ( .A(n16684), .ZN(n16686) );
  NAND2_X1 U17707 ( .A1(n19390), .A2(n17656), .ZN(n16685) );
  INV_X1 U17708 ( .A(n19453), .ZN(n17091) );
  INV_X1 U17709 ( .A(n457), .ZN(n16688) );
  XNOR2_X1 U17710 ( .A(n16689), .B(n17347), .ZN(n16692) );
  XNOR2_X1 U17711 ( .A(n16691), .B(n16690), .ZN(n17287) );
  XNOR2_X1 U17712 ( .A(n17287), .B(n16692), .ZN(n16694) );
  XNOR2_X1 U17714 ( .A(n19909), .B(n16695), .ZN(n16895) );
  XNOR2_X1 U17715 ( .A(n936), .B(n16895), .ZN(n16700) );
  XNOR2_X1 U17716 ( .A(n17339), .B(n17269), .ZN(n16698) );
  XNOR2_X1 U17717 ( .A(n16755), .B(n1386), .ZN(n16697) );
  XNOR2_X1 U17718 ( .A(n16698), .B(n16697), .ZN(n16699) );
  XNOR2_X1 U17719 ( .A(n16700), .B(n16699), .ZN(n17193) );
  XNOR2_X1 U17720 ( .A(n16844), .B(n17442), .ZN(n16879) );
  XNOR2_X1 U17721 ( .A(n17259), .B(n16879), .ZN(n16704) );
  XNOR2_X1 U17722 ( .A(n17378), .B(n106), .ZN(n16701) );
  XNOR2_X1 U17723 ( .A(n16702), .B(n16701), .ZN(n16703) );
  MUX2_X1 U17724 ( .A(n19684), .B(n935), .S(n18966), .Z(n16726) );
  XNOR2_X1 U17725 ( .A(n16705), .B(n17250), .ZN(n16710) );
  XNOR2_X1 U17726 ( .A(n16706), .B(n18006), .ZN(n16708) );
  XNOR2_X1 U17727 ( .A(n20167), .B(n16707), .ZN(n16870) );
  XNOR2_X1 U17728 ( .A(n16708), .B(n16870), .ZN(n16709) );
  XNOR2_X1 U17730 ( .A(n17276), .B(n16711), .ZN(n16712) );
  XNOR2_X1 U17731 ( .A(n16713), .B(n16712), .ZN(n16717) );
  XNOR2_X1 U17732 ( .A(n16861), .B(n17433), .ZN(n16715) );
  XNOR2_X1 U17733 ( .A(n17279), .B(n311), .ZN(n16714) );
  XNOR2_X1 U17734 ( .A(n16715), .B(n16714), .ZN(n16716) );
  XNOR2_X1 U17735 ( .A(n16717), .B(n16716), .ZN(n17695) );
  NOR2_X1 U17736 ( .A1(n18966), .A2(n17695), .ZN(n16718) );
  NAND2_X1 U17737 ( .A1(n16718), .A2(n17819), .ZN(n16724) );
  XNOR2_X1 U17738 ( .A(n17401), .B(n19720), .ZN(n16899) );
  XNOR2_X1 U17739 ( .A(n16719), .B(n16899), .ZN(n16723) );
  XNOR2_X1 U17740 ( .A(n20104), .B(n17294), .ZN(n16721) );
  XNOR2_X1 U17741 ( .A(n20125), .B(n1904), .ZN(n16720) );
  XNOR2_X1 U17742 ( .A(n16721), .B(n16720), .ZN(n16722) );
  NAND2_X1 U17744 ( .A1(n18961), .A2(n935), .ZN(n18970) );
  NAND2_X1 U17745 ( .A1(n16724), .A2(n18970), .ZN(n16725) );
  AOI22_X1 U17746 ( .A1(n20506), .A2(n17676), .B1(n17867), .B2(n20514), .ZN(
        n16727) );
  NOR2_X1 U17747 ( .A1(n16727), .A2(n19973), .ZN(n16729) );
  AND2_X1 U17748 ( .A1(n17873), .A2(n17872), .ZN(n17677) );
  NOR2_X1 U17752 ( .A1(n17840), .A2(n17835), .ZN(n17062) );
  INV_X1 U17753 ( .A(n17062), .ZN(n16732) );
  XNOR2_X1 U17755 ( .A(n17294), .B(n16900), .ZN(n16735) );
  XNOR2_X1 U17756 ( .A(n16851), .B(n16735), .ZN(n16739) );
  XNOR2_X1 U17757 ( .A(n16960), .B(n20481), .ZN(n16737) );
  XNOR2_X1 U17758 ( .A(n16854), .B(n18854), .ZN(n16736) );
  XNOR2_X1 U17759 ( .A(n16737), .B(n16736), .ZN(n16738) );
  XNOR2_X1 U17760 ( .A(n16739), .B(n16738), .ZN(n18955) );
  INV_X1 U17761 ( .A(n18955), .ZN(n16745) );
  XNOR2_X1 U17762 ( .A(n19889), .B(n16741), .ZN(n16825) );
  XNOR2_X1 U17763 ( .A(n20267), .B(n16742), .ZN(n16744) );
  NOR2_X1 U17764 ( .A1(n16745), .A2(n17831), .ZN(n16767) );
  XNOR2_X1 U17765 ( .A(n19900), .B(n20100), .ZN(n16748) );
  XNOR2_X1 U17766 ( .A(n16749), .B(n16748), .ZN(n16754) );
  XNOR2_X1 U17767 ( .A(n16840), .B(n16750), .ZN(n16752) );
  INV_X1 U17768 ( .A(n2341), .ZN(n19083) );
  XNOR2_X1 U17769 ( .A(n16996), .B(n19083), .ZN(n16751) );
  XNOR2_X1 U17770 ( .A(n16752), .B(n16751), .ZN(n16753) );
  XNOR2_X1 U17771 ( .A(n16754), .B(n16753), .ZN(n18953) );
  INV_X1 U17772 ( .A(n18953), .ZN(n17179) );
  XNOR2_X1 U17773 ( .A(n16757), .B(n16756), .ZN(n16759) );
  AOI21_X1 U17774 ( .B1(n2907), .B2(n17179), .A(n18954), .ZN(n16766) );
  XNOR2_X1 U17775 ( .A(n16761), .B(n16760), .ZN(n16860) );
  XNOR2_X1 U17776 ( .A(n16970), .B(n16971), .ZN(n16763) );
  XNOR2_X1 U17777 ( .A(n20098), .B(n2263), .ZN(n16762) );
  XNOR2_X1 U17778 ( .A(n16763), .B(n16762), .ZN(n16764) );
  XNOR2_X1 U17779 ( .A(n16765), .B(n16764), .ZN(n17180) );
  INV_X1 U17780 ( .A(n17180), .ZN(n18959) );
  MUX2_X1 U17781 ( .A(n16767), .B(n16766), .S(n18959), .Z(n16776) );
  XNOR2_X1 U17782 ( .A(n16987), .B(n2035), .ZN(n16768) );
  XNOR2_X1 U17783 ( .A(n16769), .B(n16768), .ZN(n16774) );
  XNOR2_X1 U17784 ( .A(n17291), .B(n16770), .ZN(n16771) );
  XNOR2_X1 U17785 ( .A(n16771), .B(n16772), .ZN(n16773) );
  NAND2_X1 U17786 ( .A1(n18956), .A2(n17831), .ZN(n17833) );
  INV_X1 U17787 ( .A(n17833), .ZN(n16775) );
  NOR2_X2 U17788 ( .A1(n16776), .A2(n16775), .ZN(n19134) );
  MUX2_X1 U17789 ( .A(n17079), .B(n20239), .S(n17823), .Z(n16778) );
  INV_X1 U17790 ( .A(n17825), .ZN(n17176) );
  NOR2_X1 U17791 ( .A1(n19135), .A2(n16780), .ZN(n19147) );
  INV_X1 U17792 ( .A(n19134), .ZN(n19145) );
  OR2_X1 U17794 ( .A1(n17898), .A2(n19707), .ZN(n16787) );
  NAND2_X1 U17795 ( .A1(n19910), .A2(n16025), .ZN(n16785) );
  NAND2_X1 U17796 ( .A1(n16785), .A2(n17892), .ZN(n16786) );
  AND2_X1 U17797 ( .A1(n17564), .A2(n20432), .ZN(n17161) );
  OAI21_X1 U17798 ( .B1(n17471), .B2(n20432), .A(n18539), .ZN(n16792) );
  NAND2_X1 U17799 ( .A1(n16789), .A2(n18535), .ZN(n18542) );
  NAND2_X1 U17801 ( .A1(n16790), .A2(n18538), .ZN(n16791) );
  OAI21_X1 U17802 ( .B1(n17504), .B2(n16165), .A(n1060), .ZN(n16799) );
  NAND2_X1 U17803 ( .A1(n16795), .A2(n16794), .ZN(n16796) );
  NAND2_X1 U17804 ( .A1(n16797), .A2(n16796), .ZN(n16798) );
  NAND2_X1 U17805 ( .A1(n16799), .A2(n16798), .ZN(n18545) );
  NOR2_X1 U17806 ( .A1(n17584), .A2(n18545), .ZN(n18530) );
  NOR2_X1 U17807 ( .A1(n16801), .A2(n17155), .ZN(n16804) );
  NOR2_X1 U17808 ( .A1(n18530), .A2(n19691), .ZN(n16807) );
  NAND2_X1 U17810 ( .A1(n19682), .A2(n18545), .ZN(n16806) );
  NAND2_X1 U17811 ( .A1(n16807), .A2(n16806), .ZN(n16818) );
  OAI21_X1 U17812 ( .B1(n17243), .B2(n17245), .A(n17479), .ZN(n16808) );
  NAND2_X1 U17813 ( .A1(n16809), .A2(n16808), .ZN(n18540) );
  NAND2_X1 U17814 ( .A1(n18540), .A2(n18541), .ZN(n17925) );
  NAND3_X1 U17815 ( .A1(n17923), .A2(n19682), .A3(n17925), .ZN(n16817) );
  MUX2_X1 U17816 ( .A(n18093), .B(n160), .S(n18097), .Z(n16812) );
  INV_X1 U17817 ( .A(n18093), .ZN(n17475) );
  NOR2_X1 U17818 ( .A1(n17475), .A2(n18095), .ZN(n16811) );
  MUX2_X1 U17819 ( .A(n16812), .B(n16811), .S(n18096), .Z(n16815) );
  NAND2_X1 U17820 ( .A1(n18101), .A2(n226), .ZN(n16813) );
  NOR2_X1 U17821 ( .A1(n16813), .A2(n19774), .ZN(n16814) );
  NAND3_X1 U17822 ( .A1(n16818), .A2(n16817), .A3(n16816), .ZN(n16820) );
  INV_X1 U17823 ( .A(n2337), .ZN(n16819) );
  XNOR2_X1 U17824 ( .A(n16820), .B(n16819), .ZN(Ciphertext[39]) );
  XNOR2_X1 U17825 ( .A(n16821), .B(n16742), .ZN(n16823) );
  XNOR2_X1 U17826 ( .A(n16823), .B(n16822), .ZN(n16827) );
  XNOR2_X1 U17827 ( .A(n19845), .B(n610), .ZN(n16824) );
  XOR2_X1 U17828 ( .A(n16825), .B(n16824), .Z(n16826) );
  XNOR2_X1 U17829 ( .A(n16829), .B(n16828), .ZN(n16833) );
  XNOR2_X1 U17830 ( .A(n16188), .B(n17098), .ZN(n16831) );
  XNOR2_X1 U17831 ( .A(n17288), .B(n2424), .ZN(n16830) );
  XNOR2_X1 U17832 ( .A(n16831), .B(n16830), .ZN(n16832) );
  XNOR2_X1 U17834 ( .A(n16835), .B(n16834), .ZN(n16839) );
  XNOR2_X1 U17835 ( .A(n17111), .B(n16836), .ZN(n17032) );
  XNOR2_X1 U17836 ( .A(n17110), .B(n18078), .ZN(n16837) );
  XNOR2_X1 U17837 ( .A(n17032), .B(n16837), .ZN(n16838) );
  XNOR2_X2 U17838 ( .A(n16839), .B(n16838), .ZN(n18275) );
  XNOR2_X1 U17839 ( .A(n17124), .B(n16840), .ZN(n16843) );
  XNOR2_X1 U17840 ( .A(n19704), .B(n2306), .ZN(n16842) );
  XNOR2_X1 U17841 ( .A(n16843), .B(n16842), .ZN(n16849) );
  INV_X1 U17842 ( .A(n16844), .ZN(n16845) );
  XNOR2_X1 U17843 ( .A(n16845), .B(n947), .ZN(n16846) );
  XNOR2_X1 U17844 ( .A(n16847), .B(n16846), .ZN(n16848) );
  XNOR2_X1 U17845 ( .A(n19720), .B(n17116), .ZN(n16852) );
  XNOR2_X1 U17846 ( .A(n16851), .B(n16852), .ZN(n16858) );
  XNOR2_X1 U17847 ( .A(n16853), .B(n19929), .ZN(n16856) );
  XNOR2_X1 U17848 ( .A(n16854), .B(n2233), .ZN(n16855) );
  XNOR2_X1 U17849 ( .A(n16856), .B(n16855), .ZN(n16857) );
  XNOR2_X1 U17850 ( .A(n16858), .B(n16857), .ZN(n18273) );
  INV_X1 U17851 ( .A(n18269), .ZN(n16866) );
  XNOR2_X1 U17852 ( .A(n16859), .B(n16860), .ZN(n16865) );
  XNOR2_X1 U17853 ( .A(n879), .B(n17275), .ZN(n16863) );
  XNOR2_X1 U17854 ( .A(n16861), .B(n18177), .ZN(n16862) );
  XNOR2_X1 U17855 ( .A(n16863), .B(n16862), .ZN(n16864) );
  XNOR2_X1 U17856 ( .A(n16865), .B(n16864), .ZN(n17769) );
  NAND2_X1 U17857 ( .A1(n16866), .A2(n17769), .ZN(n16867) );
  MUX2_X1 U17858 ( .A(n221), .B(n16867), .S(n18275), .Z(n16868) );
  XNOR2_X1 U17859 ( .A(n16871), .B(n16870), .ZN(n16877) );
  XNOR2_X1 U17860 ( .A(n17005), .B(n16872), .ZN(n16875) );
  XNOR2_X1 U17861 ( .A(n16873), .B(n18170), .ZN(n16874) );
  XNOR2_X1 U17862 ( .A(n16875), .B(n16874), .ZN(n16876) );
  XNOR2_X1 U17864 ( .A(n16878), .B(n16879), .ZN(n16884) );
  XNOR2_X1 U17865 ( .A(n16880), .B(n18396), .ZN(n16881) );
  XNOR2_X1 U17866 ( .A(n16882), .B(n16881), .ZN(n16883) );
  XNOR2_X1 U17867 ( .A(n16884), .B(n16883), .ZN(n18016) );
  AND2_X1 U17868 ( .A1(n20129), .A2(n18016), .ZN(n16913) );
  XNOR2_X1 U17869 ( .A(n16885), .B(n17135), .ZN(n16890) );
  XNOR2_X1 U17870 ( .A(n16886), .B(Key[63]), .ZN(n16888) );
  XNOR2_X1 U17871 ( .A(n16887), .B(n16888), .ZN(n16889) );
  XNOR2_X1 U17872 ( .A(n16892), .B(n16891), .ZN(n16897) );
  XNOR2_X1 U17873 ( .A(n16893), .B(n1840), .ZN(n16894) );
  XNOR2_X1 U17874 ( .A(n16895), .B(n16894), .ZN(n16896) );
  NAND2_X1 U17875 ( .A1(n20158), .A2(n20499), .ZN(n16912) );
  XNOR2_X1 U17876 ( .A(n16898), .B(n16899), .ZN(n16904) );
  XNOR2_X1 U17877 ( .A(n16900), .B(n19321), .ZN(n16901) );
  XNOR2_X1 U17878 ( .A(n16902), .B(n16901), .ZN(n16903) );
  NOR2_X1 U17879 ( .A1(n18976), .A2(n18975), .ZN(n18223) );
  XNOR2_X1 U17880 ( .A(n16905), .B(n16906), .ZN(n16910) );
  XNOR2_X1 U17881 ( .A(n16908), .B(n16907), .ZN(n16909) );
  XNOR2_X1 U17882 ( .A(n17379), .B(n2108), .ZN(n16915) );
  XNOR2_X1 U17883 ( .A(n16915), .B(n16914), .ZN(n16917) );
  XNOR2_X1 U17884 ( .A(n17443), .B(n955), .ZN(n16916) );
  XNOR2_X1 U17885 ( .A(n16917), .B(n16916), .ZN(n16920) );
  XNOR2_X1 U17886 ( .A(n17438), .B(n16918), .ZN(n16919) );
  XNOR2_X1 U17887 ( .A(n16920), .B(n16919), .ZN(n18042) );
  XNOR2_X1 U17888 ( .A(n19836), .B(n2323), .ZN(n16923) );
  XNOR2_X1 U17889 ( .A(n16921), .B(n19713), .ZN(n16922) );
  XNOR2_X1 U17890 ( .A(n16923), .B(n16922), .ZN(n16925) );
  XNOR2_X1 U17891 ( .A(n16988), .B(n17409), .ZN(n16924) );
  XNOR2_X1 U17892 ( .A(n16925), .B(n16924), .ZN(n18043) );
  NAND2_X1 U17893 ( .A1(n20194), .A2(n19916), .ZN(n18950) );
  XNOR2_X1 U17894 ( .A(n16927), .B(n16926), .ZN(n17432) );
  XNOR2_X1 U17895 ( .A(n16929), .B(n16928), .ZN(n16930) );
  XNOR2_X1 U17896 ( .A(n16930), .B(n17432), .ZN(n16935) );
  XNOR2_X1 U17897 ( .A(n16931), .B(n17366), .ZN(n17278) );
  XNOR2_X1 U17898 ( .A(n16932), .B(n17851), .ZN(n16933) );
  XNOR2_X1 U17899 ( .A(n17278), .B(n16933), .ZN(n16934) );
  XNOR2_X1 U17900 ( .A(n17360), .B(n16936), .ZN(n17249) );
  XNOR2_X1 U17901 ( .A(n19863), .B(n17249), .ZN(n16943) );
  XNOR2_X1 U17902 ( .A(n16938), .B(n19180), .ZN(n16941) );
  XNOR2_X1 U17903 ( .A(n16939), .B(n16181), .ZN(n16940) );
  XNOR2_X1 U17904 ( .A(n16941), .B(n16940), .ZN(n16942) );
  XNOR2_X2 U17905 ( .A(n16943), .B(n16942), .ZN(n18946) );
  XNOR2_X1 U17906 ( .A(n16945), .B(n16944), .ZN(n17403) );
  XNOR2_X1 U17907 ( .A(n17403), .B(n16946), .ZN(n16951) );
  XNOR2_X1 U17908 ( .A(n16947), .B(n17295), .ZN(n16949) );
  XNOR2_X1 U17909 ( .A(n17330), .B(n2284), .ZN(n16948) );
  XNOR2_X1 U17910 ( .A(n16949), .B(n16948), .ZN(n16950) );
  XNOR2_X1 U17911 ( .A(n16951), .B(n16950), .ZN(n18046) );
  NAND2_X1 U17913 ( .A1(n2586), .A2(n18946), .ZN(n16959) );
  XNOR2_X1 U17914 ( .A(n16952), .B(n16953), .ZN(n16958) );
  XNOR2_X1 U17915 ( .A(n16954), .B(n19706), .ZN(n16956) );
  XNOR2_X1 U17916 ( .A(n902), .B(n17932), .ZN(n16955) );
  XNOR2_X1 U17917 ( .A(n16956), .B(n16955), .ZN(n16957) );
  NAND2_X1 U17918 ( .A1(n19681), .A2(n17054), .ZN(n18891) );
  OAI21_X1 U17919 ( .B1(n19905), .B2(n18897), .A(n18891), .ZN(n17059) );
  XNOR2_X1 U17920 ( .A(n16961), .B(n16960), .ZN(n17326) );
  XNOR2_X1 U17921 ( .A(n16962), .B(n17326), .ZN(n16968) );
  XNOR2_X1 U17922 ( .A(n16964), .B(n16963), .ZN(n17118) );
  XNOR2_X1 U17923 ( .A(n20481), .B(n2384), .ZN(n16966) );
  XNOR2_X1 U17924 ( .A(n17118), .B(n16966), .ZN(n16967) );
  XNOR2_X1 U17925 ( .A(n16967), .B(n16968), .ZN(n18029) );
  INV_X1 U17926 ( .A(n18029), .ZN(n18926) );
  XNOR2_X1 U17927 ( .A(n16970), .B(n16969), .ZN(n17370) );
  XNOR2_X1 U17928 ( .A(n17133), .B(n16971), .ZN(n16972) );
  XNOR2_X1 U17929 ( .A(n17370), .B(n16972), .ZN(n16978) );
  XNOR2_X1 U17930 ( .A(n19659), .B(n16973), .ZN(n17139) );
  XNOR2_X1 U17931 ( .A(n16975), .B(n17544), .ZN(n16976) );
  XNOR2_X1 U17932 ( .A(n17139), .B(n16976), .ZN(n16977) );
  XNOR2_X1 U17933 ( .A(n16978), .B(n16977), .ZN(n18024) );
  XNOR2_X1 U17934 ( .A(n17108), .B(n16979), .ZN(n16986) );
  XNOR2_X1 U17935 ( .A(n16981), .B(n16980), .ZN(n16984) );
  XNOR2_X1 U17936 ( .A(n16982), .B(n18830), .ZN(n16983) );
  XNOR2_X1 U17937 ( .A(n16984), .B(n16983), .ZN(n16985) );
  MUX2_X1 U17939 ( .A(n18926), .B(n18024), .S(n18025), .Z(n17011) );
  XNOR2_X1 U17940 ( .A(n16988), .B(n16987), .ZN(n16989) );
  XNOR2_X1 U17941 ( .A(n16990), .B(n16989), .ZN(n16995) );
  XNOR2_X1 U17942 ( .A(n17407), .B(n19783), .ZN(n17346) );
  XNOR2_X1 U17943 ( .A(n17102), .B(n2337), .ZN(n16993) );
  XNOR2_X1 U17944 ( .A(n17346), .B(n16993), .ZN(n16994) );
  XNOR2_X1 U17945 ( .A(n16995), .B(n16994), .ZN(n18026) );
  INV_X1 U17946 ( .A(n18026), .ZN(n18931) );
  NOR2_X1 U17947 ( .A1(n18931), .A2(n18025), .ZN(n17324) );
  XNOR2_X1 U17948 ( .A(n16996), .B(n2257), .ZN(n16997) );
  XNOR2_X1 U17949 ( .A(n16998), .B(n16997), .ZN(n17001) );
  XNOR2_X1 U17950 ( .A(n17444), .B(n16999), .ZN(n17375) );
  XNOR2_X1 U17951 ( .A(n17125), .B(n17375), .ZN(n17000) );
  XNOR2_X1 U17952 ( .A(n17001), .B(n17000), .ZN(n18927) );
  NOR2_X1 U17953 ( .A1(n20207), .A2(n18927), .ZN(n17699) );
  NOR2_X1 U17954 ( .A1(n17324), .A2(n17699), .ZN(n17010) );
  XNOR2_X1 U17955 ( .A(n15935), .B(n17002), .ZN(n17004) );
  XNOR2_X1 U17956 ( .A(n17004), .B(n17003), .ZN(n17009) );
  XNOR2_X1 U17957 ( .A(n864), .B(n17355), .ZN(n17007) );
  XNOR2_X1 U17958 ( .A(n17005), .B(n2394), .ZN(n17006) );
  XNOR2_X1 U17959 ( .A(n17006), .B(n17007), .ZN(n17008) );
  INV_X1 U17961 ( .A(n18928), .ZN(n18932) );
  XNOR2_X1 U17962 ( .A(n17012), .B(n17098), .ZN(n17013) );
  XNOR2_X1 U17963 ( .A(n17345), .B(n17013), .ZN(n17018) );
  XNOR2_X1 U17964 ( .A(n17288), .B(n17347), .ZN(n17016) );
  XNOR2_X1 U17965 ( .A(n17014), .B(n1869), .ZN(n17015) );
  XNOR2_X1 U17966 ( .A(n17016), .B(n17015), .ZN(n17017) );
  XNOR2_X1 U17967 ( .A(n17019), .B(n17325), .ZN(n17023) );
  XNOR2_X1 U17968 ( .A(n17116), .B(n2382), .ZN(n17021) );
  XNOR2_X1 U17969 ( .A(n17021), .B(n17020), .ZN(n17022) );
  XNOR2_X1 U17970 ( .A(n17023), .B(n17022), .ZN(n18939) );
  NAND2_X1 U17971 ( .A1(n20501), .A2(n18939), .ZN(n18021) );
  INV_X1 U17972 ( .A(n19893), .ZN(n17025) );
  XNOR2_X1 U17973 ( .A(n17025), .B(n17024), .ZN(n17027) );
  XNOR2_X1 U17974 ( .A(n17026), .B(n17027), .ZN(n17031) );
  XNOR2_X1 U17975 ( .A(n17029), .B(n17028), .ZN(n17030) );
  XNOR2_X1 U17976 ( .A(n17031), .B(n17030), .ZN(n18936) );
  XNOR2_X1 U17979 ( .A(n17035), .B(n19336), .ZN(n17037) );
  XNOR2_X1 U17980 ( .A(n17036), .B(n17037), .ZN(n17038) );
  XNOR2_X1 U17982 ( .A(n17040), .B(n17357), .ZN(n17044) );
  XNOR2_X1 U17983 ( .A(n16181), .B(n19844), .ZN(n17042) );
  XNOR2_X1 U17984 ( .A(n17143), .B(n18848), .ZN(n17041) );
  XNOR2_X1 U17985 ( .A(n17042), .B(n17041), .ZN(n17043) );
  INV_X1 U17986 ( .A(n17187), .ZN(n18941) );
  AOI21_X1 U17987 ( .B1(n19723), .B2(n18941), .A(n18939), .ZN(n17045) );
  NAND2_X1 U17988 ( .A1(n17705), .A2(n17045), .ZN(n17053) );
  NOR2_X1 U17989 ( .A1(n20501), .A2(n17187), .ZN(n17051) );
  XNOR2_X1 U17990 ( .A(n17046), .B(n17376), .ZN(n17050) );
  XNOR2_X1 U17991 ( .A(n17378), .B(n17637), .ZN(n17047) );
  XNOR2_X1 U17992 ( .A(n17048), .B(n17047), .ZN(n17049) );
  NAND2_X1 U17993 ( .A1(n17051), .A2(n20452), .ZN(n17052) );
  OAI211_X1 U17994 ( .C1(n18021), .C2(n889), .A(n17053), .B(n17052), .ZN(
        n18916) );
  INV_X1 U17995 ( .A(n18916), .ZN(n18876) );
  AND2_X1 U17996 ( .A1(n17054), .A2(n18890), .ZN(n18874) );
  AOI22_X1 U17997 ( .A1(n19684), .A2(n935), .B1(n18966), .B2(n18961), .ZN(
        n17057) );
  NAND2_X1 U17998 ( .A1(n18966), .A2(n17818), .ZN(n17055) );
  AOI21_X1 U18000 ( .B1(n17059), .B2(n18921), .A(n17058), .ZN(n17061) );
  XNOR2_X1 U18001 ( .A(n17061), .B(n17060), .ZN(Ciphertext[106]) );
  NAND2_X1 U18002 ( .A1(n17836), .A2(n17715), .ZN(n17196) );
  OR2_X1 U18003 ( .A1(n17196), .A2(n17062), .ZN(n17065) );
  INV_X1 U18004 ( .A(n17063), .ZN(n17714) );
  NAND2_X1 U18005 ( .A1(n17714), .A2(n17840), .ZN(n17718) );
  NOR2_X1 U18006 ( .A1(n17840), .A2(n17715), .ZN(n17197) );
  NAND2_X1 U18007 ( .A1(n17197), .A2(n17838), .ZN(n17064) );
  MUX2_X1 U18008 ( .A(n17180), .B(n18955), .S(n18954), .Z(n17067) );
  INV_X1 U18009 ( .A(n18954), .ZN(n17178) );
  NAND2_X1 U18010 ( .A1(n17178), .A2(n18953), .ZN(n17066) );
  AOI21_X1 U18012 ( .B1(n854), .B2(n17181), .A(n17897), .ZN(n17070) );
  NAND2_X1 U18013 ( .A1(n17070), .A2(n17895), .ZN(n17073) );
  INV_X1 U18014 ( .A(n17896), .ZN(n17893) );
  NAND3_X1 U18015 ( .A1(n17893), .A2(n854), .A3(n17181), .ZN(n17072) );
  NAND3_X1 U18016 ( .A1(n17892), .A2(n17896), .A3(n17897), .ZN(n17071) );
  MUX2_X1 U18018 ( .A(n19163), .B(n19155), .S(n19162), .Z(n17088) );
  NAND2_X1 U18019 ( .A1(n17868), .A2(n20514), .ZN(n17076) );
  NAND2_X1 U18020 ( .A1(n19973), .A2(n17078), .ZN(n17075) );
  MUX2_X1 U18021 ( .A(n17076), .B(n17075), .S(n20506), .Z(n17077) );
  MUX2_X1 U18022 ( .A(n17823), .B(n17080), .S(n17079), .Z(n17083) );
  MUX2_X1 U18023 ( .A(n19667), .B(n17824), .S(n17825), .Z(n17082) );
  NOR2_X1 U18025 ( .A1(n19164), .A2(n19162), .ZN(n17084) );
  AOI21_X1 U18026 ( .B1(n19165), .B2(n19948), .A(n17084), .ZN(n17087) );
  OAI21_X1 U18027 ( .B1(n19947), .B2(n20185), .A(n17886), .ZN(n17085) );
  INV_X1 U18028 ( .A(n17891), .ZN(n17601) );
  XNOR2_X1 U18030 ( .A(n17090), .B(n17089), .ZN(Ciphertext[140]) );
  AND2_X1 U18031 ( .A1(n19463), .A2(n19460), .ZN(n17092) );
  MUX2_X1 U18032 ( .A(n20140), .B(n19453), .S(n20152), .Z(n17093) );
  NOR2_X1 U18033 ( .A1(n17093), .A2(n19460), .ZN(n17094) );
  NOR2_X1 U18035 ( .A1(n18111), .A2(n20114), .ZN(n17096) );
  MUX2_X1 U18036 ( .A(n19885), .B(n20488), .S(n17458), .Z(n17097) );
  XNOR2_X1 U18037 ( .A(n17099), .B(n17098), .ZN(n17100) );
  XNOR2_X1 U18038 ( .A(n17101), .B(n17100), .ZN(n17106) );
  XNOR2_X1 U18039 ( .A(n17102), .B(n573), .ZN(n17103) );
  XNOR2_X1 U18040 ( .A(n17104), .B(n17103), .ZN(n17105) );
  XNOR2_X1 U18041 ( .A(n17107), .B(n17108), .ZN(n17115) );
  XNOR2_X1 U18042 ( .A(n17109), .B(n911), .ZN(n17113) );
  XNOR2_X1 U18043 ( .A(n17111), .B(n18011), .ZN(n17112) );
  XNOR2_X1 U18044 ( .A(n17113), .B(n17112), .ZN(n17114) );
  XNOR2_X1 U18045 ( .A(n17116), .B(n2096), .ZN(n17117) );
  XNOR2_X1 U18046 ( .A(n17118), .B(n17117), .ZN(n17122) );
  XNOR2_X1 U18047 ( .A(n17120), .B(n17119), .ZN(n17121) );
  XNOR2_X1 U18048 ( .A(n17121), .B(n17122), .ZN(n17547) );
  INV_X1 U18049 ( .A(n17547), .ZN(n18229) );
  XNOR2_X1 U18050 ( .A(n17124), .B(n17123), .ZN(n17126) );
  XNOR2_X1 U18051 ( .A(n17126), .B(n17125), .ZN(n17132) );
  XNOR2_X1 U18052 ( .A(n19882), .B(n17442), .ZN(n17130) );
  XNOR2_X1 U18053 ( .A(n17128), .B(n18809), .ZN(n17129) );
  XNOR2_X1 U18054 ( .A(n17130), .B(n17129), .ZN(n17131) );
  XNOR2_X1 U18055 ( .A(n17132), .B(n17131), .ZN(n17390) );
  INV_X1 U18056 ( .A(n17390), .ZN(n18232) );
  XNOR2_X1 U18057 ( .A(n19893), .B(n17133), .ZN(n17136) );
  XNOR2_X1 U18058 ( .A(n17136), .B(n17135), .ZN(n17140) );
  XNOR2_X1 U18059 ( .A(n880), .B(n18084), .ZN(n17138) );
  XNOR2_X1 U18060 ( .A(n17142), .B(n17141), .ZN(n17147) );
  XNOR2_X1 U18061 ( .A(n864), .B(n2368), .ZN(n17145) );
  XNOR2_X1 U18062 ( .A(n17143), .B(n17416), .ZN(n17144) );
  XNOR2_X1 U18063 ( .A(n17145), .B(n17144), .ZN(n17146) );
  XNOR2_X1 U18064 ( .A(n17147), .B(n17146), .ZN(n18226) );
  OR2_X1 U18065 ( .A1(n18226), .A2(n17390), .ZN(n18121) );
  MUX2_X1 U18066 ( .A(n18121), .B(n18229), .S(n17545), .Z(n17148) );
  OAI22_X1 U18068 ( .A1(n19672), .A2(n17553), .B1(n17149), .B2(n18105), .ZN(
        n17153) );
  AND2_X1 U18069 ( .A1(n19672), .A2(n17954), .ZN(n17151) );
  NOR2_X1 U18070 ( .A1(n19737), .A2(n17959), .ZN(n17150) );
  MUX2_X1 U18073 ( .A(n17489), .B(n17154), .S(n19675), .Z(n17159) );
  INV_X1 U18074 ( .A(n17491), .ZN(n17156) );
  NOR2_X1 U18075 ( .A1(n17156), .A2(n19675), .ZN(n17157) );
  INV_X1 U18076 ( .A(n17623), .ZN(n17918) );
  NAND3_X1 U18077 ( .A1(n18596), .A2(n19669), .A3(n17918), .ZN(n17169) );
  NOR2_X1 U18078 ( .A1(n18539), .A2(n18535), .ZN(n17563) );
  INV_X1 U18079 ( .A(n17563), .ZN(n17162) );
  NAND2_X1 U18080 ( .A1(n17562), .A2(n18535), .ZN(n17160) );
  OAI21_X1 U18081 ( .B1(n18592), .B2(n18589), .A(n19665), .ZN(n17168) );
  NOR2_X1 U18082 ( .A1(n20365), .A2(n18592), .ZN(n17167) );
  MUX2_X2 U18083 ( .A(n17166), .B(n17165), .S(n160), .Z(n18597) );
  AOI22_X1 U18084 ( .A1(n17169), .A2(n17168), .B1(n17167), .B2(n18597), .ZN(
        n17171) );
  XNOR2_X1 U18085 ( .A(n17171), .B(n17170), .ZN(Ciphertext[48]) );
  OR2_X1 U18086 ( .A1(n17826), .A2(n16262), .ZN(n17177) );
  MUX2_X1 U18087 ( .A(n17825), .B(n17172), .S(n17824), .Z(n17174) );
  OR2_X1 U18088 ( .A1(n17825), .A2(n17823), .ZN(n17173) );
  MUX2_X1 U18089 ( .A(n17174), .B(n17173), .S(n17822), .Z(n17175) );
  MUX2_X1 U18090 ( .A(n17179), .B(n17178), .S(n20221), .Z(n19111) );
  OR2_X1 U18091 ( .A1(n18954), .A2(n18955), .ZN(n17832) );
  NAND2_X1 U18092 ( .A1(n18959), .A2(n18954), .ZN(n17829) );
  NAND2_X1 U18093 ( .A1(n17832), .A2(n17829), .ZN(n19106) );
  INV_X1 U18095 ( .A(n17181), .ZN(n17894) );
  AOI21_X1 U18096 ( .B1(n17894), .B2(n17893), .A(n17892), .ZN(n17186) );
  OAI21_X1 U18097 ( .B1(n17184), .B2(n17183), .A(n17182), .ZN(n17185) );
  NAND2_X1 U18098 ( .A1(n19093), .A2(n19911), .ZN(n19088) );
  INV_X1 U18099 ( .A(n18938), .ZN(n18934) );
  NOR2_X1 U18100 ( .A1(n18934), .A2(n18937), .ZN(n17707) );
  NAND2_X1 U18101 ( .A1(n17707), .A2(n18935), .ZN(n17192) );
  INV_X1 U18102 ( .A(n18019), .ZN(n18940) );
  INV_X1 U18103 ( .A(n20452), .ZN(n17188) );
  NAND3_X1 U18104 ( .A1(n18940), .A2(n17188), .A3(n889), .ZN(n17191) );
  NAND3_X1 U18105 ( .A1(n19723), .A2(n20452), .A3(n18935), .ZN(n17190) );
  INV_X1 U18106 ( .A(n18939), .ZN(n18020) );
  NAND2_X1 U18107 ( .A1(n18020), .A2(n19723), .ZN(n17189) );
  INV_X1 U18108 ( .A(n17695), .ZN(n17692) );
  NAND3_X1 U18109 ( .A1(n18961), .A2(n227), .A3(n17692), .ZN(n17195) );
  INV_X1 U18110 ( .A(n17193), .ZN(n17819) );
  OAI211_X1 U18111 ( .C1(n18966), .C2(n20127), .A(n17819), .B(n18962), .ZN(
        n17194) );
  OAI211_X1 U18112 ( .C1(n19684), .C2(n227), .A(n17195), .B(n17194), .ZN(
        n17203) );
  NAND2_X1 U18113 ( .A1(n19115), .A2(n17203), .ZN(n19085) );
  NAND2_X1 U18114 ( .A1(n19088), .A2(n19085), .ZN(n17205) );
  INV_X1 U18115 ( .A(n19093), .ZN(n19116) );
  NOR2_X1 U18116 ( .A1(n17196), .A2(n17063), .ZN(n17198) );
  NOR2_X1 U18117 ( .A1(n17198), .A2(n17197), .ZN(n17202) );
  NOR3_X1 U18118 ( .A1(n3755), .A2(n17840), .A3(n17838), .ZN(n17200) );
  AOI21_X2 U18119 ( .B1(n17202), .B2(n17201), .A(n17200), .ZN(n19098) );
  INV_X1 U18120 ( .A(n17203), .ZN(n19095) );
  OAI21_X1 U18121 ( .B1(n19098), .B2(n19095), .A(n19115), .ZN(n17204) );
  AOI22_X1 U18122 ( .A1(n19105), .A2(n17205), .B1(n19116), .B2(n17204), .ZN(
        n17206) );
  XNOR2_X1 U18123 ( .A(n17206), .B(n2216), .ZN(Ciphertext[131]) );
  AOI21_X1 U18124 ( .B1(n17211), .B2(n17208), .A(n20092), .ZN(n17209) );
  INV_X1 U18125 ( .A(n17209), .ZN(n17216) );
  AND2_X1 U18126 ( .A1(n17210), .A2(n17211), .ZN(n17212) );
  AOI22_X1 U18127 ( .A1(n17214), .A2(n17213), .B1(n16465), .B2(n17212), .ZN(
        n17215) );
  MUX2_X1 U18129 ( .A(n19383), .B(n17218), .S(n1897), .Z(n17222) );
  MUX2_X1 U18130 ( .A(n19956), .B(n17507), .S(n17512), .Z(n17230) );
  NAND2_X1 U18131 ( .A1(n3573), .A2(n17508), .ZN(n17228) );
  NAND3_X1 U18133 ( .A1(n16633), .A2(n14845), .A3(n19956), .ZN(n17227) );
  OAI21_X1 U18134 ( .B1(n19956), .B2(n17228), .A(n17227), .ZN(n17229) );
  INV_X1 U18135 ( .A(n17231), .ZN(n17232) );
  NAND2_X1 U18136 ( .A1(n17232), .A2(n19353), .ZN(n17235) );
  OAI211_X1 U18137 ( .C1(n19352), .C2(n19348), .A(n19349), .B(n20273), .ZN(
        n17233) );
  OAI21_X1 U18138 ( .B1(n17240), .B2(n19666), .A(n19372), .ZN(n17238) );
  INV_X1 U18139 ( .A(n17243), .ZN(n17241) );
  NAND2_X1 U18141 ( .A1(n17242), .A2(n20230), .ZN(n17247) );
  AOI22_X1 U18142 ( .A1(n17482), .A2(n17245), .B1(n20354), .B2(n17243), .ZN(
        n17246) );
  INV_X1 U18143 ( .A(n17249), .ZN(n17251) );
  XNOR2_X1 U18144 ( .A(n17250), .B(n17251), .ZN(n17257) );
  XNOR2_X1 U18145 ( .A(n19807), .B(n2310), .ZN(n17255) );
  XNOR2_X1 U18146 ( .A(n17253), .B(n19845), .ZN(n17254) );
  XNOR2_X1 U18147 ( .A(n17255), .B(n17254), .ZN(n17256) );
  XNOR2_X1 U18148 ( .A(n17257), .B(n17256), .ZN(n17303) );
  XNOR2_X1 U18149 ( .A(n17259), .B(n17258), .ZN(n17266) );
  XNOR2_X1 U18150 ( .A(n947), .B(n17260), .ZN(n17264) );
  XNOR2_X1 U18151 ( .A(n17264), .B(n17263), .ZN(n17265) );
  NOR2_X1 U18152 ( .A1(n17753), .A2(n18038), .ZN(n17307) );
  XNOR2_X1 U18153 ( .A(n17268), .B(n17267), .ZN(n17274) );
  XNOR2_X1 U18154 ( .A(n17269), .B(n19706), .ZN(n17272) );
  XNOR2_X1 U18155 ( .A(n17270), .B(n18146), .ZN(n17271) );
  XNOR2_X1 U18156 ( .A(n17272), .B(n17271), .ZN(n17273) );
  XNOR2_X1 U18157 ( .A(n17274), .B(n17273), .ZN(n17982) );
  XNOR2_X1 U18158 ( .A(n17275), .B(n17276), .ZN(n17277) );
  XNOR2_X1 U18159 ( .A(n17278), .B(n17277), .ZN(n17285) );
  XNOR2_X1 U18160 ( .A(n17280), .B(n17279), .ZN(n17283) );
  XNOR2_X1 U18161 ( .A(n17281), .B(n2445), .ZN(n17282) );
  XNOR2_X1 U18162 ( .A(n17283), .B(n17282), .ZN(n17284) );
  OR2_X1 U18163 ( .A1(n17982), .A2(n18238), .ZN(n18241) );
  XNOR2_X1 U18164 ( .A(n17287), .B(n17286), .ZN(n17292) );
  XNOR2_X1 U18165 ( .A(n19836), .B(n2305), .ZN(n17290) );
  INV_X1 U18166 ( .A(n17288), .ZN(n17289) );
  XNOR2_X1 U18167 ( .A(n17293), .B(n17328), .ZN(n17297) );
  XNOR2_X1 U18168 ( .A(n17294), .B(n17295), .ZN(n17296) );
  XNOR2_X1 U18169 ( .A(n17298), .B(n17299), .ZN(n17302) );
  XNOR2_X1 U18170 ( .A(n17300), .B(n17993), .ZN(n17301) );
  NAND2_X1 U18171 ( .A1(n17981), .A2(n18238), .ZN(n17983) );
  INV_X1 U18176 ( .A(n19766), .ZN(n17992) );
  INV_X1 U18177 ( .A(n18975), .ZN(n17308) );
  NAND2_X1 U18178 ( .A1(n17309), .A2(n18977), .ZN(n17313) );
  NAND2_X1 U18179 ( .A1(n18221), .A2(n20158), .ZN(n17311) );
  MUX2_X1 U18181 ( .A(n17311), .B(n17310), .S(n20499), .Z(n17312) );
  OAI21_X1 U18183 ( .B1(n19916), .B2(n18946), .A(n17315), .ZN(n17316) );
  NAND2_X1 U18184 ( .A1(n17316), .A2(n20194), .ZN(n17319) );
  NAND2_X1 U18185 ( .A1(n17317), .A2(n19916), .ZN(n17318) );
  NAND2_X1 U18187 ( .A1(n18275), .A2(n18270), .ZN(n18274) );
  OAI21_X1 U18188 ( .B1(n18269), .B2(n18270), .A(n18274), .ZN(n17320) );
  NAND2_X1 U18189 ( .A1(n20097), .A2(n19794), .ZN(n18817) );
  OAI21_X1 U18190 ( .B1(n17992), .B2(n20422), .A(n18817), .ZN(n17388) );
  OAI21_X1 U18191 ( .B1(n2120), .B2(n18928), .A(n18926), .ZN(n17323) );
  NOR2_X1 U18192 ( .A1(n20207), .A2(n18926), .ZN(n17748) );
  INV_X1 U18193 ( .A(n18024), .ZN(n18929) );
  INV_X1 U18194 ( .A(n18927), .ZN(n17700) );
  NOR2_X1 U18195 ( .A1(n18928), .A2(n17700), .ZN(n17321) );
  AOI22_X1 U18196 ( .A1(n17748), .A2(n18929), .B1(n17321), .B2(n17749), .ZN(
        n17322) );
  OAI21_X1 U18197 ( .B1(n17324), .B2(n17323), .A(n17322), .ZN(n18844) );
  INV_X1 U18198 ( .A(n18844), .ZN(n18818) );
  XNOR2_X1 U18199 ( .A(n17325), .B(n17326), .ZN(n17334) );
  XNOR2_X1 U18200 ( .A(n17328), .B(n20125), .ZN(n17332) );
  INV_X1 U18201 ( .A(n18090), .ZN(n17329) );
  XNOR2_X1 U18202 ( .A(n17330), .B(n17329), .ZN(n17331) );
  XNOR2_X1 U18203 ( .A(n17332), .B(n17331), .ZN(n17333) );
  XNOR2_X1 U18204 ( .A(n17334), .B(n17333), .ZN(n17394) );
  INV_X1 U18205 ( .A(n17394), .ZN(n18258) );
  XNOR2_X1 U18206 ( .A(n17335), .B(n20192), .ZN(n17336) );
  XNOR2_X1 U18207 ( .A(n17337), .B(n17336), .ZN(n17344) );
  XNOR2_X1 U18208 ( .A(n17339), .B(n17338), .ZN(n17342) );
  XNOR2_X1 U18209 ( .A(n19706), .B(n19052), .ZN(n17341) );
  XNOR2_X1 U18210 ( .A(n17342), .B(n17341), .ZN(n17343) );
  NOR2_X1 U18212 ( .A1(n18258), .A2(n19787), .ZN(n17976) );
  INV_X1 U18213 ( .A(n17976), .ZN(n17978) );
  XNOR2_X1 U18214 ( .A(n17345), .B(n17346), .ZN(n17353) );
  XNOR2_X1 U18215 ( .A(n19713), .B(n17347), .ZN(n17351) );
  XNOR2_X1 U18216 ( .A(n19836), .B(n20672), .ZN(n17350) );
  XNOR2_X1 U18217 ( .A(n17351), .B(n17350), .ZN(n17352) );
  XNOR2_X1 U18218 ( .A(n17353), .B(n17352), .ZN(n17374) );
  XNOR2_X1 U18219 ( .A(n15935), .B(n17355), .ZN(n17356) );
  XNOR2_X1 U18220 ( .A(n17356), .B(n17357), .ZN(n17364) );
  XNOR2_X1 U18221 ( .A(n17359), .B(n17358), .ZN(n17362) );
  XNOR2_X1 U18222 ( .A(n17360), .B(n17587), .ZN(n17361) );
  XNOR2_X1 U18223 ( .A(n17362), .B(n17361), .ZN(n17363) );
  NAND2_X1 U18224 ( .A1(n18262), .A2(n18753), .ZN(n17396) );
  XNOR2_X1 U18225 ( .A(n17366), .B(n17365), .ZN(n17368) );
  XNOR2_X1 U18226 ( .A(n17367), .B(n17368), .ZN(n17369) );
  XNOR2_X1 U18227 ( .A(n17370), .B(n17369), .ZN(n17372) );
  NAND2_X1 U18228 ( .A1(n19787), .A2(n18260), .ZN(n17373) );
  NAND3_X1 U18229 ( .A1(n17978), .A2(n17396), .A3(n17373), .ZN(n17385) );
  INV_X1 U18230 ( .A(n17374), .ZN(n17977) );
  XNOR2_X1 U18231 ( .A(n17376), .B(n17375), .ZN(n17382) );
  XNOR2_X1 U18232 ( .A(n19798), .B(n456), .ZN(n17380) );
  XNOR2_X1 U18233 ( .A(n17382), .B(n17381), .ZN(n18138) );
  INV_X1 U18234 ( .A(n18138), .ZN(n18137) );
  NAND2_X1 U18235 ( .A1(n18137), .A2(n19787), .ZN(n17383) );
  NAND2_X1 U18237 ( .A1(n18844), .A2(n20097), .ZN(n17386) );
  AOI21_X1 U18239 ( .B1(n20276), .B2(n17386), .A(n20130), .ZN(n17387) );
  AOI21_X1 U18240 ( .B1(n17388), .B2(n18818), .A(n17387), .ZN(n17389) );
  XNOR2_X1 U18241 ( .A(n17389), .B(n2055), .ZN(Ciphertext[90]) );
  INV_X1 U18242 ( .A(n18226), .ZN(n17549) );
  NOR2_X1 U18243 ( .A1(n17549), .A2(n19771), .ZN(n17392) );
  AOI21_X1 U18244 ( .B1(n18226), .B2(n17390), .A(n18233), .ZN(n17391) );
  NOR2_X1 U18245 ( .A1(n18226), .A2(n17545), .ZN(n18123) );
  NOR2_X2 U18246 ( .A1(n17393), .A2(n18123), .ZN(n18698) );
  NOR2_X1 U18247 ( .A1(n17394), .A2(n17758), .ZN(n17395) );
  INV_X1 U18248 ( .A(n18260), .ZN(n18750) );
  INV_X1 U18250 ( .A(n19751), .ZN(n17463) );
  XNOR2_X1 U18251 ( .A(n17399), .B(n17400), .ZN(n17405) );
  XNOR2_X1 U18252 ( .A(n17401), .B(n641), .ZN(n17402) );
  XNOR2_X1 U18253 ( .A(n17403), .B(n17402), .ZN(n17404) );
  XNOR2_X1 U18254 ( .A(n17407), .B(n17406), .ZN(n17408) );
  XNOR2_X1 U18255 ( .A(n17409), .B(n17408), .ZN(n17415) );
  XNOR2_X1 U18256 ( .A(n17411), .B(n17410), .ZN(n17413) );
  INV_X1 U18257 ( .A(n2417), .ZN(n19038) );
  XNOR2_X1 U18258 ( .A(n17413), .B(n17412), .ZN(n17414) );
  XNOR2_X1 U18260 ( .A(n20167), .B(n2055), .ZN(n17417) );
  XNOR2_X1 U18261 ( .A(n17418), .B(n17417), .ZN(n17422) );
  XNOR2_X1 U18262 ( .A(n17419), .B(n17420), .ZN(n17421) );
  MUX2_X1 U18263 ( .A(n18130), .B(n2475), .S(n19744), .Z(n17450) );
  XNOR2_X1 U18264 ( .A(n17424), .B(n17423), .ZN(n17430) );
  XNOR2_X1 U18265 ( .A(n19909), .B(n17425), .ZN(n17428) );
  XNOR2_X1 U18266 ( .A(n17426), .B(n345), .ZN(n17427) );
  XNOR2_X1 U18267 ( .A(n17428), .B(n17427), .ZN(n17429) );
  XNOR2_X1 U18268 ( .A(n17430), .B(n17429), .ZN(n17946) );
  XNOR2_X1 U18269 ( .A(n17431), .B(n17432), .ZN(n17437) );
  XNOR2_X1 U18270 ( .A(n17433), .B(n18284), .ZN(n17434) );
  XOR2_X1 U18271 ( .A(n17435), .B(n17434), .Z(n17436) );
  XNOR2_X1 U18274 ( .A(n17438), .B(n17439), .ZN(n17441) );
  XNOR2_X1 U18275 ( .A(n17440), .B(n17441), .ZN(n17448) );
  XNOR2_X1 U18276 ( .A(n17443), .B(n17442), .ZN(n17446) );
  XNOR2_X1 U18277 ( .A(n17444), .B(n538), .ZN(n17445) );
  XNOR2_X1 U18278 ( .A(n17446), .B(n17445), .ZN(n17447) );
  XNOR2_X1 U18279 ( .A(n17448), .B(n17447), .ZN(n18129) );
  AND2_X1 U18280 ( .A1(n17769), .A2(n18273), .ZN(n18032) );
  OAI21_X1 U18281 ( .B1(n17768), .B2(n18032), .A(n18269), .ZN(n17453) );
  INV_X1 U18282 ( .A(n17769), .ZN(n18267) );
  OAI21_X1 U18283 ( .B1(n18267), .B2(n18275), .A(n18273), .ZN(n17451) );
  INV_X1 U18284 ( .A(n18270), .ZN(n17766) );
  NAND2_X1 U18285 ( .A1(n17451), .A2(n17766), .ZN(n17452) );
  OAI21_X1 U18286 ( .B1(n18698), .B2(n17463), .A(n18706), .ZN(n17465) );
  AOI21_X1 U18288 ( .B1(n396), .B2(n18238), .A(n18240), .ZN(n17454) );
  NAND2_X1 U18289 ( .A1(n17982), .A2(n17981), .ZN(n18037) );
  MUX2_X1 U18290 ( .A(n17753), .B(n17454), .S(n18037), .Z(n17457) );
  INV_X1 U18291 ( .A(n18240), .ZN(n17455) );
  NOR3_X1 U18293 ( .A1(n17455), .A2(n19919), .A3(n17753), .ZN(n17456) );
  NOR2_X2 U18294 ( .A1(n17457), .A2(n17456), .ZN(n18072) );
  INV_X1 U18295 ( .A(n19885), .ZN(n18113) );
  INV_X1 U18296 ( .A(n17458), .ZN(n18115) );
  OAI21_X1 U18297 ( .B1(n18111), .B2(n18112), .A(n20349), .ZN(n17459) );
  NAND2_X1 U18298 ( .A1(n17460), .A2(n17459), .ZN(n17461) );
  OAI21_X1 U18299 ( .B1(n20114), .B2(n18113), .A(n17461), .ZN(n18701) );
  OAI21_X1 U18300 ( .B1(n18072), .B2(n18702), .A(n18701), .ZN(n17464) );
  AOI22_X1 U18301 ( .A1(n17465), .A2(n18072), .B1(n17464), .B2(n17463), .ZN(
        n17467) );
  XNOR2_X1 U18302 ( .A(n17467), .B(n17466), .ZN(Ciphertext[72]) );
  INV_X1 U18303 ( .A(n17564), .ZN(n17469) );
  MUX2_X1 U18304 ( .A(n17469), .B(n17468), .S(n17470), .Z(n17474) );
  NAND2_X1 U18305 ( .A1(n18539), .A2(n17565), .ZN(n17472) );
  OR2_X1 U18306 ( .A1(n17564), .A2(n17470), .ZN(n17561) );
  MUX2_X1 U18307 ( .A(n17472), .B(n17561), .S(n17471), .Z(n17473) );
  NOR2_X1 U18309 ( .A1(n18093), .A2(n226), .ZN(n17572) );
  NOR2_X1 U18310 ( .A1(n20109), .A2(n18096), .ZN(n17570) );
  OAI21_X1 U18311 ( .B1(n17572), .B2(n17570), .A(n18101), .ZN(n17478) );
  AOI21_X1 U18312 ( .B1(n18095), .B2(n18097), .A(n18096), .ZN(n17476) );
  NOR2_X1 U18314 ( .A1(n18511), .A2(n18518), .ZN(n17519) );
  NOR2_X1 U18315 ( .A1(n17482), .A2(n17481), .ZN(n17486) );
  NAND2_X1 U18316 ( .A1(n18184), .A2(n18504), .ZN(n17524) );
  OAI211_X1 U18317 ( .C1(n17505), .C2(n17504), .A(n17503), .B(n17502), .ZN(
        n17506) );
  NAND2_X1 U18319 ( .A1(n19758), .A2(n19526), .ZN(n17518) );
  OAI21_X1 U18320 ( .B1(n19956), .B2(n17508), .A(n17507), .ZN(n17516) );
  OAI21_X1 U18321 ( .B1(n19700), .B2(n17510), .A(n17509), .ZN(n17515) );
  NOR2_X1 U18322 ( .A1(n17513), .A2(n17512), .ZN(n17514) );
  NAND2_X1 U18323 ( .A1(n18519), .A2(n18512), .ZN(n17517) );
  INV_X1 U18324 ( .A(n2307), .ZN(n17522) );
  NAND3_X1 U18325 ( .A1(n17581), .A2(n2307), .A3(n18505), .ZN(n17527) );
  INV_X1 U18326 ( .A(n17519), .ZN(n17521) );
  INV_X1 U18327 ( .A(n17524), .ZN(n17520) );
  NAND3_X1 U18328 ( .A1(n17521), .A2(n17520), .A3(n2307), .ZN(n17526) );
  INV_X1 U18329 ( .A(n18505), .ZN(n17523) );
  NAND3_X1 U18330 ( .A1(n17524), .A2(n17523), .A3(n17522), .ZN(n17525) );
  AND4_X1 U18331 ( .A1(n17528), .A2(n17527), .A3(n17526), .A4(n17525), .ZN(
        Ciphertext[31]) );
  INV_X1 U18332 ( .A(n19092), .ZN(n19109) );
  INV_X1 U18335 ( .A(n19111), .ZN(n17530) );
  NAND2_X1 U18336 ( .A1(n19106), .A2(n19110), .ZN(n17529) );
  NAND2_X1 U18338 ( .A1(n19098), .A2(n17203), .ZN(n17531) );
  AOI21_X1 U18339 ( .B1(n17532), .B2(n17531), .A(n19105), .ZN(n17533) );
  AND4_X1 U18340 ( .A1(n17538), .A2(n17537), .A3(n17536), .A4(n17610), .ZN(
        n17540) );
  NAND3_X1 U18341 ( .A1(n17540), .A2(n17539), .A3(n19955), .ZN(n17541) );
  INV_X1 U18342 ( .A(n19339), .ZN(n19308) );
  NAND2_X1 U18343 ( .A1(n19308), .A2(n19340), .ZN(n17543) );
  NOR2_X1 U18344 ( .A1(n19338), .A2(n19339), .ZN(n19316) );
  INV_X1 U18345 ( .A(n17545), .ZN(n17546) );
  NOR2_X1 U18346 ( .A1(n17546), .A2(n3066), .ZN(n17548) );
  NOR3_X1 U18347 ( .A1(n17549), .A2(n17390), .A3(n19876), .ZN(n17550) );
  MUX2_X1 U18349 ( .A(n18103), .B(n18105), .S(n18107), .Z(n17555) );
  INV_X1 U18350 ( .A(n17957), .ZN(n18106) );
  MUX2_X1 U18351 ( .A(n17553), .B(n17552), .S(n18107), .Z(n17554) );
  OAI21_X1 U18354 ( .B1(n20101), .B2(n19744), .A(n17556), .ZN(n18249) );
  NAND2_X1 U18356 ( .A1(n18249), .A2(n19678), .ZN(n17557) );
  OR2_X1 U18357 ( .A1(n19673), .A2(n19679), .ZN(n17578) );
  NOR2_X1 U18358 ( .A1(n20488), .A2(n20348), .ZN(n17965) );
  INV_X1 U18359 ( .A(n17965), .ZN(n18213) );
  INV_X1 U18360 ( .A(n20349), .ZN(n18633) );
  NAND3_X1 U18361 ( .A1(n19885), .A2(n17559), .A3(n18633), .ZN(n18211) );
  OAI21_X1 U18362 ( .B1(n17565), .B2(n20432), .A(n17564), .ZN(n17566) );
  OAI21_X1 U18363 ( .B1(n18538), .B2(n17564), .A(n17566), .ZN(n17567) );
  OAI22_X1 U18364 ( .A1(n17569), .A2(n18096), .B1(n18095), .B2(n18097), .ZN(
        n17573) );
  OR3_X1 U18365 ( .A1(n17570), .A2(n18101), .A3(n160), .ZN(n17571) );
  NAND2_X1 U18367 ( .A1(n18600), .A2(n19757), .ZN(n17574) );
  OAI21_X1 U18368 ( .B1(n18625), .B2(n18600), .A(n17574), .ZN(n17575) );
  NAND2_X1 U18369 ( .A1(n17575), .A2(n19673), .ZN(n17577) );
  OAI211_X1 U18370 ( .C1(n18630), .C2(n17578), .A(n17577), .B(n17576), .ZN(
        n17580) );
  INV_X1 U18371 ( .A(n2087), .ZN(n17579) );
  XNOR2_X1 U18372 ( .A(n17580), .B(n17579), .ZN(Ciphertext[58]) );
  OAI21_X1 U18373 ( .B1(n18504), .B2(n18184), .A(n18512), .ZN(n17582) );
  XNOR2_X1 U18374 ( .A(n17583), .B(n538), .ZN(Ciphertext[35]) );
  AOI22_X1 U18377 ( .A1(n17927), .A2(n19668), .B1(n19690), .B2(n19655), .ZN(
        n17585) );
  NAND2_X1 U18378 ( .A1(n17586), .A2(n17585), .ZN(n17589) );
  INV_X1 U18379 ( .A(n17587), .ZN(n17588) );
  XNOR2_X1 U18380 ( .A(n17589), .B(n17588), .ZN(Ciphertext[36]) );
  INV_X1 U18381 ( .A(n17861), .ZN(n17864) );
  AND2_X1 U18382 ( .A1(n19360), .A2(n20212), .ZN(n17590) );
  OAI21_X1 U18383 ( .B1(n17591), .B2(n17590), .A(n17864), .ZN(n17594) );
  OAI21_X1 U18385 ( .B1(n17596), .B2(n19372), .A(n19733), .ZN(n17597) );
  NOR2_X1 U18387 ( .A1(n17600), .A2(n17599), .ZN(n17605) );
  OAI21_X1 U18388 ( .B1(n17601), .B2(n17602), .A(n17890), .ZN(n17604) );
  AND2_X1 U18389 ( .A1(n19947), .A2(n17602), .ZN(n17603) );
  OAI21_X1 U18390 ( .B1(n20364), .B2(n19292), .A(n19298), .ZN(n17617) );
  MUX2_X1 U18391 ( .A(n19402), .B(n17606), .S(n19401), .Z(n17609) );
  MUX2_X1 U18393 ( .A(n17649), .B(n17607), .S(n19401), .Z(n17608) );
  NOR2_X1 U18395 ( .A1(n20515), .A2(n19284), .ZN(n17616) );
  INV_X1 U18396 ( .A(n17610), .ZN(n17614) );
  INV_X1 U18397 ( .A(n17881), .ZN(n17613) );
  OAI211_X1 U18398 ( .C1(n17881), .C2(n196), .A(n19930), .B(n3345), .ZN(n17612) );
  OAI21_X1 U18399 ( .B1(n17613), .B2(n19832), .A(n17878), .ZN(n17611) );
  INV_X1 U18400 ( .A(n17656), .ZN(n19395) );
  AND2_X1 U18402 ( .A1(n17654), .A2(n20172), .ZN(n17618) );
  INV_X1 U18403 ( .A(n19388), .ZN(n19400) );
  AND3_X1 U18404 ( .A1(n19390), .A2(n19396), .A3(n20004), .ZN(n19282) );
  NOR3_X1 U18405 ( .A1(n19304), .A2(n19292), .A3(n20515), .ZN(n17620) );
  NOR2_X1 U18406 ( .A1(n17621), .A2(n17620), .ZN(n17622) );
  XNOR2_X1 U18407 ( .A(n17622), .B(n345), .ZN(Ciphertext[172]) );
  INV_X1 U18408 ( .A(n18589), .ZN(n17624) );
  NAND3_X1 U18409 ( .A1(n20445), .A2(n19656), .A3(n19669), .ZN(n17625) );
  OAI211_X1 U18410 ( .C1(n18597), .C2(n17627), .A(n17626), .B(n17625), .ZN(
        n17629) );
  INV_X1 U18411 ( .A(n2392), .ZN(n17628) );
  XNOR2_X1 U18412 ( .A(n17629), .B(n17628), .ZN(Ciphertext[52]) );
  NOR2_X1 U18413 ( .A1(n17630), .A2(n18701), .ZN(n17633) );
  NOR2_X1 U18414 ( .A1(n17633), .A2(n17632), .ZN(n17634) );
  XNOR2_X1 U18415 ( .A(n17634), .B(n2317), .ZN(Ciphertext[76]) );
  OAI22_X1 U18416 ( .A1(n19682), .A2(n19691), .B1(n17925), .B2(n19661), .ZN(
        n18531) );
  OAI21_X1 U18417 ( .B1(n17923), .B2(n19661), .A(n19690), .ZN(n17635) );
  AOI22_X1 U18418 ( .A1(n18531), .A2(n19668), .B1(n17635), .B2(n18546), .ZN(
        n17638) );
  XNOR2_X1 U18419 ( .A(n17638), .B(n17637), .ZN(Ciphertext[41]) );
  NAND2_X1 U18420 ( .A1(n18495), .A2(n18497), .ZN(n17914) );
  NAND2_X1 U18421 ( .A1(n18500), .A2(n17914), .ZN(n17642) );
  AOI21_X1 U18422 ( .B1(n18496), .B2(n18498), .A(n645), .ZN(n17641) );
  OAI21_X1 U18423 ( .B1(n17914), .B2(n893), .A(n645), .ZN(n17643) );
  INV_X1 U18424 ( .A(n17643), .ZN(n17646) );
  NAND2_X1 U18425 ( .A1(n18489), .A2(n18495), .ZN(n17645) );
  OAI21_X1 U18426 ( .B1(n17649), .B2(n17650), .A(n17648), .ZN(n17653) );
  MUX2_X1 U18427 ( .A(n19404), .B(n17650), .S(n17853), .Z(n17651) );
  NOR2_X1 U18428 ( .A1(n19402), .A2(n17651), .ZN(n17652) );
  NOR2_X2 U18429 ( .A1(n17653), .A2(n17652), .ZN(n19269) );
  NAND2_X1 U18431 ( .A1(n19947), .A2(n20185), .ZN(n17661) );
  NAND2_X1 U18432 ( .A1(n16261), .A2(n17663), .ZN(n17664) );
  NOR2_X1 U18433 ( .A1(n17666), .A2(n17876), .ZN(n17883) );
  NAND2_X1 U18434 ( .A1(n17883), .A2(n20162), .ZN(n19251) );
  NAND2_X1 U18435 ( .A1(n17667), .A2(n19251), .ZN(n17669) );
  NOR3_X1 U18436 ( .A1(n17879), .A2(n17668), .A3(n3345), .ZN(n19249) );
  INV_X1 U18438 ( .A(n19276), .ZN(n19271) );
  NOR2_X1 U18439 ( .A1(n19276), .A2(n19246), .ZN(n19263) );
  NOR2_X1 U18440 ( .A1(n20242), .A2(n19938), .ZN(n17670) );
  NOR2_X1 U18441 ( .A1(n17673), .A2(n17864), .ZN(n17674) );
  INV_X1 U18442 ( .A(n19278), .ZN(n19247) );
  NAND2_X1 U18443 ( .A1(n19263), .A2(n19247), .ZN(n17681) );
  AND2_X1 U18444 ( .A1(n19246), .A2(n19269), .ZN(n17685) );
  AOI22_X1 U18445 ( .A1(n1112), .A2(n20275), .B1(n20507), .B2(n20512), .ZN(
        n17679) );
  OAI21_X1 U18446 ( .B1(n17677), .B2(n17867), .A(n17676), .ZN(n17678) );
  NAND2_X1 U18447 ( .A1(n17685), .A2(n20448), .ZN(n17680) );
  OAI211_X1 U18448 ( .C1(n17682), .C2(n19271), .A(n17681), .B(n17680), .ZN(
        n17684) );
  XNOR2_X1 U18449 ( .A(n17684), .B(n17683), .ZN(Ciphertext[165]) );
  NAND2_X1 U18450 ( .A1(n19278), .A2(n19246), .ZN(n19261) );
  AND2_X1 U18451 ( .A1(n18042), .A2(n18946), .ZN(n17691) );
  NAND2_X1 U18452 ( .A1(n18047), .A2(n17687), .ZN(n17688) );
  INV_X1 U18453 ( .A(n19034), .ZN(n18061) );
  NOR2_X1 U18454 ( .A1(n18961), .A2(n17818), .ZN(n17694) );
  NOR2_X1 U18455 ( .A1(n18968), .A2(n17692), .ZN(n17693) );
  OR2_X1 U18456 ( .A1(n18968), .A2(n17695), .ZN(n17696) );
  AOI21_X1 U18457 ( .B1(n17817), .B2(n17696), .A(n227), .ZN(n17697) );
  AND2_X1 U18460 ( .A1(n18927), .A2(n18928), .ZN(n18028) );
  NAND2_X1 U18461 ( .A1(n18028), .A2(n18025), .ZN(n17703) );
  NAND2_X1 U18462 ( .A1(n17700), .A2(n18024), .ZN(n17701) );
  MUX2_X1 U18463 ( .A(n17701), .B(n18029), .S(n18025), .Z(n17702) );
  NAND2_X1 U18464 ( .A1(n18081), .A2(n19046), .ZN(n17724) );
  MUX2_X1 U18465 ( .A(n18020), .B(n889), .S(n19723), .Z(n17709) );
  NOR2_X1 U18466 ( .A1(n17707), .A2(n17706), .ZN(n17708) );
  NAND2_X1 U18467 ( .A1(n18954), .A2(n18955), .ZN(n17710) );
  OAI21_X1 U18468 ( .B1(n18959), .B2(n18955), .A(n17710), .ZN(n17713) );
  INV_X1 U18471 ( .A(n20264), .ZN(n17719) );
  OAI22_X1 U18472 ( .A1(n16731), .A2(n17719), .B1(n17714), .B2(n20423), .ZN(
        n17717) );
  INV_X1 U18473 ( .A(n17715), .ZN(n17716) );
  NAND2_X1 U18474 ( .A1(n17717), .A2(n17716), .ZN(n17722) );
  NAND2_X1 U18475 ( .A1(n17063), .A2(n16731), .ZN(n17721) );
  NAND2_X1 U18477 ( .A1(n19046), .A2(n19034), .ZN(n17723) );
  OAI21_X1 U18478 ( .B1(n20475), .B2(n19047), .A(n17723), .ZN(n18062) );
  AOI22_X1 U18479 ( .A1(n17724), .A2(n19047), .B1(n18062), .B2(n19043), .ZN(
        n17725) );
  XNOR2_X1 U18480 ( .A(n17725), .B(n642), .ZN(Ciphertext[119]) );
  NAND2_X1 U18481 ( .A1(n18453), .A2(n18468), .ZN(n17726) );
  OAI21_X1 U18485 ( .B1(n19791), .B2(n20231), .A(n18468), .ZN(n17727) );
  AOI22_X1 U18486 ( .A1(n18429), .A2(n18464), .B1(n20110), .B2(n17727), .ZN(
        n17728) );
  XNOR2_X1 U18487 ( .A(n17728), .B(n20593), .ZN(Ciphertext[23]) );
  NAND2_X1 U18488 ( .A1(n18485), .A2(n17733), .ZN(n17736) );
  NAND2_X1 U18491 ( .A1(n17731), .A2(n19816), .ZN(n17732) );
  OAI211_X1 U18492 ( .C1(n18500), .C2(n17640), .A(n17736), .B(n17732), .ZN(
        n17743) );
  XNOR2_X1 U18493 ( .A(n18498), .B(n17733), .ZN(n17734) );
  AOI21_X1 U18494 ( .B1(n17734), .B2(n17640), .A(n19816), .ZN(n17742) );
  NOR2_X1 U18495 ( .A1(n17736), .A2(n17735), .ZN(n17738) );
  NAND2_X1 U18496 ( .A1(n17738), .A2(n17739), .ZN(n17741) );
  NAND2_X1 U18499 ( .A1(n20158), .A2(n18976), .ZN(n17746) );
  OR2_X1 U18500 ( .A1(n18016), .A2(n18977), .ZN(n17745) );
  MUX2_X1 U18501 ( .A(n17746), .B(n17745), .S(n18221), .Z(n17747) );
  INV_X1 U18502 ( .A(n18807), .ZN(n18332) );
  AOI22_X1 U18503 ( .A1(n18931), .A2(n18025), .B1(n18927), .B2(n18926), .ZN(
        n17750) );
  OR2_X1 U18504 ( .A1(n18240), .A2(n19919), .ZN(n17757) );
  INV_X1 U18505 ( .A(n18237), .ZN(n17756) );
  NAND3_X1 U18507 ( .A1(n20258), .A2(n17753), .A3(n17981), .ZN(n17755) );
  INV_X1 U18508 ( .A(n18238), .ZN(n17751) );
  NAND2_X1 U18509 ( .A1(n3205), .A2(n17751), .ZN(n17752) );
  OAI211_X1 U18510 ( .C1(n17753), .C2(n18240), .A(n17982), .B(n17752), .ZN(
        n17754) );
  NAND2_X1 U18512 ( .A1(n18795), .A2(n19770), .ZN(n18335) );
  INV_X1 U18513 ( .A(n17758), .ZN(n18256) );
  NAND2_X1 U18514 ( .A1(n18256), .A2(n18138), .ZN(n17759) );
  NAND2_X1 U18515 ( .A1(n17759), .A2(n18257), .ZN(n17761) );
  NAND2_X1 U18516 ( .A1(n18754), .A2(n18256), .ZN(n17760) );
  MUX2_X1 U18517 ( .A(n17761), .B(n17760), .S(n18260), .Z(n17763) );
  NAND2_X1 U18518 ( .A1(n17763), .A2(n17762), .ZN(n17772) );
  INV_X1 U18520 ( .A(n18806), .ZN(n18800) );
  OAI21_X1 U18521 ( .B1(n18795), .B2(n19811), .A(n18800), .ZN(n17773) );
  NAND2_X1 U18522 ( .A1(n18267), .A2(n18270), .ZN(n17765) );
  MUX2_X1 U18523 ( .A(n17765), .B(n17764), .S(n18275), .Z(n17771) );
  AND2_X1 U18524 ( .A1(n18033), .A2(n18269), .ZN(n17767) );
  AOI22_X1 U18525 ( .A1(n17769), .A2(n17768), .B1(n17767), .B2(n17766), .ZN(
        n17770) );
  NOR2_X1 U18526 ( .A1(n18794), .A2(n17772), .ZN(n18333) );
  INV_X1 U18527 ( .A(n17774), .ZN(n18128) );
  AND2_X1 U18528 ( .A1(n17946), .A2(n18130), .ZN(n17776) );
  AOI21_X1 U18529 ( .B1(n18248), .B2(n18129), .A(n17776), .ZN(n17780) );
  NOR2_X1 U18530 ( .A1(n17946), .A2(n17777), .ZN(n17778) );
  NAND2_X1 U18531 ( .A1(n18129), .A2(n17778), .ZN(n17779) );
  INV_X1 U18532 ( .A(n18803), .ZN(n18331) );
  INV_X1 U18533 ( .A(n18794), .ZN(n17781) );
  NAND3_X1 U18534 ( .A1(n213), .A2(n18331), .A3(n17781), .ZN(n17782) );
  INV_X1 U18535 ( .A(n2329), .ZN(n17783) );
  NAND2_X1 U18536 ( .A1(n19302), .A2(n19292), .ZN(n19290) );
  OR2_X1 U18537 ( .A1(n19284), .A2(n19292), .ZN(n18164) );
  MUX2_X1 U18538 ( .A(n19770), .B(n19711), .S(n18807), .Z(n17786) );
  NOR2_X1 U18539 ( .A1(n19811), .A2(n18807), .ZN(n17784) );
  MUX2_X1 U18540 ( .A(n17784), .B(n18803), .S(n19711), .Z(n17785) );
  AOI21_X1 U18541 ( .B1(n18795), .B2(n17786), .A(n17785), .ZN(n17788) );
  XNOR2_X1 U18542 ( .A(n17788), .B(n17787), .ZN(Ciphertext[84]) );
  OAI22_X1 U18545 ( .A1(n17789), .A2(n17794), .B1(n2896), .B2(n17793), .ZN(
        n17795) );
  NOR3_X1 U18546 ( .A1(n17797), .A2(n17796), .A3(n17795), .ZN(Ciphertext[139])
         );
  NAND2_X1 U18547 ( .A1(n18697), .A2(n19753), .ZN(n17799) );
  OAI21_X1 U18548 ( .B1(n18698), .B2(n18701), .A(n17799), .ZN(n18695) );
  INV_X1 U18549 ( .A(n18072), .ZN(n17803) );
  INV_X1 U18550 ( .A(n18701), .ZN(n17800) );
  OAI21_X1 U18551 ( .B1(n18698), .B2(n19751), .A(n17800), .ZN(n17802) );
  AOI22_X1 U18552 ( .A1(n18695), .A2(n17803), .B1(n17802), .B2(n1055), .ZN(
        n17805) );
  XNOR2_X1 U18553 ( .A(n17805), .B(n17804), .ZN(Ciphertext[77]) );
  INV_X1 U18554 ( .A(n19143), .ZN(n19133) );
  AND2_X1 U18556 ( .A1(n20508), .A2(n19144), .ZN(n19127) );
  NAND2_X1 U18557 ( .A1(n19127), .A2(n19134), .ZN(n17809) );
  INV_X1 U18558 ( .A(n19146), .ZN(n19125) );
  NAND2_X1 U18559 ( .A1(n17807), .A2(n19125), .ZN(n17808) );
  OAI211_X1 U18560 ( .C1(n17810), .C2(n19144), .A(n17809), .B(n17808), .ZN(
        n17811) );
  XNOR2_X1 U18561 ( .A(n17811), .B(n2079), .ZN(Ciphertext[134]) );
  AND2_X1 U18562 ( .A1(n18046), .A2(n17812), .ZN(n18045) );
  INV_X1 U18563 ( .A(n18045), .ZN(n17816) );
  NAND3_X1 U18564 ( .A1(n20194), .A2(n17687), .A3(n17812), .ZN(n17815) );
  NAND4_X1 U18565 ( .A1(n17816), .A2(n17815), .A3(n17814), .A4(n17813), .ZN(
        n19059) );
  NAND2_X1 U18566 ( .A1(n17819), .A2(n18961), .ZN(n18965) );
  MUX2_X1 U18567 ( .A(n19059), .B(n19685), .S(n19060), .Z(n17850) );
  OR2_X1 U18568 ( .A1(n17836), .A2(n16731), .ZN(n17839) );
  OAI211_X1 U18569 ( .C1(n17715), .C2(n17838), .A(n17063), .B(n17839), .ZN(
        n17843) );
  INV_X1 U18570 ( .A(n17839), .ZN(n17841) );
  NAND2_X1 U18571 ( .A1(n17841), .A2(n17840), .ZN(n17842) );
  AND2_X1 U18572 ( .A1(n19060), .A2(n19067), .ZN(n19064) );
  NOR2_X1 U18573 ( .A1(n20452), .A2(n18935), .ZN(n17847) );
  OR2_X1 U18574 ( .A1(n18939), .A2(n18936), .ZN(n17845) );
  MUX2_X1 U18575 ( .A(n17845), .B(n20501), .S(n17187), .Z(n17846) );
  OAI21_X2 U18576 ( .B1(n18933), .B2(n17847), .A(n17846), .ZN(n19073) );
  NOR2_X1 U18577 ( .A1(n19060), .A2(n19073), .ZN(n17848) );
  AOI22_X1 U18578 ( .A1(n19064), .A2(n19685), .B1(n17848), .B2(n20131), .ZN(
        n17849) );
  OAI21_X1 U18579 ( .B1(n17850), .B2(n20131), .A(n17849), .ZN(n17852) );
  XNOR2_X1 U18580 ( .A(n17852), .B(n17851), .ZN(Ciphertext[122]) );
  MUX2_X1 U18581 ( .A(n19401), .B(n19402), .S(n19404), .Z(n17856) );
  INV_X1 U18582 ( .A(n19402), .ZN(n17854) );
  NOR2_X1 U18583 ( .A1(n17854), .A2(n17853), .ZN(n17855) );
  INV_X1 U18584 ( .A(n19403), .ZN(n17857) );
  NOR3_X1 U18585 ( .A1(n19401), .A2(n17857), .A3(n19402), .ZN(n17858) );
  OAI21_X1 U18586 ( .B1(n20150), .B2(n17861), .A(n17860), .ZN(n19366) );
  AOI21_X1 U18587 ( .B1(n17863), .B2(n20212), .A(n20242), .ZN(n17865) );
  OR2_X1 U18588 ( .A1(n17865), .A2(n17864), .ZN(n17866) );
  NAND2_X1 U18589 ( .A1(n19242), .A2(n20124), .ZN(n17904) );
  NAND2_X1 U18590 ( .A1(n20275), .A2(n17867), .ZN(n17869) );
  MUX2_X1 U18591 ( .A(n20507), .B(n17869), .S(n17868), .Z(n17875) );
  OAI211_X1 U18592 ( .C1(n20512), .C2(n17873), .A(n19973), .B(n1112), .ZN(
        n17874) );
  NAND2_X1 U18593 ( .A1(n17875), .A2(n17874), .ZN(n19235) );
  AND2_X1 U18595 ( .A1(n19754), .A2(n19227), .ZN(n17903) );
  AND2_X1 U18596 ( .A1(n17890), .A2(n17886), .ZN(n17888) );
  INV_X1 U18597 ( .A(n19233), .ZN(n19236) );
  AND2_X1 U18598 ( .A1(n17892), .A2(n17893), .ZN(n17902) );
  AOI21_X1 U18599 ( .B1(n17894), .B2(n17898), .A(n17893), .ZN(n17901) );
  NOR2_X1 U18600 ( .A1(n17895), .A2(n17897), .ZN(n17899) );
  INV_X1 U18601 ( .A(n19237), .ZN(n18190) );
  XNOR2_X1 U18602 ( .A(n17905), .B(n1857), .ZN(Ciphertext[157]) );
  BUF_X1 U18603 ( .A(n18287), .Z(n17936) );
  MUX2_X1 U18604 ( .A(n18357), .B(n17907), .S(n18362), .Z(n17908) );
  XNOR2_X1 U18605 ( .A(n17910), .B(n17909), .ZN(Ciphertext[1]) );
  NAND3_X1 U18606 ( .A1(n19729), .A2(n18497), .A3(n17640), .ZN(n17913) );
  INV_X1 U18607 ( .A(n19242), .ZN(n17916) );
  NAND2_X1 U18608 ( .A1(n19219), .A2(n20193), .ZN(n17915) );
  XNOR2_X1 U18609 ( .A(n17917), .B(Key[60]), .ZN(Ciphertext[161]) );
  NAND2_X1 U18610 ( .A1(n18590), .A2(n18589), .ZN(n18584) );
  NOR2_X1 U18611 ( .A1(n18589), .A2(n17918), .ZN(n18593) );
  OAI21_X1 U18612 ( .B1(n18573), .B2(n18584), .A(n17919), .ZN(n17921) );
  NOR2_X1 U18613 ( .A1(n18597), .A2(n20365), .ZN(n17920) );
  NOR2_X1 U18614 ( .A1(n17921), .A2(n17920), .ZN(n17922) );
  XNOR2_X1 U18615 ( .A(n17922), .B(n484), .ZN(Ciphertext[49]) );
  NAND3_X1 U18616 ( .A1(n17923), .A2(n19690), .A3(n19691), .ZN(n17930) );
  NAND3_X1 U18617 ( .A1(n17925), .A2(n19661), .A3(n19691), .ZN(n17929) );
  NAND4_X1 U18618 ( .A1(n17931), .A2(n17930), .A3(n17929), .A4(n17928), .ZN(
        n17934) );
  INV_X1 U18619 ( .A(n17932), .ZN(n17933) );
  XNOR2_X1 U18620 ( .A(n17934), .B(n17933), .ZN(Ciphertext[40]) );
  OAI21_X1 U18621 ( .B1(n18362), .B2(n18348), .A(n18290), .ZN(n17939) );
  INV_X1 U18622 ( .A(n17935), .ZN(n18350) );
  NAND2_X1 U18623 ( .A1(n17936), .A2(n18350), .ZN(n18364) );
  OAI211_X1 U18624 ( .C1(n18362), .C2(n18359), .A(n18364), .B(n18292), .ZN(
        n17938) );
  AOI22_X1 U18625 ( .A1(n17938), .A2(n17939), .B1(n17937), .B2(n18357), .ZN(
        n17941) );
  XNOR2_X1 U18626 ( .A(n17941), .B(n17940), .ZN(Ciphertext[2]) );
  NOR2_X1 U18627 ( .A1(n19093), .A2(n19109), .ZN(n17944) );
  OAI21_X1 U18628 ( .B1(n19095), .B2(n19112), .A(n19093), .ZN(n17943) );
  NAND2_X1 U18629 ( .A1(n19095), .A2(n19098), .ZN(n19089) );
  NAND2_X1 U18630 ( .A1(n18248), .A2(n19678), .ZN(n17953) );
  NOR2_X1 U18631 ( .A1(n19472), .A2(n18130), .ZN(n17945) );
  NOR2_X1 U18632 ( .A1(n18131), .A2(n17946), .ZN(n18251) );
  OR2_X1 U18635 ( .A1(n18251), .A2(n17950), .ZN(n17951) );
  OAI21_X1 U18637 ( .B1(n17956), .B2(n19672), .A(n17954), .ZN(n17958) );
  NAND2_X1 U18638 ( .A1(n17958), .A2(n17957), .ZN(n17963) );
  NAND3_X1 U18639 ( .A1(n17956), .A2(n17959), .A3(n18106), .ZN(n17962) );
  NAND3_X1 U18640 ( .A1(n17956), .A2(n18103), .A3(n18107), .ZN(n17961) );
  NAND2_X1 U18642 ( .A1(n17965), .A2(n18115), .ZN(n17971) );
  INV_X1 U18643 ( .A(n17966), .ZN(n17970) );
  NOR2_X1 U18644 ( .A1(n18112), .A2(n20349), .ZN(n17967) );
  OR2_X1 U18645 ( .A1(n17968), .A2(n17967), .ZN(n17969) );
  NAND2_X1 U18646 ( .A1(n18672), .A2(n18671), .ZN(n17972) );
  AOI21_X1 U18647 ( .B1(n17390), .B2(n19876), .A(n17973), .ZN(n17975) );
  NOR2_X1 U18648 ( .A1(n18229), .A2(n18233), .ZN(n18122) );
  NOR2_X1 U18649 ( .A1(n18122), .A2(n18120), .ZN(n17974) );
  MUX2_X1 U18650 ( .A(n18137), .B(n17976), .S(n18753), .Z(n17980) );
  NAND2_X1 U18651 ( .A1(n18262), .A2(n18256), .ZN(n18752) );
  AOI21_X1 U18652 ( .B1(n18258), .B2(n18260), .A(n17977), .ZN(n17979) );
  NOR2_X1 U18653 ( .A1(n18682), .A2(n19735), .ZN(n17986) );
  NAND2_X1 U18654 ( .A1(n17986), .A2(n17985), .ZN(n17987) );
  OAI21_X1 U18656 ( .B1(n17992), .B2(n20276), .A(n17991), .ZN(n18845) );
  NAND2_X1 U18657 ( .A1(n18818), .A2(n18172), .ZN(n18174) );
  AOI22_X1 U18658 ( .A1(n18845), .A2(n18817), .B1(n18811), .B2(n18174), .ZN(
        n17994) );
  XNOR2_X1 U18659 ( .A(n17994), .B(n17993), .ZN(Ciphertext[91]) );
  NAND2_X1 U18660 ( .A1(n19775), .A2(n18568), .ZN(n17996) );
  AOI21_X1 U18662 ( .B1(n17997), .B2(n17996), .A(n20169), .ZN(n17998) );
  XNOR2_X1 U18663 ( .A(n18000), .B(n17999), .ZN(Ciphertext[46]) );
  NAND2_X1 U18664 ( .A1(n18568), .A2(n18556), .ZN(n18560) );
  INV_X1 U18665 ( .A(n18559), .ZN(n18570) );
  NOR2_X1 U18666 ( .A1(n18199), .A2(n18559), .ZN(n18002) );
  INV_X1 U18667 ( .A(n18567), .ZN(n18001) );
  OAI21_X1 U18668 ( .B1(n18002), .B2(n18565), .A(n18001), .ZN(n18005) );
  OAI211_X1 U18669 ( .C1(n18560), .C2(n18570), .A(n18005), .B(n18004), .ZN(
        n18008) );
  INV_X1 U18670 ( .A(n18006), .ZN(n18007) );
  XNOR2_X1 U18671 ( .A(n18008), .B(n18007), .ZN(Ciphertext[42]) );
  MUX2_X1 U18672 ( .A(n20492), .B(n18522), .S(n18512), .Z(n18010) );
  INV_X1 U18673 ( .A(n18011), .ZN(n18012) );
  OAI21_X1 U18674 ( .B1(n19459), .B2(n19453), .A(n19460), .ZN(n18013) );
  AOI22_X1 U18675 ( .A1(n18014), .A2(n19459), .B1(n18013), .B2(n20152), .ZN(
        n18015) );
  XNOR2_X1 U18676 ( .A(n18015), .B(n2383), .ZN(Ciphertext[186]) );
  MUX2_X1 U18677 ( .A(n18016), .B(n20499), .S(n18221), .Z(n18018) );
  MUX2_X1 U18678 ( .A(n18975), .B(n18976), .S(n18978), .Z(n18017) );
  MUX2_X2 U18679 ( .A(n18018), .B(n18017), .S(n18977), .Z(n18869) );
  AOI22_X1 U18680 ( .A1(n18020), .A2(n18937), .B1(n20501), .B2(n19723), .ZN(
        n18023) );
  NAND3_X1 U18681 ( .A1(n18934), .A2(n18937), .A3(n18935), .ZN(n18022) );
  MUX2_X1 U18685 ( .A(n18270), .B(n18032), .S(n18268), .Z(n18036) );
  OAI211_X1 U18686 ( .C1(n18269), .C2(n18033), .A(n18275), .B(n18267), .ZN(
        n18034) );
  INV_X1 U18687 ( .A(n18034), .ZN(n18035) );
  MUX2_X1 U18688 ( .A(n19988), .B(n20418), .S(n18857), .Z(n18054) );
  NOR2_X1 U18689 ( .A1(n18240), .A2(n20132), .ZN(n18040) );
  NAND2_X1 U18690 ( .A1(n20258), .A2(n18038), .ZN(n18039) );
  INV_X1 U18692 ( .A(n18866), .ZN(n18850) );
  NOR2_X1 U18693 ( .A1(n20418), .A2(n18850), .ZN(n18052) );
  NOR2_X1 U18694 ( .A1(n18043), .A2(n18042), .ZN(n18044) );
  NAND2_X1 U18696 ( .A1(n18948), .A2(n2586), .ZN(n18048) );
  AOI21_X1 U18697 ( .B1(n18949), .B2(n18048), .A(n18047), .ZN(n18049) );
  INV_X1 U18701 ( .A(n19168), .ZN(n18323) );
  NAND2_X1 U18702 ( .A1(n18057), .A2(n18157), .ZN(n18058) );
  OAI21_X1 U18703 ( .B1(n20460), .B2(n18323), .A(n18058), .ZN(n18089) );
  AOI22_X1 U18704 ( .A1(n18089), .A2(n19170), .B1(n18323), .B2(n18059), .ZN(
        n18060) );
  XNOR2_X1 U18705 ( .A(n18060), .B(n2257), .ZN(Ciphertext[149]) );
  NOR2_X1 U18707 ( .A1(n20142), .A2(n19032), .ZN(n18064) );
  NAND2_X1 U18708 ( .A1(n19047), .A2(n19032), .ZN(n19031) );
  NAND2_X1 U18709 ( .A1(n18062), .A2(n19031), .ZN(n18063) );
  INV_X1 U18710 ( .A(n18065), .ZN(n18066) );
  MUX2_X1 U18711 ( .A(n19460), .B(n19463), .S(n20152), .Z(n18069) );
  MUX2_X1 U18712 ( .A(n19459), .B(n19462), .S(n20140), .Z(n18068) );
  XNOR2_X1 U18713 ( .A(n18071), .B(n18070), .ZN(Ciphertext[188]) );
  MUX2_X1 U18714 ( .A(n18072), .B(n19751), .S(n18697), .Z(n18074) );
  MUX2_X1 U18715 ( .A(n18698), .B(n18701), .S(n18703), .Z(n18073) );
  MUX2_X1 U18716 ( .A(n18074), .B(n18073), .S(n19753), .Z(n18076) );
  XNOR2_X1 U18717 ( .A(n18076), .B(n18075), .ZN(Ciphertext[74]) );
  NOR2_X1 U18719 ( .A1(n18392), .A2(n18384), .ZN(n18077) );
  NAND2_X1 U18721 ( .A1(n19992), .A2(n19046), .ZN(n18080) );
  NAND2_X1 U18722 ( .A1(n18081), .A2(n18080), .ZN(n18082) );
  MUX2_X1 U18723 ( .A(n18083), .B(n18082), .S(n19032), .Z(n18086) );
  INV_X1 U18724 ( .A(n18084), .ZN(n18085) );
  XNOR2_X1 U18725 ( .A(n18086), .B(n18085), .ZN(Ciphertext[116]) );
  INV_X1 U18726 ( .A(n18327), .ZN(n19174) );
  INV_X1 U18727 ( .A(n19169), .ZN(n18087) );
  AOI22_X1 U18728 ( .A1(n18089), .A2(n18088), .B1(n18161), .B2(n18087), .ZN(
        n18091) );
  XNOR2_X1 U18729 ( .A(n18091), .B(n18090), .ZN(Ciphertext[145]) );
  AOI22_X1 U18730 ( .A1(n18095), .A2(n18094), .B1(n19774), .B2(n160), .ZN(
        n18102) );
  INV_X1 U18731 ( .A(n18096), .ZN(n18098) );
  OAI21_X1 U18732 ( .B1(n18099), .B2(n18098), .A(n18097), .ZN(n18100) );
  INV_X1 U18734 ( .A(n18651), .ZN(n18119) );
  NAND2_X1 U18735 ( .A1(n19737), .A2(n18107), .ZN(n18104) );
  OAI211_X1 U18736 ( .C1(n19658), .C2(n18107), .A(n18106), .B(n18105), .ZN(
        n18109) );
  MUX2_X1 U18738 ( .A(n18113), .B(n18112), .S(n18111), .Z(n18636) );
  AND2_X1 U18739 ( .A1(n18115), .A2(n19885), .ZN(n18117) );
  MUX2_X2 U18740 ( .A(n18636), .B(n18634), .S(n20349), .Z(n18656) );
  AOI21_X1 U18742 ( .B1(n18119), .B2(n18648), .A(n19624), .ZN(n18145) );
  AOI22_X1 U18743 ( .A1(n18123), .A2(n3066), .B1(n18122), .B2(n18226), .ZN(
        n18124) );
  NAND2_X1 U18744 ( .A1(n18125), .A2(n18124), .ZN(n18644) );
  AND2_X1 U18745 ( .A1(n18644), .A2(n18651), .ZN(n18144) );
  INV_X1 U18746 ( .A(n18144), .ZN(n18641) );
  AOI21_X1 U18747 ( .B1(n18128), .B2(n18127), .A(n18126), .ZN(n18136) );
  NOR2_X1 U18748 ( .A1(n18129), .A2(n19472), .ZN(n18134) );
  NOR2_X1 U18749 ( .A1(n18131), .A2(n18130), .ZN(n18133) );
  MUX2_X1 U18750 ( .A(n18134), .B(n18133), .S(n20101), .Z(n18135) );
  NOR2_X1 U18752 ( .A1(n18656), .A2(n18650), .ZN(n18143) );
  AOI21_X1 U18753 ( .B1(n18137), .B2(n18754), .A(n18262), .ZN(n18142) );
  NAND2_X1 U18754 ( .A1(n18257), .A2(n18138), .ZN(n18139) );
  AOI21_X1 U18755 ( .B1(n18139), .B2(n18260), .A(n18258), .ZN(n18141) );
  INV_X1 U18756 ( .A(n19757), .ZN(n18626) );
  NAND3_X1 U18758 ( .A1(n18625), .A2(n19673), .A3(n18626), .ZN(n18147) );
  INV_X1 U18759 ( .A(n2221), .ZN(n18148) );
  NOR2_X1 U18760 ( .A1(n19685), .A2(n19073), .ZN(n18150) );
  INV_X1 U18761 ( .A(n19059), .ZN(n19075) );
  AND2_X1 U18762 ( .A1(n19075), .A2(n19060), .ZN(n18149) );
  INV_X1 U18763 ( .A(n19074), .ZN(n19058) );
  MUX2_X1 U18764 ( .A(n18150), .B(n18149), .S(n19058), .Z(n18154) );
  INV_X1 U18765 ( .A(n18151), .ZN(n19069) );
  NAND2_X1 U18767 ( .A1(n19079), .A2(n19073), .ZN(n18152) );
  OAI21_X1 U18768 ( .B1(n19055), .B2(n19067), .A(n18152), .ZN(n18153) );
  NOR2_X1 U18769 ( .A1(n18154), .A2(n18153), .ZN(n18155) );
  XNOR2_X1 U18770 ( .A(n18155), .B(n1869), .ZN(Ciphertext[123]) );
  OAI21_X1 U18771 ( .B1(n18156), .B2(n20460), .A(n18320), .ZN(n18160) );
  INV_X1 U18772 ( .A(n18157), .ZN(n18318) );
  OAI21_X1 U18773 ( .B1(n18318), .B2(n18319), .A(n18158), .ZN(n18159) );
  AOI22_X1 U18774 ( .A1(n18161), .A2(n18160), .B1(n18159), .B2(n18323), .ZN(
        n18162) );
  XNOR2_X1 U18775 ( .A(n18162), .B(n1840), .ZN(Ciphertext[148]) );
  NAND2_X1 U18776 ( .A1(n20434), .A2(n19284), .ZN(n18163) );
  OAI21_X1 U18777 ( .B1(n19298), .B2(n19284), .A(n18163), .ZN(n18165) );
  NAND2_X1 U18779 ( .A1(n18688), .A2(n19735), .ZN(n18679) );
  OAI21_X1 U18780 ( .B1(n18672), .B2(n18666), .A(n18679), .ZN(n18169) );
  OAI21_X1 U18782 ( .B1(n18682), .B2(n19510), .A(n18671), .ZN(n18168) );
  AOI22_X1 U18783 ( .A1(n18169), .A2(n18682), .B1(n18666), .B2(n18168), .ZN(
        n18171) );
  XNOR2_X1 U18784 ( .A(n18171), .B(n18170), .ZN(Ciphertext[66]) );
  OR2_X1 U18785 ( .A1(n18831), .A2(n18172), .ZN(n18827) );
  OAI22_X1 U18786 ( .A1(n18827), .A2(n18834), .B1(n18813), .B2(n20097), .ZN(
        n18176) );
  NAND2_X1 U18787 ( .A1(n20422), .A2(n19766), .ZN(n18841) );
  OAI21_X1 U18788 ( .B1(n20130), .B2(n20097), .A(n18841), .ZN(n18175) );
  OAI22_X1 U18789 ( .A1(n18176), .A2(n18175), .B1(n18813), .B2(n18174), .ZN(
        n18178) );
  XNOR2_X1 U18790 ( .A(n18178), .B(n18177), .ZN(Ciphertext[92]) );
  NAND2_X1 U18791 ( .A1(n18630), .A2(n18600), .ZN(n18181) );
  INV_X1 U18792 ( .A(n18625), .ZN(n18619) );
  AOI22_X1 U18795 ( .A1(n18181), .A2(n18180), .B1(n18179), .B2(n18630), .ZN(
        n18182) );
  XNOR2_X1 U18796 ( .A(n18182), .B(n2100), .ZN(Ciphertext[54]) );
  MUX2_X1 U18797 ( .A(n18522), .B(n18511), .S(n19773), .Z(n18186) );
  NAND2_X1 U18798 ( .A1(n18504), .A2(n18512), .ZN(n18183) );
  OAI21_X1 U18799 ( .B1(n18504), .B2(n18184), .A(n18183), .ZN(n18185) );
  MUX2_X1 U18800 ( .A(n18186), .B(n18185), .S(n19758), .Z(n18188) );
  INV_X1 U18801 ( .A(n2375), .ZN(n18187) );
  XNOR2_X1 U18802 ( .A(n18188), .B(n18187), .ZN(Ciphertext[32]) );
  INV_X1 U18803 ( .A(n19227), .ZN(n19239) );
  OAI21_X1 U18804 ( .B1(n19754), .B2(n19239), .A(n19229), .ZN(n18193) );
  NAND2_X1 U18805 ( .A1(n19242), .A2(n18190), .ZN(n18192) );
  NOR2_X1 U18806 ( .A1(n19237), .A2(n19238), .ZN(n19225) );
  NOR2_X1 U18807 ( .A1(n19225), .A2(n19227), .ZN(n18191) );
  AOI22_X1 U18808 ( .A1(n18193), .A2(n19242), .B1(n18192), .B2(n18191), .ZN(
        n18194) );
  XNOR2_X1 U18809 ( .A(n18194), .B(n2296), .ZN(Ciphertext[156]) );
  INV_X1 U18810 ( .A(n18644), .ZN(n18654) );
  INV_X1 U18811 ( .A(n18648), .ZN(n18642) );
  OAI21_X1 U18812 ( .B1(n18654), .B2(n18642), .A(n18651), .ZN(n18197) );
  NAND2_X1 U18813 ( .A1(n18648), .A2(n18651), .ZN(n18195) );
  OAI21_X1 U18814 ( .B1(n18656), .B2(n19935), .A(n18195), .ZN(n18647) );
  INV_X1 U18815 ( .A(n19745), .ZN(n18196) );
  AOI22_X1 U18816 ( .A1(n18197), .A2(n18656), .B1(n18647), .B2(n18196), .ZN(
        n18198) );
  XNOR2_X1 U18817 ( .A(n18198), .B(n2306), .ZN(Ciphertext[65]) );
  NAND2_X1 U18818 ( .A1(n18555), .A2(n18565), .ZN(n18200) );
  NAND2_X1 U18819 ( .A1(n18561), .A2(n18200), .ZN(n18571) );
  INV_X1 U18820 ( .A(n18555), .ZN(n18566) );
  AND2_X1 U18821 ( .A1(n19775), .A2(n18566), .ZN(n18202) );
  AOI22_X1 U18822 ( .A1(n18571), .A2(n18560), .B1(n18202), .B2(n18201), .ZN(
        n18204) );
  XNOR2_X1 U18823 ( .A(n18204), .B(n18203), .ZN(Ciphertext[43]) );
  OAI21_X1 U18824 ( .B1(n20142), .B2(n18061), .A(n19992), .ZN(n18205) );
  OAI21_X1 U18825 ( .B1(n19993), .B2(n19046), .A(n18205), .ZN(n18207) );
  NAND3_X1 U18826 ( .A1(n938), .A2(n20142), .A3(n19032), .ZN(n18206) );
  INV_X1 U18828 ( .A(n18208), .ZN(n18209) );
  INV_X1 U18831 ( .A(n18211), .ZN(n18212) );
  AOI21_X1 U18832 ( .B1(n18214), .B2(n18213), .A(n18212), .ZN(n18215) );
  AND2_X1 U18833 ( .A1(n18622), .A2(n19509), .ZN(n18218) );
  NAND2_X1 U18834 ( .A1(n18218), .A2(n18630), .ZN(n18217) );
  OAI21_X1 U18835 ( .B1(n18219), .B2(n18218), .A(n18217), .ZN(n18220) );
  XNOR2_X1 U18836 ( .A(n18220), .B(n2420), .ZN(Ciphertext[56]) );
  NOR2_X1 U18837 ( .A1(n20158), .A2(n18978), .ZN(n18225) );
  OAI21_X1 U18838 ( .B1(n18225), .B2(n18976), .A(n224), .ZN(n18722) );
  NAND2_X1 U18839 ( .A1(n18721), .A2(n18722), .ZN(n18709) );
  INV_X1 U18840 ( .A(n18709), .ZN(n18763) );
  NOR2_X1 U18841 ( .A1(n18232), .A2(n18226), .ZN(n18227) );
  NAND2_X1 U18842 ( .A1(n19876), .A2(n18227), .ZN(n18236) );
  INV_X1 U18843 ( .A(n18233), .ZN(n18228) );
  NAND3_X1 U18844 ( .A1(n18228), .A2(n17390), .A3(n3066), .ZN(n18231) );
  NAND2_X1 U18845 ( .A1(n18229), .A2(n18233), .ZN(n18230) );
  AND2_X1 U18846 ( .A1(n18231), .A2(n18230), .ZN(n18235) );
  NAND3_X1 U18847 ( .A1(n17549), .A2(n18233), .A3(n18232), .ZN(n18234) );
  INV_X1 U18848 ( .A(n18762), .ZN(n18772) );
  NAND3_X1 U18851 ( .A1(n20258), .A2(n396), .A3(n20132), .ZN(n18245) );
  INV_X1 U18854 ( .A(n18248), .ZN(n18250) );
  OAI21_X1 U18855 ( .B1(n19678), .B2(n19472), .A(n18251), .ZN(n18254) );
  OAI21_X1 U18856 ( .B1(n18762), .B2(n19803), .A(n18255), .ZN(n18266) );
  NAND2_X1 U18857 ( .A1(n18258), .A2(n18257), .ZN(n18259) );
  OAI211_X1 U18858 ( .C1(n18260), .C2(n19787), .A(n18259), .B(n18753), .ZN(
        n18261) );
  OAI21_X1 U18859 ( .B1(n18263), .B2(n18262), .A(n18261), .ZN(n18265) );
  NOR2_X1 U18860 ( .A1(n18752), .A2(n18264), .ZN(n18758) );
  NOR2_X2 U18861 ( .A1(n18265), .A2(n18758), .ZN(n18741) );
  INV_X1 U18862 ( .A(n18741), .ZN(n18783) );
  NAND2_X1 U18863 ( .A1(n18266), .A2(n18783), .ZN(n18277) );
  NAND2_X1 U18864 ( .A1(n221), .A2(n18267), .ZN(n18272) );
  NAND2_X1 U18865 ( .A1(n18269), .A2(n18268), .ZN(n18271) );
  MUX2_X1 U18866 ( .A(n18272), .B(n18271), .S(n18270), .Z(n18719) );
  OAI211_X1 U18867 ( .C1(n18275), .C2(n18033), .A(n18274), .B(n18273), .ZN(
        n18720) );
  NAND2_X1 U18868 ( .A1(n18719), .A2(n18720), .ZN(n18775) );
  AND2_X1 U18869 ( .A1(n18775), .A2(n18741), .ZN(n18782) );
  NAND2_X1 U18870 ( .A1(n18782), .A2(n18763), .ZN(n18276) );
  INV_X1 U18871 ( .A(n18278), .ZN(n18279) );
  MUX2_X1 U18872 ( .A(n18656), .B(n18651), .S(n19934), .Z(n18283) );
  NAND3_X1 U18873 ( .A1(n18644), .A2(n18642), .A3(n19934), .ZN(n18281) );
  OAI211_X1 U18874 ( .C1(n18283), .C2(n18644), .A(n18282), .B(n18281), .ZN(
        n18285) );
  XNOR2_X1 U18875 ( .A(n18285), .B(n18284), .ZN(Ciphertext[62]) );
  INV_X1 U18876 ( .A(n18286), .ZN(n18293) );
  OAI21_X1 U18877 ( .B1(n18289), .B2(n18288), .A(n18365), .ZN(n18291) );
  NAND2_X1 U18878 ( .A1(n18290), .A2(n18359), .ZN(n18360) );
  OAI211_X1 U18879 ( .C1(n18293), .C2(n18292), .A(n18291), .B(n18360), .ZN(
        n18295) );
  XNOR2_X1 U18880 ( .A(n18295), .B(n18294), .ZN(Ciphertext[0]) );
  INV_X1 U18881 ( .A(n19163), .ZN(n19154) );
  NOR2_X1 U18882 ( .A1(n19948), .A2(n19154), .ZN(n18296) );
  NOR2_X1 U18883 ( .A1(n18296), .A2(n19683), .ZN(n18303) );
  INV_X1 U18884 ( .A(n19165), .ZN(n18297) );
  NAND2_X1 U18885 ( .A1(n19948), .A2(n18297), .ZN(n18302) );
  INV_X1 U18886 ( .A(n19162), .ZN(n18298) );
  NAND2_X1 U18887 ( .A1(n18298), .A2(n19163), .ZN(n18300) );
  NAND3_X1 U18888 ( .A1(n19155), .A2(n19708), .A3(n18306), .ZN(n18299) );
  OAI21_X1 U18889 ( .B1(n19948), .B2(n18300), .A(n18299), .ZN(n18301) );
  AOI21_X1 U18890 ( .B1(n18303), .B2(n18302), .A(n18301), .ZN(n18305) );
  XNOR2_X1 U18891 ( .A(n18305), .B(n18304), .ZN(Ciphertext[141]) );
  NOR2_X1 U18892 ( .A1(n19708), .A2(n19692), .ZN(n18307) );
  NAND2_X1 U18893 ( .A1(n19340), .A2(n19339), .ZN(n19311) );
  INV_X1 U18894 ( .A(n19338), .ZN(n19309) );
  NAND2_X1 U18895 ( .A1(n19329), .A2(n19339), .ZN(n18309) );
  NAND3_X1 U18898 ( .A1(n19333), .A2(n19324), .A3(n19308), .ZN(n18314) );
  NAND3_X1 U18900 ( .A1(n16544), .A2(n19749), .A3(n19334), .ZN(n18313) );
  INV_X1 U18901 ( .A(n2323), .ZN(n18316) );
  NAND2_X1 U18902 ( .A1(n18318), .A2(n18317), .ZN(n19175) );
  NAND3_X1 U18903 ( .A1(n18324), .A2(n20460), .A3(n18323), .ZN(n18325) );
  OAI211_X1 U18904 ( .C1(n20460), .C2(n19175), .A(n18326), .B(n18325), .ZN(
        n18328) );
  XNOR2_X1 U18905 ( .A(n18328), .B(n2445), .ZN(Ciphertext[146]) );
  NAND2_X1 U18906 ( .A1(n18800), .A2(n18795), .ZN(n18329) );
  OAI21_X1 U18907 ( .B1(n18331), .B2(n19811), .A(n18329), .ZN(n18808) );
  AOI22_X1 U18908 ( .A1(n18808), .A2(n18335), .B1(n18334), .B2(n18333), .ZN(
        n18336) );
  XNOR2_X1 U18909 ( .A(n18336), .B(n2454), .ZN(Ciphertext[85]) );
  NOR2_X1 U18910 ( .A1(n19134), .A2(n870), .ZN(n19148) );
  INV_X1 U18911 ( .A(n18338), .ZN(n18339) );
  INV_X1 U18913 ( .A(n18341), .ZN(n18343) );
  NOR2_X1 U18914 ( .A1(n18343), .A2(n18342), .ZN(n18346) );
  INV_X1 U18915 ( .A(n18359), .ZN(n18345) );
  NAND4_X1 U18916 ( .A1(n20234), .A2(n18346), .A3(n18345), .A4(n18344), .ZN(
        n18353) );
  NAND2_X1 U18917 ( .A1(n17936), .A2(n18348), .ZN(n18351) );
  NAND3_X1 U18918 ( .A1(n18351), .A2(n18350), .A3(n18349), .ZN(n18352) );
  OAI211_X1 U18919 ( .C1(n18365), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        n18356) );
  XNOR2_X1 U18920 ( .A(n18356), .B(n18355), .ZN(Ciphertext[3]) );
  OAI21_X1 U18921 ( .B1(n18359), .B2(n18358), .A(n18357), .ZN(n18361) );
  INV_X1 U18924 ( .A(n18366), .ZN(n18367) );
  XNOR2_X1 U18925 ( .A(n18368), .B(n18367), .ZN(Ciphertext[4]) );
  NOR2_X1 U18926 ( .A1(n20361), .A2(n18382), .ZN(n18369) );
  OAI21_X1 U18927 ( .B1(n18392), .B2(n19763), .A(n19501), .ZN(n18371) );
  NAND2_X1 U18928 ( .A1(n18371), .A2(n20361), .ZN(n18372) );
  NAND2_X1 U18929 ( .A1(n18373), .A2(n18372), .ZN(n18375) );
  INV_X1 U18930 ( .A(n2413), .ZN(n18374) );
  XNOR2_X1 U18931 ( .A(n18375), .B(n18374), .ZN(Ciphertext[6]) );
  INV_X1 U18933 ( .A(n18392), .ZN(n18383) );
  OAI21_X1 U18934 ( .B1(n18383), .B2(n18384), .A(n18381), .ZN(n18378) );
  NOR2_X1 U18936 ( .A1(n20361), .A2(n18384), .ZN(n18385) );
  NAND2_X1 U18937 ( .A1(n18385), .A2(n20437), .ZN(n18386) );
  AOI21_X1 U18938 ( .B1(n20611), .B2(n20361), .A(n20437), .ZN(n18395) );
  OAI22_X1 U18939 ( .A1(n18395), .A2(n18394), .B1(n18393), .B2(n18392), .ZN(
        n18398) );
  INV_X1 U18940 ( .A(n18396), .ZN(n18397) );
  XNOR2_X1 U18941 ( .A(n18398), .B(n18397), .ZN(Ciphertext[11]) );
  NOR2_X1 U18942 ( .A1(n20003), .A2(n15529), .ZN(n18417) );
  NAND2_X1 U18943 ( .A1(n18417), .A2(n18407), .ZN(n18403) );
  NAND2_X1 U18945 ( .A1(n19702), .A2(n18423), .ZN(n18399) );
  INV_X1 U18947 ( .A(n2394), .ZN(n18405) );
  INV_X1 U18948 ( .A(n18423), .ZN(n18416) );
  INV_X1 U18949 ( .A(n2382), .ZN(n18410) );
  XNOR2_X1 U18950 ( .A(n18411), .B(n18410), .ZN(Ciphertext[13]) );
  AND2_X1 U18951 ( .A1(n18423), .A2(n18412), .ZN(n18413) );
  NOR2_X1 U18952 ( .A1(n18414), .A2(n18413), .ZN(n18419) );
  AOI22_X1 U18953 ( .A1(n18417), .A2(n18416), .B1(n18415), .B2(n18425), .ZN(
        n18418) );
  OAI21_X1 U18954 ( .B1(n18419), .B2(n18425), .A(n18418), .ZN(n18422) );
  INV_X1 U18955 ( .A(n18420), .ZN(n18421) );
  XNOR2_X1 U18956 ( .A(n18422), .B(n18421), .ZN(Ciphertext[16]) );
  NOR2_X1 U18957 ( .A1(n18424), .A2(n18423), .ZN(n18426) );
  INV_X1 U18958 ( .A(n2280), .ZN(n18428) );
  OAI211_X1 U18961 ( .C1(n18464), .C2(n18465), .A(n19791), .B(n20232), .ZN(
        n18430) );
  INV_X1 U18963 ( .A(n18433), .ZN(n18434) );
  XNOR2_X1 U18964 ( .A(n18435), .B(n18434), .ZN(Ciphertext[19]) );
  INV_X1 U18965 ( .A(n18464), .ZN(n18436) );
  NAND2_X1 U18966 ( .A1(n18469), .A2(n18453), .ZN(n18440) );
  OAI21_X1 U18967 ( .B1(n18442), .B2(n18436), .A(n18440), .ZN(n18451) );
  INV_X1 U18968 ( .A(n18441), .ZN(n18438) );
  NAND3_X1 U18969 ( .A1(n18465), .A2(n18466), .A3(n20148), .ZN(n18437) );
  OAI211_X1 U18970 ( .C1(n18438), .C2(n18466), .A(n18439), .B(n18437), .ZN(
        n18450) );
  OR2_X1 U18971 ( .A1(n18440), .A2(n18439), .ZN(n18449) );
  OAI21_X1 U18972 ( .B1(n20139), .B2(n18468), .A(n18443), .ZN(n18444) );
  NAND3_X1 U18973 ( .A1(n19825), .A2(n18446), .A3(n18445), .ZN(n18448) );
  OAI211_X1 U18974 ( .C1(n18451), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        Ciphertext[20]) );
  OAI21_X1 U18975 ( .B1(n18461), .B2(n18464), .A(n18465), .ZN(n18458) );
  NOR2_X1 U18976 ( .A1(n20110), .A2(n18453), .ZN(n18457) );
  OR3_X1 U18977 ( .A1(n20110), .A2(n20232), .A3(n18453), .ZN(n18456) );
  INV_X1 U18978 ( .A(n18468), .ZN(n18463) );
  NAND3_X1 U18979 ( .A1(n18466), .A2(n18463), .A3(n20139), .ZN(n18455) );
  OAI211_X1 U18980 ( .C1(n18458), .C2(n18457), .A(n18456), .B(n18455), .ZN(
        n18460) );
  INV_X1 U18981 ( .A(n347), .ZN(n18459) );
  XNOR2_X1 U18982 ( .A(n18460), .B(n18459), .ZN(Ciphertext[21]) );
  AOI21_X1 U18983 ( .B1(n18463), .B2(n19791), .A(n18461), .ZN(n18472) );
  AOI21_X1 U18984 ( .B1(n20139), .B2(n18464), .A(n20110), .ZN(n18471) );
  NAND2_X1 U18985 ( .A1(n18469), .A2(n20148), .ZN(n18470) );
  XNOR2_X1 U18986 ( .A(n18474), .B(n18473), .ZN(Ciphertext[22]) );
  NOR3_X1 U18987 ( .A1(n18485), .A2(n18500), .A3(n18478), .ZN(n18475) );
  OAI21_X1 U18988 ( .B1(n18497), .B2(n18498), .A(n18475), .ZN(n18477) );
  INV_X1 U18989 ( .A(n18478), .ZN(n18481) );
  NOR2_X1 U18990 ( .A1(n18498), .A2(n18481), .ZN(n18486) );
  NAND2_X1 U18991 ( .A1(n18486), .A2(n19816), .ZN(n18476) );
  NAND2_X1 U18992 ( .A1(n18477), .A2(n18476), .ZN(n18494) );
  NAND3_X1 U18993 ( .A1(n18500), .A2(n18478), .A3(n17640), .ZN(n18484) );
  OR2_X1 U18994 ( .A1(n18498), .A2(n18478), .ZN(n18487) );
  NAND3_X1 U18995 ( .A1(n18495), .A2(n18478), .A3(n18498), .ZN(n18479) );
  NAND2_X1 U18996 ( .A1(n18487), .A2(n18479), .ZN(n18480) );
  NAND2_X1 U18997 ( .A1(n18480), .A2(n893), .ZN(n18483) );
  NAND3_X1 U18998 ( .A1(n18496), .A2(n893), .A3(n18481), .ZN(n18482) );
  NAND3_X1 U18999 ( .A1(n18484), .A2(n18483), .A3(n18482), .ZN(n18493) );
  NAND3_X1 U19000 ( .A1(n18486), .A2(n18501), .A3(n893), .ZN(n18492) );
  INV_X1 U19001 ( .A(n18487), .ZN(n18488) );
  NAND3_X1 U19002 ( .A1(n19729), .A2(n19816), .A3(n18488), .ZN(n18491) );
  OAI211_X1 U19003 ( .C1(n18494), .C2(n18493), .A(n18492), .B(n18491), .ZN(
        Ciphertext[25]) );
  AOI22_X1 U19004 ( .A1(n18500), .A2(n17640), .B1(n18495), .B2(n18498), .ZN(
        n18502) );
  OAI21_X1 U19005 ( .B1(n214), .B2(n18517), .A(n18518), .ZN(n18528) );
  NAND2_X1 U19006 ( .A1(n19773), .A2(n18517), .ZN(n18510) );
  NAND2_X1 U19007 ( .A1(n20492), .A2(n18517), .ZN(n18507) );
  NAND2_X1 U19008 ( .A1(n19526), .A2(n18507), .ZN(n18509) );
  OAI21_X1 U19009 ( .B1(n20433), .B2(n18510), .A(n18509), .ZN(n18527) );
  NAND2_X1 U19010 ( .A1(n19758), .A2(Key[124]), .ZN(n18514) );
  OR2_X1 U19011 ( .A1(n19773), .A2(n20492), .ZN(n18523) );
  XNOR2_X1 U19012 ( .A(n18512), .B(n18517), .ZN(n18513) );
  OAI22_X1 U19013 ( .A1(n18514), .A2(n18523), .B1(n18513), .B2(n19758), .ZN(
        n18515) );
  NAND2_X1 U19014 ( .A1(n18515), .A2(n18504), .ZN(n18526) );
  OR2_X1 U19015 ( .A1(n19773), .A2(Key[124]), .ZN(n18520) );
  INV_X1 U19016 ( .A(n18520), .ZN(n18524) );
  OAI22_X1 U19017 ( .A1(n18520), .A2(n20492), .B1(n19758), .B2(n18517), .ZN(
        n18521) );
  OAI211_X1 U19018 ( .C1(n18524), .C2(n18523), .A(n18522), .B(n18521), .ZN(
        n18525) );
  OAI211_X1 U19019 ( .C1(n18528), .C2(n18527), .A(n18526), .B(n18525), .ZN(
        Ciphertext[33]) );
  NAND2_X1 U19020 ( .A1(n18529), .A2(n19682), .ZN(n18553) );
  AOI22_X1 U19021 ( .A1(n18532), .A2(n18531), .B1(n18553), .B2(n18530), .ZN(
        n18533) );
  XNOR2_X1 U19022 ( .A(n18533), .B(n2233), .ZN(Ciphertext[37]) );
  MUX2_X1 U19023 ( .A(n18535), .B(n17564), .S(n20432), .Z(n18536) );
  NAND2_X1 U19024 ( .A1(n18539), .A2(n18536), .ZN(n18537) );
  OAI21_X1 U19025 ( .B1(n18539), .B2(n18538), .A(n18537), .ZN(n18543) );
  NAND4_X1 U19026 ( .A1(n18543), .A2(n18542), .A3(n18541), .A4(n18540), .ZN(
        n18549) );
  NAND2_X1 U19027 ( .A1(n18543), .A2(n18542), .ZN(n18544) );
  OAI21_X1 U19028 ( .B1(n19682), .B2(n18545), .A(n18544), .ZN(n18548) );
  NAND2_X1 U19029 ( .A1(n19682), .A2(n19691), .ZN(n18547) );
  OAI211_X1 U19030 ( .C1(n19682), .C2(n18549), .A(n18548), .B(n18547), .ZN(
        n18551) );
  OAI21_X1 U19031 ( .B1(n18553), .B2(n18552), .A(n18551), .ZN(n18554) );
  XNOR2_X1 U19032 ( .A(n18554), .B(Key[63]), .ZN(Ciphertext[38]) );
  NOR2_X1 U19033 ( .A1(n18555), .A2(n18568), .ZN(n18558) );
  NOR2_X1 U19034 ( .A1(n18565), .A2(n18556), .ZN(n18557) );
  MUX2_X1 U19035 ( .A(n18558), .B(n18557), .S(n18567), .Z(n18563) );
  OAI22_X1 U19036 ( .A1(n18561), .A2(n18566), .B1(n18560), .B2(n18559), .ZN(
        n18562) );
  NOR2_X1 U19037 ( .A1(n18563), .A2(n18562), .ZN(n18564) );
  XNOR2_X1 U19038 ( .A(n18564), .B(n404), .ZN(Ciphertext[45]) );
  OAI21_X1 U19039 ( .B1(n19775), .B2(n18566), .A(n18565), .ZN(n18569) );
  AOI22_X1 U19040 ( .A1(n18571), .A2(n18570), .B1(n18569), .B2(n18568), .ZN(
        n18572) );
  XNOR2_X1 U19041 ( .A(n18572), .B(n2349), .ZN(Ciphertext[47]) );
  NAND2_X1 U19042 ( .A1(n18573), .A2(n18597), .ZN(n18579) );
  NOR2_X1 U19043 ( .A1(n20445), .A2(n18597), .ZN(n18576) );
  NOR2_X1 U19044 ( .A1(n20365), .A2(n19656), .ZN(n18575) );
  NAND3_X1 U19045 ( .A1(n20445), .A2(n18589), .A3(n19669), .ZN(n18578) );
  XNOR2_X1 U19046 ( .A(n18580), .B(n2344), .ZN(Ciphertext[50]) );
  INV_X1 U19047 ( .A(n18597), .ZN(n18583) );
  NOR2_X1 U19048 ( .A1(n20445), .A2(n19656), .ZN(n18581) );
  NAND2_X1 U19049 ( .A1(n18581), .A2(n19665), .ZN(n18582) );
  OAI211_X1 U19050 ( .C1(n18589), .C2(n20445), .A(n18584), .B(n18583), .ZN(
        n18586) );
  OAI21_X1 U19051 ( .B1(n18590), .B2(n18589), .A(n19656), .ZN(n18591) );
  NAND2_X1 U19052 ( .A1(n18597), .A2(n18591), .ZN(n18595) );
  NAND2_X1 U19053 ( .A1(n18593), .A2(n18592), .ZN(n18594) );
  OAI211_X1 U19054 ( .C1(n18597), .C2(n18596), .A(n18595), .B(n18594), .ZN(
        n18599) );
  XNOR2_X1 U19055 ( .A(n18599), .B(n18598), .ZN(Ciphertext[53]) );
  NAND2_X1 U19056 ( .A1(n19679), .A2(n2248), .ZN(n18606) );
  INV_X1 U19057 ( .A(n2248), .ZN(n18610) );
  AND3_X1 U19058 ( .A1(n18622), .A2(n18610), .A3(n19679), .ZN(n18607) );
  OR2_X1 U19059 ( .A1(n18620), .A2(n18610), .ZN(n18612) );
  NOR2_X1 U19060 ( .A1(n18612), .A2(n18600), .ZN(n18601) );
  OAI21_X1 U19061 ( .B1(n18607), .B2(n18601), .A(n18626), .ZN(n18605) );
  NAND3_X1 U19062 ( .A1(n18603), .A2(n19509), .A3(n18610), .ZN(n18604) );
  OAI211_X1 U19063 ( .C1(n19673), .C2(n18606), .A(n18605), .B(n18604), .ZN(
        n18618) );
  INV_X1 U19064 ( .A(n18607), .ZN(n18609) );
  NAND3_X1 U19065 ( .A1(n18619), .A2(n2248), .A3(n18613), .ZN(n18608) );
  OAI21_X1 U19066 ( .B1(n18619), .B2(n18609), .A(n18608), .ZN(n18617) );
  NAND4_X1 U19068 ( .A1(n19877), .A2(n18619), .A3(n18610), .A4(n18613), .ZN(
        n18616) );
  INV_X1 U19069 ( .A(n18612), .ZN(n18614) );
  NAND3_X1 U19070 ( .A1(n20188), .A2(n18614), .A3(n18613), .ZN(n18615) );
  OAI211_X1 U19071 ( .C1(n18618), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        Ciphertext[55]) );
  NOR2_X1 U19072 ( .A1(n18621), .A2(n19679), .ZN(n18623) );
  NOR2_X1 U19073 ( .A1(n18623), .A2(n18622), .ZN(n18624) );
  OAI21_X1 U19074 ( .B1(n18626), .B2(n18625), .A(n18624), .ZN(n18627) );
  OAI211_X1 U19075 ( .C1(n20188), .C2(n18629), .A(n18628), .B(n18627), .ZN(
        n18632) );
  XNOR2_X1 U19076 ( .A(n18632), .B(n18631), .ZN(Ciphertext[57]) );
  NOR2_X1 U19078 ( .A1(n18634), .A2(n18633), .ZN(n18638) );
  NOR2_X1 U19079 ( .A1(n18636), .A2(n20349), .ZN(n18637) );
  OAI211_X1 U19080 ( .C1(n18644), .C2(n19745), .A(n18639), .B(n19934), .ZN(
        n18640) );
  NOR2_X1 U19081 ( .A1(n18644), .A2(n18648), .ZN(n18659) );
  NAND2_X1 U19082 ( .A1(n18656), .A2(n19934), .ZN(n18646) );
  NOR2_X1 U19085 ( .A1(n19935), .A2(n18650), .ZN(n18655) );
  NOR2_X1 U19086 ( .A1(n19934), .A2(n18651), .ZN(n18653) );
  XNOR2_X1 U19089 ( .A(n18661), .B(n18660), .ZN(Ciphertext[63]) );
  INV_X1 U19090 ( .A(n18679), .ZN(n18663) );
  NOR2_X1 U19091 ( .A1(n18672), .A2(n18671), .ZN(n18684) );
  NOR2_X1 U19092 ( .A1(n18684), .A2(n19735), .ZN(n18662) );
  NAND2_X1 U19093 ( .A1(n18686), .A2(n18672), .ZN(n18675) );
  OAI22_X1 U19094 ( .A1(n18663), .A2(n18662), .B1(n18669), .B2(n18675), .ZN(
        n18665) );
  XNOR2_X1 U19095 ( .A(n18665), .B(n18664), .ZN(Ciphertext[67]) );
  NOR2_X1 U19096 ( .A1(n18688), .A2(n18666), .ZN(n18668) );
  NAND3_X1 U19097 ( .A1(n19510), .A2(n18671), .A3(n18686), .ZN(n18678) );
  NOR2_X1 U19098 ( .A1(n18673), .A2(n18672), .ZN(n18674) );
  NOR2_X1 U19099 ( .A1(n18688), .A2(n18674), .ZN(n18676) );
  NAND2_X1 U19100 ( .A1(n18676), .A2(n18675), .ZN(n18677) );
  OAI211_X1 U19101 ( .C1(n18682), .C2(n18679), .A(n18678), .B(n18677), .ZN(
        n18680) );
  XNOR2_X1 U19102 ( .A(n18680), .B(n1781), .ZN(Ciphertext[69]) );
  NOR2_X1 U19103 ( .A1(n18688), .A2(n19510), .ZN(n18685) );
  INV_X1 U19104 ( .A(n18682), .ZN(n18683) );
  OAI21_X1 U19105 ( .B1(n18685), .B2(n18684), .A(n18683), .ZN(n18690) );
  OAI21_X1 U19106 ( .B1(n18686), .B2(n18672), .A(n17964), .ZN(n18687) );
  NAND2_X1 U19107 ( .A1(n18688), .A2(n18687), .ZN(n18689) );
  NAND2_X1 U19108 ( .A1(n18690), .A2(n18689), .ZN(n18693) );
  XNOR2_X1 U19110 ( .A(n18693), .B(n19640), .ZN(Ciphertext[71]) );
  AND2_X1 U19111 ( .A1(n18698), .A2(n18703), .ZN(n18699) );
  NAND2_X1 U19112 ( .A1(n18072), .A2(n18702), .ZN(n18694) );
  AOI22_X1 U19113 ( .A1(n18695), .A2(n18706), .B1(n18699), .B2(n18694), .ZN(
        n18696) );
  XNOR2_X1 U19114 ( .A(n18696), .B(n2222), .ZN(Ciphertext[73]) );
  OAI21_X1 U19115 ( .B1(n18698), .B2(n19753), .A(n18697), .ZN(n18700) );
  NAND3_X1 U19116 ( .A1(n19751), .A2(n18702), .A3(n18701), .ZN(n18704) );
  OAI211_X1 U19117 ( .C1(n18072), .C2(n18706), .A(n18705), .B(n18704), .ZN(
        n18708) );
  INV_X1 U19118 ( .A(n2376), .ZN(n18707) );
  XNOR2_X1 U19119 ( .A(n18708), .B(n18707), .ZN(Ciphertext[75]) );
  AND2_X1 U19120 ( .A1(n18775), .A2(n18709), .ZN(n18761) );
  NAND2_X1 U19121 ( .A1(n18761), .A2(n19803), .ZN(n18715) );
  NAND2_X1 U19123 ( .A1(n18746), .A2(n18781), .ZN(n18714) );
  INV_X1 U19124 ( .A(n18775), .ZN(n18711) );
  INV_X1 U19127 ( .A(n18716), .ZN(n18717) );
  NOR2_X1 U19129 ( .A1(n18774), .A2(n18762), .ZN(n18771) );
  NAND2_X1 U19130 ( .A1(n18771), .A2(n18763), .ZN(n18725) );
  AND2_X1 U19131 ( .A1(n18781), .A2(n18741), .ZN(n18776) );
  INV_X1 U19132 ( .A(n18776), .ZN(n18724) );
  NAND4_X1 U19133 ( .A1(n18719), .A2(n18722), .A3(n18721), .A4(n18720), .ZN(
        n18728) );
  NAND3_X1 U19134 ( .A1(n18774), .A2(n18773), .A3(n18728), .ZN(n18723) );
  NAND4_X1 U19135 ( .A1(n18725), .A2(n18726), .A3(n18724), .A4(n18723), .ZN(
        n18732) );
  INV_X1 U19136 ( .A(n18726), .ZN(n18727) );
  NAND2_X1 U19137 ( .A1(n18776), .A2(n18727), .ZN(n18731) );
  NAND4_X1 U19138 ( .A1(n18763), .A2(n18772), .A3(n18727), .A4(n18749), .ZN(
        n18730) );
  NAND4_X1 U19139 ( .A1(n18728), .A2(n18774), .A3(n18773), .A4(n18727), .ZN(
        n18729) );
  NAND4_X1 U19140 ( .A1(n18732), .A2(n18731), .A3(n18730), .A4(n18729), .ZN(
        Ciphertext[79]) );
  INV_X1 U19141 ( .A(n2381), .ZN(n18743) );
  AND2_X1 U19142 ( .A1(n18773), .A2(n18743), .ZN(n18733) );
  NAND3_X1 U19143 ( .A1(n18733), .A2(n18781), .A3(n18772), .ZN(n18737) );
  NAND3_X1 U19146 ( .A1(n18762), .A2(n18773), .A3(n2381), .ZN(n18735) );
  NAND2_X1 U19151 ( .A1(n18741), .A2(n18773), .ZN(n18742) );
  NAND3_X1 U19152 ( .A1(n18763), .A2(n2381), .A3(n18742), .ZN(n18745) );
  NAND3_X1 U19153 ( .A1(n18746), .A2(n18763), .A3(n18743), .ZN(n18744) );
  OAI21_X1 U19154 ( .B1(n18746), .B2(n18745), .A(n18744), .ZN(n18747) );
  NAND2_X1 U19156 ( .A1(n18750), .A2(n18753), .ZN(n18751) );
  NAND2_X1 U19157 ( .A1(n18752), .A2(n18751), .ZN(n18757) );
  NAND2_X1 U19158 ( .A1(n18754), .A2(n18753), .ZN(n18756) );
  MUX2_X1 U19159 ( .A(n18757), .B(n18756), .S(n20438), .Z(n18760) );
  INV_X1 U19160 ( .A(n18758), .ZN(n18759) );
  NAND2_X1 U19161 ( .A1(n18760), .A2(n18759), .ZN(n18766) );
  NAND2_X1 U19162 ( .A1(n18766), .A2(n18761), .ZN(n18765) );
  NAND3_X1 U19163 ( .A1(n18763), .A2(n18773), .A3(n18762), .ZN(n18764) );
  OAI211_X1 U19164 ( .C1(n18767), .C2(n18766), .A(n18765), .B(n18764), .ZN(
        n18770) );
  INV_X1 U19165 ( .A(n18768), .ZN(n18769) );
  XNOR2_X1 U19166 ( .A(n18770), .B(n18769), .ZN(Ciphertext[81]) );
  NAND2_X1 U19167 ( .A1(n18771), .A2(n18775), .ZN(n18780) );
  OAI21_X1 U19168 ( .B1(n18774), .B2(n18773), .A(n18772), .ZN(n18785) );
  NAND2_X1 U19169 ( .A1(n18785), .A2(n18783), .ZN(n18778) );
  NAND2_X1 U19170 ( .A1(n18776), .A2(n18775), .ZN(n18777) );
  NAND4_X1 U19171 ( .A1(n18780), .A2(n18779), .A3(n18778), .A4(n18777), .ZN(
        n18789) );
  OR2_X1 U19172 ( .A1(n18780), .A2(n18779), .ZN(n18788) );
  NAND3_X1 U19173 ( .A1(n18782), .A2(n18784), .A3(n18781), .ZN(n18787) );
  NAND3_X1 U19174 ( .A1(n18785), .A2(n18784), .A3(n18783), .ZN(n18786) );
  NAND4_X1 U19175 ( .A1(n18789), .A2(n18788), .A3(n18787), .A4(n18786), .ZN(
        Ciphertext[83]) );
  MUX2_X1 U19176 ( .A(n18794), .B(n18807), .S(n19770), .Z(n18791) );
  NAND2_X1 U19177 ( .A1(n18794), .A2(n17772), .ZN(n18804) );
  OAI21_X1 U19178 ( .B1(n19711), .B2(n18331), .A(n18804), .ZN(n18790) );
  MUX2_X1 U19179 ( .A(n18791), .B(n18790), .S(n18795), .Z(n18793) );
  XNOR2_X1 U19180 ( .A(n18793), .B(n18792), .ZN(Ciphertext[86]) );
  MUX2_X1 U19181 ( .A(n17772), .B(n19711), .S(n18803), .Z(n18799) );
  NAND2_X1 U19182 ( .A1(n18807), .A2(n18800), .ZN(n18797) );
  NAND2_X1 U19183 ( .A1(n18794), .A2(n18803), .ZN(n18796) );
  OAI21_X1 U19184 ( .B1(n18800), .B2(n18799), .A(n18798), .ZN(n18802) );
  XNOR2_X1 U19185 ( .A(n18802), .B(n296), .ZN(Ciphertext[88]) );
  NAND2_X1 U19186 ( .A1(n18804), .A2(n18803), .ZN(n18805) );
  AOI22_X1 U19187 ( .A1(n18808), .A2(n18807), .B1(n19770), .B2(n18805), .ZN(
        n18810) );
  XNOR2_X1 U19188 ( .A(n18810), .B(n18809), .ZN(Ciphertext[89]) );
  NAND3_X1 U19189 ( .A1(n20130), .A2(n18172), .A3(n20276), .ZN(n18816) );
  NAND3_X1 U19190 ( .A1(n18814), .A2(n18813), .A3(n18812), .ZN(n18815) );
  OAI211_X1 U19191 ( .C1(n18818), .C2(n18817), .A(n18815), .B(n18816), .ZN(
        n18820) );
  XNOR2_X1 U19192 ( .A(n18820), .B(n1783), .ZN(Ciphertext[93]) );
  XNOR2_X1 U19193 ( .A(n19766), .B(n18830), .ZN(n18822) );
  NAND3_X1 U19194 ( .A1(n18822), .A2(n20276), .A3(n19794), .ZN(n18839) );
  AND2_X1 U19195 ( .A1(n18172), .A2(n18830), .ZN(n18829) );
  NOR2_X1 U19196 ( .A1(n19890), .A2(n18830), .ZN(n18823) );
  AOI21_X1 U19197 ( .B1(n18829), .B2(n19890), .A(n18823), .ZN(n18826) );
  NOR2_X1 U19198 ( .A1(n18172), .A2(n18830), .ZN(n18835) );
  NOR2_X1 U19199 ( .A1(n19794), .A2(n18835), .ZN(n18825) );
  OAI211_X1 U19200 ( .C1(n20130), .C2(n18827), .A(n18826), .B(n18825), .ZN(
        n18838) );
  NOR2_X1 U19201 ( .A1(n20422), .A2(n18830), .ZN(n18832) );
  INV_X1 U19202 ( .A(n18831), .ZN(n18840) );
  OAI211_X1 U19203 ( .C1(n18833), .C2(n18832), .A(n18840), .B(n19794), .ZN(
        n18837) );
  NAND3_X1 U19204 ( .A1(n18840), .A2(n18835), .A3(n18834), .ZN(n18836) );
  NAND4_X1 U19205 ( .A1(n18839), .A2(n18838), .A3(n18837), .A4(n18836), .ZN(
        Ciphertext[94]) );
  NAND2_X1 U19206 ( .A1(n18841), .A2(n18840), .ZN(n18843) );
  AOI22_X1 U19207 ( .A1(n18845), .A2(n19890), .B1(n18843), .B2(n19794), .ZN(
        n18846) );
  XNOR2_X1 U19208 ( .A(n18846), .B(n2108), .ZN(Ciphertext[95]) );
  AOI21_X1 U19210 ( .B1(n19917), .B2(n19988), .A(n18850), .ZN(n18847) );
  INV_X1 U19211 ( .A(n18848), .ZN(n18849) );
  OAI21_X1 U19212 ( .B1(n18871), .B2(n18853), .A(n18852), .ZN(n18856) );
  INV_X1 U19213 ( .A(n18854), .ZN(n18855) );
  XNOR2_X1 U19214 ( .A(n18856), .B(n18855), .ZN(Ciphertext[97]) );
  NAND2_X1 U19215 ( .A1(n18857), .A2(n20259), .ZN(n18860) );
  OR2_X1 U19216 ( .A1(n3030), .A2(n19988), .ZN(n18859) );
  OAI21_X1 U19217 ( .B1(n18862), .B2(n20259), .A(n18861), .ZN(n18865) );
  INV_X1 U19218 ( .A(n18863), .ZN(n18864) );
  XNOR2_X1 U19219 ( .A(n18865), .B(n18864), .ZN(Ciphertext[100]) );
  AOI21_X1 U19220 ( .B1(n20418), .B2(n20117), .A(n20259), .ZN(n18870) );
  OAI22_X1 U19221 ( .A1(n18871), .A2(n3030), .B1(n18870), .B2(n18869), .ZN(
        n18873) );
  INV_X1 U19222 ( .A(n2164), .ZN(n18872) );
  XNOR2_X1 U19223 ( .A(n18873), .B(n18872), .ZN(Ciphertext[101]) );
  INV_X1 U19224 ( .A(n18921), .ZN(n18898) );
  NAND2_X1 U19225 ( .A1(n19874), .A2(n18876), .ZN(n18879) );
  NAND2_X1 U19226 ( .A1(n18899), .A2(n18916), .ZN(n18901) );
  NOR2_X1 U19227 ( .A1(n18901), .A2(n19681), .ZN(n18875) );
  NOR2_X1 U19228 ( .A1(n18875), .A2(n18874), .ZN(n18878) );
  NAND3_X1 U19229 ( .A1(n18897), .A2(n19681), .A3(n18876), .ZN(n18877) );
  OAI211_X1 U19230 ( .C1(n18898), .C2(n18879), .A(n18878), .B(n18877), .ZN(
        n18881) );
  XNOR2_X1 U19231 ( .A(n18881), .B(n18880), .ZN(Ciphertext[102]) );
  INV_X1 U19232 ( .A(n18899), .ZN(n18882) );
  INV_X1 U19233 ( .A(n18918), .ZN(n18886) );
  AND2_X1 U19234 ( .A1(n17054), .A2(n18897), .ZN(n18917) );
  NAND2_X1 U19235 ( .A1(n18917), .A2(n18882), .ZN(n18885) );
  INV_X1 U19236 ( .A(n18897), .ZN(n18883) );
  OAI211_X1 U19237 ( .C1(n19664), .C2(n19874), .A(n18883), .B(n19681), .ZN(
        n18884) );
  NAND3_X1 U19238 ( .A1(n18886), .A2(n18885), .A3(n18884), .ZN(n18889) );
  INV_X1 U19239 ( .A(n18887), .ZN(n18888) );
  XNOR2_X1 U19240 ( .A(n18889), .B(n18888), .ZN(Ciphertext[103]) );
  MUX2_X1 U19241 ( .A(n18890), .B(n18916), .S(n18921), .Z(n18893) );
  NAND2_X1 U19242 ( .A1(n18897), .A2(n18890), .ZN(n18919) );
  NAND2_X1 U19243 ( .A1(n18919), .A2(n18891), .ZN(n18892) );
  MUX2_X1 U19244 ( .A(n18893), .B(n18892), .S(n19874), .Z(n18895) );
  INV_X1 U19245 ( .A(n2446), .ZN(n18894) );
  XNOR2_X1 U19246 ( .A(n18895), .B(n18894), .ZN(Ciphertext[104]) );
  NAND2_X1 U19247 ( .A1(n19874), .A2(n18897), .ZN(n18896) );
  OAI21_X1 U19248 ( .B1(n19681), .B2(n18897), .A(n18896), .ZN(n18911) );
  NAND2_X1 U19249 ( .A1(n18898), .A2(n18911), .ZN(n18904) );
  NOR2_X1 U19250 ( .A1(n19905), .A2(n19874), .ZN(n18907) );
  AOI21_X1 U19251 ( .B1(n18907), .B2(n19681), .A(n18909), .ZN(n18903) );
  INV_X1 U19252 ( .A(n18901), .ZN(n18902) );
  NAND2_X1 U19253 ( .A1(n18921), .A2(n18902), .ZN(n18905) );
  NAND3_X1 U19254 ( .A1(n18904), .A2(n18903), .A3(n18905), .ZN(n18915) );
  INV_X1 U19255 ( .A(n18905), .ZN(n18910) );
  NOR2_X1 U19256 ( .A1(n18890), .A2(n2203), .ZN(n18908) );
  AOI22_X1 U19257 ( .A1(n18910), .A2(n18909), .B1(n18908), .B2(n18907), .ZN(
        n18914) );
  NOR2_X1 U19258 ( .A1(n18921), .A2(n2203), .ZN(n18912) );
  NAND2_X1 U19259 ( .A1(n18912), .A2(n18911), .ZN(n18913) );
  NAND3_X1 U19260 ( .A1(n18915), .A2(n18914), .A3(n18913), .ZN(Ciphertext[105]) );
  OAI21_X1 U19261 ( .B1(n18918), .B2(n18917), .A(n19664), .ZN(n18923) );
  NAND2_X1 U19262 ( .A1(n18919), .A2(n19905), .ZN(n18920) );
  XNOR2_X1 U19263 ( .A(n18925), .B(n18924), .ZN(Ciphertext[107]) );
  NAND2_X1 U19264 ( .A1(n18932), .A2(n18926), .ZN(n18930) );
  NAND2_X1 U19265 ( .A1(n20501), .A2(n18937), .ZN(n18943) );
  NAND2_X1 U19266 ( .A1(n18940), .A2(n18939), .ZN(n18942) );
  MUX2_X1 U19267 ( .A(n18943), .B(n18942), .S(n18941), .Z(n18944) );
  NOR2_X1 U19268 ( .A1(n2058), .A2(n19654), .ZN(n18974) );
  MUX2_X1 U19269 ( .A(n18948), .B(n19916), .S(n18946), .Z(n18952) );
  MUX2_X1 U19270 ( .A(n18950), .B(n18949), .S(n17687), .Z(n18951) );
  AOI22_X1 U19271 ( .A1(n219), .A2(n18954), .B1(n18955), .B2(n18953), .ZN(
        n18960) );
  OR2_X1 U19272 ( .A1(n20221), .A2(n18955), .ZN(n18958) );
  INV_X1 U19274 ( .A(n18961), .ZN(n18963) );
  NAND2_X1 U19275 ( .A1(n18963), .A2(n18962), .ZN(n18964) );
  AND2_X1 U19276 ( .A1(n18965), .A2(n18964), .ZN(n18973) );
  INV_X1 U19277 ( .A(n18966), .ZN(n18967) );
  OR2_X1 U19278 ( .A1(n19684), .A2(n18967), .ZN(n18971) );
  MUX2_X1 U19279 ( .A(n18971), .B(n18970), .S(n20127), .Z(n18972) );
  OAI21_X1 U19280 ( .B1(n18973), .B2(n220), .A(n18972), .ZN(n19011) );
  INV_X1 U19281 ( .A(n19680), .ZN(n19025) );
  OAI21_X1 U19282 ( .B1(n18974), .B2(n19004), .A(n19025), .ZN(n18983) );
  MUX2_X1 U19283 ( .A(n18976), .B(n20158), .S(n18978), .Z(n18981) );
  AOI21_X1 U19284 ( .B1(n18981), .B2(n18980), .A(n18979), .ZN(n19002) );
  AND2_X1 U19285 ( .A1(n19001), .A2(n19002), .ZN(n19010) );
  INV_X1 U19286 ( .A(n19010), .ZN(n19015) );
  INV_X1 U19288 ( .A(n18984), .ZN(n18985) );
  NOR2_X1 U19289 ( .A1(n19011), .A2(n19687), .ZN(n18995) );
  NAND2_X1 U19291 ( .A1(n2058), .A2(n19724), .ZN(n18987) );
  INV_X1 U19292 ( .A(n19021), .ZN(n18986) );
  AOI22_X1 U19293 ( .A1(n18986), .A2(n19687), .B1(n19013), .B2(n19002), .ZN(
        n19026) );
  OAI22_X1 U19294 ( .A1(n18995), .A2(n18987), .B1(n19026), .B2(n19004), .ZN(
        n18990) );
  INV_X1 U19295 ( .A(n18988), .ZN(n18989) );
  XNOR2_X1 U19296 ( .A(n18990), .B(n18989), .ZN(Ciphertext[109]) );
  INV_X1 U19297 ( .A(n19023), .ZN(n18994) );
  INV_X1 U19298 ( .A(n19009), .ZN(n18999) );
  NAND2_X1 U19299 ( .A1(n18999), .A2(n19654), .ZN(n18993) );
  NAND2_X1 U19300 ( .A1(n18999), .A2(n19867), .ZN(n18991) );
  NAND2_X1 U19301 ( .A1(n18995), .A2(n19866), .ZN(n18996) );
  XNOR2_X1 U19302 ( .A(n18998), .B(n18997), .ZN(Ciphertext[110]) );
  NOR2_X1 U19303 ( .A1(n19687), .A2(n19654), .ZN(n19003) );
  INV_X1 U19304 ( .A(n19002), .ZN(n19022) );
  AOI22_X1 U19305 ( .A1(n19004), .A2(n19680), .B1(n19003), .B2(n19022), .ZN(
        n19005) );
  OAI21_X1 U19306 ( .B1(n19006), .B2(n19866), .A(n19005), .ZN(n19008) );
  XNOR2_X1 U19307 ( .A(n19008), .B(n19007), .ZN(Ciphertext[111]) );
  NOR2_X1 U19308 ( .A1(n19687), .A2(n19866), .ZN(n19012) );
  AOI22_X1 U19309 ( .A1(n19012), .A2(n19680), .B1(n19010), .B2(n19687), .ZN(
        n19017) );
  NAND2_X1 U19310 ( .A1(n19013), .A2(n19022), .ZN(n19014) );
  NAND3_X1 U19311 ( .A1(n19015), .A2(n19014), .A3(n19867), .ZN(n19016) );
  NAND2_X1 U19312 ( .A1(n19017), .A2(n19016), .ZN(n19020) );
  INV_X1 U19313 ( .A(n19018), .ZN(n19019) );
  XNOR2_X1 U19314 ( .A(n19020), .B(n19019), .ZN(Ciphertext[112]) );
  OAI21_X1 U19315 ( .B1(n19023), .B2(n19022), .A(n19867), .ZN(n19024) );
  OAI21_X1 U19316 ( .B1(n19026), .B2(n19025), .A(n19024), .ZN(n19029) );
  INV_X1 U19317 ( .A(n19027), .ZN(n19028) );
  XNOR2_X1 U19318 ( .A(n19029), .B(n19028), .ZN(Ciphertext[113]) );
  NOR2_X1 U19320 ( .A1(n19046), .A2(n19032), .ZN(n19033) );
  AOI21_X1 U19321 ( .B1(n20475), .B2(n19034), .A(n19047), .ZN(n19036) );
  NAND2_X1 U19322 ( .A1(n19036), .A2(n19035), .ZN(n19037) );
  XNOR2_X1 U19323 ( .A(n19039), .B(n19038), .ZN(Ciphertext[117]) );
  NOR2_X1 U19324 ( .A1(n20475), .A2(n19993), .ZN(n19042) );
  AND2_X1 U19325 ( .A1(n19992), .A2(n19047), .ZN(n19041) );
  OAI21_X1 U19326 ( .B1(n19042), .B2(n19041), .A(n19046), .ZN(n19051) );
  INV_X1 U19327 ( .A(n19047), .ZN(n19045) );
  NAND3_X1 U19328 ( .A1(n19045), .A2(n20475), .A3(n20142), .ZN(n19050) );
  INV_X1 U19329 ( .A(n19046), .ZN(n19048) );
  NAND3_X1 U19330 ( .A1(n19048), .A2(n18061), .A3(n19047), .ZN(n19049) );
  NAND3_X1 U19331 ( .A1(n19051), .A2(n19050), .A3(n19049), .ZN(n19054) );
  INV_X1 U19332 ( .A(n19052), .ZN(n19053) );
  XNOR2_X1 U19333 ( .A(n19054), .B(n19053), .ZN(Ciphertext[118]) );
  INV_X1 U19334 ( .A(n19073), .ZN(n19076) );
  OAI21_X1 U19335 ( .B1(n19076), .B2(n20131), .A(n19055), .ZN(n19057) );
  INV_X1 U19336 ( .A(n19067), .ZN(n19077) );
  NAND3_X1 U19337 ( .A1(n19069), .A2(n20131), .A3(n19077), .ZN(n19056) );
  NAND2_X1 U19338 ( .A1(n19058), .A2(n19076), .ZN(n19063) );
  INV_X1 U19339 ( .A(n19079), .ZN(n19062) );
  NAND3_X1 U19340 ( .A1(n19653), .A2(n19073), .A3(n19059), .ZN(n19061) );
  OAI211_X1 U19341 ( .C1(n19064), .C2(n19063), .A(n19062), .B(n19061), .ZN(
        n19066) );
  INV_X1 U19342 ( .A(n2384), .ZN(n19065) );
  XNOR2_X1 U19343 ( .A(n19066), .B(n19065), .ZN(Ciphertext[121]) );
  INV_X1 U19344 ( .A(n19068), .ZN(n19082) );
  AOI21_X1 U19345 ( .B1(n19075), .B2(n19073), .A(n19082), .ZN(n19072) );
  NOR2_X1 U19346 ( .A1(n19685), .A2(n19067), .ZN(n19070) );
  AOI21_X1 U19347 ( .B1(n20131), .B2(n19073), .A(n19075), .ZN(n19081) );
  NOR2_X1 U19348 ( .A1(n19076), .A2(n19075), .ZN(n19078) );
  OAI21_X1 U19349 ( .B1(n19079), .B2(n19078), .A(n19077), .ZN(n19080) );
  XNOR2_X1 U19350 ( .A(n19084), .B(n19083), .ZN(Ciphertext[125]) );
  NOR2_X1 U19351 ( .A1(n19105), .A2(n19112), .ZN(n19090) );
  INV_X1 U19352 ( .A(n19085), .ZN(n19086) );
  XNOR2_X1 U19353 ( .A(n19091), .B(n304), .ZN(Ciphertext[127]) );
  NOR2_X1 U19354 ( .A1(n19093), .A2(n19911), .ZN(n19101) );
  INV_X1 U19355 ( .A(n19094), .ZN(n19097) );
  NAND2_X1 U19356 ( .A1(n19112), .A2(n19095), .ZN(n19096) );
  NAND2_X1 U19357 ( .A1(n19097), .A2(n19096), .ZN(n19100) );
  AND2_X1 U19358 ( .A1(n19115), .A2(n19098), .ZN(n19118) );
  INV_X1 U19361 ( .A(n19102), .ZN(n19103) );
  INV_X1 U19363 ( .A(n19105), .ZN(n19122) );
  INV_X1 U19364 ( .A(n19106), .ZN(n19107) );
  NAND2_X1 U19365 ( .A1(n19107), .A2(n19110), .ZN(n19108) );
  OAI211_X1 U19366 ( .C1(n19111), .C2(n19110), .A(n19109), .B(n19108), .ZN(
        n19121) );
  NOR2_X1 U19367 ( .A1(n19115), .A2(n17203), .ZN(n19117) );
  OAI21_X1 U19368 ( .B1(n19118), .B2(n19117), .A(n19116), .ZN(n19119) );
  OAI211_X1 U19369 ( .C1(n19122), .C2(n19121), .A(n19120), .B(n19119), .ZN(
        n19124) );
  XNOR2_X1 U19370 ( .A(n19124), .B(n19123), .ZN(Ciphertext[130]) );
  NOR2_X1 U19371 ( .A1(n19144), .A2(n19134), .ZN(n19126) );
  AOI22_X1 U19372 ( .A1(n19126), .A2(n19125), .B1(n19133), .B2(n19144), .ZN(
        n19129) );
  NAND2_X1 U19373 ( .A1(n19127), .A2(n19146), .ZN(n19128) );
  OAI211_X1 U19374 ( .C1(n19130), .C2(n833), .A(n19129), .B(n19128), .ZN(
        n19131) );
  XNOR2_X1 U19375 ( .A(n19131), .B(n293), .ZN(Ciphertext[132]) );
  NAND2_X1 U19376 ( .A1(n19144), .A2(n16780), .ZN(n19132) );
  OAI211_X1 U19377 ( .C1(n19135), .C2(n19144), .A(n19133), .B(n19132), .ZN(
        n19139) );
  NAND3_X1 U19378 ( .A1(n19135), .A2(n19134), .A3(n870), .ZN(n19138) );
  NAND3_X1 U19379 ( .A1(n19146), .A2(n16780), .A3(n19151), .ZN(n19137) );
  NAND3_X1 U19380 ( .A1(n19139), .A2(n19138), .A3(n19137), .ZN(n19142) );
  INV_X1 U19381 ( .A(n19140), .ZN(n19141) );
  XNOR2_X1 U19382 ( .A(n19142), .B(n19141), .ZN(Ciphertext[136]) );
  AOI21_X1 U19383 ( .B1(n19145), .B2(n19144), .A(n870), .ZN(n19150) );
  OAI21_X1 U19384 ( .B1(n19148), .B2(n19147), .A(n19146), .ZN(n19149) );
  OAI21_X1 U19385 ( .B1(n19151), .B2(n19150), .A(n19149), .ZN(n19153) );
  XNOR2_X1 U19386 ( .A(n19153), .B(n19152), .ZN(Ciphertext[137]) );
  INV_X1 U19387 ( .A(n19155), .ZN(n19161) );
  AOI21_X1 U19388 ( .B1(n2918), .B2(n19165), .A(n19161), .ZN(n19156) );
  OAI22_X1 U19389 ( .A1(n19157), .A2(n19165), .B1(n19708), .B2(n19156), .ZN(
        n19160) );
  INV_X1 U19390 ( .A(n19158), .ZN(n19159) );
  XNOR2_X1 U19391 ( .A(n19160), .B(n19159), .ZN(Ciphertext[138]) );
  XNOR2_X1 U19392 ( .A(n19167), .B(n875), .ZN(Ciphertext[143]) );
  NAND2_X1 U19393 ( .A1(n19171), .A2(n19170), .ZN(n19172) );
  OAI211_X1 U19394 ( .C1(n19175), .C2(n19174), .A(n19173), .B(n19172), .ZN(
        n19177) );
  INV_X1 U19395 ( .A(n2424), .ZN(n19176) );
  XNOR2_X1 U19396 ( .A(n19177), .B(n19176), .ZN(Ciphertext[147]) );
  INV_X1 U19397 ( .A(n19182), .ZN(n19201) );
  OAI21_X1 U19399 ( .B1(n19197), .B2(n19208), .A(n19193), .ZN(n19179) );
  OAI21_X1 U19400 ( .B1(n19210), .B2(n19189), .A(n19209), .ZN(n19178) );
  AOI22_X1 U19401 ( .A1(n19179), .A2(n19210), .B1(n19197), .B2(n19178), .ZN(
        n19181) );
  XNOR2_X1 U19402 ( .A(n19181), .B(n19180), .ZN(Ciphertext[150]) );
  AND2_X1 U19403 ( .A1(n19190), .A2(n19208), .ZN(n19187) );
  AOI21_X1 U19404 ( .B1(n19212), .B2(n19193), .A(n19187), .ZN(n19185) );
  NAND2_X1 U19405 ( .A1(n19210), .A2(n19189), .ZN(n19183) );
  XNOR2_X1 U19408 ( .A(n19186), .B(n1904), .ZN(Ciphertext[151]) );
  INV_X1 U19409 ( .A(n19187), .ZN(n19188) );
  INV_X1 U19410 ( .A(n19196), .ZN(n19198) );
  OAI211_X1 U19411 ( .C1(n19208), .C2(n19201), .A(n19188), .B(n19198), .ZN(
        n19192) );
  NAND3_X1 U19412 ( .A1(n19209), .A2(n19190), .A3(n19189), .ZN(n19191) );
  OAI211_X1 U19413 ( .C1(n19210), .C2(n19193), .A(n19192), .B(n19191), .ZN(
        n19195) );
  INV_X1 U19414 ( .A(n1996), .ZN(n19194) );
  XNOR2_X1 U19415 ( .A(n19195), .B(n19194), .ZN(Ciphertext[153]) );
  OAI21_X1 U19416 ( .B1(n19197), .B2(n19209), .A(n19842), .ZN(n19215) );
  AND2_X1 U19417 ( .A1(n19208), .A2(n19209), .ZN(n19200) );
  OAI21_X1 U19418 ( .B1(n19210), .B2(n19201), .A(n19198), .ZN(n19199) );
  OAI21_X1 U19419 ( .B1(n19215), .B2(n19200), .A(n19199), .ZN(n19204) );
  NAND3_X1 U19420 ( .A1(n19202), .A2(n19197), .A3(n19201), .ZN(n19203) );
  NAND2_X1 U19421 ( .A1(n19204), .A2(n19203), .ZN(n19207) );
  INV_X1 U19422 ( .A(n19205), .ZN(n19206) );
  XNOR2_X1 U19423 ( .A(n19207), .B(n19206), .ZN(Ciphertext[154]) );
  NOR2_X1 U19424 ( .A1(n2943), .A2(n19209), .ZN(n19214) );
  INV_X1 U19425 ( .A(n19210), .ZN(n19211) );
  NAND2_X1 U19426 ( .A1(n19212), .A2(n19211), .ZN(n19213) );
  OAI21_X1 U19427 ( .B1(n19215), .B2(n19214), .A(n19213), .ZN(n19218) );
  INV_X1 U19428 ( .A(n19216), .ZN(n19217) );
  XNOR2_X1 U19429 ( .A(n19218), .B(n19217), .ZN(Ciphertext[155]) );
  MUX2_X1 U19430 ( .A(n19242), .B(n19227), .S(n19233), .Z(n19221) );
  AND2_X1 U19431 ( .A1(n19238), .A2(n19234), .ZN(n19220) );
  AOI22_X1 U19432 ( .A1(n19221), .A2(n20124), .B1(n19220), .B2(n19219), .ZN(
        n19224) );
  INV_X1 U19433 ( .A(n19222), .ZN(n19223) );
  XNOR2_X1 U19434 ( .A(n19224), .B(n19223), .ZN(Ciphertext[158]) );
  INV_X1 U19435 ( .A(n19225), .ZN(n19230) );
  OAI222_X1 U19436 ( .A1(n19239), .A2(n19230), .B1(n19229), .B2(n19242), .C1(
        n19236), .C2(n19228), .ZN(n19232) );
  INV_X1 U19437 ( .A(n632), .ZN(n19231) );
  XNOR2_X1 U19438 ( .A(n19232), .B(n19231), .ZN(Ciphertext[159]) );
  NAND2_X1 U19439 ( .A1(n19233), .A2(n20124), .ZN(n19241) );
  NAND3_X1 U19440 ( .A1(n19239), .A2(n19238), .A3(n20193), .ZN(n19240) );
  INV_X1 U19441 ( .A(n19243), .ZN(n19244) );
  XNOR2_X1 U19442 ( .A(n19245), .B(n19244), .ZN(Ciphertext[160]) );
  NOR2_X1 U19443 ( .A1(n19269), .A2(n19274), .ZN(n19268) );
  INV_X1 U19444 ( .A(n19268), .ZN(n19258) );
  INV_X1 U19445 ( .A(n19269), .ZN(n19275) );
  INV_X1 U19446 ( .A(n19246), .ZN(n19267) );
  NAND3_X1 U19447 ( .A1(n19275), .A2(n19247), .A3(n19267), .ZN(n19257) );
  INV_X1 U19448 ( .A(n19248), .ZN(n19253) );
  INV_X1 U19449 ( .A(n19249), .ZN(n19250) );
  OAI211_X1 U19450 ( .C1(n19253), .C2(n20162), .A(n19251), .B(n19250), .ZN(
        n19254) );
  NAND3_X1 U19451 ( .A1(n19278), .A2(n19254), .A3(n19267), .ZN(n19255) );
  NAND4_X1 U19452 ( .A1(n19258), .A2(n19257), .A3(n19256), .A4(n19255), .ZN(
        n19260) );
  XNOR2_X1 U19453 ( .A(n19260), .B(n19259), .ZN(Ciphertext[162]) );
  NAND3_X1 U19454 ( .A1(n19261), .A2(n19269), .A3(n2816), .ZN(n19262) );
  OAI21_X1 U19455 ( .B1(n19279), .B2(n19263), .A(n19262), .ZN(n19265) );
  XNOR2_X1 U19456 ( .A(n19265), .B(n19264), .ZN(Ciphertext[163]) );
  NOR2_X1 U19457 ( .A1(n19278), .A2(n19267), .ZN(n19266) );
  INV_X1 U19458 ( .A(n2123), .ZN(n19273) );
  OAI22_X1 U19459 ( .A1(n19279), .A2(n19278), .B1(n19277), .B2(n20444), .ZN(
        n19281) );
  XNOR2_X1 U19460 ( .A(n19281), .B(n19280), .ZN(Ciphertext[167]) );
  OAI21_X1 U19461 ( .B1(n20434), .B2(n19284), .A(n19290), .ZN(n19288) );
  NOR3_X1 U19462 ( .A1(n19298), .A2(n19283), .A3(n19282), .ZN(n19286) );
  OAI21_X1 U19463 ( .B1(n19298), .B2(n19292), .A(n19284), .ZN(n19285) );
  INV_X1 U19467 ( .A(n19290), .ZN(n19295) );
  INV_X1 U19468 ( .A(n19299), .ZN(n19291) );
  AOI22_X1 U19469 ( .A1(n1773), .A2(n19292), .B1(n19298), .B2(n19291), .ZN(
        n19305) );
  NAND2_X1 U19470 ( .A1(n20510), .A2(n20218), .ZN(n19293) );
  OAI22_X1 U19471 ( .A1(n19305), .A2(n19295), .B1(n19294), .B2(n19293), .ZN(
        n19297) );
  XNOR2_X1 U19472 ( .A(n19297), .B(n19296), .ZN(Ciphertext[169]) );
  OAI21_X1 U19473 ( .B1(n20364), .B2(n20218), .A(n19298), .ZN(n19301) );
  OAI21_X1 U19475 ( .B1(n19305), .B2(n19304), .A(n19303), .ZN(n19307) );
  INV_X1 U19476 ( .A(n456), .ZN(n19306) );
  XNOR2_X1 U19477 ( .A(n19307), .B(n19306), .ZN(Ciphertext[173]) );
  OAI21_X1 U19478 ( .B1(n19309), .B2(n19308), .A(n19333), .ZN(n19313) );
  AOI21_X1 U19479 ( .B1(n19311), .B2(n19310), .A(n19338), .ZN(n19312) );
  AOI21_X1 U19480 ( .B1(n19334), .B2(n19313), .A(n19312), .ZN(n19314) );
  XNOR2_X1 U19481 ( .A(n19314), .B(n2310), .ZN(Ciphertext[174]) );
  INV_X1 U19482 ( .A(n19315), .ZN(n19320) );
  INV_X1 U19483 ( .A(n19316), .ZN(n19317) );
  NAND3_X1 U19484 ( .A1(n19317), .A2(n19324), .A3(n19749), .ZN(n19319) );
  INV_X1 U19485 ( .A(n19333), .ZN(n19327) );
  NAND3_X1 U19486 ( .A1(n19327), .A2(n19308), .A3(n19329), .ZN(n19318) );
  INV_X1 U19488 ( .A(n19321), .ZN(n19322) );
  NOR2_X1 U19490 ( .A1(n19333), .A2(n19324), .ZN(n19326) );
  OAI21_X1 U19491 ( .B1(n19326), .B2(n19340), .A(n19336), .ZN(n19325) );
  OAI211_X1 U19492 ( .C1(n19336), .C2(n19326), .A(n19325), .B(n19955), .ZN(
        n19346) );
  OAI21_X1 U19493 ( .B1(n19334), .B2(n19336), .A(n19327), .ZN(n19332) );
  NAND2_X1 U19494 ( .A1(n19749), .A2(n19336), .ZN(n19331) );
  NAND3_X1 U19495 ( .A1(n19333), .A2(n19329), .A3(n19337), .ZN(n19330) );
  NAND4_X1 U19496 ( .A1(n19340), .A2(n19332), .A3(n19331), .A4(n19330), .ZN(
        n19345) );
  NOR2_X1 U19497 ( .A1(n19333), .A2(n19955), .ZN(n19335) );
  NAND4_X1 U19498 ( .A1(n19340), .A2(n19336), .A3(n19335), .A4(n19334), .ZN(
        n19344) );
  XNOR2_X1 U19499 ( .A(n19338), .B(n19337), .ZN(n19342) );
  NOR2_X1 U19500 ( .A1(n19340), .A2(n19955), .ZN(n19341) );
  NAND2_X1 U19501 ( .A1(n19342), .A2(n19341), .ZN(n19343) );
  NAND4_X1 U19502 ( .A1(n19346), .A2(n19345), .A3(n19344), .A4(n19343), .ZN(
        Ciphertext[178]) );
  AND2_X1 U19503 ( .A1(n20240), .A2(n19349), .ZN(n19359) );
  OAI21_X1 U19504 ( .B1(n20244), .B2(n19348), .A(n19347), .ZN(n19358) );
  NAND2_X1 U19505 ( .A1(n19351), .A2(n20273), .ZN(n19356) );
  NAND2_X1 U19506 ( .A1(n19353), .A2(n19352), .ZN(n19355) );
  MUX2_X1 U19507 ( .A(n19356), .B(n19355), .S(n20240), .Z(n19357) );
  OAI21_X1 U19508 ( .B1(n19359), .B2(n19358), .A(n19357), .ZN(n19444) );
  INV_X1 U19509 ( .A(n19444), .ZN(n19409) );
  NOR2_X1 U19510 ( .A1(n19361), .A2(n19360), .ZN(n19369) );
  INV_X1 U19511 ( .A(n20212), .ZN(n19364) );
  NAND2_X1 U19512 ( .A1(n19364), .A2(n19938), .ZN(n19368) );
  NAND2_X1 U19513 ( .A1(n19366), .A2(n19365), .ZN(n19367) );
  OAI21_X1 U19514 ( .B1(n19369), .B2(n19368), .A(n19367), .ZN(n19440) );
  INV_X1 U19515 ( .A(n19440), .ZN(n19381) );
  MUX2_X1 U19516 ( .A(n19373), .B(n19666), .S(n19370), .Z(n19379) );
  NAND2_X1 U19517 ( .A1(n19373), .A2(n19372), .ZN(n19377) );
  OAI21_X1 U19521 ( .B1(n1897), .B2(n20463), .A(n19382), .ZN(n19384) );
  NOR2_X1 U19522 ( .A1(n19388), .A2(n20004), .ZN(n19393) );
  NOR2_X1 U19523 ( .A1(n19390), .A2(n20172), .ZN(n19392) );
  OAI21_X1 U19524 ( .B1(n19393), .B2(n19392), .A(n19391), .ZN(n19398) );
  NAND3_X1 U19525 ( .A1(n19396), .A2(n19395), .A3(n20004), .ZN(n19397) );
  NAND2_X1 U19526 ( .A1(n3827), .A2(n19425), .ZN(n19408) );
  OAI21_X1 U19527 ( .B1(n19402), .B2(n19403), .A(n19401), .ZN(n19406) );
  OAI21_X1 U19529 ( .B1(n19409), .B2(n19442), .A(n19418), .ZN(n19407) );
  AOI22_X1 U19530 ( .A1(n19409), .A2(n19408), .B1(n19407), .B2(n19439), .ZN(
        n19411) );
  XNOR2_X1 U19531 ( .A(n19411), .B(n19410), .ZN(Ciphertext[180]) );
  INV_X1 U19532 ( .A(n19442), .ZN(n19434) );
  NOR2_X1 U19533 ( .A1(n19439), .A2(n19440), .ZN(n19430) );
  OAI21_X1 U19534 ( .B1(n19444), .B2(n19434), .A(n19430), .ZN(n19413) );
  AND2_X1 U19535 ( .A1(n19440), .A2(n19432), .ZN(n19445) );
  OAI21_X1 U19536 ( .B1(n19445), .B2(n19434), .A(n19425), .ZN(n19412) );
  NAND2_X1 U19537 ( .A1(n19413), .A2(n19412), .ZN(n19415) );
  INV_X1 U19538 ( .A(n2298), .ZN(n19414) );
  XNOR2_X1 U19539 ( .A(n19415), .B(n19414), .ZN(Ciphertext[181]) );
  MUX2_X1 U19540 ( .A(n19444), .B(n19439), .S(n19441), .Z(n19416) );
  NAND2_X1 U19541 ( .A1(n19416), .A2(n19442), .ZN(n19421) );
  XNOR2_X1 U19546 ( .A(n19423), .B(n19422), .ZN(Ciphertext[182]) );
  NAND2_X1 U19547 ( .A1(n19442), .A2(n19440), .ZN(n19424) );
  NAND2_X1 U19548 ( .A1(n19424), .A2(n19448), .ZN(n19429) );
  INV_X1 U19549 ( .A(n19439), .ZN(n19426) );
  NAND3_X1 U19550 ( .A1(n19426), .A2(n19442), .A3(n19418), .ZN(n19427) );
  OAI211_X1 U19551 ( .C1(n19430), .C2(n19429), .A(n19428), .B(n19427), .ZN(
        n19431) );
  XNOR2_X1 U19552 ( .A(n19431), .B(n2709), .ZN(Ciphertext[183]) );
  MUX2_X1 U19553 ( .A(n19440), .B(n19439), .S(n19432), .Z(n19435) );
  NAND2_X1 U19554 ( .A1(n19439), .A2(n19432), .ZN(n19433) );
  INV_X1 U19555 ( .A(n19436), .ZN(n19437) );
  XNOR2_X1 U19556 ( .A(n19438), .B(n19437), .ZN(Ciphertext[184]) );
  AOI21_X1 U19557 ( .B1(n19440), .B2(n19439), .A(n19418), .ZN(n19449) );
  INV_X1 U19558 ( .A(n19441), .ZN(n19443) );
  NOR2_X1 U19559 ( .A1(n19443), .A2(n19442), .ZN(n19446) );
  OAI21_X1 U19560 ( .B1(n19446), .B2(n19445), .A(n19444), .ZN(n19447) );
  OAI21_X1 U19561 ( .B1(n19449), .B2(n19448), .A(n19447), .ZN(n19451) );
  INV_X1 U19562 ( .A(n620), .ZN(n19450) );
  XNOR2_X1 U19563 ( .A(n19451), .B(n19450), .ZN(Ciphertext[185]) );
  OAI22_X1 U19564 ( .A1(n212), .A2(n19453), .B1(n19463), .B2(n19460), .ZN(
        n19466) );
  NAND2_X1 U19565 ( .A1(n19453), .A2(n19459), .ZN(n19454) );
  AOI22_X1 U19566 ( .A1(n19466), .A2(n19456), .B1(n19738), .B2(n19454), .ZN(
        n19458) );
  XNOR2_X1 U19567 ( .A(n19458), .B(n19457), .ZN(Ciphertext[187]) );
  INV_X1 U19568 ( .A(n19459), .ZN(n19465) );
  INV_X1 U19569 ( .A(n19460), .ZN(n19461) );
  OAI21_X1 U19570 ( .B1(n19463), .B2(n19462), .A(n19461), .ZN(n19464) );
  AOI22_X1 U19571 ( .A1(n19466), .A2(n19465), .B1(n19464), .B2(n212), .ZN(
        n19468) );
  XNOR2_X1 U19572 ( .A(n19468), .B(n19467), .ZN(Ciphertext[191]) );
  NAND3_X2 U8160 ( .A1(n3556), .A2(n3553), .A3(n3552), .ZN(n9635) );
  NOR2_X2 U1007 ( .A1(n8164), .A2(n8163), .ZN(n9070) );
  MUX2_X2 U1001 ( .A(n11878), .B(n11877), .S(n12577), .Z(n13848) );
  XNOR2_X2 U4182 ( .A(n5166), .B(n5165), .ZN(n2792) );
  INV_X1 U281 ( .A(n15479), .ZN(n17909) );
  MUX2_X2 U68 ( .A(n4195), .B(n4194), .S(n4370), .Z(n5424) );
  NOR2_X2 U257 ( .A1(n11542), .A2(n11543), .ZN(n12029) );
  OR2_X2 U1842 ( .A1(n2876), .A2(n2880), .ZN(n7202) );
  NOR2_X1 U851 ( .A1(n12223), .A2(n10925), .ZN(n12121) );
  AOI21_X1 U1550 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n11830) );
  BUF_X2 U1449 ( .A(n14626), .Z(n954) );
  BUF_X1 U1116 ( .A(n5762), .Z(n8205) );
  BUF_X2 U8440 ( .A(n16673), .Z(n19349) );
  BUF_X1 U1649 ( .A(n11389), .Z(n11870) );
  INV_X1 U739 ( .A(n9391), .ZN(n10594) );
  OR2_X2 U1763 ( .A1(n427), .A2(n3625), .ZN(n9029) );
  NAND2_X1 U79 ( .A1(n615), .A2(n446), .ZN(n6782) );
  NAND3_X2 U10038 ( .A1(n5549), .A2(n5547), .A3(n5548), .ZN(n7155) );
  CLKBUF_X1 U2021 ( .A(Key[117]), .Z(n19102) );
  XNOR2_X1 U981 ( .A(Key[155]), .B(Plaintext[155]), .ZN(n4567) );
  XNOR2_X1 U2030 ( .A(Plaintext[136]), .B(Key[136]), .ZN(n4271) );
  CLKBUF_X1 U2014 ( .A(Key[6]), .Z(n18691) );
  XNOR2_X1 U512 ( .A(Key[30]), .B(Plaintext[30]), .ZN(n4911) );
  XNOR2_X1 U436 ( .A(Key[26]), .B(Plaintext[26]), .ZN(n4945) );
  XNOR2_X1 U1981 ( .A(Key[25]), .B(Plaintext[25]), .ZN(n4940) );
  BUF_X1 U8874 ( .A(n4518), .Z(n4523) );
  XNOR2_X1 U539 ( .A(n3857), .B(Key[90]), .ZN(n5095) );
  AND2_X1 U9103 ( .A1(n4940), .A2(n4118), .ZN(n4886) );
  XNOR2_X1 U955 ( .A(n3971), .B(Key[40]), .ZN(n4962) );
  XNOR2_X1 U154 ( .A(n3844), .B(Key[82]), .ZN(n5115) );
  BUF_X1 U3464 ( .A(n4152), .Z(n4546) );
  OAI211_X1 U121 ( .C1(n4290), .C2(n4018), .A(n4017), .B(n4627), .ZN(n5322) );
  OR2_X1 U1946 ( .A1(n4041), .A2(n4769), .ZN(n5034) );
  OR2_X1 U1914 ( .A1(n3886), .A2(n3885), .ZN(n1776) );
  AND2_X1 U5819 ( .A1(n3550), .A2(n3549), .ZN(n1807) );
  AND2_X1 U416 ( .A1(n4086), .A2(n4085), .ZN(n6000) );
  NAND2_X1 U546 ( .A1(n643), .A2(n664), .ZN(n5803) );
  MUX2_X1 U557 ( .A(n3955), .B(n3954), .S(n4609), .Z(n5573) );
  INV_X1 U8512 ( .A(n5148), .ZN(n5582) );
  NAND2_X1 U244 ( .A1(n1985), .A2(n4292), .ZN(n5628) );
  INV_X1 U466 ( .A(n5264), .ZN(n6143) );
  NAND2_X1 U510 ( .A1(n3262), .A2(n5522), .ZN(n5973) );
  OR2_X1 U630 ( .A1(n4183), .A2(n4184), .ZN(n6708) );
  INV_X1 U420 ( .A(n7188), .ZN(n6427) );
  OAI21_X1 U5974 ( .B1(n5566), .B2(n1895), .A(n1894), .ZN(n7382) );
  OR2_X1 U6480 ( .A1(n5131), .A2(n5130), .ZN(n7144) );
  OAI21_X1 U745 ( .B1(n6063), .B2(n6064), .A(n6062), .ZN(n7017) );
  XNOR2_X1 U10555 ( .A(n6477), .B(n7253), .ZN(n6660) );
  NAND3_X1 U1831 ( .A1(n2396), .A2(n2099), .A3(n2098), .ZN(n7151) );
  XNOR2_X1 U818 ( .A(n7322), .B(n7321), .ZN(n8325) );
  XNOR2_X1 U11019 ( .A(n6930), .B(n6929), .ZN(n8165) );
  XNOR2_X1 U864 ( .A(n6006), .B(n6005), .ZN(n8197) );
  XNOR2_X1 U10975 ( .A(n6870), .B(n6869), .ZN(n8352) );
  BUF_X1 U349 ( .A(n7877), .Z(n8044) );
  OAI211_X1 U10917 ( .C1(n8385), .C2(n6800), .A(n6799), .B(n7685), .ZN(n9310)
         );
  OAI21_X1 U11588 ( .B1(n7694), .B2(n7693), .A(n7692), .ZN(n8904) );
  OR2_X1 U10816 ( .A1(n6654), .A2(n6653), .ZN(n9189) );
  NAND4_X2 U282 ( .A1(n3719), .A2(n5299), .A3(n3718), .A4(n5298), .ZN(n1037)
         );
  NAND3_X1 U1112 ( .A1(n3311), .A2(n8255), .A3(n769), .ZN(n9130) );
  INV_X1 U3832 ( .A(n8797), .ZN(n9112) );
  INV_X1 U1710 ( .A(n670), .ZN(n9256) );
  OR2_X1 U1713 ( .A1(n8611), .A2(n7537), .ZN(n8698) );
  OR3_X1 U3524 ( .A1(n8649), .A2(n8991), .A3(n20265), .ZN(n2887) );
  NAND3_X1 U6214 ( .A1(n2015), .A2(n8629), .A3(n2014), .ZN(n10582) );
  OAI211_X1 U870 ( .C1(n2651), .C2(n2650), .A(n8412), .B(n2652), .ZN(n10425)
         );
  INV_X1 U1673 ( .A(n10237), .ZN(n9994) );
  XNOR2_X1 U2595 ( .A(n20156), .B(n10046), .ZN(n10347) );
  XNOR2_X1 U849 ( .A(n9522), .B(n9521), .ZN(n10960) );
  XNOR2_X1 U12608 ( .A(n9474), .B(n9473), .ZN(n11148) );
  XNOR2_X1 U8115 ( .A(n9907), .B(n9906), .ZN(n3507) );
  BUF_X1 U814 ( .A(n11087), .Z(n11454) );
  NAND3_X1 U615 ( .A1(n576), .A2(n9199), .A3(n9200), .ZN(n12354) );
  NAND2_X1 U604 ( .A1(n11288), .A2(n19972), .ZN(n12811) );
  NAND2_X1 U2177 ( .A1(n3489), .A2(n10949), .ZN(n12126) );
  NAND3_X1 U2087 ( .A1(n9485), .A2(n3381), .A3(n2045), .ZN(n12180) );
  OAI21_X1 U14040 ( .B1(n11434), .B2(n11433), .A(n11432), .ZN(n12167) );
  OAI211_X1 U7470 ( .C1(n11250), .C2(n11383), .A(n11249), .B(n11384), .ZN(
        n12372) );
  NAND3_X1 U1547 ( .A1(n1278), .A2(n766), .A3(n765), .ZN(n11942) );
  OR2_X1 U415 ( .A1(n11995), .A2(n11997), .ZN(n12322) );
  OR2_X1 U115 ( .A1(n12534), .A2(n12532), .ZN(n12293) );
  OR2_X1 U3010 ( .A1(n12492), .A2(n253), .ZN(n12813) );
  NOR2_X1 U14580 ( .A1(n12327), .A2(n12514), .ZN(n13269) );
  AND3_X1 U2716 ( .A1(n1828), .A2(n1827), .A3(n609), .ZN(n13427) );
  NAND3_X1 U609 ( .A1(n2148), .A2(n12144), .A3(n2147), .ZN(n13644) );
  XNOR2_X1 U135 ( .A(n12626), .B(n12625), .ZN(n14791) );
  XNOR2_X1 U904 ( .A(n13548), .B(n13547), .ZN(n14482) );
  XNOR2_X1 U7204 ( .A(n2624), .B(n2623), .ZN(n14236) );
  XNOR2_X1 U189 ( .A(n13516), .B(n13515), .ZN(n14487) );
  XNOR2_X1 U338 ( .A(n1973), .B(n13349), .ZN(n14693) );
  XNOR2_X1 U15104 ( .A(n13024), .B(n13023), .ZN(n14506) );
  OR2_X1 U611 ( .A1(n14693), .A2(n200), .ZN(n14696) );
  NAND4_X1 U15972 ( .A1(n14253), .A2(n14254), .A3(n14255), .A4(n14252), .ZN(
        n15531) );
  AOI21_X1 U927 ( .B1(n14301), .B2(n14508), .A(n14300), .ZN(n14902) );
  OAI21_X1 U471 ( .B1(n13671), .B2(n14247), .A(n14246), .ZN(n15921) );
  NOR2_X1 U6095 ( .A1(n15458), .A2(n20173), .ZN(n15239) );
  NOR2_X1 U16897 ( .A1(n230), .A2(n868), .ZN(n15851) );
  AND2_X1 U4890 ( .A1(n1217), .A2(n1220), .ZN(n17328) );
  AND4_X1 U4152 ( .A1(n15668), .A2(n1018), .A3(n15669), .A4(n15670), .ZN(n955)
         );
  XNOR2_X1 U6147 ( .A(n16958), .B(n16957), .ZN(n17812) );
  XNOR2_X1 U6801 ( .A(n16218), .B(n16217), .ZN(n17489) );
  XNOR2_X1 U111 ( .A(n14634), .B(n14633), .ZN(n17508) );
  BUF_X1 U834 ( .A(n18092), .Z(n160) );
  BUF_X1 U317 ( .A(n16263), .Z(n17079) );
  XNOR2_X1 U140 ( .A(n16235), .B(n16234), .ZN(n17492) );
  CLKBUF_X1 U116 ( .A(n16805), .Z(n17959) );
  AOI21_X1 U3674 ( .B1(n2335), .B2(n17510), .A(n16634), .ZN(n18342) );
  AOI22_X1 U18029 ( .A1(n17086), .A2(n17602), .B1(n17085), .B2(n17601), .ZN(
        n18306) );
  AND3_X1 U18017 ( .A1(n17073), .A2(n17072), .A3(n17071), .ZN(n19162) );
  NOR2_X1 U6415 ( .A1(n16815), .A2(n16814), .ZN(n18529) );
  OR2_X1 U17153 ( .A1(n16114), .A2(n16113), .ZN(n19170) );
  AOI21_X1 U81 ( .B1(n17230), .B2(n17510), .A(n17229), .ZN(n18392) );
  XNOR2_X1 U283 ( .A(Key[61]), .B(Plaintext[61]), .ZN(n4651) );
  CLKBUF_X1 U567 ( .A(Key[186]), .Z(n106) );
  CLKBUF_X1 U1199 ( .A(Key[156]), .Z(n2306) );
  XNOR2_X1 U2368 ( .A(n3908), .B(Key[156]), .ZN(n4571) );
  INV_X1 U6122 ( .A(n5107), .ZN(n3259) );
  XNOR2_X1 U5154 ( .A(n6797), .B(n6798), .ZN(n8386) );
  INV_X1 U9776 ( .A(n8301), .ZN(n8046) );
  NAND2_X1 U6706 ( .A1(n7871), .A2(n7615), .ZN(n7618) );
  AND2_X1 U6895 ( .A1(n7888), .A2(n7887), .ZN(n9275) );
  INV_X1 U13968 ( .A(n12021), .ZN(n12369) );
  NAND2_X1 U1003 ( .A1(n11809), .A2(n11810), .ZN(n12212) );
  AOI21_X2 U10 ( .B1(n14259), .B2(n15421), .A(n14258), .ZN(n16836) );
  XNOR2_X2 U16959 ( .A(n15942), .B(n15941), .ZN(n17823) );
  BUF_X2 U4245 ( .A(n14000), .Z(n14620) );
  XNOR2_X2 U826 ( .A(n4035), .B(Key[132]), .ZN(n4095) );
  NAND2_X2 U907 ( .A1(n597), .A2(n599), .ZN(n10349) );
  NAND4_X2 U1872 ( .A1(n5609), .A2(n5607), .A3(n5608), .A4(n5606), .ZN(n6558)
         );
  AND4_X2 U1684 ( .A1(n8788), .A2(n8787), .A3(n3466), .A4(n3465), .ZN(n9771)
         );
  NAND2_X2 U2350 ( .A1(n445), .A2(n1483), .ZN(n7333) );
  AND3_X2 U117 ( .A1(n344), .A2(n11369), .A3(n11368), .ZN(n12312) );
  NAND3_X2 U7799 ( .A1(n3191), .A2(n4672), .A3(n3192), .ZN(n6171) );
  MUX2_X2 U6207 ( .A(n8406), .B(n8405), .S(n9164), .Z(n9794) );
  MUX2_X2 U1679 ( .A(n7806), .B(n7805), .S(n2243), .Z(n10262) );
  AND2_X2 U1743 ( .A1(n2259), .A2(n2258), .ZN(n9159) );
  AND2_X2 U184 ( .A1(n7698), .A2(n7697), .ZN(n8720) );
  OAI21_X2 U771 ( .B1(n4751), .B2(n4750), .A(n4749), .ZN(n5172) );
  BUF_X2 U1650 ( .A(n9492), .Z(n10649) );
  AND2_X2 U253 ( .A1(n9497), .A2(n9496), .ZN(n11673) );
  NOR2_X2 U7979 ( .A1(n14786), .A2(n14785), .ZN(n15582) );
  OAI211_X2 U2865 ( .C1(n2888), .C2(n9278), .A(n2887), .B(n702), .ZN(n10185)
         );
  AND3_X2 U1492 ( .A1(n3531), .A2(n1641), .A3(n1020), .ZN(n12713) );
  NOR2_X2 U580 ( .A1(n9047), .A2(n9048), .ZN(n9289) );
  BUF_X2 U14 ( .A(n12658), .Z(n15766) );
  OAI211_X2 U702 ( .C1(n15264), .C2(n15265), .A(n15263), .B(n15262), .ZN(
        n16987) );
  OR3_X1 U8469 ( .A1(n14599), .A2(n14603), .A3(n19918), .ZN(n3815) );
  AND3_X1 U3 ( .A1(n17065), .A2(n17718), .A3(n17064), .ZN(n19163) );
  AOI211_X1 U4 ( .C1(n14449), .C2(n14453), .A(n13927), .B(n14452), .ZN(n12929)
         );
  XNOR2_X1 U7 ( .A(n10184), .B(n10183), .ZN(n19830) );
  NOR2_X2 U120 ( .A1(n11811), .A2(n11638), .ZN(n12207) );
  OAI211_X2 U137 ( .C1(n7682), .C2(n8166), .A(n7681), .B(n7680), .ZN(n19941)
         );
  OAI22_X1 U151 ( .A1(n14342), .A2(n13931), .B1(n14335), .B2(n12879), .ZN(
        n14050) );
  NOR2_X1 U153 ( .A1(n18741), .A2(n18775), .ZN(n18746) );
  INV_X1 U155 ( .A(n16665), .ZN(n1897) );
  INV_X1 U187 ( .A(n2684), .ZN(n3223) );
  XOR2_X1 U198 ( .A(n17422), .B(n17421), .Z(n19472) );
  BUF_X2 U201 ( .A(n14325), .Z(n14352) );
  XNOR2_X1 U226 ( .A(n6210), .B(n3805), .ZN(n8195) );
  BUF_X1 U245 ( .A(n6381), .Z(n19476) );
  AOI21_X1 U252 ( .B1(n4718), .B2(n4717), .A(n4716), .ZN(n6381) );
  XNOR2_X2 U264 ( .A(n12853), .B(n12852), .ZN(n14449) );
  BUF_X1 U293 ( .A(n16921), .Z(n19860) );
  AND3_X2 U325 ( .A1(n3324), .A2(n3325), .A3(n3566), .ZN(n12506) );
  XNOR2_X1 U363 ( .A(n9511), .B(n9510), .ZN(n11144) );
  NOR2_X2 U365 ( .A1(n3677), .A2(n7467), .ZN(n8550) );
  AND3_X2 U381 ( .A1(n11916), .A2(n3161), .A3(n3160), .ZN(n12470) );
  XNOR2_X2 U422 ( .A(n10308), .B(n10307), .ZN(n11255) );
  XNOR2_X1 U484 ( .A(n12779), .B(n12778), .ZN(n12800) );
  XNOR2_X2 U507 ( .A(Key[98]), .B(Plaintext[98]), .ZN(n5075) );
  NAND2_X2 U520 ( .A1(n3622), .A2(n393), .ZN(n5668) );
  XNOR2_X2 U533 ( .A(Key[51]), .B(Plaintext[51]), .ZN(n4856) );
  XNOR2_X2 U579 ( .A(n3923), .B(Key[170]), .ZN(n4343) );
  OAI211_X2 U623 ( .C1(n705), .C2(n708), .A(n706), .B(n704), .ZN(n10506) );
  XNOR2_X2 U625 ( .A(n11936), .B(n11935), .ZN(n19875) );
  AND3_X2 U652 ( .A1(n1673), .A2(n1710), .A3(n1711), .ZN(n11586) );
  OAI211_X1 U665 ( .C1(n7840), .C2(n8910), .A(n7839), .B(n7838), .ZN(n9009) );
  BUF_X2 U674 ( .A(n16321), .Z(n18539) );
  XNOR2_X2 U675 ( .A(n3921), .B(Key[169]), .ZN(n4517) );
  CLKBUF_X1 U685 ( .A(n10575), .Z(n11499) );
  XNOR2_X2 U716 ( .A(Key[111]), .B(Plaintext[111]), .ZN(n5087) );
  INV_X1 U724 ( .A(n5095), .ZN(n4788) );
  XNOR2_X2 U751 ( .A(Key[152]), .B(Plaintext[152]), .ZN(n4752) );
  NAND2_X2 U754 ( .A1(n5157), .A2(n499), .ZN(n7364) );
  XNOR2_X2 U822 ( .A(n10479), .B(n10478), .ZN(n11034) );
  XNOR2_X2 U839 ( .A(n1285), .B(n9599), .ZN(n11292) );
  OAI211_X2 U847 ( .C1(n2846), .C2(n11160), .A(n2842), .B(n19570), .ZN(n1508)
         );
  XNOR2_X2 U862 ( .A(Key[146]), .B(Plaintext[146]), .ZN(n4744) );
  OAI211_X2 U871 ( .C1(n5831), .C2(n6018), .A(n5830), .B(n5829), .ZN(n7154) );
  OAI21_X2 U876 ( .B1(n11268), .B2(n11336), .A(n602), .ZN(n12374) );
  XNOR2_X1 U893 ( .A(n12743), .B(n12744), .ZN(n14347) );
  XNOR2_X2 U906 ( .A(n3153), .B(Key[143]), .ZN(n4555) );
  OAI21_X2 U919 ( .B1(n15151), .B2(n15150), .A(n15149), .ZN(n16900) );
  XNOR2_X2 U920 ( .A(n4028), .B(Key[114]), .ZN(n4697) );
  INV_X1 U944 ( .A(n18376), .ZN(n19501) );
  NAND2_X1 U949 ( .A1(n1844), .A2(n16255), .ZN(n18495) );
  NOR2_X1 U953 ( .A1(n16658), .A2(n17208), .ZN(n17217) );
  OR2_X1 U958 ( .A1(n15400), .A2(n15892), .ZN(n14285) );
  INV_X1 U961 ( .A(n14700), .ZN(n19503) );
  INV_X1 U969 ( .A(n12372), .ZN(n19504) );
  INV_X1 U976 ( .A(n4970), .ZN(n19507) );
  OR2_X1 U1011 ( .A1(n16249), .A2(n16248), .ZN(n19729) );
  NOR2_X1 U1013 ( .A1(n20214), .A2(n19098), .ZN(n19113) );
  NOR2_X1 U1016 ( .A1(n18781), .A2(n18741), .ZN(n19551) );
  AND4_X1 U1026 ( .A1(n3548), .A2(n3544), .A3(n3545), .A4(n3547), .ZN(n19681)
         );
  NOR2_X2 U1037 ( .A1(n16441), .A2(n16440), .ZN(n19775) );
  AND3_X1 U1053 ( .A1(n17073), .A2(n17072), .A3(n17071), .ZN(n19708) );
  NOR2_X1 U1059 ( .A1(n18136), .A2(n18135), .ZN(n19745) );
  INV_X1 U1073 ( .A(n18673), .ZN(n19510) );
  INV_X1 U1088 ( .A(n19390), .ZN(n19511) );
  XNOR2_X1 U1128 ( .A(n16204), .B(n16203), .ZN(n18534) );
  XNOR2_X1 U1268 ( .A(n17377), .B(n19640), .ZN(n16119) );
  INV_X1 U1282 ( .A(n15852), .ZN(n17433) );
  MUX2_X1 U1302 ( .A(n12936), .B(n12935), .S(n15380), .Z(n17104) );
  CLKBUF_X1 U1310 ( .A(n15502), .Z(n19813) );
  NAND2_X1 U1325 ( .A1(n19537), .A2(n14368), .ZN(n15905) );
  INV_X1 U1328 ( .A(n15502), .ZN(n19512) );
  OAI21_X1 U1330 ( .B1(n14365), .B2(n14364), .A(n19538), .ZN(n19537) );
  INV_X1 U1346 ( .A(n15709), .ZN(n19514) );
  OR2_X1 U1349 ( .A1(n2314), .A2(n14599), .ZN(n13855) );
  OR2_X1 U1352 ( .A1(n20513), .A2(n14599), .ZN(n14600) );
  AND2_X1 U1380 ( .A1(n11473), .A2(n11472), .ZN(n924) );
  OR2_X1 U1396 ( .A1(n8402), .A2(n8401), .ZN(n19769) );
  XNOR2_X1 U1402 ( .A(n10014), .B(n10015), .ZN(n11573) );
  OAI21_X1 U1424 ( .B1(n9564), .B2(n19590), .A(n2169), .ZN(n8415) );
  AND2_X1 U1453 ( .A1(n9249), .A2(n8974), .ZN(n3356) );
  AND2_X1 U1454 ( .A1(n477), .A2(n19550), .ZN(n8499) );
  AND2_X1 U1474 ( .A1(n8602), .A2(n8743), .ZN(n8483) );
  INV_X1 U1486 ( .A(n9106), .ZN(n19515) );
  INV_X1 U1498 ( .A(n8974), .ZN(n19516) );
  OR2_X1 U1500 ( .A1(n5965), .A2(n19579), .ZN(n19577) );
  INV_X1 U1502 ( .A(n8772), .ZN(n19517) );
  BUF_X2 U1508 ( .A(n8735), .Z(n19518) );
  INV_X1 U1517 ( .A(n8828), .ZN(n19519) );
  INV_X1 U1618 ( .A(n8384), .ZN(n19589) );
  INV_X1 U1621 ( .A(n7500), .ZN(n19651) );
  INV_X1 U1626 ( .A(n8316), .ZN(n19520) );
  INV_X1 U1629 ( .A(n7903), .ZN(n19521) );
  INV_X1 U1641 ( .A(n5410), .ZN(n5681) );
  INV_X1 U1645 ( .A(n5704), .ZN(n5996) );
  INV_X1 U1652 ( .A(n5382), .ZN(n6194) );
  INV_X1 U1663 ( .A(n6206), .ZN(n19522) );
  AND2_X1 U1746 ( .A1(n4609), .A2(n4177), .ZN(n19963) );
  XNOR2_X1 U1754 ( .A(n3870), .B(Key[34]), .ZN(n4952) );
  OR2_X1 U1755 ( .A1(n4319), .A2(n4324), .ZN(n4146) );
  INV_X1 U1765 ( .A(n4651), .ZN(n19523) );
  XNOR2_X1 U1766 ( .A(Key[135]), .B(Plaintext[135]), .ZN(n19788) );
  AND2_X1 U1768 ( .A1(n4467), .A2(n4887), .ZN(n4889) );
  BUF_X1 U1803 ( .A(n4041), .Z(n5032) );
  OR2_X1 U1832 ( .A1(n4204), .A2(n5010), .ZN(n19540) );
  CLKBUF_X1 U1848 ( .A(n4094), .Z(n5029) );
  XNOR2_X1 U1851 ( .A(Key[168]), .B(Plaintext[168]), .ZN(n4187) );
  AND2_X1 U1852 ( .A1(n6050), .A2(n3351), .ZN(n3665) );
  OR2_X1 U1855 ( .A1(n3959), .A2(n5405), .ZN(n5316) );
  OR2_X1 U1887 ( .A1(n5291), .A2(n5645), .ZN(n2321) );
  INV_X1 U1939 ( .A(n3351), .ZN(n6052) );
  OR2_X1 U1958 ( .A1(n5158), .A2(n5429), .ZN(n499) );
  XNOR2_X1 U2029 ( .A(n7230), .B(n7151), .ZN(n6495) );
  XNOR2_X1 U2048 ( .A(n7304), .B(n6348), .ZN(n6961) );
  XNOR2_X1 U2051 ( .A(n6789), .B(n6788), .ZN(n8132) );
  OR2_X1 U2088 ( .A1(n7932), .A2(n7931), .ZN(n1453) );
  OR2_X1 U2107 ( .A1(n7648), .A2(n8079), .ZN(n19622) );
  OR2_X1 U2108 ( .A1(n9242), .A2(n9189), .ZN(n431) );
  AND2_X1 U2109 ( .A1(n8304), .A2(n2792), .ZN(n1244) );
  CLKBUF_X1 U2116 ( .A(n8221), .Z(n19809) );
  AOI21_X1 U2135 ( .B1(n8382), .B2(n8381), .A(n19589), .ZN(n8391) );
  OAI211_X1 U2150 ( .C1(n7902), .C2(n7909), .A(n19582), .B(n7754), .ZN(n2251)
         );
  INV_X1 U2156 ( .A(n803), .ZN(n9211) );
  NOR3_X1 U2231 ( .A1(n9130), .A2(n9129), .A3(n9201), .ZN(n9131) );
  XNOR2_X1 U2232 ( .A(n9391), .B(n9392), .ZN(n10454) );
  NAND2_X1 U2235 ( .A1(n1398), .A2(n8425), .ZN(n694) );
  AND2_X1 U2267 ( .A1(n19878), .A2(n11174), .ZN(n19614) );
  CLKBUF_X1 U2282 ( .A(n11884), .Z(n909) );
  OR2_X1 U2283 ( .A1(n10945), .A2(n1654), .ZN(n19571) );
  AOI22_X1 U2317 ( .A1(n10828), .A2(n10827), .B1(n10826), .B2(n11041), .ZN(
        n12202) );
  OR2_X1 U2334 ( .A1(n12380), .A2(n12381), .ZN(n19592) );
  AOI21_X1 U2344 ( .B1(n10452), .B2(n10451), .A(n2656), .ZN(n10471) );
  BUF_X1 U2362 ( .A(n11769), .Z(n12528) );
  OAI21_X1 U2388 ( .B1(n11684), .B2(n11685), .A(n19585), .ZN(n19584) );
  INV_X1 U2421 ( .A(n2220), .ZN(n19535) );
  XNOR2_X1 U2424 ( .A(n13539), .B(n13716), .ZN(n13771) );
  XNOR2_X1 U2425 ( .A(n13312), .B(n13791), .ZN(n13483) );
  INV_X1 U2432 ( .A(n2684), .ZN(n19598) );
  BUF_X1 U2438 ( .A(n14490), .Z(n14753) );
  INV_X1 U2439 ( .A(n14369), .ZN(n19538) );
  CLKBUF_X1 U2440 ( .A(n14779), .Z(n877) );
  XOR2_X1 U2446 ( .A(n13334), .B(n13333), .Z(n19895) );
  INV_X1 U2452 ( .A(n19634), .ZN(n19600) );
  AND2_X1 U2488 ( .A1(n3431), .A2(n15606), .ZN(n19542) );
  NAND2_X1 U2514 ( .A1(n13978), .A2(n2353), .ZN(n15874) );
  AND2_X1 U2515 ( .A1(n2288), .A2(n15503), .ZN(n3019) );
  OR2_X1 U2519 ( .A1(n14786), .A2(n14785), .ZN(n19958) );
  BUF_X1 U2525 ( .A(n15746), .Z(n15182) );
  OR2_X1 U2544 ( .A1(n14961), .A2(n15287), .ZN(n19573) );
  AND2_X1 U2613 ( .A1(n15875), .A2(n15714), .ZN(n15146) );
  OR3_X1 U2668 ( .A1(n19888), .A2(n19583), .A3(n15470), .ZN(n1075) );
  OR2_X1 U2714 ( .A1(n15467), .A2(n15470), .ZN(n2358) );
  BUF_X1 U2747 ( .A(n17127), .Z(n19882) );
  CLKBUF_X1 U2762 ( .A(n17547), .Z(n19771) );
  NOR2_X1 U2764 ( .A1(n19974), .A2(n19744), .ZN(n18248) );
  XNOR2_X1 U2770 ( .A(n16710), .B(n16709), .ZN(n17818) );
  MUX2_X1 U2772 ( .A(n15269), .B(n15268), .S(n15846), .Z(n16691) );
  XNOR2_X1 U2778 ( .A(n16352), .B(n16351), .ZN(n18111) );
  OR2_X1 U2786 ( .A1(n17830), .A2(n219), .ZN(n18957) );
  AND2_X1 U2819 ( .A1(n17855), .A2(n17), .ZN(n15) );
  NAND2_X1 U2853 ( .A1(n17247), .A2(n17246), .ZN(n18384) );
  AND2_X1 U2858 ( .A1(n17452), .A2(n17453), .ZN(n18702) );
  OR2_X1 U2877 ( .A1(n17750), .A2(n18929), .ZN(n19574) );
  OR2_X1 U2901 ( .A1(n18064), .A2(n19035), .ZN(n2399) );
  OR2_X1 U2932 ( .A1(n18709), .A2(n18733), .ZN(n18736) );
  OAI21_X1 U3018 ( .B1(n17177), .B2(n17176), .A(n17175), .ZN(n19105) );
  OAI211_X1 U3064 ( .C1(n18381), .C2(n2274), .A(n18387), .B(n18386), .ZN(
        n19969) );
  CLKBUF_X1 U3101 ( .A(Key[39]), .Z(n18284) );
  CLKBUF_X1 U3109 ( .A(Key[123]), .Z(n18075) );
  CLKBUF_X1 U3117 ( .A(Key[75]), .Z(n17851) );
  XOR2_X1 U3122 ( .A(n18749), .B(n2381), .Z(n19525) );
  AND3_X1 U3137 ( .A1(n3085), .A2(n975), .A3(n17506), .ZN(n19526) );
  NAND3_X1 U3146 ( .A1(n12525), .A2(n3256), .A3(n182), .ZN(n19527) );
  INV_X1 U3166 ( .A(n9837), .ZN(n19606) );
  AND2_X1 U3168 ( .A1(n4500), .A2(n409), .ZN(n5841) );
  INV_X1 U3180 ( .A(n5841), .ZN(n19968) );
  AOI22_X1 U3239 ( .A1(n4139), .A2(n4962), .B1(n4377), .B2(n4138), .ZN(n5524)
         );
  AND2_X1 U3256 ( .A1(n7528), .A2(n7908), .ZN(n19528) );
  INV_X1 U3267 ( .A(n5435), .ZN(n19562) );
  INV_X1 U3277 ( .A(n5798), .ZN(n5429) );
  INV_X1 U3296 ( .A(n9780), .ZN(n19553) );
  INV_X1 U3315 ( .A(n7788), .ZN(n19579) );
  AND2_X1 U3328 ( .A1(n7562), .A2(n6705), .ZN(n19529) );
  XOR2_X1 U3330 ( .A(n13112), .B(n13113), .Z(n19530) );
  XNOR2_X1 U3342 ( .A(n12954), .B(n12953), .ZN(n14641) );
  XOR2_X1 U3380 ( .A(n12712), .B(n13457), .Z(n19531) );
  AND2_X1 U3392 ( .A1(n20221), .A2(n18953), .ZN(n19532) );
  INV_X1 U3434 ( .A(n18656), .ZN(n19624) );
  AND3_X1 U3469 ( .A1(n18737), .A2(n18736), .A3(n18735), .ZN(n19533) );
  OR2_X1 U3527 ( .A1(n19286), .A2(n19285), .ZN(n19534) );
  NAND2_X1 U3583 ( .A1(n19536), .A2(n19535), .ZN(n12914) );
  NAND2_X1 U3702 ( .A1(n12297), .A2(n12296), .ZN(n19536) );
  NAND2_X1 U3709 ( .A1(n4248), .A2(n19540), .ZN(n19539) );
  NAND2_X1 U3722 ( .A1(n17217), .A2(n19541), .ZN(n16467) );
  NAND2_X1 U3756 ( .A1(n20135), .A2(n17211), .ZN(n19541) );
  NOR2_X1 U3769 ( .A1(n19542), .A2(n20007), .ZN(n14976) );
  NAND2_X1 U3870 ( .A1(n4570), .A2(n4370), .ZN(n4509) );
  NAND2_X1 U3892 ( .A1(n12569), .A2(n12570), .ZN(n12571) );
  OAI211_X1 U3916 ( .C1(n14227), .C2(n20376), .A(n19543), .B(n14412), .ZN(
        n2903) );
  NAND2_X1 U3949 ( .A1(n13403), .A2(n14408), .ZN(n19543) );
  NAND3_X1 U4009 ( .A1(n20464), .A2(n4697), .A3(n5040), .ZN(n19544) );
  NOR2_X1 U4053 ( .A1(n20535), .A2(n18869), .ZN(n18853) );
  NAND2_X1 U4119 ( .A1(n2891), .A2(n14703), .ZN(n14380) );
  XNOR2_X1 U4122 ( .A(n17366), .B(n18308), .ZN(n16145) );
  XNOR2_X1 U4183 ( .A(n10286), .B(n9802), .ZN(n9756) );
  NAND2_X1 U4191 ( .A1(n7577), .A2(n7576), .ZN(n9802) );
  NAND2_X1 U4342 ( .A1(n19740), .A2(n192), .ZN(n15705) );
  NAND2_X1 U4369 ( .A1(n2659), .A2(n17149), .ZN(n3235) );
  NAND3_X1 U4370 ( .A1(n2782), .A2(n2781), .A3(n2989), .ZN(n19638) );
  NAND3_X1 U4404 ( .A1(n233), .A2(n15815), .A3(n228), .ZN(n3374) );
  NAND2_X1 U4407 ( .A1(n19547), .A2(n19546), .ZN(n10700) );
  NAND2_X1 U4452 ( .A1(n11292), .A2(n10697), .ZN(n19546) );
  NAND2_X1 U4453 ( .A1(n10696), .A2(n10978), .ZN(n19547) );
  NAND2_X1 U4456 ( .A1(n19549), .A2(n19548), .ZN(n15852) );
  NAND2_X1 U4483 ( .A1(n15408), .A2(n15407), .ZN(n19548) );
  NAND2_X1 U4518 ( .A1(n2791), .A2(n15616), .ZN(n19549) );
  NOR2_X1 U4533 ( .A1(n19528), .A2(n7531), .ZN(n19550) );
  AOI21_X1 U4566 ( .B1(n19525), .B2(n19803), .A(n19551), .ZN(n19650) );
  INV_X1 U4665 ( .A(n4144), .ZN(n4398) );
  NAND2_X1 U4676 ( .A1(n4144), .A2(n4141), .ZN(n4143) );
  NAND2_X1 U4683 ( .A1(n4914), .A2(n4140), .ZN(n4144) );
  NAND2_X1 U4689 ( .A1(n14828), .A2(n3223), .ZN(n2685) );
  NAND2_X1 U4690 ( .A1(n11348), .A2(n11349), .ZN(n11352) );
  NAND2_X1 U4698 ( .A1(n19554), .A2(n19552), .ZN(n8666) );
  NAND2_X1 U4734 ( .A1(n9782), .A2(n19553), .ZN(n19552) );
  NAND2_X1 U4737 ( .A1(n9779), .A2(n9780), .ZN(n19554) );
  NAND2_X1 U4742 ( .A1(n12151), .A2(n20618), .ZN(n19555) );
  NOR2_X1 U4745 ( .A1(n12157), .A2(n19558), .ZN(n19557) );
  NAND2_X1 U4768 ( .A1(n9068), .A2(n2504), .ZN(n2502) );
  NAND2_X1 U4819 ( .A1(n5014), .A2(n4555), .ZN(n4737) );
  NAND2_X1 U4914 ( .A1(n19562), .A2(n5704), .ZN(n19561) );
  OR2_X2 U4941 ( .A1(n4078), .A2(n4079), .ZN(n5704) );
  OAI21_X1 U4942 ( .B1(n20479), .B2(n19564), .A(n19563), .ZN(n10648) );
  NAND2_X1 U4945 ( .A1(n10968), .A2(n11559), .ZN(n19563) );
  NAND2_X1 U5040 ( .A1(n9274), .A2(n20265), .ZN(n19565) );
  NAND2_X1 U5072 ( .A1(n6166), .A2(n6172), .ZN(n6170) );
  NAND2_X1 U5092 ( .A1(n19568), .A2(n19566), .ZN(n10647) );
  NAND2_X1 U5108 ( .A1(n10646), .A2(n19567), .ZN(n19566) );
  INV_X1 U5139 ( .A(n10968), .ZN(n19567) );
  NAND2_X1 U5167 ( .A1(n11553), .A2(n9017), .ZN(n10646) );
  NAND2_X1 U5170 ( .A1(n10645), .A2(n10968), .ZN(n19568) );
  NAND2_X1 U5173 ( .A1(n19569), .A2(n4570), .ZN(n4259) );
  NAND2_X1 U5177 ( .A1(n4573), .A2(n4507), .ZN(n19569) );
  NAND3_X1 U5235 ( .A1(n607), .A2(n11160), .A3(n19571), .ZN(n19570) );
  NAND2_X1 U5300 ( .A1(n20012), .A2(n8282), .ZN(n7601) );
  NAND2_X1 U5313 ( .A1(n328), .A2(n3704), .ZN(n15081) );
  NAND2_X1 U5324 ( .A1(n2768), .A2(n2766), .ZN(n328) );
  NAND2_X1 U5359 ( .A1(n2414), .A2(n17866), .ZN(n19238) );
  OR2_X1 U5360 ( .A1(n10246), .A2(n11886), .ZN(n2130) );
  NAND2_X1 U5361 ( .A1(n9018), .A2(n9295), .ZN(n9299) );
  OR2_X2 U5392 ( .A1(n3261), .A2(n8514), .ZN(n8676) );
  NAND2_X1 U5408 ( .A1(n16782), .A2(n16783), .ZN(n1559) );
  NAND2_X1 U5447 ( .A1(n17069), .A2(n17896), .ZN(n16783) );
  NAND2_X1 U5546 ( .A1(n213), .A2(n18797), .ZN(n2179) );
  MUX2_X1 U5549 ( .A(n6195), .B(n6196), .S(n5382), .Z(n6197) );
  NAND2_X1 U5592 ( .A1(n14287), .A2(n241), .ZN(n1976) );
  NAND3_X1 U5678 ( .A1(n114), .A2(n20128), .A3(n18037), .ZN(n19575) );
  OR2_X2 U5745 ( .A1(n4316), .A2(n19576), .ZN(n5633) );
  NAND2_X1 U5751 ( .A1(n4314), .A2(n4362), .ZN(n19576) );
  NAND2_X1 U5761 ( .A1(n12203), .A2(n125), .ZN(n1190) );
  AND2_X1 U5774 ( .A1(n14032), .A2(n14637), .ZN(n13985) );
  NAND2_X1 U5832 ( .A1(n19579), .A2(n8299), .ZN(n19578) );
  NAND2_X1 U5837 ( .A1(n885), .A2(n8990), .ZN(n9272) );
  NAND2_X1 U5865 ( .A1(n2539), .A2(n2538), .ZN(n19580) );
  NAND2_X1 U5869 ( .A1(n4441), .A2(n2670), .ZN(n1922) );
  NAND2_X1 U5928 ( .A1(n4160), .A2(n4524), .ZN(n19581) );
  INV_X1 U5949 ( .A(n15468), .ZN(n19583) );
  NAND2_X1 U5953 ( .A1(n19584), .A2(n11688), .ZN(n13622) );
  INV_X1 U5990 ( .A(n12576), .ZN(n19585) );
  NOR2_X1 U6016 ( .A1(n19601), .A2(n19600), .ZN(n13973) );
  OAI211_X2 U6017 ( .C1(n16778), .C2(n17176), .A(n19587), .B(n19586), .ZN(
        n19144) );
  NAND2_X1 U6034 ( .A1(n3293), .A2(n20239), .ZN(n19586) );
  NAND2_X1 U6073 ( .A1(n16777), .A2(n19667), .ZN(n19587) );
  NAND2_X1 U6109 ( .A1(n1471), .A2(n11831), .ZN(n13843) );
  NAND2_X1 U6139 ( .A1(n824), .A2(n823), .ZN(n8419) );
  NAND2_X1 U6193 ( .A1(n8003), .A2(n7591), .ZN(n7477) );
  XNOR2_X1 U6208 ( .A(n19588), .B(n19410), .ZN(n7217) );
  NAND2_X1 U6209 ( .A1(n5245), .A2(n5244), .ZN(n19588) );
  INV_X1 U6224 ( .A(n352), .ZN(n19590) );
  NAND3_X1 U6232 ( .A1(n771), .A2(n772), .A3(n8665), .ZN(n419) );
  OAI211_X1 U6248 ( .C1(n8354), .C2(n8359), .A(n19591), .B(n7504), .ZN(n6902)
         );
  NAND2_X1 U6287 ( .A1(n19651), .A2(n8354), .ZN(n19591) );
  NAND3_X1 U6289 ( .A1(n12379), .A2(n12378), .A3(n19592), .ZN(n13600) );
  NAND2_X1 U6342 ( .A1(n2333), .A2(n2332), .ZN(n12378) );
  NAND2_X1 U6356 ( .A1(n3560), .A2(n19593), .ZN(n1720) );
  NOR2_X1 U6382 ( .A1(n4865), .A2(n19523), .ZN(n19593) );
  XNOR2_X1 U6393 ( .A(n19594), .B(n18848), .ZN(n9761) );
  NAND3_X1 U6396 ( .A1(n8170), .A2(n8168), .A3(n8169), .ZN(n19594) );
  NAND2_X1 U6397 ( .A1(n9832), .A2(n11263), .ZN(n1132) );
  NAND2_X1 U6405 ( .A1(n755), .A2(n756), .ZN(n9832) );
  NAND2_X1 U6427 ( .A1(n20129), .A2(n18976), .ZN(n17310) );
  NAND2_X1 U6441 ( .A1(n8659), .A2(n8658), .ZN(n19595) );
  NAND2_X1 U6458 ( .A1(n3519), .A2(n8660), .ZN(n19596) );
  NAND2_X1 U6487 ( .A1(n8134), .A2(n8135), .ZN(n8136) );
  NOR2_X2 U6513 ( .A1(n2776), .A2(n8570), .ZN(n10254) );
  OAI22_X1 U6555 ( .A1(n20468), .A2(n12101), .B1(n11271), .B2(n10684), .ZN(
        n9659) );
  NOR2_X1 U6560 ( .A1(n19984), .A2(n19598), .ZN(n19597) );
  OAI21_X2 U6562 ( .B1(n3961), .B2(n5408), .A(n1182), .ZN(n7304) );
  OAI21_X2 U6592 ( .B1(n9933), .B2(n11522), .A(n9932), .ZN(n12004) );
  OR2_X1 U6607 ( .A1(n15179), .A2(n15181), .ZN(n19599) );
  OAI21_X1 U6610 ( .B1(n6020), .B2(n6021), .A(n19660), .ZN(n445) );
  NAND2_X1 U6626 ( .A1(n3246), .A2(n14522), .ZN(n19601) );
  NAND2_X1 U6645 ( .A1(n2529), .A2(n2530), .ZN(n2528) );
  NAND2_X1 U6670 ( .A1(n19602), .A2(n12641), .ZN(n12643) );
  NAND2_X1 U6686 ( .A1(n389), .A2(n12640), .ZN(n19602) );
  NAND2_X1 U6699 ( .A1(n2387), .A2(n2386), .ZN(n7624) );
  NAND2_X1 U6703 ( .A1(n12569), .A2(n12258), .ZN(n19603) );
  NAND2_X1 U6730 ( .A1(n2065), .A2(n8602), .ZN(n19604) );
  NAND2_X1 U6745 ( .A1(n3328), .A2(n348), .ZN(n3327) );
  NAND2_X1 U6754 ( .A1(n20504), .A2(n8064), .ZN(n1433) );
  OR2_X1 U6765 ( .A1(n14098), .A2(n14338), .ZN(n19607) );
  OAI21_X1 U6766 ( .B1(n14096), .B2(n14095), .A(n14094), .ZN(n19608) );
  OR2_X1 U6789 ( .A1(n14103), .A2(n14787), .ZN(n14063) );
  XNOR2_X1 U6803 ( .A(n19609), .B(n13135), .ZN(n3364) );
  XNOR2_X1 U6807 ( .A(n3365), .B(n13651), .ZN(n19609) );
  XNOR2_X1 U6822 ( .A(n19610), .B(n19103), .ZN(Ciphertext[128]) );
  NOR2_X2 U6844 ( .A1(n19611), .A2(n15640), .ZN(n16412) );
  NAND3_X1 U6860 ( .A1(n6055), .A2(n5785), .A3(n5891), .ZN(n3865) );
  NAND3_X1 U6863 ( .A1(n3838), .A2(n1137), .A3(n19612), .ZN(n5782) );
  NAND2_X1 U6890 ( .A1(n14223), .A2(n14224), .ZN(n14225) );
  NAND2_X1 U6904 ( .A1(n9063), .A2(n19805), .ZN(n2300) );
  NAND2_X1 U6917 ( .A1(n3072), .A2(n1765), .ZN(n9063) );
  NAND3_X1 U6924 ( .A1(n12572), .A2(n12017), .A3(n242), .ZN(n12019) );
  MUX2_X1 U6986 ( .A(n14823), .B(n14822), .S(n14821), .Z(n19613) );
  AOI21_X1 U7026 ( .B1(n10912), .B2(n9487), .A(n19614), .ZN(n9490) );
  NAND3_X1 U7028 ( .A1(n19615), .A2(n1009), .A3(n12562), .ZN(n11895) );
  NAND2_X1 U7030 ( .A1(n3733), .A2(n12262), .ZN(n19615) );
  OAI22_X1 U7039 ( .A1(n15817), .A2(n19958), .B1(n15816), .B2(n15815), .ZN(
        n2114) );
  NAND2_X1 U7058 ( .A1(n19617), .A2(n19616), .ZN(n5410) );
  NAND2_X1 U7065 ( .A1(n4889), .A2(n4888), .ZN(n19616) );
  NAND2_X1 U7098 ( .A1(n4891), .A2(n4890), .ZN(n19617) );
  NAND2_X1 U7103 ( .A1(n11951), .A2(n11598), .ZN(n11957) );
  NAND2_X1 U7109 ( .A1(n20367), .A2(n7480), .ZN(n7483) );
  XNOR2_X1 U7111 ( .A(n13768), .B(n13600), .ZN(n13282) );
  NOR2_X1 U7138 ( .A1(n10830), .A2(n11421), .ZN(n10831) );
  NAND2_X1 U7141 ( .A1(n385), .A2(n5893), .ZN(n7258) );
  OAI21_X1 U7160 ( .B1(n2120), .B2(n18024), .A(n19618), .ZN(n18027) );
  NAND2_X1 U7169 ( .A1(n18928), .A2(n18024), .ZN(n19618) );
  NAND2_X1 U7170 ( .A1(n7674), .A2(n8365), .ZN(n7510) );
  XNOR2_X2 U7171 ( .A(n6395), .B(n6394), .ZN(n7674) );
  NAND2_X1 U7172 ( .A1(n11604), .A2(n12416), .ZN(n11608) );
  NAND2_X1 U7179 ( .A1(n11603), .A2(n20350), .ZN(n11604) );
  MUX2_X1 U7242 ( .A(n4304), .B(n4303), .S(n4982), .Z(n19619) );
  OAI21_X1 U7244 ( .B1(n19110), .B2(n19532), .A(n19620), .ZN(n17712) );
  NAND2_X1 U7245 ( .A1(n19110), .A2(n17710), .ZN(n19620) );
  NAND3_X1 U7258 ( .A1(n3028), .A2(n3030), .A3(n20117), .ZN(n3027) );
  NAND3_X1 U7265 ( .A1(n19621), .A2(n3701), .A3(n2482), .ZN(n3700) );
  NAND3_X1 U7266 ( .A1(n286), .A2(n5746), .A3(n5745), .ZN(n19621) );
  NAND2_X1 U7275 ( .A1(n19623), .A2(n19622), .ZN(n3791) );
  NAND2_X1 U7280 ( .A1(n3793), .A2(n3795), .ZN(n19623) );
  NAND2_X1 U7288 ( .A1(n19625), .A2(n19624), .ZN(n18658) );
  NAND2_X1 U7289 ( .A1(n18648), .A2(n19935), .ZN(n19625) );
  XNOR2_X1 U7311 ( .A(n19627), .B(n19626), .ZN(Ciphertext[168]) );
  INV_X1 U7352 ( .A(n2455), .ZN(n19626) );
  NAND2_X1 U7363 ( .A1(n19633), .A2(n19629), .ZN(n19283) );
  INV_X1 U7372 ( .A(n19630), .ZN(n19629) );
  AOI21_X1 U7382 ( .B1(n19632), .B2(n19631), .A(n19400), .ZN(n19630) );
  NAND2_X1 U7448 ( .A1(n19391), .A2(n19390), .ZN(n19632) );
  NAND2_X1 U7462 ( .A1(n17618), .A2(n19400), .ZN(n19633) );
  INV_X1 U7468 ( .A(n951), .ZN(n19634) );
  XNOR2_X1 U7482 ( .A(n19635), .B(n3460), .ZN(n13007) );
  XNOR2_X1 U7487 ( .A(n13703), .B(n19796), .ZN(n19635) );
  XNOR2_X2 U7488 ( .A(n19637), .B(n19636), .ZN(n11234) );
  XNOR2_X1 U7492 ( .A(n10158), .B(n9864), .ZN(n19636) );
  XNOR2_X1 U7497 ( .A(n9992), .B(n9863), .ZN(n19637) );
  NAND2_X1 U7559 ( .A1(n332), .A2(n333), .ZN(n11345) );
  NAND3_X2 U7668 ( .A1(n19638), .A2(n6959), .A3(n6958), .ZN(n10249) );
  NAND2_X1 U7678 ( .A1(n19639), .A2(n1616), .ZN(n8977) );
  OAI21_X1 U7695 ( .B1(n8970), .B2(n1618), .A(n9252), .ZN(n19639) );
  OR2_X1 U7708 ( .A1(n11866), .A2(n11870), .ZN(n9776) );
  INV_X1 U7774 ( .A(n18691), .ZN(n19640) );
  NAND2_X1 U7796 ( .A1(n7820), .A2(n278), .ZN(n7521) );
  NAND2_X1 U7817 ( .A1(n19641), .A2(n7755), .ZN(n2259) );
  OAI22_X1 U7825 ( .A1(n7909), .A2(n6904), .B1(n19521), .B2(n7754), .ZN(n19641) );
  OAI21_X1 U7859 ( .B1(n249), .B2(n12354), .A(n12174), .ZN(n11656) );
  NAND2_X1 U7889 ( .A1(n12354), .A2(n12352), .ZN(n12174) );
  NAND2_X1 U7890 ( .A1(n7831), .A2(n7832), .ZN(n9007) );
  NAND2_X1 U7918 ( .A1(n19643), .A2(n19642), .ZN(n13743) );
  NAND2_X1 U7944 ( .A1(n13730), .A2(n14381), .ZN(n19642) );
  NAND2_X1 U7945 ( .A1(n13731), .A2(n19644), .ZN(n19643) );
  INV_X1 U7946 ( .A(n14381), .ZN(n19644) );
  OAI21_X1 U7953 ( .B1(n635), .B2(n19645), .A(n634), .ZN(n16580) );
  OAI21_X1 U7959 ( .B1(n20436), .B2(n19372), .A(n19646), .ZN(n19645) );
  INV_X1 U8004 ( .A(n19370), .ZN(n19647) );
  AOI21_X1 U8017 ( .B1(n19648), .B2(n11109), .A(n11106), .ZN(n10772) );
  NAND2_X1 U8041 ( .A1(n11429), .A2(n11041), .ZN(n19648) );
  OR2_X2 U8042 ( .A1(n9231), .A2(n9230), .ZN(n9987) );
  NAND3_X1 U8043 ( .A1(n19649), .A2(n18241), .A3(n18240), .ZN(n18246) );
  NAND2_X1 U8046 ( .A1(n20132), .A2(n18238), .ZN(n19649) );
  AOI21_X1 U8068 ( .B1(n19650), .B2(n19533), .A(n18747), .ZN(Ciphertext[80])
         );
  NAND3_X1 U8069 ( .A1(n2174), .A2(n9331), .A3(n8866), .ZN(n8867) );
  NAND2_X1 U8133 ( .A1(n19057), .A2(n19067), .ZN(n71) );
  NAND3_X1 U8141 ( .A1(n1812), .A2(n11113), .A3(n11452), .ZN(n1804) );
  BUF_X2 U8178 ( .A(n18287), .Z(n18362) );
  AND2_X1 U8196 ( .A1(n19163), .A2(n19162), .ZN(n17790) );
  XNOR2_X1 U8223 ( .A(n13112), .B(n13113), .ZN(n19652) );
  INV_X1 U8262 ( .A(n19069), .ZN(n19653) );
  NAND2_X1 U8281 ( .A1(n18944), .A2(n2062), .ZN(n19654) );
  OAI211_X2 U8361 ( .C1(n18633), .C2(n959), .A(n1069), .B(n1013), .ZN(n18592)
         );
  OAI211_X1 U8366 ( .C1(n17161), .C2(n16792), .A(n16791), .B(n18542), .ZN(
        n19655) );
  XOR2_X1 U8373 ( .A(n9842), .B(n10299), .Z(n8509) );
  XNOR2_X1 U8377 ( .A(n13057), .B(n13018), .ZN(n13457) );
  XNOR2_X1 U8385 ( .A(n12712), .B(n13457), .ZN(n19657) );
  XOR2_X1 U8405 ( .A(n9503), .B(n8548), .Z(n8567) );
  NAND2_X1 U8422 ( .A1(n18944), .A2(n2062), .ZN(n19001) );
  OAI21_X1 U8430 ( .B1(n3576), .B2(n13943), .A(n13942), .ZN(n19659) );
  OAI21_X1 U8434 ( .B1(n3576), .B2(n13943), .A(n13942), .ZN(n16974) );
  OR2_X1 U8444 ( .A1(n3569), .A2(n5823), .ZN(n19660) );
  AND2_X1 U8503 ( .A1(n16799), .A2(n16798), .ZN(n19661) );
  AOI22_X1 U8514 ( .A1(n14084), .A2(n20500), .B1(n14081), .B2(n14082), .ZN(
        n15515) );
  OR2_X1 U8562 ( .A1(n9241), .A2(n9240), .ZN(n19663) );
  CLKBUF_X1 U8597 ( .A(n18916), .Z(n19664) );
  NOR2_X1 U8652 ( .A1(n17153), .A2(n17152), .ZN(n19665) );
  NOR2_X1 U8654 ( .A1(n17153), .A2(n17152), .ZN(n18590) );
  OR2_X1 U8661 ( .A1(n12003), .A2(n1637), .ZN(n3239) );
  XNOR2_X1 U8664 ( .A(n16559), .B(n16558), .ZN(n19371) );
  XNOR2_X1 U8676 ( .A(n16065), .B(n16064), .ZN(n16308) );
  XOR2_X1 U8716 ( .A(n15953), .B(n15954), .Z(n19667) );
  CLKBUF_X1 U8737 ( .A(Key[173]), .Z(n19140) );
  OR2_X1 U8772 ( .A1(n17153), .A2(n17152), .ZN(n19669) );
  NOR2_X1 U8798 ( .A1(n19010), .A2(n19670), .ZN(n2050) );
  AND3_X1 U8810 ( .A1(n19011), .A2(n19654), .A3(n19687), .ZN(n19670) );
  XNOR2_X1 U8857 ( .A(n16399), .B(n16400), .ZN(n19672) );
  OAI21_X1 U8877 ( .B1(n17555), .B2(n18106), .A(n17554), .ZN(n19673) );
  XNOR2_X1 U8995 ( .A(n16223), .B(n16222), .ZN(n19675) );
  XNOR2_X1 U8998 ( .A(n16223), .B(n16222), .ZN(n17494) );
  OAI211_X1 U9068 ( .C1(n15807), .C2(n15808), .A(n15805), .B(n19966), .ZN(
        n16982) );
  INV_X1 U9122 ( .A(n15420), .ZN(n19676) );
  XNOR2_X1 U9125 ( .A(n16230), .B(n16229), .ZN(n17493) );
  XOR2_X1 U9224 ( .A(n17448), .B(n17447), .Z(n19678) );
  NAND2_X1 U9225 ( .A1(n17557), .A2(n2797), .ZN(n19679) );
  OAI21_X1 U9262 ( .B1(n18973), .B2(n220), .A(n18972), .ZN(n19680) );
  CLKBUF_X1 U9382 ( .A(n18306), .Z(n19683) );
  XNOR2_X1 U9444 ( .A(n16694), .B(n16693), .ZN(n19684) );
  NAND2_X1 U9497 ( .A1(n102), .A2(n17820), .ZN(n19685) );
  XNOR2_X1 U9595 ( .A(n16694), .B(n16693), .ZN(n18968) );
  BUF_X1 U9791 ( .A(n7443), .Z(n19686) );
  XNOR2_X1 U9967 ( .A(n5423), .B(n5422), .ZN(n7443) );
  OAI211_X1 U10006 ( .C1(n18960), .C2(n18959), .A(n18958), .B(n18957), .ZN(
        n19687) );
  OAI211_X1 U10071 ( .C1(n18960), .C2(n18959), .A(n18958), .B(n18957), .ZN(
        n19009) );
  XNOR2_X2 U10097 ( .A(n3851), .B(Key[77]), .ZN(n19688) );
  OAI21_X1 U10107 ( .B1(n922), .B2(n12457), .A(n12456), .ZN(n19689) );
  XNOR2_X1 U10196 ( .A(n3851), .B(Key[77]), .ZN(n5258) );
  OAI21_X1 U10261 ( .B1(n922), .B2(n12457), .A(n12456), .ZN(n13584) );
  AND2_X1 U10351 ( .A1(n18540), .A2(n18541), .ZN(n19690) );
  OAI21_X1 U10360 ( .B1(n2691), .B2(n16804), .A(n16803), .ZN(n19691) );
  OAI21_X1 U10453 ( .B1(n2691), .B2(n16804), .A(n16803), .ZN(n18546) );
  INV_X1 U10788 ( .A(n12332), .ZN(n12335) );
  OR2_X1 U10970 ( .A1(n15879), .A2(n15153), .ZN(n14924) );
  OAI21_X1 U10979 ( .B1(n17068), .B2(n17067), .A(n17066), .ZN(n19692) );
  OAI21_X1 U10994 ( .B1(n17068), .B2(n17067), .A(n17066), .ZN(n19155) );
  NAND4_X2 U11000 ( .A1(n1207), .A2(n1573), .A3(n968), .A4(n1209), .ZN(n15714)
         );
  AND2_X1 U11192 ( .A1(n15750), .A2(n25), .ZN(n16044) );
  INV_X1 U11236 ( .A(n14350), .ZN(n19693) );
  XNOR2_X1 U11403 ( .A(n12806), .B(n12805), .ZN(n14327) );
  AND2_X1 U11453 ( .A1(n2647), .A2(n12122), .ZN(n19694) );
  OR2_X1 U11471 ( .A1(n13896), .A2(n13895), .ZN(n28) );
  OR2_X1 U11512 ( .A1(n17495), .A2(n17492), .ZN(n19695) );
  OR2_X1 U11618 ( .A1(n15313), .A2(n14620), .ZN(n1266) );
  AND3_X1 U11724 ( .A1(n3528), .A2(n5685), .A3(n3527), .ZN(n19698) );
  AND3_X1 U11728 ( .A1(n3528), .A2(n5685), .A3(n3527), .ZN(n19699) );
  OAI21_X1 U11806 ( .B1(n5326), .B2(n5327), .A(n5325), .ZN(n7041) );
  XNOR2_X1 U11881 ( .A(n14376), .B(n14375), .ZN(n19700) );
  INV_X1 U11906 ( .A(n20003), .ZN(n19702) );
  OAI21_X1 U11922 ( .B1(n14848), .B2(n16172), .A(n14847), .ZN(n18400) );
  XOR2_X1 U11955 ( .A(n12953), .B(n12954), .Z(n19703) );
  OAI211_X1 U11970 ( .C1(n14838), .C2(n14534), .A(n14533), .B(n14532), .ZN(
        n19704) );
  OAI211_X1 U11982 ( .C1(n14838), .C2(n14534), .A(n14533), .B(n14532), .ZN(
        n19705) );
  NAND2_X1 U12026 ( .A1(n14881), .A2(n1490), .ZN(n19706) );
  NAND2_X1 U12029 ( .A1(n14881), .A2(n1490), .ZN(n17340) );
  OAI21_X1 U12095 ( .B1(n10843), .B2(n1812), .A(n10842), .ZN(n12589) );
  AND2_X1 U12139 ( .A1(n14154), .A2(n14393), .ZN(n19709) );
  XOR2_X1 U12151 ( .A(n10552), .B(n10582), .Z(n9760) );
  AND2_X1 U12159 ( .A1(n7849), .A2(n7850), .ZN(n19710) );
  NAND2_X1 U12163 ( .A1(n17771), .A2(n17770), .ZN(n19711) );
  NAND2_X1 U12210 ( .A1(n17771), .A2(n17770), .ZN(n18794) );
  NOR2_X1 U12272 ( .A1(n17669), .A2(n19249), .ZN(n19276) );
  AOI21_X2 U12275 ( .B1(n15578), .B2(n693), .A(n692), .ZN(n19713) );
  AOI21_X1 U12347 ( .B1(n15578), .B2(n693), .A(n692), .ZN(n17348) );
  NOR2_X1 U12389 ( .A1(n6206), .A2(n19492), .ZN(n5839) );
  XNOR2_X1 U12401 ( .A(n10189), .B(n10190), .ZN(n11430) );
  NAND2_X1 U12596 ( .A1(n102), .A2(n17820), .ZN(n19068) );
  AND2_X1 U12625 ( .A1(n737), .A2(n7509), .ZN(n19715) );
  NAND4_X1 U12668 ( .A1(n9281), .A2(n9279), .A3(n9282), .A4(n9280), .ZN(n19717) );
  NAND4_X1 U12767 ( .A1(n9281), .A2(n9279), .A3(n9282), .A4(n9280), .ZN(n19718) );
  XNOR2_X1 U12875 ( .A(n10585), .B(n10586), .ZN(n19719) );
  NAND4_X1 U12877 ( .A1(n9281), .A2(n9279), .A3(n9282), .A4(n9280), .ZN(n10490) );
  NOR2_X1 U12903 ( .A1(n15469), .A2(n15465), .ZN(n15234) );
  OAI21_X1 U12916 ( .B1(n12171), .B2(n12172), .A(n12170), .ZN(n19721) );
  OR2_X1 U12917 ( .A1(n14291), .A2(n129), .ZN(n19722) );
  OAI21_X1 U12972 ( .B1(n12171), .B2(n12172), .A(n12170), .ZN(n13721) );
  XNOR2_X1 U12975 ( .A(n17039), .B(n17038), .ZN(n19723) );
  AND2_X1 U13093 ( .A1(n18944), .A2(n2062), .ZN(n19724) );
  XNOR2_X1 U13099 ( .A(n17039), .B(n17038), .ZN(n18019) );
  XNOR2_X1 U13253 ( .A(n10111), .B(n10110), .ZN(n19725) );
  OAI211_X1 U13273 ( .C1(n10817), .C2(n19949), .A(n1357), .B(n1356), .ZN(
        n19726) );
  OAI211_X1 U13503 ( .C1(n10817), .C2(n19949), .A(n1357), .B(n1356), .ZN(n948)
         );
  XNOR2_X1 U13535 ( .A(n13478), .B(n13477), .ZN(n19727) );
  XNOR2_X1 U13536 ( .A(n13478), .B(n13477), .ZN(n19728) );
  XNOR2_X1 U13547 ( .A(n13477), .B(n13478), .ZN(n14746) );
  XNOR2_X1 U13580 ( .A(n6966), .B(n7211), .ZN(n6883) );
  NAND2_X1 U13630 ( .A1(n5261), .A2(n2175), .ZN(n19730) );
  NAND2_X1 U13643 ( .A1(n5261), .A2(n2175), .ZN(n6867) );
  BUF_X1 U13692 ( .A(n8828), .Z(n19896) );
  XNOR2_X1 U13697 ( .A(n13627), .B(n13628), .ZN(n19731) );
  XNOR2_X1 U13743 ( .A(n13627), .B(n13628), .ZN(n14393) );
  NOR2_X1 U13779 ( .A1(n19763), .A2(n18394), .ZN(n1296) );
  XNOR2_X1 U14010 ( .A(n20519), .B(n16576), .ZN(n19733) );
  XNOR2_X1 U14108 ( .A(n16577), .B(n16576), .ZN(n19380) );
  BUF_X1 U14109 ( .A(n13029), .Z(n19734) );
  OAI21_X1 U14149 ( .B1(n19919), .B2(n17983), .A(n3206), .ZN(n19735) );
  OAI21_X1 U14157 ( .B1(n19919), .B2(n17983), .A(n3206), .ZN(n18673) );
  XOR2_X1 U14178 ( .A(n9428), .B(n9944), .Z(n19736) );
  XNOR2_X1 U14209 ( .A(n16387), .B(n16693), .ZN(n19737) );
  AND2_X1 U14281 ( .A1(n19462), .A2(n19463), .ZN(n19738) );
  AND3_X1 U14365 ( .A1(n13958), .A2(n13956), .A3(n402), .ZN(n19740) );
  XOR2_X1 U14494 ( .A(n7288), .B(n6410), .Z(n19741) );
  XOR2_X1 U14495 ( .A(n13024), .B(n13023), .Z(n19742) );
  NOR2_X1 U14500 ( .A1(n15360), .A2(n15359), .ZN(n19743) );
  NOR2_X1 U14503 ( .A1(n15360), .A2(n15359), .ZN(n16359) );
  XNOR2_X1 U14512 ( .A(n17106), .B(n17105), .ZN(n19876) );
  XNOR2_X1 U14550 ( .A(n17421), .B(n17422), .ZN(n19744) );
  NOR2_X1 U14581 ( .A1(n18136), .A2(n18135), .ZN(n18650) );
  NAND2_X1 U14599 ( .A1(n8922), .A2(n2301), .ZN(n19746) );
  BUF_X1 U14698 ( .A(n14548), .Z(n19748) );
  NAND2_X1 U14787 ( .A1(n16501), .A2(n16500), .ZN(n19749) );
  XNOR2_X1 U14788 ( .A(n9758), .B(n9757), .ZN(n19750) );
  NOR2_X1 U14789 ( .A1(n17397), .A2(n17398), .ZN(n19751) );
  XNOR2_X1 U14790 ( .A(n9758), .B(n9757), .ZN(n11390) );
  NOR2_X1 U14861 ( .A1(n17398), .A2(n17397), .ZN(n18703) );
  AND2_X1 U14930 ( .A1(n328), .A2(n3704), .ZN(n19752) );
  NAND2_X1 U14983 ( .A1(n17452), .A2(n17453), .ZN(n19753) );
  AND2_X1 U14984 ( .A1(n17875), .A2(n17874), .ZN(n19754) );
  OAI21_X1 U15028 ( .B1(n10853), .B2(n11367), .A(n11365), .ZN(n19755) );
  NAND2_X1 U15048 ( .A1(n1590), .A2(n10873), .ZN(n19756) );
  OAI21_X1 U15085 ( .B1(n10853), .B2(n11367), .A(n11365), .ZN(n1590) );
  NAND2_X1 U15125 ( .A1(n1590), .A2(n10873), .ZN(n12242) );
  OAI21_X1 U15132 ( .B1(n20429), .B2(n17573), .A(n17571), .ZN(n19757) );
  OAI21_X1 U15337 ( .B1(n20429), .B2(n17573), .A(n17571), .ZN(n18621) );
  OAI211_X1 U15377 ( .C1(n12884), .C2(n2039), .A(n12883), .B(n12882), .ZN(
        n12888) );
  NAND2_X1 U15466 ( .A1(n17478), .A2(n17477), .ZN(n19758) );
  NAND2_X1 U15485 ( .A1(n17478), .A2(n17477), .ZN(n18518) );
  BUF_X1 U15486 ( .A(n15349), .Z(n19759) );
  AOI21_X1 U15518 ( .B1(n14501), .B2(n13509), .A(n13508), .ZN(n15349) );
  OAI211_X1 U15520 ( .C1(n9451), .C2(n6442), .A(n6441), .B(n6440), .ZN(n19760)
         );
  XOR2_X1 U15523 ( .A(n13614), .B(n13613), .Z(n19761) );
  XNOR2_X1 U15544 ( .A(n15978), .B(n15977), .ZN(n17873) );
  AND2_X1 U15601 ( .A1(n17247), .A2(n17246), .ZN(n19763) );
  OAI21_X1 U15759 ( .B1(n17307), .B2(n18241), .A(n20093), .ZN(n19766) );
  NOR2_X1 U15781 ( .A1(n7738), .A2(n7737), .ZN(n19767) );
  OR2_X1 U15818 ( .A1(n8402), .A2(n8401), .ZN(n19768) );
  NOR2_X1 U15837 ( .A1(n7738), .A2(n7737), .ZN(n9792) );
  OR2_X1 U15851 ( .A1(n8402), .A2(n8401), .ZN(n12353) );
  OAI211_X1 U15930 ( .C1(n17757), .C2(n17756), .A(n17755), .B(n17754), .ZN(
        n19770) );
  OAI211_X1 U15958 ( .C1(n17757), .C2(n17756), .A(n17755), .B(n17754), .ZN(
        n18806) );
  XOR2_X1 U16103 ( .A(n13595), .B(n13598), .Z(n13606) );
  NAND2_X1 U16249 ( .A1(n15498), .A2(n15500), .ZN(n460) );
  NAND4_X2 U16260 ( .A1(n15478), .A2(n15476), .A3(n15477), .A4(n375), .ZN(
        n17401) );
  XNOR2_X1 U16272 ( .A(n16422), .B(n16519), .ZN(n19774) );
  XNOR2_X1 U16336 ( .A(n16422), .B(n16519), .ZN(n18093) );
  XNOR2_X1 U16373 ( .A(n4030), .B(Key[113]), .ZN(n19776) );
  XNOR2_X1 U16390 ( .A(n4030), .B(Key[113]), .ZN(n19777) );
  XNOR2_X1 U16467 ( .A(n4030), .B(Key[113]), .ZN(n4701) );
  XNOR2_X1 U16521 ( .A(n9406), .B(n9405), .ZN(n19779) );
  XNOR2_X1 U16523 ( .A(n9406), .B(n9405), .ZN(n10694) );
  OAI21_X1 U16583 ( .B1(n5857), .B2(n6159), .A(n2795), .ZN(n19780) );
  OAI21_X1 U16597 ( .B1(n5857), .B2(n6159), .A(n2795), .ZN(n7137) );
  XNOR2_X1 U16642 ( .A(n11625), .B(n11626), .ZN(n19781) );
  OAI21_X1 U16692 ( .B1(n14918), .B2(n14917), .A(n148), .ZN(n19782) );
  OAI21_X1 U16746 ( .B1(n14918), .B2(n14917), .A(n148), .ZN(n19783) );
  XNOR2_X1 U16807 ( .A(n11625), .B(n11626), .ZN(n14810) );
  BUF_X1 U16881 ( .A(n12617), .Z(n19784) );
  XOR2_X1 U16900 ( .A(n16981), .B(n17035), .Z(n17337) );
  XNOR2_X1 U16924 ( .A(n17344), .B(n17343), .ZN(n18257) );
  OAI211_X1 U16945 ( .C1(n8958), .C2(n8505), .A(n8504), .B(n8503), .ZN(n19785)
         );
  OAI211_X1 U17058 ( .C1(n8958), .C2(n8505), .A(n8504), .B(n8503), .ZN(n19786)
         );
  XNOR2_X1 U17083 ( .A(n17344), .B(n17343), .ZN(n19787) );
  XNOR2_X1 U17105 ( .A(Key[135]), .B(Plaintext[135]), .ZN(n5023) );
  OAI21_X1 U17113 ( .B1(n5011), .B2(n5010), .A(n5009), .ZN(n19789) );
  OAI21_X1 U17159 ( .B1(n5011), .B2(n5010), .A(n5009), .ZN(n19790) );
  OAI21_X1 U17181 ( .B1(n5011), .B2(n5010), .A(n5009), .ZN(n6031) );
  AND2_X1 U17200 ( .A1(n16467), .A2(n60), .ZN(n19791) );
  NOR2_X1 U17290 ( .A1(n11596), .A2(n11597), .ZN(n19792) );
  NOR2_X1 U17304 ( .A1(n11596), .A2(n11597), .ZN(n12861) );
  BUF_X1 U17409 ( .A(n18842), .Z(n19794) );
  OAI21_X1 U17410 ( .B1(n17320), .B2(n18033), .A(n3691), .ZN(n18842) );
  AOI21_X1 U17480 ( .B1(n12329), .B2(n12328), .A(n13269), .ZN(n19797) );
  NAND4_X1 U17488 ( .A1(n15689), .A2(n15691), .A3(n15690), .A4(n93), .ZN(
        n19798) );
  NAND4_X1 U17500 ( .A1(n15689), .A2(n15691), .A3(n15690), .A4(n93), .ZN(
        n19799) );
  NAND4_X1 U17576 ( .A1(n15689), .A2(n15691), .A3(n15690), .A4(n93), .ZN(
        n17379) );
  INV_X1 U17643 ( .A(n8196), .ZN(n19802) );
  NAND3_X1 U17667 ( .A1(n18247), .A2(n18246), .A3(n18245), .ZN(n19803) );
  BUF_X1 U17713 ( .A(n5524), .Z(n19804) );
  INV_X1 U17729 ( .A(n8830), .ZN(n19805) );
  BUF_X1 U17809 ( .A(n10199), .Z(n19806) );
  AOI22_X1 U17912 ( .A1(n8679), .A2(n8830), .B1(n8678), .B2(n9060), .ZN(n10199) );
  OAI211_X1 U17960 ( .C1(n15332), .C2(n15866), .A(n15331), .B(n15330), .ZN(
        n19807) );
  OAI211_X1 U17981 ( .C1(n15332), .C2(n15866), .A(n15331), .B(n15330), .ZN(
        n17252) );
  NOR2_X1 U18024 ( .A1(n6049), .A2(n6048), .ZN(n5330) );
  XNOR2_X1 U18071 ( .A(n6448), .B(n6447), .ZN(n8221) );
  OAI21_X1 U18072 ( .B1(n2326), .B2(n2325), .A(n2324), .ZN(n7405) );
  BUF_X1 U18180 ( .A(n8098), .Z(n8238) );
  XNOR2_X2 U18211 ( .A(n1693), .B(n6841), .ZN(n8157) );
  NAND3_X2 U18249 ( .A1(n601), .A2(n17594), .A3(n17593), .ZN(n19284) );
  XOR2_X1 U18273 ( .A(n13776), .B(n13369), .Z(n2521) );
  AND2_X1 U18287 ( .A1(n17763), .A2(n17762), .ZN(n19811) );
  XOR2_X1 U18292 ( .A(n6289), .B(n6288), .Z(n19812) );
  OAI211_X1 U18313 ( .C1(n20206), .C2(n13867), .A(n1790), .B(n1789), .ZN(
        n15502) );
  CLKBUF_X1 U18318 ( .A(n17497), .Z(n19814) );
  INV_X1 U18348 ( .A(n18497), .ZN(n19816) );
  XNOR2_X1 U18352 ( .A(n15526), .B(n15525), .ZN(n17497) );
  XOR2_X1 U18355 ( .A(n9409), .B(n9410), .Z(n19817) );
  OAI21_X1 U18366 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n19818) );
  XNOR2_X1 U18375 ( .A(n12719), .B(n12718), .ZN(n19819) );
  XNOR2_X1 U18437 ( .A(n2488), .B(Key[17]), .ZN(n19822) );
  XNOR2_X1 U18469 ( .A(n2488), .B(Key[17]), .ZN(n4302) );
  XNOR2_X1 U18470 ( .A(n15137), .B(n15136), .ZN(n19823) );
  XNOR2_X1 U18484 ( .A(n15137), .B(n15136), .ZN(n1718) );
  XOR2_X1 U18511 ( .A(n13534), .B(n19887), .Z(n19824) );
  OR2_X1 U18519 ( .A1(n20231), .A2(n20139), .ZN(n19825) );
  XNOR2_X1 U18594 ( .A(n6524), .B(n6523), .ZN(n19826) );
  AOI21_X1 U18718 ( .B1(n7792), .B2(n7791), .A(n7790), .ZN(n8985) );
  AOI21_X1 U18741 ( .B1(n14538), .B2(n2676), .A(n14537), .ZN(n19828) );
  XOR2_X1 U18757 ( .A(n12990), .B(n12989), .Z(n19831) );
  XNOR2_X1 U18781 ( .A(n10184), .B(n10183), .ZN(n11431) );
  XOR2_X1 U18849 ( .A(n16065), .B(n16064), .Z(n19832) );
  NAND3_X1 U18852 ( .A1(n11185), .A2(n2948), .A3(n2949), .ZN(n19833) );
  NAND3_X1 U19067 ( .A1(n2006), .A2(n3137), .A3(n3136), .ZN(n17349) );
  BUF_X1 U19083 ( .A(n11132), .Z(n19837) );
  OR2_X1 U19084 ( .A1(n14278), .A2(n1409), .ZN(n19838) );
  AOI22_X1 U19122 ( .A1(n8643), .A2(n8929), .B1(n8598), .B2(n8933), .ZN(n10179) );
  OAI211_X1 U19144 ( .C1(n3603), .C2(n3604), .A(n5814), .B(n3602), .ZN(n19840)
         );
  OAI211_X1 U19145 ( .C1(n3603), .C2(n3604), .A(n5814), .B(n3602), .ZN(n19841)
         );
  OAI21_X1 U19147 ( .B1(n16317), .B2(n1112), .A(n16316), .ZN(n19842) );
  OAI211_X1 U19148 ( .C1(n3603), .C2(n3604), .A(n5814), .B(n3602), .ZN(n7231)
         );
  OAI21_X1 U19149 ( .B1(n16317), .B2(n1112), .A(n16316), .ZN(n19196) );
  XNOR2_X1 U19150 ( .A(n10585), .B(n10586), .ZN(n11491) );
  NOR2_X1 U19155 ( .A1(n14139), .A2(n14138), .ZN(n19844) );
  NOR2_X1 U19273 ( .A1(n14139), .A2(n14138), .ZN(n19845) );
  XNOR2_X1 U19287 ( .A(n3419), .B(n13654), .ZN(n14722) );
  NOR2_X1 U19290 ( .A1(n14139), .A2(n14138), .ZN(n15936) );
  XOR2_X1 U19360 ( .A(n13446), .B(n13644), .Z(n12159) );
  XOR2_X1 U19362 ( .A(n16951), .B(n16950), .Z(n19846) );
  XOR2_X1 U19464 ( .A(n7122), .B(n7081), .Z(n19847) );
  XNOR2_X1 U19465 ( .A(n14963), .B(n16969), .ZN(n19849) );
  OAI21_X1 U19466 ( .B1(n14505), .B2(n14506), .A(n14504), .ZN(n15284) );
  CLKBUF_X1 U19573 ( .A(n6754), .Z(n19850) );
  XNOR2_X1 U19574 ( .A(n9425), .B(n9424), .ZN(n19851) );
  XNOR2_X1 U19575 ( .A(n9425), .B(n9424), .ZN(n11000) );
  XOR2_X1 U19576 ( .A(n7317), .B(n7091), .Z(n19852) );
  OAI211_X1 U19577 ( .C1(n3494), .C2(n19941), .A(n3495), .B(n3492), .ZN(n19853) );
  OAI211_X1 U19578 ( .C1(n3494), .C2(n19941), .A(n3495), .B(n3492), .ZN(n9669)
         );
  NAND3_X2 U19582 ( .A1(n2847), .A2(n2850), .A3(n838), .ZN(n10126) );
  XNOR2_X1 U19583 ( .A(n7293), .B(n7292), .ZN(n19856) );
  NOR2_X1 U19586 ( .A1(n8512), .A2(n8513), .ZN(n8510) );
  XOR2_X1 U19587 ( .A(n12732), .B(n12733), .Z(n19859) );
  BUF_X1 U19588 ( .A(n12636), .Z(n19861) );
  OAI211_X2 U19590 ( .C1(n9128), .C2(n9127), .A(n9126), .B(n9125), .ZN(n10079)
         );
  XNOR2_X1 U19591 ( .A(n17359), .B(n16429), .ZN(n19863) );
  XNOR2_X1 U19592 ( .A(n10006), .B(n10005), .ZN(n19864) );
  XNOR2_X1 U19593 ( .A(n10006), .B(n10005), .ZN(n11514) );
  XNOR2_X1 U19594 ( .A(n5270), .B(n5269), .ZN(n19865) );
  XNOR2_X1 U19595 ( .A(n5270), .B(n5269), .ZN(n3748) );
  OAI21_X1 U19596 ( .B1(n18952), .B2(n2590), .A(n18951), .ZN(n19866) );
  OAI21_X1 U19597 ( .B1(n18952), .B2(n2590), .A(n18951), .ZN(n19867) );
  OAI21_X1 U19598 ( .B1(n18952), .B2(n2590), .A(n18951), .ZN(n19021) );
  XOR2_X1 U19599 ( .A(Key[101]), .B(Plaintext[101]), .Z(n19868) );
  OAI211_X1 U19600 ( .C1(n12235), .C2(n12236), .A(n12234), .B(n12233), .ZN(
        n19869) );
  OAI211_X1 U19602 ( .C1(n12235), .C2(n12236), .A(n12234), .B(n12233), .ZN(
        n13511) );
  CLKBUF_X1 U19603 ( .A(n10299), .Z(n19871) );
  XOR2_X1 U19604 ( .A(n1524), .B(n1523), .Z(n19872) );
  OAI21_X1 U19606 ( .B1(n18962), .B2(n17057), .A(n17056), .ZN(n19874) );
  OAI21_X1 U19607 ( .B1(n18962), .B2(n17057), .A(n17056), .ZN(n18899) );
  XNOR2_X1 U19608 ( .A(n11936), .B(n11935), .ZN(n14619) );
  OR2_X1 U19609 ( .A1(n17551), .A2(n17550), .ZN(n19877) );
  XNOR2_X1 U19610 ( .A(n17106), .B(n17105), .ZN(n17545) );
  XOR2_X1 U19611 ( .A(n9350), .B(n9349), .Z(n19878) );
  NOR2_X1 U19612 ( .A1(n13318), .A2(n478), .ZN(n19879) );
  OAI21_X1 U19613 ( .B1(n7846), .B2(n20251), .A(n1236), .ZN(n19880) );
  OAI21_X1 U19614 ( .B1(n7846), .B2(n20251), .A(n1236), .ZN(n9271) );
  XNOR2_X1 U19615 ( .A(n638), .B(n6732), .ZN(n19881) );
  OAI211_X1 U19617 ( .C1(n13264), .C2(n14738), .A(n13263), .B(n1849), .ZN(
        n19884) );
  AOI21_X1 U19618 ( .B1(n12276), .B2(n12300), .A(n1872), .ZN(n12945) );
  OAI211_X1 U19619 ( .C1(n13264), .C2(n14738), .A(n13263), .B(n1849), .ZN(
        n15667) );
  XNOR2_X1 U19620 ( .A(n16340), .B(n16339), .ZN(n19885) );
  XNOR2_X1 U19621 ( .A(n16340), .B(n16339), .ZN(n18114) );
  XNOR2_X1 U19622 ( .A(n16758), .B(n15827), .ZN(n16673) );
  XOR2_X1 U19623 ( .A(n10285), .B(n10284), .Z(n19886) );
  OAI211_X1 U19624 ( .C1(n12333), .C2(n11974), .A(n11973), .B(n11972), .ZN(
        n19887) );
  CLKBUF_X1 U19627 ( .A(n18844), .Z(n19890) );
  OAI21_X1 U19628 ( .B1(n14567), .B2(n14566), .A(n14565), .ZN(n19891) );
  OAI21_X1 U19630 ( .B1(n15765), .B2(n15248), .A(n15247), .ZN(n19894) );
  OAI211_X1 U19631 ( .C1(n11807), .C2(n12537), .A(n11806), .B(n11805), .ZN(
        n13519) );
  XNOR2_X1 U19633 ( .A(n10042), .B(n10041), .ZN(n19897) );
  OAI211_X1 U19634 ( .C1(n7696), .C2(n7504), .A(n7503), .B(n7502), .ZN(n8828)
         );
  XNOR2_X1 U19635 ( .A(n10042), .B(n10041), .ZN(n11211) );
  XNOR2_X1 U19636 ( .A(n15483), .B(n15482), .ZN(n19898) );
  XOR2_X1 U19637 ( .A(n13762), .B(n13616), .Z(n19899) );
  OAI211_X1 U19639 ( .C1(n15208), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        n19900) );
  OAI211_X1 U19640 ( .C1(n15208), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        n16747) );
  INV_X1 U19641 ( .A(n18497), .ZN(n18489) );
  INV_X1 U19642 ( .A(n10726), .ZN(n11093) );
  XNOR2_X1 U19643 ( .A(n6623), .B(n6622), .ZN(n19901) );
  XNOR2_X1 U19644 ( .A(n6623), .B(n6622), .ZN(n8175) );
  OAI21_X1 U19645 ( .B1(n17713), .B2(n20221), .A(n17712), .ZN(n19043) );
  XNOR2_X1 U19646 ( .A(n13992), .B(n16566), .ZN(n19903) );
  OAI211_X1 U19647 ( .C1(n12381), .C2(n12380), .A(n12379), .B(n12378), .ZN(
        n19904) );
  CLKBUF_X1 U19648 ( .A(n17054), .Z(n19905) );
  XNOR2_X1 U19649 ( .A(n2520), .B(n2519), .ZN(n19906) );
  XNOR2_X1 U19650 ( .A(n13766), .B(n13765), .ZN(n19907) );
  XNOR2_X1 U19651 ( .A(n13766), .B(n13765), .ZN(n19908) );
  OAI211_X1 U19652 ( .C1(n15514), .C2(n15513), .A(n15512), .B(n519), .ZN(
        n19909) );
  OAI211_X1 U19653 ( .C1(n15514), .C2(n15513), .A(n15512), .B(n519), .ZN(
        n16082) );
  XNOR2_X1 U19654 ( .A(n16033), .B(n17371), .ZN(n19910) );
  MUX2_X2 U19656 ( .A(n17011), .B(n17010), .S(n18932), .Z(n18921) );
  INV_X1 U19657 ( .A(n12609), .ZN(n19971) );
  OAI211_X1 U19658 ( .C1(n3896), .C2(n4947), .A(n3895), .B(n3894), .ZN(n19912)
         );
  XOR2_X1 U19659 ( .A(n10593), .B(n10592), .Z(n19913) );
  XOR2_X1 U19660 ( .A(n6878), .B(n6877), .Z(n19914) );
  XOR2_X1 U19661 ( .A(n8821), .B(n8822), .Z(n19915) );
  XNOR2_X1 U19662 ( .A(n16925), .B(n16924), .ZN(n19916) );
  OR2_X1 U19663 ( .A1(n18050), .A2(n18049), .ZN(n19917) );
  XNOR2_X1 U19664 ( .A(n13821), .B(n13822), .ZN(n19918) );
  XOR2_X1 U19665 ( .A(n17266), .B(n17265), .Z(n19919) );
  XNOR2_X1 U19666 ( .A(n13821), .B(n13822), .ZN(n14250) );
  XNOR2_X1 U19667 ( .A(n10429), .B(n10428), .ZN(n19920) );
  BUF_X1 U19668 ( .A(n14692), .Z(n19921) );
  XNOR2_X1 U19669 ( .A(n10429), .B(n10428), .ZN(n11443) );
  XNOR2_X1 U19670 ( .A(n5727), .B(n5726), .ZN(n19922) );
  NOR2_X1 U19671 ( .A1(n12190), .A2(n2426), .ZN(n19923) );
  NOR2_X1 U19672 ( .A1(n12190), .A2(n2426), .ZN(n13383) );
  XOR2_X1 U19673 ( .A(n15483), .B(n15482), .Z(n19924) );
  XNOR2_X1 U19674 ( .A(n2211), .B(n6772), .ZN(n19925) );
  NOR2_X1 U19676 ( .A1(n14862), .A2(n1489), .ZN(n19927) );
  NOR2_X1 U19677 ( .A1(n14862), .A2(n1489), .ZN(n19928) );
  NOR2_X1 U19678 ( .A1(n14862), .A2(n1489), .ZN(n17425) );
  XNOR2_X1 U19680 ( .A(n16049), .B(n16048), .ZN(n19930) );
  XNOR2_X1 U19681 ( .A(n16049), .B(n16048), .ZN(n17666) );
  OAI21_X1 U19682 ( .B1(n14578), .B2(n20187), .A(n14577), .ZN(n19931) );
  OAI21_X1 U19683 ( .B1(n14578), .B2(n20187), .A(n14577), .ZN(n15828) );
  XOR2_X1 U19685 ( .A(n16935), .B(n16934), .Z(n19933) );
  INV_X1 U19686 ( .A(n18652), .ZN(n19935) );
  OAI21_X1 U19687 ( .B1(n18142), .B2(n18141), .A(n18140), .ZN(n18652) );
  XOR2_X1 U19688 ( .A(n16532), .B(n16531), .Z(n19936) );
  OAI211_X1 U19689 ( .C1(n12428), .C2(n3649), .A(n12098), .B(n12097), .ZN(
        n19937) );
  XNOR2_X1 U19690 ( .A(n1436), .B(n16509), .ZN(n19938) );
  XOR2_X1 U19691 ( .A(n13046), .B(n13045), .Z(n19940) );
  OAI211_X1 U19692 ( .C1(n7682), .C2(n8166), .A(n7681), .B(n7680), .ZN(n9354)
         );
  XOR2_X1 U19694 ( .A(n16352), .B(n16351), .Z(n19943) );
  OAI211_X1 U19695 ( .C1(n5225), .C2(n5768), .A(n5224), .B(n5223), .ZN(n19944)
         );
  OAI211_X1 U19696 ( .C1(n5225), .C2(n5768), .A(n5224), .B(n5223), .ZN(n7187)
         );
  AOI21_X1 U19697 ( .B1(n9133), .B2(n9132), .A(n9131), .ZN(n10077) );
  AOI21_X1 U19698 ( .B1(n12297), .B2(n12296), .A(n2220), .ZN(n19946) );
  XNOR2_X1 U19699 ( .A(n16087), .B(n16086), .ZN(n19947) );
  XNOR2_X1 U19700 ( .A(n16087), .B(n16086), .ZN(n17887) );
  MUX2_X1 U19701 ( .A(n17083), .B(n17082), .S(n20239), .Z(n19948) );
  MUX2_X1 U19702 ( .A(n17083), .B(n17082), .S(n20239), .Z(n19164) );
  XNOR2_X2 U19708 ( .A(n13326), .B(n13327), .ZN(n14385) );
  AOI22_X1 U19709 ( .A1(n6160), .A2(n5614), .B1(n5613), .B2(n5612), .ZN(n19953) );
  NAND2_X1 U19711 ( .A1(n565), .A2(n1154), .ZN(n19954) );
  OAI21_X1 U19712 ( .B1(n20240), .B2(n16543), .A(n16542), .ZN(n19955) );
  XNOR2_X1 U19714 ( .A(n3575), .B(n3574), .ZN(n19956) );
  XNOR2_X1 U19715 ( .A(n3575), .B(n3574), .ZN(n17223) );
  XOR2_X1 U19716 ( .A(n9096), .B(n9097), .Z(n19957) );
  OR2_X1 U19717 ( .A1(n11349), .A2(n11347), .ZN(n11060) );
  XOR2_X1 U19719 ( .A(n10408), .B(n10407), .Z(n19959) );
  NAND2_X1 U19720 ( .A1(n9308), .A2(n9313), .ZN(n1128) );
  AND2_X2 U19721 ( .A1(n19960), .A2(n19529), .ZN(n9313) );
  NAND2_X1 U19722 ( .A1(n1584), .A2(n8113), .ZN(n19960) );
  NAND2_X1 U19723 ( .A1(n19962), .A2(n18042), .ZN(n17814) );
  NOR2_X1 U19724 ( .A1(n18948), .A2(n17812), .ZN(n19962) );
  NAND2_X1 U19725 ( .A1(n19963), .A2(n4330), .ZN(n3110) );
  NAND2_X1 U19726 ( .A1(n4177), .A2(n4613), .ZN(n4330) );
  OAI21_X2 U19727 ( .B1(n15548), .B2(n2803), .A(n1100), .ZN(n16872) );
  NOR3_X1 U19728 ( .A1(n11953), .A2(n11829), .A3(n11952), .ZN(n2562) );
  NAND4_X1 U19729 ( .A1(n11822), .A2(n19964), .A3(n11821), .A4(n13270), .ZN(
        n11823) );
  NAND2_X1 U19730 ( .A1(n12325), .A2(n11997), .ZN(n19964) );
  NAND2_X1 U19732 ( .A1(n15802), .A2(n15801), .ZN(n19966) );
  NAND2_X1 U19733 ( .A1(n5840), .A2(n19967), .ZN(n7143) );
  NAND2_X1 U19734 ( .A1(n19522), .A2(n19968), .ZN(n19967) );
  NAND2_X1 U19735 ( .A1(n1293), .A2(n15402), .ZN(n15069) );
  XNOR2_X1 U19736 ( .A(n19969), .B(n18389), .ZN(Ciphertext[9]) );
  OAI21_X1 U19737 ( .B1(n12610), .B2(n19971), .A(n19970), .ZN(n12239) );
  NAND2_X1 U19738 ( .A1(n12610), .A2(n12237), .ZN(n19970) );
  NAND2_X1 U19740 ( .A1(n7980), .A2(n7767), .ZN(n7769) );
  NAND2_X1 U19741 ( .A1(n19517), .A2(n7752), .ZN(n3554) );
  NAND2_X1 U19742 ( .A1(n15108), .A2(n14947), .ZN(n16329) );
  NAND2_X1 U19743 ( .A1(n14944), .A2(n15292), .ZN(n14946) );
  OR2_X1 U19746 ( .A1(n11289), .A2(n9559), .ZN(n19972) );
  XNOR2_X1 U19747 ( .A(n13261), .B(n13262), .ZN(n14736) );
  OAI211_X1 U19748 ( .C1(n12333), .C2(n11974), .A(n11973), .B(n11972), .ZN(
        n12997) );
  AND3_X2 U1521 ( .A1(n11994), .A2(n11993), .A3(n12333), .ZN(n13481) );
  BUF_X1 U1416 ( .A(n16011), .Z(n901) );
  NAND2_X2 U915 ( .A1(n14118), .A2(n14117), .ZN(n16126) );
  XNOR2_X2 U2647 ( .A(n6561), .B(n6560), .ZN(n8100) );
  MUX2_X2 U891 ( .A(n14075), .B(n14074), .S(n3223), .Z(n15748) );
  AND2_X2 U2961 ( .A1(n13182), .A2(n13181), .ZN(n785) );
  BUF_X2 U14440 ( .A(n12061), .Z(n12595) );
  INV_X1 U17527 ( .A(n17650), .ZN(n19401) );
  NAND2_X2 U1744 ( .A1(n3750), .A2(n970), .ZN(n9105) );
  BUF_X2 U8534 ( .A(n7457), .Z(n8196) );
  BUF_X1 U1619 ( .A(n11147), .Z(n11016) );
  BUF_X1 U1315 ( .A(n15310), .Z(n19662) );
  OAI21_X2 U6746 ( .B1(n7869), .B2(n7870), .A(n7868), .ZN(n10264) );
  XNOR2_X1 U555 ( .A(n9690), .B(n9689), .ZN(n11377) );
  OAI22_X2 U1092 ( .A1(n9933), .A2(n10635), .B1(n10923), .B2(n2469), .ZN(
        n12352) );
  OAI211_X2 U6737 ( .C1(n5373), .C2(n5398), .A(n5372), .B(n5371), .ZN(n7316)
         );
  XNOR2_X1 U2601 ( .A(n5940), .B(n5939), .ZN(n8300) );
  NAND2_X2 U1915 ( .A1(n3350), .A2(n3349), .ZN(n6050) );
  INV_X1 U15140 ( .A(n19336), .ZN(n19337) );
  NAND3_X2 U848 ( .A1(n2898), .A2(n2899), .A3(n2897), .ZN(n3305) );
  BUF_X1 U8972 ( .A(n16982), .Z(n19674) );
  BUF_X1 U224 ( .A(n8195), .Z(n19474) );
  OR3_X1 U4696 ( .A1(n8652), .A2(n9262), .A3(n7866), .ZN(n8655) );
  NOR2_X2 U6176 ( .A1(n3213), .A2(n3215), .ZN(n19190) );
  NOR2_X2 U19584 ( .A1(n8512), .A2(n8513), .ZN(n19857) );
  XNOR2_X1 U8825 ( .A(Key[144]), .B(Plaintext[144]), .ZN(n4750) );
  CLKBUF_X1 U1247 ( .A(Key[175]), .Z(n2100) );
  XNOR2_X1 U8855 ( .A(Key[165]), .B(Plaintext[165]), .ZN(n3948) );
  XNOR2_X1 U9023 ( .A(n4045), .B(Key[106]), .ZN(n5101) );
  AND2_X1 U6816 ( .A1(n4351), .A2(n4352), .ZN(n5717) );
  AND3_X1 U1935 ( .A1(n5505), .A2(n5504), .A3(n5510), .ZN(n6007) );
  OAI211_X1 U73 ( .C1(n4608), .C2(n4607), .A(n4606), .B(n4605), .ZN(n5745) );
  AND2_X1 U5550 ( .A1(n4579), .A2(n4580), .ZN(n5382) );
  NAND2_X1 U554 ( .A1(n4267), .A2(n4266), .ZN(n6129) );
  AND3_X1 U6032 ( .A1(n3008), .A2(n3009), .A3(n4735), .ZN(n6113) );
  AND2_X1 U1901 ( .A1(n4918), .A2(n4917), .ZN(n5476) );
  AND2_X1 U56 ( .A1(n3640), .A2(n5226), .ZN(n6220) );
  OR2_X1 U9641 ( .A1(n4995), .A2(n5138), .ZN(n4997) );
  NAND2_X1 U897 ( .A1(n5123), .A2(n1978), .ZN(n7046) );
  NAND2_X1 U924 ( .A1(n1708), .A2(n1705), .ZN(n7392) );
  OAI211_X1 U439 ( .C1(n5275), .C2(n19562), .A(n5274), .B(n5273), .ZN(n6850)
         );
  NAND2_X1 U4748 ( .A1(n1886), .A2(n1885), .ZN(n7267) );
  OAI211_X1 U10333 ( .C1(n6160), .C2(n6159), .A(n6158), .B(n6157), .ZN(n7348)
         );
  BUF_X1 U470 ( .A(n5984), .Z(n7272) );
  BUF_X1 U941 ( .A(n7009), .Z(n179) );
  XNOR2_X1 U10260 ( .A(n5962), .B(n5961), .ZN(n8299) );
  XNOR2_X1 U11101 ( .A(n7029), .B(n7030), .ZN(n7836) );
  BUF_X1 U692 ( .A(n6510), .Z(n7560) );
  NAND2_X1 U547 ( .A1(n7498), .A2(n3377), .ZN(n9291) );
  INV_X1 U4861 ( .A(n8722), .ZN(n9358) );
  OR2_X1 U1737 ( .A1(n8223), .A2(n8224), .ZN(n8797) );
  AND2_X1 U7666 ( .A1(n3075), .A2(n3073), .ZN(n9031) );
  NAND2_X1 U7995 ( .A1(n3384), .A2(n3383), .ZN(n8527) );
  INV_X1 U1470 ( .A(n8419), .ZN(n9209) );
  AND2_X1 U5581 ( .A1(n7804), .A2(n7803), .ZN(n8987) );
  OAI211_X1 U914 ( .C1(n8611), .C2(n7540), .A(n7539), .B(n7538), .ZN(n9947) );
  OAI21_X1 U6707 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n9817) );
  NAND2_X1 U3538 ( .A1(n8519), .A2(n8518), .ZN(n10461) );
  NAND2_X1 U4864 ( .A1(n1202), .A2(n1200), .ZN(n10436) );
  AND3_X1 U1671 ( .A1(n8626), .A2(n8625), .A3(n8624), .ZN(n10002) );
  AND2_X1 U3871 ( .A1(n9323), .A2(n9838), .ZN(n9960) );
  XNOR2_X1 U859 ( .A(n9823), .B(n9822), .ZN(n11263) );
  XNOR2_X1 U1633 ( .A(n1823), .B(n9316), .ZN(n11177) );
  XNOR2_X1 U3241 ( .A(n2496), .B(n2495), .ZN(n11192) );
  XNOR2_X1 U7367 ( .A(n8590), .B(n8591), .ZN(n10926) );
  XNOR2_X1 U1642 ( .A(n10147), .B(n10146), .ZN(n11057) );
  XNOR2_X1 U592 ( .A(n9929), .B(n9928), .ZN(n11076) );
  INV_X1 U179 ( .A(n10513), .ZN(n11440) );
  BUF_X1 U731 ( .A(n10112), .Z(n10813) );
  NAND3_X1 U13717 ( .A1(n202), .A2(n2861), .A3(n11376), .ZN(n10858) );
  INV_X1 U13393 ( .A(n10724), .ZN(n11051) );
  OR2_X1 U3259 ( .A1(n9546), .A2(n9547), .ZN(n3176) );
  OR2_X1 U1572 ( .A1(n9490), .A2(n9489), .ZN(n9491) );
  INV_X1 U1557 ( .A(n9491), .ZN(n12179) );
  MUX2_X1 U13621 ( .A(n10744), .B(n10743), .S(n10936), .Z(n12754) );
  OAI21_X1 U827 ( .B1(n10648), .B2(n11556), .A(n10647), .ZN(n12421) );
  OAI211_X1 U3938 ( .C1(n11050), .C2(n11459), .A(n2130), .B(n10260), .ZN(
        n12339) );
  OR2_X1 U2295 ( .A1(n12590), .A2(n12200), .ZN(n1252) );
  NOR2_X1 U3413 ( .A1(n10659), .A2(n10658), .ZN(n13088) );
  MUX2_X1 U14164 ( .A(n11663), .B(n11662), .S(n11661), .Z(n13651) );
  AOI22_X1 U614 ( .A1(n13144), .A2(n13146), .B1(n11099), .B2(n11098), .ZN(
        n13280) );
  AND3_X1 U129 ( .A1(n1981), .A2(n10850), .A3(n1980), .ZN(n12709) );
  NAND3_X1 U4719 ( .A1(n12112), .A2(n12113), .A3(n12111), .ZN(n13398) );
  AND2_X1 U763 ( .A1(n12447), .A2(n12446), .ZN(n13697) );
  NAND2_X1 U266 ( .A1(n11919), .A2(n40), .ZN(n13453) );
  INV_X1 U3615 ( .A(n14249), .ZN(n1262) );
  XNOR2_X1 U1468 ( .A(n13663), .B(n13662), .ZN(n14717) );
  XNOR2_X1 U14960 ( .A(n12858), .B(n12857), .ZN(n14451) );
  BUF_X1 U124 ( .A(n14420), .Z(n19939) );
  XNOR2_X1 U909 ( .A(n11103), .B(n11102), .ZN(n14780) );
  XNOR2_X1 U946 ( .A(n12943), .B(n12942), .ZN(n14644) );
  MUX2_X1 U6806 ( .A(n13630), .B(n13629), .S(n19731), .Z(n15682) );
  MUX2_X2 U15881 ( .A(n14110), .B(n14109), .S(n14723), .Z(n15495) );
  NAND2_X1 U995 ( .A1(n13949), .A2(n2952), .ZN(n16016) );
  NAND2_X1 U15063 ( .A1(n12975), .A2(n12976), .ZN(n15777) );
  NOR2_X1 U164 ( .A1(n14756), .A2(n14755), .ZN(n15503) );
  BUF_X1 U959 ( .A(n15515), .Z(n19502) );
  AND2_X1 U397 ( .A1(n14616), .A2(n14615), .ZN(n15276) );
  OR2_X1 U1063 ( .A1(n15567), .A2(n15566), .ZN(n14954) );
  AND2_X1 U5473 ( .A1(n2564), .A2(n2565), .ZN(n15870) );
  XNOR2_X1 U544 ( .A(n15889), .B(n15888), .ZN(n19352) );
  CLKBUF_X1 U1336 ( .A(n18026), .Z(n17749) );
  INV_X1 U17439 ( .A(n17955), .ZN(n18107) );
  MUX2_X1 U18695 ( .A(n18045), .B(n18044), .S(n18946), .Z(n18050) );
  OAI211_X1 U843 ( .C1(n2819), .C2(n17664), .A(n2818), .B(n2817), .ZN(n2816)
         );
  AOI22_X1 U5765 ( .A1(n17614), .A2(n17613), .B1(n17612), .B2(n17611), .ZN(
        n19299) );
  OAI21_X1 U8402 ( .B1(n16913), .B2(n16912), .A(n16911), .ZN(n18897) );
  AND3_X1 U196 ( .A1(n18247), .A2(n18246), .A3(n18245), .ZN(n18773) );
  NAND2_X1 U2062 ( .A1(n17747), .A2(n319), .ZN(n18807) );
  OAI211_X1 U2093 ( .C1(n20648), .C2(n16797), .A(n2633), .B(n16168), .ZN(
        n18497) );
  OR2_X1 U1039 ( .A1(n15965), .A2(n15964), .ZN(n18057) );
  OR2_X1 U650 ( .A1(n20124), .A2(n19233), .ZN(n19229) );
  INV_X1 U9292 ( .A(n5717), .ZN(n5714) );
  INV_X1 U1015 ( .A(n5349), .ZN(n6156) );
  CLKBUF_X1 U3720 ( .A(n3855), .Z(n5785) );
  NAND2_X2 U161 ( .A1(n3658), .A2(n1807), .ZN(n5605) );
  MUX2_X1 U5895 ( .A(n5890), .B(n5889), .S(n5888), .Z(n6761) );
  OAI211_X1 U431 ( .C1(n5654), .C2(n5653), .A(n5652), .B(n5651), .ZN(n6912) );
  INV_X1 U3791 ( .A(n7470), .ZN(n8293) );
  AND2_X1 U1686 ( .A1(n1103), .A2(n1102), .ZN(n9414) );
  XNOR2_X1 U6090 ( .A(n9156), .B(n9155), .ZN(n11556) );
  INV_X1 U3911 ( .A(n9351), .ZN(n11178) );
  NAND2_X1 U1495 ( .A1(n3277), .A2(n3276), .ZN(n13572) );
  NAND3_X1 U2594 ( .A1(n11861), .A2(n542), .A3(n541), .ZN(n13064) );
  OR2_X1 U2700 ( .A1(n14022), .A2(n14021), .ZN(n14288) );
  BUF_X1 U1071 ( .A(n13946), .Z(n14688) );
  OAI211_X1 U6010 ( .C1(n12695), .C2(n14419), .A(n3635), .B(n3636), .ZN(n15341) );
  AOI22_X1 U550 ( .A1(n15605), .A2(n15604), .B1(n15603), .B2(n15602), .ZN(
        n16970) );
  MUX2_X1 U38 ( .A(n16315), .B(n16314), .S(n20512), .Z(n16316) );
  CLKBUF_X1 U11616 ( .A(n18009), .Z(n18522) );
  MUX2_X2 U1136 ( .A(n4661), .B(n4660), .S(n4841), .Z(n6168) );
  NAND3_X2 U289 ( .A1(n7435), .A2(n7434), .A3(n7433), .ZN(n9295) );
  NOR2_X2 U4569 ( .A1(n14331), .A2(n14330), .ZN(n15470) );
  AND2_X2 U5326 ( .A1(n3594), .A2(n3595), .ZN(n9204) );
  NOR2_X2 U5119 ( .A1(n11669), .A2(n11668), .ZN(n12940) );
  BUF_X2 U1750 ( .A(n8103), .Z(n9328) );
  XNOR2_X2 U12894 ( .A(n10503), .B(n9770), .ZN(n11866) );
  AND3_X2 U777 ( .A1(n822), .A2(n3585), .A3(n3584), .ZN(n953) );
  NOR2_X2 U141 ( .A1(n6188), .A2(n6187), .ZN(n19778) );
  AOI22_X2 U2761 ( .A1(n15039), .A2(n15698), .B1(n15702), .B2(n15040), .ZN(
        n17143) );
  NAND3_X2 U255 ( .A1(n6179), .A2(n6177), .A3(n6178), .ZN(n7032) );
  MUX2_X2 U6882 ( .A(n6086), .B(n6085), .S(n3529), .Z(n7354) );
  MUX2_X2 U10348 ( .A(n8554), .B(n8553), .S(n8814), .Z(n10421) );
  NAND2_X2 U2639 ( .A1(n3135), .A2(n3296), .ZN(n12686) );
  OR2_X2 U753 ( .A1(n8246), .A2(n8253), .ZN(n900) );
  AND2_X2 U657 ( .A1(n14816), .A2(n14815), .ZN(n15813) );
  BUF_X1 U1289 ( .A(n18667), .Z(n18666) );
  XNOR2_X2 U11221 ( .A(n7200), .B(n7199), .ZN(n8313) );
  OR2_X2 U559 ( .A1(n104), .A2(n11450), .ZN(n12523) );
  AND2_X2 U472 ( .A1(n2077), .A2(n2076), .ZN(n5401) );
  MUX2_X1 U4538 ( .A(n5561), .B(n5560), .S(n5559), .Z(n7080) );
  BUF_X2 U892 ( .A(n7568), .Z(n7864) );
  AOI22_X1 U1510 ( .A1(n12064), .A2(n12063), .B1(n12201), .B2(n12062), .ZN(
        n13027) );
  BUF_X2 U841 ( .A(n14425), .Z(n14424) );
  AOI21_X1 U26 ( .B1(n8692), .B2(n8691), .A(n8690), .ZN(n12349) );
  OAI22_X1 U31 ( .A1(n3220), .A2(n3221), .B1(n7311), .B2(n7343), .ZN(n8928) );
  BUF_X1 U75 ( .A(n13468), .Z(n13818) );
  BUF_X1 U84 ( .A(n10179), .Z(n19839) );
  BUF_X1 U97 ( .A(n14829), .Z(n19986) );
  BUF_X1 U105 ( .A(n18858), .Z(n19989) );
  XNOR2_X1 U112 ( .A(n2991), .B(n2992), .ZN(n17831) );
  NAND2_X1 U122 ( .A1(n16467), .A2(n60), .ZN(n18453) );
  OR2_X2 U127 ( .A1(n3791), .A2(n3794), .ZN(n8846) );
  NOR2_X2 U136 ( .A1(n11128), .A2(n2029), .ZN(n12382) );
  OAI21_X2 U142 ( .B1(n10878), .B2(n10879), .A(n10877), .ZN(n19854) );
  XNOR2_X2 U165 ( .A(n13007), .B(n13006), .ZN(n14648) );
  AOI21_X2 U167 ( .B1(n10888), .B2(n10887), .A(n10886), .ZN(n12609) );
  NAND2_X2 U185 ( .A1(n13915), .A2(n3222), .ZN(n15864) );
  OAI211_X2 U197 ( .C1(n14093), .C2(n14094), .A(n12802), .B(n12801), .ZN(
        n15469) );
  XOR2_X1 U203 ( .A(n15969), .B(n15968), .Z(n19973) );
  XOR2_X1 U217 ( .A(n14942), .B(n14943), .Z(n19975) );
  MUX2_X2 U259 ( .A(n8009), .B(n8008), .S(n8314), .Z(n8831) );
  XNOR2_X2 U306 ( .A(n17285), .B(n17284), .ZN(n18238) );
  AOI21_X2 U309 ( .B1(n13990), .B2(n13991), .A(n15303), .ZN(n16566) );
  NAND3_X2 U340 ( .A1(n14212), .A2(n14211), .A3(n3274), .ZN(n15618) );
  AND3_X2 U353 ( .A1(n2823), .A2(n16265), .A3(n2822), .ZN(n19209) );
  NAND3_X2 U373 ( .A1(n1095), .A2(n5287), .A3(n5288), .ZN(n7266) );
  BUF_X1 U382 ( .A(n5589), .Z(n19980) );
  OAI211_X1 U388 ( .C1(n5091), .C2(n5090), .A(n1360), .B(n5089), .ZN(n5589) );
  BUF_X2 U395 ( .A(n12800), .Z(n19485) );
  XNOR2_X2 U418 ( .A(n16208), .B(n16207), .ZN(n17564) );
  XNOR2_X2 U423 ( .A(n12753), .B(n12752), .ZN(n14828) );
  NAND4_X2 U425 ( .A1(n15786), .A2(n15785), .A3(n15787), .A4(n15784), .ZN(
        n16278) );
  NOR2_X2 U427 ( .A1(n15623), .A2(n15624), .ZN(n16960) );
  NAND3_X2 U428 ( .A1(n5994), .A2(n5993), .A3(n5992), .ZN(n7050) );
  XNOR2_X2 U456 ( .A(n12319), .B(n12318), .ZN(n14796) );
  NAND3_X2 U468 ( .A1(n2346), .A2(n11017), .A3(n2345), .ZN(n13767) );
  XNOR2_X1 U491 ( .A(n13214), .B(n13213), .ZN(n14022) );
  NAND2_X2 U508 ( .A1(n1380), .A2(n3707), .ZN(n13048) );
  AND3_X2 U509 ( .A1(n6847), .A2(n6846), .A3(n6845), .ZN(n9307) );
  AND2_X2 U514 ( .A1(n20342), .A2(n20341), .ZN(n17355) );
  XNOR2_X2 U521 ( .A(n17009), .B(n17008), .ZN(n18928) );
  NAND3_X2 U522 ( .A1(n12220), .A2(n3360), .A3(n3359), .ZN(n12230) );
  MUX2_X2 U541 ( .A(n5427), .B(n5426), .S(n5668), .Z(n7116) );
  NAND3_X2 U545 ( .A1(n9237), .A2(n3060), .A3(n3059), .ZN(n10484) );
  BUF_X2 U549 ( .A(n16320), .Z(n17471) );
  OAI21_X2 U576 ( .B1(n10692), .B2(n19851), .A(n10691), .ZN(n12631) );
  NAND2_X2 U584 ( .A1(n19608), .A2(n19607), .ZN(n15741) );
  OR2_X1 U585 ( .A1(n8301), .A2(n2792), .ZN(n8047) );
  XNOR2_X2 U586 ( .A(n5214), .B(n5213), .ZN(n8301) );
  XNOR2_X2 U626 ( .A(n16536), .B(n16537), .ZN(n19360) );
  OAI21_X2 U627 ( .B1(n13094), .B2(n15120), .A(n13093), .ZN(n15686) );
  INV_X1 U628 ( .A(n9017), .ZN(n19564) );
  XNOR2_X2 U641 ( .A(n3947), .B(Key[180]), .ZN(n4548) );
  NOR2_X2 U647 ( .A1(n16631), .A2(n16630), .ZN(n18365) );
  XNOR2_X2 U656 ( .A(n8719), .B(n8718), .ZN(n11168) );
  NOR2_X2 U677 ( .A1(n5731), .A2(n1476), .ZN(n6743) );
  BUF_X1 U700 ( .A(n11191), .Z(n19983) );
  XNOR2_X1 U707 ( .A(n10547), .B(n10546), .ZN(n11191) );
  NOR2_X2 U721 ( .A1(n8666), .A2(n9781), .ZN(n10595) );
  OAI21_X2 U723 ( .B1(n2988), .B2(n15170), .A(n13993), .ZN(n16926) );
  NAND2_X2 U725 ( .A1(n5982), .A2(n5981), .ZN(n7047) );
  OAI21_X2 U737 ( .B1(n8110), .B2(n8151), .A(n8109), .ZN(n9330) );
  BUF_X1 U743 ( .A(n14829), .Z(n19985) );
  XNOR2_X1 U757 ( .A(n12739), .B(n12738), .ZN(n14829) );
  XNOR2_X2 U764 ( .A(n3858), .B(Key[91]), .ZN(n4405) );
  OR2_X2 U775 ( .A1(n5503), .A2(n5508), .ZN(n5914) );
  NAND2_X2 U778 ( .A1(n15415), .A2(n15414), .ZN(n17133) );
  AND3_X2 U809 ( .A1(n2249), .A2(n3443), .A3(n3442), .ZN(n15636) );
  OAI21_X2 U823 ( .B1(n12076), .B2(n12075), .A(n3269), .ZN(n13659) );
  AND3_X2 U824 ( .A1(n1619), .A2(n1621), .A3(n1622), .ZN(n6966) );
  BUF_X1 U837 ( .A(n18858), .Z(n19988) );
  OAI211_X1 U850 ( .C1(n18023), .C2(n18936), .A(n18022), .B(n18021), .ZN(
        n18858) );
  XNOR2_X2 U866 ( .A(n7398), .B(n7399), .ZN(n8026) );
  OAI21_X2 U880 ( .B1(n745), .B2(n9578), .A(n744), .ZN(n10261) );
  OAI21_X2 U887 ( .B1(n5912), .B2(n4876), .A(n4875), .ZN(n7184) );
  OAI21_X2 U899 ( .B1(n7859), .B2(n7556), .A(n6550), .ZN(n9241) );
  BUF_X2 U902 ( .A(n11129), .Z(n11418) );
  OAI21_X2 U912 ( .B1(n4958), .B2(n4959), .A(n20339), .ZN(n5569) );
  OAI211_X2 U922 ( .C1(n11977), .C2(n11800), .A(n11799), .B(n11798), .ZN(
        n13810) );
  OAI22_X2 U923 ( .A1(n1268), .A2(n1267), .B1(n7654), .B2(n7653), .ZN(n10456)
         );
  NAND3_X2 U926 ( .A1(n2054), .A2(n12058), .A3(n2052), .ZN(n13658) );
  NOR2_X2 U929 ( .A1(n3670), .A2(n11146), .ZN(n12281) );
  BUF_X1 U939 ( .A(n19040), .Z(n19992) );
  CLKBUF_X1 U940 ( .A(n19040), .Z(n19993) );
  NOR2_X1 U942 ( .A1(n17698), .A2(n17697), .ZN(n19040) );
  OAI211_X2 U945 ( .C1(n9226), .C2(n9053), .A(n1759), .B(n9227), .ZN(n10087)
         );
  XNOR2_X2 U947 ( .A(n6628), .B(n6629), .ZN(n8178) );
  XNOR2_X2 U948 ( .A(n6310), .B(n6311), .ZN(n7984) );
  NOR2_X2 U966 ( .A1(n3502), .A2(n3501), .ZN(n10296) );
  NOR2_X2 U972 ( .A1(n1175), .A2(n9791), .ZN(n12508) );
  OAI21_X2 U974 ( .B1(n11983), .B2(n11635), .A(n11634), .ZN(n13734) );
  XNOR2_X2 U988 ( .A(Key[86]), .B(Plaintext[86]), .ZN(n4410) );
  OAI211_X2 U998 ( .C1(n18128), .C2(n18129), .A(n17780), .B(n17779), .ZN(
        n18803) );
  XNOR2_X2 U999 ( .A(n547), .B(Key[188]), .ZN(n4365) );
  XNOR2_X2 U1056 ( .A(Key[163]), .B(Plaintext[163]), .ZN(n4350) );
  OAI21_X2 U1070 ( .B1(n5003), .B2(n4253), .A(n99), .ZN(n6133) );
  AOI21_X2 U1089 ( .B1(n11895), .B2(n11894), .A(n11893), .ZN(n13422) );
  OR2_X1 U1110 ( .A1(n18847), .A2(n3028), .ZN(n20041) );
  BUF_X1 U1114 ( .A(n18454), .Z(n18466) );
  INV_X1 U1118 ( .A(n15529), .ZN(n19997) );
  NAND2_X1 U1145 ( .A1(n16472), .A2(n16473), .ZN(n18465) );
  XNOR2_X1 U1234 ( .A(n3093), .B(n3090), .ZN(n16306) );
  XNOR2_X1 U1266 ( .A(n16069), .B(n16068), .ZN(n17881) );
  OR2_X1 U1279 ( .A1(n12930), .A2(n12929), .ZN(n231) );
  OAI211_X1 U1295 ( .C1(n922), .C2(n11946), .A(n10792), .B(n10791), .ZN(n13336) );
  INV_X1 U1296 ( .A(n11192), .ZN(n19998) );
  INV_X1 U1301 ( .A(n11526), .ZN(n19999) );
  INV_X1 U1303 ( .A(n1449), .ZN(n20000) );
  BUF_X1 U1304 ( .A(n9310), .Z(n20011) );
  INV_X1 U1327 ( .A(n8100), .ZN(n8112) );
  INV_X1 U1333 ( .A(n3748), .ZN(n20001) );
  INV_X1 U1347 ( .A(n5081), .ZN(n20002) );
  CLKBUF_X1 U1353 ( .A(Key[57]), .Z(n18177) );
  CLKBUF_X1 U1368 ( .A(Key[185]), .Z(n645) );
  OR2_X1 U1384 ( .A1(n19130), .A2(n19125), .ZN(n3142) );
  OAI21_X1 U1410 ( .B1(n17499), .B2(n16480), .A(n16479), .ZN(n18464) );
  OR2_X1 U1423 ( .A1(n18157), .A2(n18057), .ZN(n18158) );
  BUF_X2 U1426 ( .A(n18652), .Z(n19934) );
  OAI21_X1 U1451 ( .B1(n17385), .B2(n17384), .A(n17383), .ZN(n20276) );
  AND2_X1 U1455 ( .A1(n17319), .A2(n17318), .ZN(n18172) );
  INV_X1 U1488 ( .A(n18400), .ZN(n20003) );
  OR2_X1 U1518 ( .A1(n16543), .A2(n20240), .ZN(n20065) );
  OAI211_X1 U1525 ( .C1(n16677), .C2(n16676), .A(n16675), .B(n2206), .ZN(
        n20152) );
  XNOR2_X1 U1606 ( .A(n16774), .B(n16773), .ZN(n20221) );
  XNOR2_X1 U1624 ( .A(n17018), .B(n17017), .ZN(n18938) );
  XNOR2_X1 U1630 ( .A(n17405), .B(n17404), .ZN(n18130) );
  INV_X1 U1639 ( .A(n19389), .ZN(n20004) );
  NAND3_X1 U1648 ( .A1(n20022), .A2(n1757), .A3(n1610), .ZN(n16562) );
  INV_X1 U1691 ( .A(n15696), .ZN(n20005) );
  INV_X1 U1724 ( .A(n231), .ZN(n15166) );
  INV_X1 U1725 ( .A(n15898), .ZN(n20006) );
  INV_X1 U1738 ( .A(n16128), .ZN(n20007) );
  NAND2_X1 U1762 ( .A1(n20284), .A2(n20283), .ZN(n15657) );
  CLKBUF_X1 U1798 ( .A(n11717), .Z(n20215) );
  NAND2_X1 U1804 ( .A1(n8903), .A2(n3279), .ZN(n12002) );
  NAND2_X1 U1805 ( .A1(n11280), .A2(n11279), .ZN(n12488) );
  INV_X1 U1822 ( .A(n3667), .ZN(n20297) );
  NAND3_X1 U1874 ( .A1(n1750), .A2(n529), .A3(n1753), .ZN(n10274) );
  OR2_X1 U1900 ( .A1(n9188), .A2(n268), .ZN(n2014) );
  INV_X1 U1916 ( .A(n9328), .ZN(n20008) );
  INV_X1 U1978 ( .A(n8276), .ZN(n20009) );
  OR2_X1 U2047 ( .A1(n7898), .A2(n2703), .ZN(n20315) );
  OR2_X1 U2065 ( .A1(n8083), .A2(n20107), .ZN(n20086) );
  XNOR2_X1 U2077 ( .A(n3020), .B(n6994), .ZN(n7922) );
  XNOR2_X1 U2095 ( .A(n6304), .B(n6305), .ZN(n7921) );
  INV_X1 U2100 ( .A(n7600), .ZN(n20012) );
  XNOR2_X1 U2113 ( .A(n6233), .B(n6232), .ZN(n7932) );
  XNOR2_X1 U2148 ( .A(n5454), .B(n5453), .ZN(n8286) );
  NAND2_X1 U2160 ( .A1(n804), .A2(n1082), .ZN(n1081) );
  AND2_X1 U2194 ( .A1(n4600), .A2(n30), .ZN(n20203) );
  AND3_X1 U2218 ( .A1(n4998), .A2(n4996), .A3(n4999), .ZN(n20028) );
  NAND4_X1 U2219 ( .A1(n5771), .A2(n5772), .A3(n5774), .A4(n5773), .ZN(n6927)
         );
  INV_X1 U2236 ( .A(n5767), .ZN(n5734) );
  BUF_X1 U2269 ( .A(n4501), .Z(n6204) );
  INV_X1 U2275 ( .A(n5719), .ZN(n5604) );
  NAND2_X1 U2276 ( .A1(n19619), .A2(n4309), .ZN(n4598) );
  INV_X1 U2284 ( .A(n4860), .ZN(n20085) );
  OR2_X1 U2291 ( .A1(n4793), .A2(n5108), .ZN(n5104) );
  CLKBUF_X1 U2292 ( .A(n5112), .Z(n20256) );
  BUF_X1 U2316 ( .A(n4317), .Z(n4325) );
  INV_X1 U2339 ( .A(n5717), .ZN(n20034) );
  OR2_X1 U2345 ( .A1(n4489), .A2(n4488), .ZN(n4501) );
  MUX2_X1 U2373 ( .A(n4226), .B(n4224), .S(n3996), .Z(n3997) );
  OAI211_X1 U2383 ( .C1(n4557), .C2(n4750), .A(n3915), .B(n3914), .ZN(n6049)
         );
  XNOR2_X1 U2396 ( .A(Key[112]), .B(Plaintext[112]), .ZN(n5083) );
  OR2_X1 U2404 ( .A1(n6379), .A2(n5728), .ZN(n1746) );
  AND2_X1 U2419 ( .A1(n20034), .A2(n5719), .ZN(n4368) );
  OR2_X1 U2420 ( .A1(n5328), .A2(n6048), .ZN(n2081) );
  AND2_X1 U2447 ( .A1(n5063), .A2(n5064), .ZN(n20036) );
  INV_X1 U2460 ( .A(n5643), .ZN(n5645) );
  OR2_X1 U2472 ( .A1(n5002), .A2(n5571), .ZN(n20282) );
  CLKBUF_X1 U2473 ( .A(n5276), .Z(n5818) );
  OR2_X1 U2474 ( .A1(n7674), .A2(n8365), .ZN(n8362) );
  INV_X1 U2481 ( .A(n6523), .ZN(n20314) );
  BUF_X1 U2496 ( .A(n6345), .Z(n7504) );
  INV_X1 U2500 ( .A(n9114), .ZN(n20346) );
  INV_X1 U2504 ( .A(n9239), .ZN(n20322) );
  CLKBUF_X1 U2530 ( .A(n8087), .Z(n20254) );
  INV_X1 U2604 ( .A(n9329), .ZN(n20313) );
  AND2_X1 U2605 ( .A1(n9003), .A2(n2883), .ZN(n20037) );
  NAND2_X1 U2609 ( .A1(n7565), .A2(n7566), .ZN(n9362) );
  AND3_X1 U2660 ( .A1(n3311), .A2(n8255), .A3(n769), .ZN(n20146) );
  CLKBUF_X1 U2662 ( .A(n8985), .Z(n19827) );
  OR2_X1 U2705 ( .A1(n9122), .A2(n8812), .ZN(n8457) );
  XNOR2_X1 U2723 ( .A(n10602), .B(n20324), .ZN(n19505) );
  OR2_X1 U2724 ( .A1(n20366), .A2(n11142), .ZN(n10961) );
  AOI22_X1 U2735 ( .A1(n12107), .A2(n12104), .B1(n3186), .B2(n3601), .ZN(
        n11633) );
  INV_X1 U2741 ( .A(n12008), .ZN(n12507) );
  XNOR2_X1 U2787 ( .A(n13047), .B(n20053), .ZN(n12676) );
  INV_X1 U2790 ( .A(n12258), .ZN(n13146) );
  XNOR2_X1 U2799 ( .A(n2189), .B(n13252), .ZN(n14268) );
  OAI21_X1 U2848 ( .B1(n12655), .B2(n14788), .A(n14790), .ZN(n20284) );
  XNOR2_X1 U2861 ( .A(n12587), .B(n12588), .ZN(n14787) );
  CLKBUF_X1 U2862 ( .A(n14679), .Z(n20120) );
  INV_X1 U2908 ( .A(n15505), .ZN(n20288) );
  INV_X1 U2949 ( .A(n15221), .ZN(n15665) );
  NOR2_X1 U2972 ( .A1(n15204), .A2(n15756), .ZN(n15208) );
  INV_X1 U3011 ( .A(n16129), .ZN(n747) );
  NAND4_X1 U3079 ( .A1(n2815), .A2(n15758), .A3(n15757), .A4(n15760), .ZN(n66)
         );
  OR2_X1 U3102 ( .A1(n15540), .A2(n20006), .ZN(n14911) );
  AND2_X1 U3127 ( .A1(n15661), .A2(n15662), .ZN(n20021) );
  INV_X1 U3128 ( .A(n16295), .ZN(n16880) );
  OAI21_X1 U3157 ( .B1(n15765), .B2(n15248), .A(n15247), .ZN(n19893) );
  XNOR2_X1 U3164 ( .A(n16964), .B(n14987), .ZN(n16284) );
  XNOR2_X1 U3169 ( .A(n16044), .B(n17407), .ZN(n16769) );
  OR2_X1 U3186 ( .A1(n17690), .A2(n17691), .ZN(n20307) );
  XNOR2_X1 U3232 ( .A(n963), .B(n17140), .ZN(n3066) );
  INV_X1 U3253 ( .A(n18620), .ZN(n19509) );
  OR2_X1 U3394 ( .A1(n16155), .A2(n18057), .ZN(n19169) );
  CLKBUF_X1 U3422 ( .A(Key[159]), .Z(n2079) );
  CLKBUF_X1 U3442 ( .A(Key[93]), .Z(n2263) );
  CLKBUF_X1 U3460 ( .A(Key[41]), .Z(n345) );
  NAND3_X1 U3532 ( .A1(n13950), .A2(n14690), .A3(n14688), .ZN(n20014) );
  NAND2_X1 U3558 ( .A1(n4855), .A2(n4907), .ZN(n20015) );
  XOR2_X1 U3644 ( .A(Key[108]), .B(Plaintext[108]), .Z(n20016) );
  INV_X1 U3680 ( .A(n5859), .ZN(n20334) );
  OR2_X1 U3710 ( .A1(n4714), .A2(n4788), .ZN(n20017) );
  INV_X1 U3753 ( .A(n4501), .ZN(n6218) );
  INV_X1 U3790 ( .A(n2792), .ZN(n20057) );
  INV_X1 U3845 ( .A(n12514), .ZN(n20073) );
  XOR2_X1 U3849 ( .A(n13778), .B(n13266), .Z(n20018) );
  INV_X1 U3860 ( .A(n19043), .ZN(n20074) );
  XOR2_X1 U3901 ( .A(n16092), .B(n16093), .Z(n20019) );
  NAND2_X1 U4044 ( .A1(n1354), .A2(n8208), .ZN(n20020) );
  XNOR2_X1 U4063 ( .A(n16295), .B(n20100), .ZN(n16297) );
  NAND2_X1 U4074 ( .A1(n5610), .A2(n6152), .ZN(n6160) );
  NAND2_X1 U4086 ( .A1(n659), .A2(n2533), .ZN(n19270) );
  NAND2_X1 U4091 ( .A1(n20015), .A2(n4499), .ZN(n3706) );
  NAND3_X1 U4105 ( .A1(n1613), .A2(n1615), .A3(n1758), .ZN(n20022) );
  AND2_X2 U4150 ( .A1(n20023), .A2(n2969), .ZN(n17002) );
  OAI21_X1 U4156 ( .B1(n15399), .B2(n2968), .A(n197), .ZN(n20023) );
  NOR2_X1 U4201 ( .A1(n276), .A2(n20024), .ZN(n3076) );
  NAND2_X1 U4320 ( .A1(n8001), .A2(n2548), .ZN(n20024) );
  INV_X1 U4326 ( .A(n6871), .ZN(n8140) );
  XNOR2_X1 U4335 ( .A(n6862), .B(n6861), .ZN(n6871) );
  NAND3_X1 U4338 ( .A1(n19662), .A2(n15061), .A3(n15309), .ZN(n14989) );
  NAND3_X1 U4387 ( .A1(n20025), .A2(n15637), .A3(n15638), .ZN(n19611) );
  NAND3_X1 U4443 ( .A1(n20063), .A2(n230), .A3(n15843), .ZN(n20025) );
  XNOR2_X1 U4526 ( .A(n13108), .B(n13711), .ZN(n12923) );
  NOR2_X2 U4528 ( .A1(n11847), .A2(n11848), .ZN(n13711) );
  NAND2_X1 U4619 ( .A1(n12095), .A2(n12429), .ZN(n11611) );
  NAND2_X1 U4701 ( .A1(n3046), .A2(n3295), .ZN(n20026) );
  INV_X1 U4711 ( .A(n10725), .ZN(n20027) );
  NAND2_X1 U4722 ( .A1(n5442), .A2(n5641), .ZN(n4165) );
  OAI21_X1 U4741 ( .B1(n8327), .B2(n9104), .A(n8326), .ZN(n10048) );
  NAND2_X1 U4750 ( .A1(n7800), .A2(n7799), .ZN(n2627) );
  NAND2_X2 U4777 ( .A1(n4997), .A2(n20028), .ZN(n7318) );
  OAI21_X1 U4786 ( .B1(n3806), .B2(n9304), .A(n9298), .ZN(n20029) );
  OAI211_X1 U4787 ( .C1(n17943), .C2(n3038), .A(n1450), .B(n3036), .ZN(n3035)
         );
  INV_X1 U4801 ( .A(n10329), .ZN(n10327) );
  NAND2_X1 U4829 ( .A1(n2451), .A2(n13939), .ZN(n20030) );
  INV_X1 U4850 ( .A(n20031), .ZN(Ciphertext[26]) );
  OAI211_X1 U4928 ( .C1(n17743), .C2(n17742), .A(n17740), .B(n17741), .ZN(
        n20031) );
  NAND3_X1 U4985 ( .A1(n7703), .A2(n7542), .A3(n19881), .ZN(n7544) );
  NOR2_X1 U4998 ( .A1(n10505), .A2(n10836), .ZN(n10523) );
  OAI21_X1 U5019 ( .B1(n300), .B2(n18495), .A(n20033), .ZN(n17731) );
  NAND3_X1 U5047 ( .A1(n18495), .A2(n300), .A3(n17729), .ZN(n20033) );
  NAND3_X1 U5088 ( .A1(n9303), .A2(n9302), .A3(n3788), .ZN(n10598) );
  NAND2_X1 U5117 ( .A1(n19922), .A2(n7871), .ZN(n7422) );
  NAND2_X1 U5141 ( .A1(n5595), .A2(n5519), .ZN(n3409) );
  AOI21_X2 U5143 ( .B1(n9557), .B2(n9558), .A(n9556), .ZN(n11659) );
  NOR2_X2 U5185 ( .A1(n61), .A2(n4346), .ZN(n5719) );
  NAND3_X1 U5208 ( .A1(n20035), .A2(n7618), .A3(n586), .ZN(n2097) );
  NAND2_X1 U5255 ( .A1(n11387), .A2(n11386), .ZN(n11393) );
  NAND2_X1 U5264 ( .A1(n20038), .A2(n4943), .ZN(n4949) );
  NAND2_X1 U5284 ( .A1(n4941), .A2(n4940), .ZN(n20038) );
  NOR2_X1 U5288 ( .A1(n18630), .A2(n19509), .ZN(n20039) );
  AND2_X1 U5304 ( .A1(n14819), .A2(n14818), .ZN(n20040) );
  NAND2_X1 U5320 ( .A1(n15241), .A2(n15242), .ZN(n17279) );
  NAND2_X1 U5323 ( .A1(n12260), .A2(n19603), .ZN(n13762) );
  NAND3_X1 U5348 ( .A1(n3027), .A2(n20042), .A3(n20041), .ZN(n1374) );
  NAND2_X1 U5352 ( .A1(n18853), .A2(n3030), .ZN(n20042) );
  NAND2_X1 U5377 ( .A1(n8377), .A2(n8370), .ZN(n7541) );
  NAND2_X1 U5437 ( .A1(n4764), .A2(n4269), .ZN(n20043) );
  NOR2_X1 U5472 ( .A1(n4737), .A2(n20044), .ZN(n19559) );
  INV_X1 U5474 ( .A(n4732), .ZN(n20044) );
  NAND2_X1 U5494 ( .A1(n4734), .A2(n4277), .ZN(n4732) );
  NAND3_X1 U5571 ( .A1(n14419), .A2(n14418), .A3(n14359), .ZN(n3636) );
  NAND2_X1 U5637 ( .A1(n20047), .A2(n20045), .ZN(n15253) );
  NAND2_X1 U5661 ( .A1(n20046), .A2(n17243), .ZN(n20045) );
  NAND2_X1 U5675 ( .A1(n17480), .A2(n20353), .ZN(n20046) );
  NAND2_X1 U5772 ( .A1(n15252), .A2(n17241), .ZN(n20047) );
  NAND2_X1 U5790 ( .A1(n20048), .A2(n18399), .ZN(n18402) );
  OAI21_X1 U5793 ( .B1(n18407), .B2(n18412), .A(n20003), .ZN(n20048) );
  XNOR2_X1 U5798 ( .A(n20050), .B(n20049), .ZN(Ciphertext[99]) );
  INV_X1 U5854 ( .A(n18055), .ZN(n20049) );
  NAND2_X1 U5874 ( .A1(n20052), .A2(n20051), .ZN(n20050) );
  NAND2_X1 U5890 ( .A1(n18054), .A2(n18869), .ZN(n20051) );
  INV_X1 U5902 ( .A(n2222), .ZN(n20053) );
  NAND2_X1 U5912 ( .A1(n12178), .A2(n2260), .ZN(n13047) );
  NAND3_X1 U5921 ( .A1(n18648), .A2(n19745), .A3(n18654), .ZN(n582) );
  NOR2_X2 U5924 ( .A1(n12314), .A2(n2338), .ZN(n13309) );
  NAND2_X1 U5937 ( .A1(n63), .A2(n20054), .ZN(n10151) );
  NAND2_X1 U5951 ( .A1(n369), .A2(n257), .ZN(n11607) );
  AND2_X2 U5963 ( .A1(n8147), .A2(n8148), .ZN(n9346) );
  NAND3_X1 U5983 ( .A1(n20056), .A2(n8301), .A3(n20055), .ZN(n7452) );
  NAND2_X1 U5984 ( .A1(n8304), .A2(n2792), .ZN(n20055) );
  NAND2_X1 U6035 ( .A1(n20057), .A2(n8305), .ZN(n20056) );
  INV_X1 U6096 ( .A(n20059), .ZN(n20058) );
  OAI21_X1 U6104 ( .B1(n4951), .B2(n4911), .A(n4477), .ZN(n20059) );
  NAND2_X1 U6116 ( .A1(n4476), .A2(n4958), .ZN(n20060) );
  NAND2_X1 U6123 ( .A1(n15400), .A2(n15892), .ZN(n15540) );
  NAND2_X1 U6161 ( .A1(n15442), .A2(n15676), .ZN(n15678) );
  XNOR2_X1 U6181 ( .A(n20061), .B(n18084), .ZN(n8776) );
  NAND2_X1 U6195 ( .A1(n8775), .A2(n2882), .ZN(n20061) );
  NAND2_X1 U6225 ( .A1(n1792), .A2(n3592), .ZN(n3591) );
  NAND2_X1 U6230 ( .A1(n397), .A2(n8295), .ZN(n9100) );
  XNOR2_X1 U6235 ( .A(n13233), .B(n20018), .ZN(n13235) );
  NAND3_X1 U6242 ( .A1(n20062), .A2(n4286), .A3(n4287), .ZN(n1985) );
  NAND2_X1 U6250 ( .A1(n4288), .A2(n4623), .ZN(n20062) );
  OR2_X1 U6328 ( .A1(n7848), .A2(n8079), .ZN(n7849) );
  NAND2_X1 U6338 ( .A1(n19354), .A2(n16540), .ZN(n17234) );
  INV_X1 U6343 ( .A(n15845), .ZN(n20063) );
  NAND2_X1 U6346 ( .A1(n4913), .A2(n4914), .ZN(n4915) );
  NAND2_X1 U6348 ( .A1(n16542), .A2(n20065), .ZN(n19339) );
  NAND2_X1 U6353 ( .A1(n16541), .A2(n19352), .ZN(n16542) );
  NAND2_X1 U6392 ( .A1(n20014), .A2(n20066), .ZN(n15221) );
  NAND2_X1 U6443 ( .A1(n13365), .A2(n14696), .ZN(n20066) );
  NAND2_X1 U6448 ( .A1(n20068), .A2(n20067), .ZN(n5612) );
  NAND3_X1 U6455 ( .A1(n4392), .A2(n4681), .A3(n4486), .ZN(n20067) );
  NAND2_X1 U6462 ( .A1(n4390), .A2(n4389), .ZN(n20068) );
  NAND2_X1 U6463 ( .A1(n19347), .A2(n16673), .ZN(n16635) );
  OAI211_X1 U6472 ( .C1(n18365), .C2(n18364), .A(n20070), .B(n20069), .ZN(
        n18368) );
  OR2_X1 U6481 ( .A1(n18360), .A2(n17936), .ZN(n20069) );
  NAND2_X1 U6491 ( .A1(n20071), .A2(n18360), .ZN(n20070) );
  INV_X1 U6500 ( .A(n18361), .ZN(n20071) );
  NAND2_X1 U6509 ( .A1(n19956), .A2(n17508), .ZN(n20072) );
  NOR2_X1 U6519 ( .A1(n12323), .A2(n20073), .ZN(n2658) );
  NAND2_X1 U6520 ( .A1(n12326), .A2(n11997), .ZN(n12323) );
  OAI22_X1 U6539 ( .A1(n19045), .A2(n20074), .B1(n19047), .B2(n19992), .ZN(
        n18083) );
  NAND3_X2 U6547 ( .A1(n15869), .A2(n20077), .A3(n20076), .ZN(n17124) );
  NAND2_X1 U6549 ( .A1(n15865), .A2(n15864), .ZN(n20076) );
  NAND2_X1 U6564 ( .A1(n15867), .A2(n15866), .ZN(n20077) );
  NAND2_X2 U6586 ( .A1(n28), .A2(n20079), .ZN(n15720) );
  NAND2_X1 U6634 ( .A1(n1350), .A2(n1352), .ZN(n20079) );
  AND3_X2 U6660 ( .A1(n3417), .A2(n1012), .A3(n3416), .ZN(n10430) );
  OAI21_X2 U6673 ( .B1(n11775), .B2(n11180), .A(n11181), .ZN(n13833) );
  NAND2_X1 U6732 ( .A1(n7459), .A2(n2021), .ZN(n1567) );
  INV_X1 U6735 ( .A(n5861), .ZN(n5615) );
  NAND2_X1 U6741 ( .A1(n5859), .A2(n3188), .ZN(n5861) );
  NAND2_X1 U6772 ( .A1(n15078), .A2(n2723), .ZN(n14479) );
  OR3_X1 U6797 ( .A1(n17676), .A2(n20512), .A3(n17867), .ZN(n16000) );
  NAND3_X1 U6830 ( .A1(n3283), .A2(n3285), .A3(n16734), .ZN(n19135) );
  NAND3_X1 U6851 ( .A1(n16733), .A2(n3287), .A3(n16732), .ZN(n16734) );
  NAND2_X1 U6889 ( .A1(n20080), .A2(n2089), .ZN(n7896) );
  NAND2_X1 U6905 ( .A1(n20082), .A2(n20504), .ZN(n20080) );
  OAI21_X1 U6918 ( .B1(n8184), .B2(n8059), .A(n7892), .ZN(n20082) );
  OAI21_X1 U6948 ( .B1(n18613), .B2(n18625), .A(n18629), .ZN(n18179) );
  NAND2_X1 U6949 ( .A1(n18622), .A2(n19679), .ZN(n18629) );
  NAND3_X1 U7002 ( .A1(n3085), .A2(n17506), .A3(n975), .ZN(n19773) );
  NAND2_X1 U7007 ( .A1(n339), .A2(n16480), .ZN(n3085) );
  NAND2_X1 U7022 ( .A1(n3252), .A2(n14468), .ZN(n13924) );
  XNOR2_X2 U7115 ( .A(n12706), .B(n12705), .ZN(n14468) );
  NAND2_X2 U7116 ( .A1(n20084), .A2(n20083), .ZN(n6068) );
  NAND3_X1 U7124 ( .A1(n3989), .A2(n4860), .A3(n4498), .ZN(n20083) );
  NAND2_X1 U7135 ( .A1(n3991), .A2(n20085), .ZN(n20084) );
  NAND2_X1 U7140 ( .A1(n12508), .A2(n12008), .ZN(n126) );
  AND2_X2 U7153 ( .A1(n12362), .A2(n12363), .ZN(n12008) );
  NAND2_X1 U7188 ( .A1(n2188), .A2(n20086), .ZN(n8089) );
  OAI21_X1 U7233 ( .B1(n1211), .B2(n8705), .A(n20087), .ZN(n2776) );
  NAND2_X1 U7264 ( .A1(n2777), .A2(n1211), .ZN(n20087) );
  NAND3_X1 U7378 ( .A1(n20088), .A2(n5075), .A3(n5076), .ZN(n448) );
  NAND2_X1 U7405 ( .A1(n5074), .A2(n5080), .ZN(n20088) );
  NOR2_X2 U7406 ( .A1(n11705), .A2(n20089), .ZN(n13623) );
  AOI21_X1 U7424 ( .B1(n11702), .B2(n11703), .A(n11701), .ZN(n20089) );
  NAND2_X1 U7425 ( .A1(n17557), .A2(n2797), .ZN(n18620) );
  INV_X1 U7471 ( .A(n20090), .ZN(n18315) );
  OAI22_X1 U7472 ( .A1(n18309), .A2(n19340), .B1(n19309), .B2(n19311), .ZN(
        n20090) );
  XOR2_X1 U7554 ( .A(n17034), .B(n17032), .Z(n17039) );
  OR2_X1 U7562 ( .A1(n20091), .A2(n19758), .ZN(n3579) );
  NAND2_X1 U7570 ( .A1(n19526), .A2(n18511), .ZN(n20091) );
  INV_X1 U7592 ( .A(n18057), .ZN(n1035) );
  XOR2_X1 U7606 ( .A(n13097), .B(n13400), .Z(n13102) );
  XNOR2_X1 U7629 ( .A(n14942), .B(n14943), .ZN(n20092) );
  OAI21_X1 U7644 ( .B1(n20330), .B2(n14352), .A(n20329), .ZN(n14329) );
  MUX2_X1 U7657 ( .A(n17455), .B(n17983), .S(n20132), .Z(n20093) );
  NAND2_X1 U7684 ( .A1(n17313), .A2(n17312), .ZN(n18834) );
  OR2_X1 U7686 ( .A1(n17790), .A2(n17791), .ZN(n17794) );
  BUF_X1 U7717 ( .A(n15876), .Z(n20094) );
  OAI22_X1 U7720 ( .A1(n2675), .A2(n3366), .B1(n2678), .B2(n2677), .ZN(n15876)
         );
  XNOR2_X1 U7738 ( .A(n9673), .B(n9672), .ZN(n20095) );
  AOI21_X1 U7790 ( .B1(n3116), .B2(n19667), .A(n3115), .ZN(n18151) );
  NAND2_X1 U7826 ( .A1(n17319), .A2(n17318), .ZN(n20097) );
  XNOR2_X1 U7835 ( .A(n9604), .B(n9603), .ZN(n11290) );
  BUF_X1 U7836 ( .A(n17281), .Z(n20098) );
  OAI211_X1 U7840 ( .C1(n15885), .C2(n16012), .A(n13970), .B(n13969), .ZN(
        n17281) );
  MUX2_X2 U7851 ( .A(n19111), .B(n19106), .S(n19110), .Z(n19093) );
  XNOR2_X1 U7852 ( .A(n10097), .B(n10096), .ZN(n20099) );
  XNOR2_X1 U7880 ( .A(n10097), .B(n10096), .ZN(n11360) );
  AOI22_X2 U7931 ( .A1(n12092), .A2(n12091), .B1(n12090), .B2(n12089), .ZN(
        n13462) );
  CLKBUF_X1 U7934 ( .A(n14112), .Z(n15423) );
  AOI22_X1 U7948 ( .A1(n15197), .A2(n15198), .B1(n15500), .B2(n15196), .ZN(
        n20100) );
  AOI22_X1 U7961 ( .A1(n15197), .A2(n15198), .B1(n15500), .B2(n15196), .ZN(
        n16746) );
  XNOR2_X1 U7962 ( .A(n17415), .B(n17414), .ZN(n20101) );
  XNOR2_X1 U7978 ( .A(n15764), .B(n15763), .ZN(n20240) );
  NAND3_X2 U7982 ( .A1(n11941), .A2(n11940), .A3(n1400), .ZN(n13390) );
  AOI21_X1 U8002 ( .B1(n15725), .B2(n15724), .A(n15723), .ZN(n20102) );
  AOI21_X1 U8020 ( .B1(n15725), .B2(n15724), .A(n15723), .ZN(n16407) );
  INV_X1 U8030 ( .A(n15165), .ZN(n20103) );
  BUF_X1 U8063 ( .A(n12888), .Z(n19513) );
  NAND3_X1 U8065 ( .A1(n2007), .A2(n15161), .A3(n2293), .ZN(n20104) );
  NAND3_X1 U8096 ( .A1(n2007), .A2(n15161), .A3(n2293), .ZN(n17299) );
  XNOR2_X1 U8098 ( .A(n3831), .B(Key[70]), .ZN(n20105) );
  BUF_X1 U8108 ( .A(n11515), .Z(n20106) );
  XNOR2_X1 U8161 ( .A(n3831), .B(Key[70]), .ZN(n4420) );
  XNOR2_X1 U8164 ( .A(n9982), .B(n9981), .ZN(n11515) );
  XNOR2_X1 U8177 ( .A(n6549), .B(n6548), .ZN(n20107) );
  XNOR2_X1 U8180 ( .A(n6549), .B(n6548), .ZN(n20108) );
  XNOR2_X1 U8197 ( .A(n16428), .B(n16427), .ZN(n20109) );
  OAI21_X1 U8225 ( .B1(n3081), .B2(n17507), .A(n3080), .ZN(n20110) );
  OAI21_X2 U8362 ( .B1(n15052), .B2(n15053), .A(n15051), .ZN(n16873) );
  NAND2_X1 U8368 ( .A1(n1106), .A2(n3388), .ZN(n20111) );
  NAND2_X1 U8372 ( .A1(n14616), .A2(n14615), .ZN(n20112) );
  BUF_X1 U8376 ( .A(n2748), .Z(n20113) );
  XOR2_X1 U8382 ( .A(n16361), .B(n16362), .Z(n20114) );
  OAI21_X1 U8400 ( .B1(n7984), .B2(n7921), .A(n1726), .ZN(n502) );
  NOR2_X1 U8404 ( .A1(n8948), .A2(n528), .ZN(n20115) );
  NOR2_X1 U8429 ( .A1(n8948), .A2(n528), .ZN(n10527) );
  OR2_X1 U8441 ( .A1(n18036), .A2(n18035), .ZN(n20117) );
  OR2_X1 U8449 ( .A1(n15733), .A2(n3431), .ZN(n15736) );
  OR2_X1 U8450 ( .A1(n11360), .A2(n10112), .ZN(n11358) );
  NAND3_X1 U8647 ( .A1(n1469), .A2(n13960), .A3(n13959), .ZN(n15879) );
  NOR2_X1 U8653 ( .A1(n15098), .A2(n15099), .ZN(n20121) );
  XNOR2_X1 U8720 ( .A(n13420), .B(n13421), .ZN(n14679) );
  NOR2_X1 U8727 ( .A1(n15098), .A2(n15099), .ZN(n2542) );
  OAI211_X2 U8792 ( .C1(n12346), .C2(n12497), .A(n12006), .B(n2901), .ZN(
        n13677) );
  NAND2_X1 U8906 ( .A1(n11737), .A2(n11736), .ZN(n20123) );
  AND2_X1 U8909 ( .A1(n2414), .A2(n17866), .ZN(n20124) );
  NAND2_X1 U8921 ( .A1(n11737), .A2(n11736), .ZN(n13695) );
  AOI21_X1 U8949 ( .B1(n15715), .B2(n15716), .A(n20094), .ZN(n73) );
  OAI21_X1 U8950 ( .B1(n14976), .B2(n14977), .A(n14975), .ZN(n20125) );
  OAI21_X1 U8956 ( .B1(n14976), .B2(n14977), .A(n14975), .ZN(n20126) );
  OAI21_X1 U8959 ( .B1(n14976), .B2(n14977), .A(n14975), .ZN(n17327) );
  XNOR2_X1 U9082 ( .A(n16710), .B(n16709), .ZN(n20127) );
  NAND2_X1 U9141 ( .A1(n3205), .A2(n18038), .ZN(n20128) );
  XOR2_X1 U9239 ( .A(n16877), .B(n16876), .Z(n20129) );
  AND2_X1 U9251 ( .A1(n17313), .A2(n17312), .ZN(n20130) );
  NAND2_X1 U9293 ( .A1(n2268), .A2(n17834), .ZN(n20131) );
  NAND2_X1 U9294 ( .A1(n2268), .A2(n17834), .ZN(n19074) );
  XNOR2_X1 U9310 ( .A(n17257), .B(n17256), .ZN(n20132) );
  BUF_X1 U9311 ( .A(n15697), .Z(n20133) );
  AOI22_X1 U9320 ( .A1(n14014), .A2(n14013), .B1(n19488), .B2(n14012), .ZN(
        n15697) );
  AND2_X1 U9322 ( .A1(n8775), .A2(n2882), .ZN(n20134) );
  AOI21_X1 U9372 ( .B1(n12511), .B2(n1609), .A(n12510), .ZN(n12512) );
  INV_X1 U9389 ( .A(n14261), .ZN(n20311) );
  OAI211_X1 U9601 ( .C1(n14227), .C2(n14731), .A(n14226), .B(n14225), .ZN(
        n15422) );
  OR2_X1 U9621 ( .A1(n12657), .A2(n14791), .ZN(n20283) );
  XNOR2_X1 U9622 ( .A(n14915), .B(n15953), .ZN(n20135) );
  OAI21_X1 U9887 ( .B1(n17216), .B2(n17217), .A(n17215), .ZN(n18377) );
  INV_X1 U10070 ( .A(n15619), .ZN(n20138) );
  OR2_X1 U10074 ( .A1(n15309), .A2(n15059), .ZN(n15396) );
  OAI21_X1 U10135 ( .B1(n17596), .B2(n16657), .A(n16656), .ZN(n20140) );
  INV_X1 U10138 ( .A(n14792), .ZN(n20141) );
  OAI21_X1 U10232 ( .B1(n17713), .B2(n20221), .A(n17712), .ZN(n20142) );
  XNOR2_X1 U10284 ( .A(Key[5]), .B(Plaintext[5]), .ZN(n20143) );
  XNOR2_X1 U10490 ( .A(Key[5]), .B(Plaintext[5]), .ZN(n4622) );
  INV_X1 U10523 ( .A(n19942), .ZN(n20144) );
  BUF_X1 U10721 ( .A(n7475), .Z(n19942) );
  INV_X1 U10869 ( .A(n15696), .ZN(n20145) );
  BUF_X1 U10875 ( .A(n18468), .Z(n20148) );
  OAI21_X1 U10965 ( .B1(n1897), .B2(n16483), .A(n16482), .ZN(n18468) );
  OR2_X1 U10966 ( .A1(n11105), .A2(n11104), .ZN(n20300) );
  NAND3_X1 U10995 ( .A1(n5904), .A2(n5903), .A3(n4847), .ZN(n20149) );
  NAND3_X1 U11107 ( .A1(n5904), .A2(n5903), .A3(n4847), .ZN(n6090) );
  OAI21_X1 U11343 ( .B1(n4843), .B2(n4842), .A(n3978), .ZN(n5904) );
  XOR2_X1 U11347 ( .A(n16536), .B(n16537), .Z(n20150) );
  OR2_X1 U11361 ( .A1(n16128), .A2(n15607), .ZN(n15733) );
  BUF_X1 U11374 ( .A(n15671), .Z(n20151) );
  AOI22_X1 U11375 ( .A1(n13459), .A2(n14678), .B1(n13458), .B2(n14550), .ZN(
        n15671) );
  OAI211_X1 U11406 ( .C1(n16677), .C2(n16676), .A(n16675), .B(n2206), .ZN(
        n18067) );
  MUX2_X1 U11492 ( .A(n8970), .B(n7727), .S(n9256), .Z(n7738) );
  OAI21_X1 U11568 ( .B1(n11075), .B2(n11486), .A(n11074), .ZN(n20153) );
  OAI21_X1 U11577 ( .B1(n11075), .B2(n11486), .A(n11074), .ZN(n12253) );
  XNOR2_X1 U11578 ( .A(n7069), .B(n7068), .ZN(n20154) );
  XNOR2_X1 U11590 ( .A(n7069), .B(n7068), .ZN(n7991) );
  OAI211_X1 U11591 ( .C1(n11927), .C2(n11926), .A(n11924), .B(n11925), .ZN(
        n13702) );
  OR2_X1 U11598 ( .A1(n8468), .A2(n8467), .ZN(n20156) );
  INV_X1 U11633 ( .A(n14571), .ZN(n20157) );
  XNOR2_X2 U11647 ( .A(n13229), .B(n13228), .ZN(n14571) );
  OAI211_X2 U11708 ( .C1(n15748), .C2(n19502), .A(n15597), .B(n15596), .ZN(
        n16886) );
  XNOR2_X1 U11760 ( .A(n16890), .B(n16889), .ZN(n20158) );
  XNOR2_X1 U11764 ( .A(n16890), .B(n16889), .ZN(n18975) );
  NAND2_X2 U11867 ( .A1(n19580), .A2(n12395), .ZN(n13259) );
  OR2_X1 U11887 ( .A1(n11174), .A2(n10962), .ZN(n20317) );
  CLKBUF_X1 U11905 ( .A(n2984), .Z(n20159) );
  NOR2_X1 U12004 ( .A1(n17221), .A2(n16639), .ZN(n16641) );
  BUF_X1 U12005 ( .A(n11871), .Z(n20160) );
  BUF_X1 U12119 ( .A(n10332), .Z(n20161) );
  XNOR2_X1 U12141 ( .A(n16074), .B(n16073), .ZN(n20162) );
  NAND3_X1 U12142 ( .A1(n3343), .A2(n3344), .A3(n113), .ZN(n20163) );
  AND2_X1 U12216 ( .A1(n558), .A2(n559), .ZN(n20164) );
  XNOR2_X1 U12364 ( .A(n7012), .B(n7011), .ZN(n20165) );
  XNOR2_X1 U12380 ( .A(n7012), .B(n7011), .ZN(n7833) );
  XNOR2_X1 U12385 ( .A(n6261), .B(n6262), .ZN(n20166) );
  OAI211_X1 U12400 ( .C1(n15325), .C2(n1491), .A(n15324), .B(n15323), .ZN(
        n20167) );
  OAI211_X1 U12455 ( .C1(n15325), .C2(n1491), .A(n15324), .B(n15323), .ZN(
        n17416) );
  XOR2_X1 U12690 ( .A(n15436), .B(n15435), .Z(n20168) );
  NAND2_X1 U12691 ( .A1(n2959), .A2(n16445), .ZN(n20169) );
  NOR2_X1 U12752 ( .A1(n3565), .A2(n12512), .ZN(n13619) );
  XOR2_X1 U12862 ( .A(n13593), .B(n13594), .Z(n20171) );
  XNOR2_X1 U13005 ( .A(n16597), .B(n16598), .ZN(n20172) );
  NAND2_X1 U13267 ( .A1(n13505), .A2(n2138), .ZN(n20173) );
  NAND2_X1 U13268 ( .A1(n13505), .A2(n2138), .ZN(n15457) );
  CLKBUF_X1 U13269 ( .A(n8220), .Z(n20174) );
  XNOR2_X1 U13343 ( .A(n6473), .B(n6472), .ZN(n8220) );
  NOR2_X2 U13458 ( .A1(n7670), .A2(n7669), .ZN(n20176) );
  NOR2_X1 U13544 ( .A1(n7670), .A2(n7669), .ZN(n10200) );
  XNOR2_X1 U13545 ( .A(n6797), .B(n6798), .ZN(n20177) );
  AOI22_X1 U13599 ( .A1(n13975), .A2(n19940), .B1(n13974), .B2(n14499), .ZN(
        n20178) );
  AOI22_X1 U13632 ( .A1(n13975), .A2(n19940), .B1(n13974), .B2(n14499), .ZN(
        n15709) );
  XOR2_X1 U13668 ( .A(n963), .B(n17140), .Z(n20179) );
  XNOR2_X1 U13790 ( .A(n6455), .B(n6454), .ZN(n20180) );
  XNOR2_X1 U13873 ( .A(n13847), .B(n2679), .ZN(n20181) );
  XNOR2_X1 U13900 ( .A(n13847), .B(n2679), .ZN(n14603) );
  NOR2_X1 U13981 ( .A1(n14735), .A2(n14734), .ZN(n20182) );
  NOR2_X1 U14024 ( .A1(n14735), .A2(n14734), .ZN(n20183) );
  AOI22_X2 U14113 ( .A1(n14955), .A2(n15043), .B1(n15802), .B2(n14954), .ZN(
        n16711) );
  XNOR2_X1 U14196 ( .A(n16092), .B(n16093), .ZN(n20185) );
  INV_X1 U14197 ( .A(n12312), .ZN(n20186) );
  AND2_X1 U14402 ( .A1(n14573), .A2(n14572), .ZN(n20187) );
  INV_X1 U14403 ( .A(n19877), .ZN(n20188) );
  INV_X1 U14462 ( .A(n20235), .ZN(n11404) );
  XNOR2_X1 U14587 ( .A(n7359), .B(n7358), .ZN(n20189) );
  INV_X1 U14646 ( .A(n10601), .ZN(n20324) );
  XNOR2_X1 U14686 ( .A(n3908), .B(Key[156]), .ZN(n20190) );
  AOI22_X1 U14725 ( .A1(n11242), .A2(n11349), .B1(n11241), .B2(n11350), .ZN(
        n12021) );
  NOR2_X1 U14745 ( .A1(n15718), .A2(n73), .ZN(n20192) );
  CLKBUF_X1 U14746 ( .A(n19237), .Z(n20193) );
  NOR2_X1 U14824 ( .A1(n15718), .A2(n73), .ZN(n16027) );
  OAI21_X1 U15015 ( .B1(n17902), .B2(n17901), .A(n17900), .ZN(n19237) );
  XOR2_X1 U15022 ( .A(n16920), .B(n16919), .Z(n20194) );
  XNOR2_X1 U15059 ( .A(n6223), .B(n6224), .ZN(n20195) );
  OAI22_X1 U15154 ( .A1(n19519), .A2(n9579), .B1(n8577), .B2(n19715), .ZN(
        n20196) );
  XNOR2_X1 U15165 ( .A(n6223), .B(n6224), .ZN(n7935) );
  AND2_X1 U15166 ( .A1(n1640), .A2(n15310), .ZN(n15397) );
  XNOR2_X1 U15361 ( .A(n6079), .B(n6078), .ZN(n20198) );
  OAI211_X1 U15362 ( .C1(n12570), .C2(n13146), .A(n12019), .B(n12018), .ZN(
        n20199) );
  XNOR2_X1 U15363 ( .A(n6079), .B(n6078), .ZN(n8055) );
  OAI211_X1 U15385 ( .C1(n12570), .C2(n13146), .A(n12019), .B(n12018), .ZN(
        n13059) );
  XNOR2_X1 U15421 ( .A(n6885), .B(n6884), .ZN(n20200) );
  OAI22_X1 U15440 ( .A1(n11673), .A2(n12179), .B1(n11650), .B2(n11670), .ZN(
        n20201) );
  XNOR2_X1 U15479 ( .A(Key[108]), .B(Plaintext[108]), .ZN(n20202) );
  XNOR2_X1 U15500 ( .A(n13692), .B(n13691), .ZN(n20204) );
  XNOR2_X1 U15501 ( .A(n13692), .B(n13691), .ZN(n14378) );
  INV_X1 U15534 ( .A(n4136), .ZN(n20205) );
  XOR2_X1 U15535 ( .A(n13061), .B(n13062), .Z(n20206) );
  XNOR2_X1 U15536 ( .A(n16995), .B(n16994), .ZN(n20207) );
  XNOR2_X1 U15562 ( .A(n5321), .B(n7134), .ZN(n20208) );
  XNOR2_X1 U15583 ( .A(n6819), .B(n7218), .ZN(n20209) );
  INV_X1 U15584 ( .A(n912), .ZN(n20330) );
  OAI211_X1 U15772 ( .C1(n8784), .C2(n8783), .A(n3807), .B(n8782), .ZN(n20210)
         );
  OAI211_X1 U15813 ( .C1(n8784), .C2(n8783), .A(n3807), .B(n8782), .ZN(n20211)
         );
  OR2_X1 U15817 ( .A1(n8780), .A2(n9107), .ZN(n3807) );
  XNOR2_X1 U15842 ( .A(n16526), .B(n16525), .ZN(n20212) );
  XNOR2_X1 U15872 ( .A(n16526), .B(n16525), .ZN(n19362) );
  OR2_X1 U16014 ( .A1(n5941), .A2(n20243), .ZN(n8295) );
  XOR2_X1 U16031 ( .A(n13663), .B(n13662), .Z(n20213) );
  XNOR2_X2 U16085 ( .A(n2772), .B(n2771), .ZN(n10980) );
  AND4_X1 U16154 ( .A1(n17192), .A2(n17191), .A3(n17190), .A4(n17189), .ZN(
        n20214) );
  INV_X1 U16158 ( .A(n8103), .ZN(n9326) );
  OAI211_X1 U16244 ( .C1(n4404), .C2(n5856), .A(n4403), .B(n4402), .ZN(n20216)
         );
  OAI211_X1 U16246 ( .C1(n4404), .C2(n5856), .A(n4403), .B(n4402), .ZN(n2571)
         );
  XOR2_X1 U16312 ( .A(n16060), .B(n16061), .Z(n20217) );
  AOI22_X1 U16315 ( .A1(n17614), .A2(n17613), .B1(n17612), .B2(n17611), .ZN(
        n20218) );
  XNOR2_X1 U16316 ( .A(n17355), .B(n16181), .ZN(n20219) );
  XNOR2_X1 U16389 ( .A(n16774), .B(n16773), .ZN(n18956) );
  NAND2_X1 U16404 ( .A1(n11963), .A2(n3396), .ZN(n20222) );
  NAND2_X1 U16419 ( .A1(n11963), .A2(n3396), .ZN(n20223) );
  OAI211_X1 U16496 ( .C1(n262), .C2(n9328), .A(n1408), .B(n20313), .ZN(n2173)
         );
  NAND4_X1 U16499 ( .A1(n5738), .A2(n5740), .A3(n5737), .A4(n5739), .ZN(n20224) );
  NAND4_X1 U16598 ( .A1(n5738), .A2(n5740), .A3(n5737), .A4(n5739), .ZN(n20225) );
  NAND4_X1 U16600 ( .A1(n5738), .A2(n5740), .A3(n5737), .A4(n5739), .ZN(n6767)
         );
  OAI211_X1 U16620 ( .C1(n5823), .C2(n5448), .A(n3567), .B(n3568), .ZN(n20227)
         );
  XOR2_X1 U16663 ( .A(n9799), .B(n9462), .Z(n20228) );
  OAI211_X1 U16702 ( .C1(n5823), .C2(n5448), .A(n3567), .B(n3568), .ZN(n7121)
         );
  XNOR2_X1 U16718 ( .A(Key[140]), .B(Plaintext[140]), .ZN(n20229) );
  XNOR2_X1 U16727 ( .A(n10584), .B(n20491), .ZN(n10218) );
  XNOR2_X1 U16742 ( .A(Key[140]), .B(Plaintext[140]), .ZN(n5017) );
  XOR2_X1 U16743 ( .A(n15250), .B(n15968), .Z(n20230) );
  NOR2_X1 U16751 ( .A1(n16464), .A2(n2297), .ZN(n20231) );
  NOR2_X1 U16761 ( .A1(n16464), .A2(n2297), .ZN(n20232) );
  NOR2_X1 U16783 ( .A1(n16464), .A2(n2297), .ZN(n18454) );
  XNOR2_X1 U16803 ( .A(n10065), .B(n10064), .ZN(n20233) );
  XNOR2_X1 U16865 ( .A(n10065), .B(n10064), .ZN(n10897) );
  OR2_X1 U16870 ( .A1(n16632), .A2(n17513), .ZN(n20234) );
  OAI211_X2 U16909 ( .C1(n15105), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n16695) );
  XNOR2_X2 U16953 ( .A(n20236), .B(n9575), .ZN(n20235) );
  XOR2_X1 U16993 ( .A(n9692), .B(n9573), .Z(n20236) );
  XOR2_X1 U17032 ( .A(n12906), .B(n13848), .Z(n20237) );
  XNOR2_X1 U17203 ( .A(n15937), .B(n15938), .ZN(n20239) );
  XNOR2_X1 U17204 ( .A(n15937), .B(n15938), .ZN(n17172) );
  NAND4_X1 U17292 ( .A1(n17192), .A2(n17191), .A3(n17190), .A4(n17189), .ZN(
        n19115) );
  XNOR2_X1 U17339 ( .A(n15764), .B(n15763), .ZN(n19354) );
  BUF_X1 U17354 ( .A(n5563), .Z(n20241) );
  XNOR2_X1 U17424 ( .A(n16532), .B(n16531), .ZN(n20242) );
  XOR2_X1 U17433 ( .A(n5962), .B(n5961), .Z(n20243) );
  NAND2_X2 U17571 ( .A1(n2591), .A2(n14345), .ZN(n15906) );
  XNOR2_X1 U17575 ( .A(n4065), .B(n4064), .ZN(n20247) );
  XNOR2_X1 U17605 ( .A(n20248), .B(n20249), .ZN(n14410) );
  XNOR2_X1 U17658 ( .A(n13388), .B(n13389), .ZN(n20248) );
  XOR2_X1 U17743 ( .A(n13393), .B(n13392), .Z(n20249) );
  NOR2_X2 U17754 ( .A1(n9084), .A2(n9083), .ZN(n9986) );
  BUF_X1 U17863 ( .A(n6919), .Z(n20250) );
  XOR2_X1 U17938 ( .A(n1074), .B(n1073), .Z(n20251) );
  XNOR2_X1 U17977 ( .A(n6741), .B(n6740), .ZN(n20252) );
  OAI211_X1 U17978 ( .C1(n874), .C2(n12622), .A(n12621), .B(n12620), .ZN(
        n20253) );
  XNOR2_X1 U18011 ( .A(n6741), .B(n6740), .ZN(n8376) );
  OAI211_X1 U18034 ( .C1(n874), .C2(n12622), .A(n12621), .B(n12620), .ZN(
        n13585) );
  OAI21_X1 U18132 ( .B1(n11483), .B2(n11215), .A(n11214), .ZN(n12479) );
  XNOR2_X1 U18140 ( .A(n2738), .B(Key[79]), .ZN(n5112) );
  XNOR2_X1 U18172 ( .A(n5940), .B(n5939), .ZN(n20257) );
  XOR2_X1 U18173 ( .A(n17274), .B(n17273), .Z(n20258) );
  BUF_X1 U18174 ( .A(n18866), .Z(n20259) );
  OAI21_X1 U18175 ( .B1(n19575), .B2(n18040), .A(n18039), .ZN(n18866) );
  OAI21_X1 U18182 ( .B1(n11983), .B2(n12619), .A(n11982), .ZN(n20260) );
  INV_X1 U18186 ( .A(n19598), .ZN(n20261) );
  INV_X1 U18236 ( .A(n8370), .ZN(n20294) );
  XNOR2_X1 U18238 ( .A(n12903), .B(n12904), .ZN(n20262) );
  XNOR2_X1 U18259 ( .A(n12903), .B(n12904), .ZN(n701) );
  NOR2_X1 U18333 ( .A1(n19068), .A2(n18151), .ZN(n19079) );
  XOR2_X1 U18334 ( .A(n13532), .B(n13531), .Z(n20263) );
  XNOR2_X1 U18384 ( .A(n16121), .B(n16120), .ZN(n20264) );
  AND3_X2 U18430 ( .A1(n3428), .A2(n3432), .A3(n3426), .ZN(n16980) );
  OAI21_X1 U18458 ( .B1(n1244), .B2(n1243), .A(n1242), .ZN(n20265) );
  OAI21_X1 U18483 ( .B1(n1244), .B2(n1243), .A(n1242), .ZN(n8990) );
  XNOR2_X1 U18498 ( .A(n10219), .B(n19818), .ZN(n20268) );
  XNOR2_X1 U18506 ( .A(n16406), .B(n16027), .ZN(n20269) );
  XNOR2_X1 U18543 ( .A(n7280), .B(n7281), .ZN(n20270) );
  XNOR2_X1 U18544 ( .A(n6524), .B(n20314), .ZN(n8083) );
  XNOR2_X1 U18661 ( .A(n14017), .B(n14018), .ZN(n20271) );
  XOR2_X1 U18682 ( .A(n13069), .B(n13068), .Z(n20272) );
  XOR2_X1 U18691 ( .A(n15854), .B(n15855), .Z(n20273) );
  XOR2_X1 U18699 ( .A(n6930), .B(n6929), .Z(n20274) );
  XNOR2_X1 U18700 ( .A(n15969), .B(n15968), .ZN(n20275) );
  OAI21_X1 U18720 ( .B1(n17385), .B2(n17384), .A(n17383), .ZN(n18831) );
  OAI211_X2 U18793 ( .C1(n3118), .C2(n8341), .A(n3119), .B(n20277), .ZN(n9563)
         );
  NAND2_X1 U18794 ( .A1(n3122), .A2(n3121), .ZN(n20277) );
  NAND2_X1 U18896 ( .A1(n7685), .A2(n8381), .ZN(n7716) );
  NAND2_X1 U18897 ( .A1(n19561), .A2(n4080), .ZN(n5707) );
  AOI22_X2 U18912 ( .A1(n15169), .A2(n15168), .B1(n15378), .B2(n15170), .ZN(
        n16615) );
  NAND2_X1 U18922 ( .A1(n20279), .A2(n20278), .ZN(n10758) );
  NAND2_X1 U18923 ( .A1(n11526), .A2(n11521), .ZN(n20278) );
  XNOR2_X1 U18946 ( .A(n20123), .B(n12769), .ZN(n13698) );
  NAND3_X1 U18960 ( .A1(n12227), .A2(n10941), .A3(n12229), .ZN(n10942) );
  NAND2_X2 U19319 ( .A1(n20281), .A2(n738), .ZN(n9576) );
  NAND2_X1 U19359 ( .A1(n7512), .A2(n7511), .ZN(n20281) );
  NAND2_X1 U19489 ( .A1(n7852), .A2(n8159), .ZN(n2840) );
  NAND2_X1 U19545 ( .A1(n1865), .A2(n1868), .ZN(n2630) );
  NAND2_X1 U19579 ( .A1(n5001), .A2(n20282), .ZN(n7088) );
  NAND3_X1 U19580 ( .A1(n5770), .A2(n5545), .A3(n5734), .ZN(n5740) );
  NAND2_X1 U19581 ( .A1(n15473), .A2(n15767), .ZN(n15478) );
  NAND3_X1 U19585 ( .A1(n5147), .A2(n5146), .A3(n5572), .ZN(n5152) );
  XNOR2_X1 U19629 ( .A(n13465), .B(n13464), .ZN(n20285) );
  NAND2_X1 U19632 ( .A1(n4515), .A2(n4514), .ZN(n5767) );
  NAND3_X1 U19638 ( .A1(n338), .A2(n1383), .A3(n12663), .ZN(n16347) );
  NAND3_X1 U19693 ( .A1(n1478), .A2(n1477), .A3(n9361), .ZN(n8964) );
  OR2_X1 U19705 ( .A1(n15657), .A2(n12658), .ZN(n12659) );
  OAI21_X2 U19706 ( .B1(n488), .B2(n11657), .A(n487), .ZN(n13134) );
  NAND2_X1 U19707 ( .A1(n19112), .A2(n19105), .ZN(n20286) );
  NAND3_X1 U19718 ( .A1(n7813), .A2(n7814), .A3(n7479), .ZN(n465) );
  NAND2_X1 U19731 ( .A1(n15275), .A2(n15270), .ZN(n15272) );
  NAND2_X1 U19749 ( .A1(n14935), .A2(n20288), .ZN(n1613) );
  INV_X1 U19751 ( .A(n13615), .ZN(n14597) );
  NAND2_X1 U19752 ( .A1(n19647), .A2(n19372), .ZN(n19646) );
  NAND2_X1 U19753 ( .A1(n18216), .A2(n1194), .ZN(n1193) );
  NAND2_X1 U19754 ( .A1(n20005), .A2(n15702), .ZN(n15141) );
  XNOR2_X1 U19755 ( .A(n20290), .B(n19322), .ZN(Ciphertext[175]) );
  NAND3_X1 U19756 ( .A1(n19319), .A2(n19320), .A3(n19318), .ZN(n20290) );
  OAI22_X1 U19757 ( .A1(n19514), .A2(n13989), .B1(n15714), .B2(n15148), .ZN(
        n13990) );
  NOR2_X1 U19758 ( .A1(n16170), .A2(n20291), .ZN(n16632) );
  NOR2_X1 U19759 ( .A1(n14845), .A2(n16633), .ZN(n20291) );
  NAND2_X1 U19760 ( .A1(n7726), .A2(n7856), .ZN(n20292) );
  OAI211_X1 U19761 ( .C1(n8376), .C2(n19881), .A(n20295), .B(n20294), .ZN(
        n20293) );
  NAND2_X1 U19762 ( .A1(n8373), .A2(n19881), .ZN(n20295) );
  INV_X1 U19763 ( .A(n4926), .ZN(n4385) );
  NAND2_X1 U19764 ( .A1(n3967), .A2(n4921), .ZN(n4926) );
  NAND2_X1 U19765 ( .A1(n20298), .A2(n20297), .ZN(n12313) );
  NAND2_X1 U19766 ( .A1(n11362), .A2(n11361), .ZN(n20298) );
  NAND2_X1 U19768 ( .A1(n10768), .A2(n11104), .ZN(n20299) );
  NAND2_X1 U19770 ( .A1(n3862), .A2(n3861), .ZN(n20301) );
  XNOR2_X1 U19771 ( .A(n20302), .B(n16599), .ZN(n16385) );
  XNOR2_X1 U19772 ( .A(n19782), .B(n2329), .ZN(n20302) );
  NAND2_X1 U19773 ( .A1(n20305), .A2(n20303), .ZN(n12486) );
  NAND2_X1 U19774 ( .A1(n12476), .A2(n20304), .ZN(n20303) );
  INV_X1 U19775 ( .A(n19833), .ZN(n20304) );
  NAND2_X1 U19776 ( .A1(n12475), .A2(n19833), .ZN(n20305) );
  NAND2_X1 U19778 ( .A1(n689), .A2(n18946), .ZN(n20306) );
  OAI211_X1 U19779 ( .C1(n8672), .C2(n8674), .A(n20309), .B(n20308), .ZN(n8519) );
  NAND2_X1 U19780 ( .A1(n19857), .A2(n9023), .ZN(n20308) );
  NAND2_X1 U19781 ( .A1(n9022), .A2(n8672), .ZN(n20309) );
  OAI21_X1 U19782 ( .B1(n14260), .B2(n20311), .A(n20310), .ZN(n14019) );
  NAND2_X1 U19783 ( .A1(n14260), .A2(n13981), .ZN(n20310) );
  NAND2_X1 U19784 ( .A1(n2889), .A2(n14702), .ZN(n15370) );
  NAND2_X1 U19785 ( .A1(n2890), .A2(n14230), .ZN(n2889) );
  OR2_X2 U19786 ( .A1(n3957), .A2(n20312), .ZN(n3959) );
  NOR2_X1 U19787 ( .A1(n3956), .A2(n4291), .ZN(n20312) );
  NAND2_X1 U19788 ( .A1(n7686), .A2(n8385), .ZN(n8131) );
  NAND3_X1 U19789 ( .A1(n2702), .A2(n1006), .A3(n20315), .ZN(n8993) );
  OR3_X1 U19791 ( .A1(n11528), .A2(n11527), .A3(n11521), .ZN(n12221) );
  NAND2_X1 U19792 ( .A1(n19761), .A2(n14396), .ZN(n13615) );
  NAND2_X1 U19793 ( .A1(n20316), .A2(n19421), .ZN(n19423) );
  NAND3_X1 U19795 ( .A1(n20318), .A2(n20317), .A3(n11176), .ZN(n10656) );
  NAND2_X1 U19796 ( .A1(n11178), .A2(n10962), .ZN(n20318) );
  NOR2_X1 U19797 ( .A1(n14637), .A2(n20319), .ZN(n12974) );
  OR2_X1 U19798 ( .A1(n19703), .A2(n14032), .ZN(n20319) );
  NAND2_X1 U19799 ( .A1(n20320), .A2(n210), .ZN(n4896) );
  NAND2_X1 U19800 ( .A1(n3231), .A2(n4136), .ZN(n20320) );
  NAND3_X1 U19801 ( .A1(n8053), .A2(n19474), .A3(n8193), .ZN(n7626) );
  NAND2_X1 U19802 ( .A1(n20322), .A2(n20321), .ZN(n2637) );
  NAND2_X1 U19803 ( .A1(n9241), .A2(n9240), .ZN(n20321) );
  OAI21_X1 U19804 ( .B1(n19606), .B2(n20505), .A(n20323), .ZN(n8543) );
  NAND2_X1 U19805 ( .A1(n20505), .A2(n20476), .ZN(n20323) );
  OAI21_X1 U19808 ( .B1(n19100), .B2(n19101), .A(n20326), .ZN(n19610) );
  AOI22_X1 U19809 ( .A1(n19101), .A2(n19105), .B1(n19112), .B2(n19118), .ZN(
        n20326) );
  INV_X1 U19810 ( .A(n7688), .ZN(n20327) );
  NAND2_X1 U19811 ( .A1(n7685), .A2(n20327), .ZN(n1422) );
  OR3_X1 U19812 ( .A1(n9354), .A2(n8720), .A3(n9528), .ZN(n592) );
  OAI21_X1 U19813 ( .B1(n2685), .B2(n2697), .A(n20328), .ZN(n14047) );
  NAND2_X1 U19814 ( .A1(n19597), .A2(n14827), .ZN(n20328) );
  NOR2_X1 U19815 ( .A1(n5142), .A2(n5143), .ZN(n6494) );
  NAND2_X1 U19816 ( .A1(n14352), .A2(n14326), .ZN(n20329) );
  NAND2_X1 U19817 ( .A1(n3519), .A2(n2883), .ZN(n2882) );
  NAND2_X1 U19818 ( .A1(n2884), .A2(n1401), .ZN(n3519) );
  OAI211_X1 U19820 ( .C1(n17524), .C2(n17519), .A(n17522), .B(n20331), .ZN(
        n17528) );
  INV_X1 U19821 ( .A(n17581), .ZN(n20331) );
  INV_X1 U19822 ( .A(n699), .ZN(n698) );
  NOR2_X1 U19824 ( .A1(n14435), .A2(n14171), .ZN(n14431) );
  NAND2_X1 U19826 ( .A1(n20333), .A2(n20332), .ZN(n4464) );
  NAND2_X1 U19827 ( .A1(n6141), .A2(n5859), .ZN(n20332) );
  AND2_X2 U19829 ( .A1(n20335), .A2(n20337), .ZN(n16335) );
  INV_X1 U19830 ( .A(n20336), .ZN(n20335) );
  OAI21_X1 U19831 ( .B1(n15519), .B2(n3821), .A(n15518), .ZN(n20336) );
  NAND2_X1 U19832 ( .A1(n15522), .A2(n15521), .ZN(n20337) );
  NAND2_X1 U19833 ( .A1(n12490), .A2(n11912), .ZN(n12492) );
  NAND2_X1 U19834 ( .A1(n14090), .A2(n939), .ZN(n15516) );
  OAI22_X1 U19836 ( .A1(n3601), .A2(n11275), .B1(n11271), .B2(n11381), .ZN(
        n20338) );
  OR2_X2 U19837 ( .A1(n4149), .A2(n4150), .ZN(n5643) );
  OAI22_X1 U19838 ( .A1(n15112), .A2(n15113), .B1(n15114), .B2(n15604), .ZN(
        n15118) );
  NAND2_X1 U19839 ( .A1(n20112), .A2(n15275), .ZN(n15113) );
  NAND2_X1 U19841 ( .A1(n15370), .A2(n15371), .ZN(n15565) );
  NAND2_X1 U19842 ( .A1(n75), .A2(n78), .ZN(n20339) );
  AND2_X2 U19843 ( .A1(n1592), .A2(n1189), .ZN(n12208) );
  NAND2_X1 U19844 ( .A1(n19979), .A2(n5914), .ZN(n5915) );
  NAND2_X1 U19846 ( .A1(n10833), .A2(n11037), .ZN(n20340) );
  NAND2_X1 U19847 ( .A1(n15534), .A2(n15921), .ZN(n20341) );
  NAND2_X1 U19848 ( .A1(n20343), .A2(n2974), .ZN(n20342) );
  NAND2_X1 U19849 ( .A1(n15532), .A2(n15531), .ZN(n20343) );
  NAND2_X1 U19850 ( .A1(n20345), .A2(n20344), .ZN(n8669) );
  NAND2_X1 U19851 ( .A1(n9112), .A2(n9114), .ZN(n20344) );
  OAI21_X1 U19852 ( .B1(n1602), .B2(n9217), .A(n20346), .ZN(n20345) );
  AOI21_X2 U19853 ( .B1(n11362), .B2(n11361), .A(n3667), .ZN(n19952) );
  AOI21_X2 U19854 ( .B1(n12329), .B2(n12328), .A(n13269), .ZN(n19796) );
  AOI22_X2 U19855 ( .A1(n1419), .A2(n12293), .B1(n11772), .B2(n12533), .ZN(
        n19697) );
  OAI211_X2 U19857 ( .C1(n12267), .C2(n12565), .A(n976), .B(n1043), .ZN(n13703) );
  NAND2_X2 U6130 ( .A1(n2159), .A2(n1975), .ZN(n13725) );
  MUX2_X2 U1841 ( .A(n6103), .B(n6102), .S(n6101), .Z(n7218) );
  BUF_X2 U720 ( .A(n4268), .Z(n5024) );
  OAI211_X2 U705 ( .C1(n5103), .C2(n1421), .A(n5110), .B(n1420), .ZN(n6010) );
  NOR2_X2 U17999 ( .A1(n14583), .A2(n14582), .ZN(n16750) );
  BUF_X1 U379 ( .A(n5589), .Z(n19979) );
  NAND2_X2 U1860 ( .A1(n3194), .A2(n1745), .ZN(n7248) );
  NOR2_X2 U12692 ( .A1(n3565), .A2(n12512), .ZN(n20170) );
  OR2_X2 U2249 ( .A1(n4164), .A2(n4163), .ZN(n5442) );
  BUF_X1 U2696 ( .A(n15284), .Z(n19848) );
  BUF_X1 U740 ( .A(n14829), .Z(n19984) );
  XNOR2_X2 U62 ( .A(Key[10]), .B(Plaintext[10]), .ZN(n4125) );
  BUF_X2 U820 ( .A(n5031), .Z(n153) );
  OAI22_X2 U772 ( .A1(n3259), .A2(n4694), .B1(n5107), .B2(n4695), .ZN(n6183)
         );
  BUF_X1 U231 ( .A(n3846), .Z(n5116) );
  XNOR2_X2 U658 ( .A(n3945), .B(Key[181]), .ZN(n4313) );
  BUF_X1 U561 ( .A(n14120), .Z(n14703) );
  XNOR2_X2 U440 ( .A(Key[9]), .B(Plaintext[9]), .ZN(n4319) );
  OR2_X2 U1677 ( .A1(n7175), .A2(n7174), .ZN(n9842) );
  NOR2_X2 U852 ( .A1(n11728), .A2(n682), .ZN(n13248) );
  AND3_X2 U2893 ( .A1(n728), .A2(n14546), .A3(n14545), .ZN(n15645) );
  NAND2_X2 U173 ( .A1(n1586), .A2(n4218), .ZN(n6016) );
  AND3_X2 U2318 ( .A1(n1815), .A2(n1816), .A3(n1818), .ZN(n15979) );
  BUF_X2 U957 ( .A(n17831), .Z(n19110) );
  BUF_X1 U371 ( .A(n6404), .Z(n6707) );
  NOR2_X1 U2532 ( .A1(n14278), .A2(n1409), .ZN(n15536) );
  BUF_X2 U689 ( .A(n13316), .Z(n14705) );
  MUX2_X2 U6855 ( .A(n17975), .B(n17974), .S(n17549), .Z(n18688) );
  AND2_X2 U717 ( .A1(n8320), .A2(n8319), .ZN(n8872) );
  NAND2_X2 U166 ( .A1(n15901), .A2(n15902), .ZN(n16283) );
  AND3_X2 U9269 ( .A1(n6212), .A2(n7628), .A3(n6211), .ZN(n8708) );
  BUF_X2 U2909 ( .A(n14849), .Z(n15474) );
  OR2_X2 U1008 ( .A1(n2303), .A2(n7858), .ZN(n9266) );
  AND3_X2 U1680 ( .A1(n16050), .A2(n3147), .A3(n3146), .ZN(n16373) );
  XNOR2_X2 U408 ( .A(n4053), .B(Key[129]), .ZN(n4100) );
  AND2_X2 U1393 ( .A1(n20163), .A2(n20164), .ZN(n19227) );
  BUF_X2 U168 ( .A(n13563), .Z(n15121) );
  BUF_X1 U1281 ( .A(n13227), .Z(n20226) );
  NAND3_X2 U8331 ( .A1(n1877), .A2(n1997), .A3(n1998), .ZN(n17335) );
  XNOR2_X2 U1835 ( .A(n10135), .B(n10136), .ZN(n11349) );
  OR2_X2 U207 ( .A1(n8128), .A2(n6438), .ZN(n8129) );
  NAND2_X2 U568 ( .A1(n2635), .A2(n7452), .ZN(n8672) );
  BUF_X1 U310 ( .A(n10882), .Z(n11569) );
  BUF_X2 U1097 ( .A(n17374), .Z(n18262) );
  XNOR2_X2 U687 ( .A(Key[116]), .B(Plaintext[116]), .ZN(n5046) );
  NAND3_X2 U3679 ( .A1(n3598), .A2(n3453), .A3(n4451), .ZN(n5859) );
  NAND3_X2 U2314 ( .A1(n1455), .A2(n1454), .A3(n6001), .ZN(n6982) );
  OAI22_X2 U1678 ( .A1(n8336), .A2(n8335), .B1(n8334), .B2(n8333), .ZN(n9648)
         );
  OR2_X2 U501 ( .A1(n15426), .A2(n14243), .ZN(n15421) );
  BUF_X1 U18376 ( .A(n16690), .Z(n19820) );
  OAI21_X2 U18733 ( .B1(n18102), .B2(n18101), .A(n18100), .ZN(n18651) );
  NAND2_X2 U4237 ( .A1(n2789), .A2(n3275), .ZN(n15546) );
  OAI22_X2 U6938 ( .A1(n2973), .A2(n15553), .B1(n15552), .B2(n15551), .ZN(
        n17359) );
  XNOR2_X2 U2720 ( .A(n16848), .B(n16849), .ZN(n18269) );
  AND3_X2 U877 ( .A1(n715), .A2(n2380), .A3(n714), .ZN(n17438) );
  OR2_X2 U2955 ( .A1(n7987), .A2(n7986), .ZN(n9166) );
  NAND2_X2 U6265 ( .A1(n8120), .A2(n900), .ZN(n9331) );
  XNOR2_X2 U1461 ( .A(n11852), .B(n11851), .ZN(n15313) );
  AND2_X2 U6898 ( .A1(n3248), .A2(n18254), .ZN(n18774) );
  BUF_X1 U1839 ( .A(n7133), .Z(n899) );
  MUX2_X2 U9825 ( .A(n5263), .B(n5262), .S(n5691), .Z(n6520) );
  BUF_X1 U225 ( .A(n15777), .Z(n19977) );
  INV_X1 U368 ( .A(n13937), .ZN(n14419) );
  XNOR2_X2 U13323 ( .A(n10292), .B(n10293), .ZN(n11257) );
  AOI22_X2 U387 ( .A1(n15367), .A2(n15366), .B1(n15369), .B2(n15368), .ZN(
        n17127) );
  NAND2_X2 U5587 ( .A1(n780), .A2(n19574), .ZN(n18795) );
  OAI21_X2 U1568 ( .B1(n11355), .B2(n11354), .A(n11353), .ZN(n3260) );
  AND3_X2 U1499 ( .A1(n3464), .A2(n1008), .A3(n11758), .ZN(n13717) );
  BUF_X2 U746 ( .A(n5782), .Z(n6055) );
  NAND2_X2 U18737 ( .A1(n18110), .A2(n18109), .ZN(n18648) );
  OAI21_X2 U19 ( .B1(n4159), .B2(n4158), .A(n4157), .ZN(n5641) );
  OR2_X2 U410 ( .A1(n623), .A2(n3833), .ZN(n3855) );
  XNOR2_X2 U7843 ( .A(n7085), .B(n7084), .ZN(n8014) );
  BUF_X1 U13645 ( .A(n19092), .Z(n19112) );
  XNOR2_X2 U885 ( .A(n10386), .B(n10385), .ZN(n11131) );
  BUF_X1 U19679 ( .A(n17300), .Z(n19929) );
  NAND3_X2 U679 ( .A1(n5306), .A2(n5307), .A3(n5305), .ZN(n6687) );
  MUX2_X2 U15436 ( .A(n13461), .B(n13460), .S(n15666), .Z(n17291) );
  BUF_X2 U653 ( .A(n9009), .Z(n19490) );
  BUF_X1 U447 ( .A(n5264), .Z(n6139) );
  XNOR2_X2 U1108 ( .A(n17292), .B(n3207), .ZN(n18240) );
  AOI22_X2 U6588 ( .A1(n2680), .A2(n10895), .B1(n10893), .B2(n10894), .ZN(
        n12600) );
  NOR2_X2 U11987 ( .A1(n8491), .A2(n8490), .ZN(n10442) );
  CLKBUF_X3 U51 ( .A(n6871), .Z(n8272) );
  XNOR2_X2 U622 ( .A(n7947), .B(n7946), .ZN(n11161) );
  OAI21_X2 U15269 ( .B1(n15311), .B2(n14992), .A(n14991), .ZN(n16227) );
  AND2_X2 U1849 ( .A1(n1323), .A2(n1322), .ZN(n9799) );
  NAND2_X2 U2655 ( .A1(n579), .A2(n14835), .ZN(n17295) );
  OAI211_X2 U12023 ( .C1(n14813), .C2(n2808), .A(n14592), .B(n14591), .ZN(
        n15601) );
  AOI21_X2 U7950 ( .B1(n14521), .B2(n13565), .A(n13564), .ZN(n15052) );
  BUF_X1 U232 ( .A(n15777), .Z(n19978) );
  NAND3_X2 U1740 ( .A1(n4798), .A2(n2699), .A3(n19544), .ZN(n5990) );
  NAND4_X2 U284 ( .A1(n14141), .A2(n14140), .A3(n3006), .A4(n3005), .ZN(n15510) );
  XNOR2_X1 U1075 ( .A(n12995), .B(n12994), .ZN(n951) );
  NOR2_X2 U4800 ( .A1(n8082), .A2(n8081), .ZN(n8866) );
  AND3_X2 U24 ( .A1(n12613), .A2(n12612), .A3(n12611), .ZN(n13518) );
  BUF_X1 U240 ( .A(n6381), .Z(n19475) );
  NAND2_X2 U1856 ( .A1(n5702), .A2(n5701), .ZN(n7332) );
  XNOR2_X2 U6385 ( .A(n16826), .B(n16827), .ZN(n18033) );
  NAND2_X2 U9565 ( .A1(n350), .A2(n349), .ZN(n16330) );
  OR2_X2 U6697 ( .A1(n8463), .A2(n8462), .ZN(n9329) );
  INV_X1 U11377 ( .A(n7453), .ZN(n8297) );
  NAND3_X2 U1064 ( .A1(n1824), .A2(n14606), .A3(n14607), .ZN(n15274) );
  AND2_X1 U1397 ( .A1(n15311), .A2(n360), .ZN(n15399) );
  MUX2_X2 U5362 ( .A(n15027), .B(n15026), .S(n16629), .Z(n18425) );
  BUF_X2 U889 ( .A(n14347), .Z(n19496) );
  XNOR2_X2 U11912 ( .A(n8397), .B(n8398), .ZN(n11159) );
  OAI21_X2 U868 ( .B1(n1554), .B2(n15561), .A(n1553), .ZN(n17407) );
  NAND2_X2 U526 ( .A1(n11780), .A2(n11779), .ZN(n13601) );
  XNOR2_X2 U287 ( .A(n10278), .B(n10277), .ZN(n11253) );
  BUF_X1 U8146 ( .A(n18151), .Z(n19060) );
  XNOR2_X2 U1824 ( .A(n7001), .B(n7000), .ZN(n7974) );
  BUF_X2 U1052 ( .A(n16447), .Z(n17155) );
  BUF_X1 U1795 ( .A(n7571), .Z(n8151) );
  BUF_X2 U463 ( .A(n6578), .Z(n8239) );
  AOI21_X2 U1307 ( .B1(n16726), .B2(n20127), .A(n16725), .ZN(n870) );
  BUF_X1 U17460 ( .A(n16673), .Z(n20244) );
  CLKBUF_X1 U1192 ( .A(Key[144]), .Z(n456) );
  XNOR2_X1 U828 ( .A(Key[121]), .B(Plaintext[121]), .ZN(n4769) );
  CLKBUF_X1 U1223 ( .A(Key[82]), .Z(n2023) );
  XNOR2_X1 U8741 ( .A(Key[20]), .B(Plaintext[20]), .ZN(n4928) );
  XNOR2_X1 U8912 ( .A(Key[43]), .B(Plaintext[43]), .ZN(n4968) );
  XNOR2_X1 U8918 ( .A(Key[46]), .B(Plaintext[46]), .ZN(n4965) );
  XNOR2_X1 U921 ( .A(Key[14]), .B(Plaintext[14]), .ZN(n4306) );
  CLKBUF_X1 U1376 ( .A(Key[69]), .Z(n17544) );
  CLKBUF_X1 U1370 ( .A(Key[103]), .Z(n17535) );
  XNOR2_X1 U101 ( .A(Key[154]), .B(Plaintext[154]), .ZN(n4756) );
  CLKBUF_X1 U1371 ( .A(Key[30]), .Z(n2349) );
  CLKBUF_X1 U1357 ( .A(Key[167]), .Z(n17095) );
  CLKBUF_X1 U1355 ( .A(Key[88]), .Z(n20064) );
  XNOR2_X1 U971 ( .A(Key[118]), .B(Plaintext[118]), .ZN(n5045) );
  BUF_X1 U605 ( .A(n4638), .Z(n19524) );
  XNOR2_X1 U8871 ( .A(n3939), .B(Key[178]), .ZN(n4185) );
  BUF_X1 U322 ( .A(n4056), .Z(n5058) );
  BUF_X1 U8499 ( .A(n4100), .Z(n5060) );
  AND2_X1 U1717 ( .A1(n1390), .A2(n1389), .ZN(n3351) );
  AND2_X1 U445 ( .A1(n3891), .A2(n3890), .ZN(n5300) );
  OR2_X1 U1925 ( .A1(n4374), .A2(n4373), .ZN(n5715) );
  AND2_X1 U433 ( .A1(n614), .A2(n4639), .ZN(n5743) );
  OR2_X1 U1138 ( .A1(n3976), .A2(n3975), .ZN(n6072) );
  OR2_X1 U6578 ( .A1(n4448), .A2(n4447), .ZN(n5860) );
  NAND2_X1 U1934 ( .A1(n3853), .A2(n306), .ZN(n6057) );
  MUX2_X1 U9650 ( .A(n5008), .B(n5007), .S(n5006), .Z(n5009) );
  AND2_X1 U1924 ( .A1(n5051), .A2(n5050), .ZN(n5926) );
  NAND2_X1 U9643 ( .A1(n2480), .A2(n3641), .ZN(n5226) );
  OR2_X1 U438 ( .A1(n4074), .A2(n4075), .ZN(n5434) );
  AND3_X1 U1929 ( .A1(n4024), .A2(n4023), .A3(n4022), .ZN(n5251) );
  NAND2_X1 U9134 ( .A1(n4155), .A2(n4154), .ZN(n5443) );
  AND2_X1 U479 ( .A1(n4991), .A2(n4990), .ZN(n5562) );
  NAND2_X1 U683 ( .A1(n3399), .A2(n964), .ZN(n5279) );
  NAND2_X1 U682 ( .A1(n2739), .A2(n5015), .ZN(n5328) );
  AND2_X1 U1920 ( .A1(n4774), .A2(n4773), .ZN(n6107) );
  OR2_X1 U1899 ( .A1(n4934), .A2(n4933), .ZN(n5683) );
  NAND2_X1 U861 ( .A1(n1942), .A2(n4906), .ZN(n5684) );
  NAND2_X1 U19769 ( .A1(n20301), .A2(n20017), .ZN(n6059) );
  NAND3_X1 U357 ( .A1(n4014), .A2(n1534), .A3(n1533), .ZN(n5393) );
  OAI211_X1 U9056 ( .C1(n4712), .C2(n4783), .A(n4070), .B(n4069), .ZN(n5997)
         );
  AND2_X1 U9781 ( .A1(n5220), .A2(n5219), .ZN(n5945) );
  BUF_X1 U910 ( .A(n6167), .Z(n170) );
  BUF_X1 U9672 ( .A(n5914), .Z(n5916) );
  AND2_X1 U8273 ( .A1(n3684), .A2(n4386), .ZN(n6150) );
  NAND2_X1 U2436 ( .A1(n4068), .A2(n4067), .ZN(n5998) );
  NAND2_X1 U218 ( .A1(n1768), .A2(n1769), .ZN(n3569) );
  BUF_X1 U1986 ( .A(n5304), .Z(n5891) );
  INV_X1 U1882 ( .A(n5622), .ZN(n5621) );
  MUX2_X1 U10105 ( .A(n5672), .B(n5671), .S(n5670), .Z(n5679) );
  OAI211_X1 U261 ( .C1(n6014), .C2(n6013), .A(n6012), .B(n6011), .ZN(n6990) );
  NAND3_X1 U2196 ( .A1(n5066), .A2(n5065), .A3(n20036), .ZN(n7373) );
  OR2_X1 U6935 ( .A1(n5198), .A2(n5197), .ZN(n6641) );
  AOI22_X1 U19710 ( .A1(n6160), .A2(n5614), .B1(n5613), .B2(n5612), .ZN(n7297)
         );
  NAND2_X1 U1998 ( .A1(n1435), .A2(n1170), .ZN(n7196) );
  NAND3_X1 U5200 ( .A1(n1871), .A2(n1870), .A3(n5451), .ZN(n7289) );
  NAND3_X1 U1863 ( .A1(n2639), .A2(n6053), .A3(n2638), .ZN(n7018) );
  OAI21_X1 U727 ( .B1(n4779), .B2(n5640), .A(n4778), .ZN(n7336) );
  OAI211_X1 U1868 ( .C1(n5462), .C2(n1867), .A(n5461), .B(n5460), .ZN(n7160)
         );
  OR2_X1 U1343 ( .A1(n5195), .A2(n5194), .ZN(n6776) );
  XNOR2_X1 U10304 ( .A(n7116), .B(n7354), .ZN(n6718) );
  NAND2_X1 U1843 ( .A1(n5482), .A2(n5481), .ZN(n7306) );
  AOI21_X1 U4673 ( .B1(n5183), .B2(n5182), .A(n5181), .ZN(n7273) );
  XNOR2_X1 U6805 ( .A(n5134), .B(n5133), .ZN(n8184) );
  XNOR2_X1 U854 ( .A(n6332), .B(n6331), .ZN(n7739) );
  XNOR2_X1 U791 ( .A(n7037), .B(n7038), .ZN(n7958) );
  XNOR2_X1 U7402 ( .A(n2825), .B(n2824), .ZN(n8370) );
  XNOR2_X1 U9506 ( .A(n4728), .B(n4729), .ZN(n8190) );
  BUF_X1 U1792 ( .A(n6837), .Z(n7852) );
  INV_X1 U11473 ( .A(n7542), .ZN(n8372) );
  BUF_X1 U663 ( .A(n7684), .Z(n8381) );
  XNOR2_X1 U2104 ( .A(n5491), .B(n5490), .ZN(n8034) );
  XNOR2_X1 U504 ( .A(n6357), .B(n6356), .ZN(n7500) );
  CLKBUF_X1 U50 ( .A(n7481), .Z(n7949) );
  BUF_X1 U1782 ( .A(n7493), .Z(n7679) );
  BUF_X1 U773 ( .A(n7487), .Z(n7968) );
  XNOR2_X1 U898 ( .A(n5377), .B(n5376), .ZN(n7445) );
  BUF_X1 U18094 ( .A(n7621), .Z(n8069) );
  OAI211_X1 U540 ( .C1(n2875), .C2(n7893), .A(n7892), .B(n7607), .ZN(n8729) );
  OAI211_X1 U89 ( .C1(n1411), .C2(n1010), .A(n7617), .B(n1410), .ZN(n8743) );
  OAI22_X1 U2559 ( .A1(n7468), .A2(n8289), .B1(n8024), .B2(n8292), .ZN(n8294)
         );
  OAI211_X1 U8530 ( .C1(n7835), .C2(n7773), .A(n7772), .B(n7771), .ZN(n8997)
         );
  NOR2_X1 U916 ( .A1(n6909), .A2(n6910), .ZN(n8611) );
  NAND2_X1 U1739 ( .A1(n6901), .A2(n6902), .ZN(n9158) );
  OAI211_X1 U451 ( .C1(n8050), .C2(n8309), .A(n8049), .B(n8048), .ZN(n9066) );
  INV_X1 U6587 ( .A(n8542), .ZN(n9836) );
  BUF_X1 U234 ( .A(n8748), .Z(n8931) );
  OAI21_X1 U100 ( .B1(n7784), .B2(n7783), .A(n7782), .ZN(n9177) );
  AND3_X1 U46 ( .A1(n2251), .A2(n2252), .A3(n1784), .ZN(n9149) );
  NAND2_X1 U441 ( .A1(n8275), .A2(n8274), .ZN(n9129) );
  NAND3_X1 U1111 ( .A1(n2190), .A2(n2191), .A3(n6586), .ZN(n6587) );
  AND2_X1 U280 ( .A1(n7437), .A2(n2986), .ZN(n9296) );
  AND2_X1 U1704 ( .A1(n1657), .A2(n7810), .ZN(n9006) );
  BUF_X1 U1718 ( .A(n8500), .Z(n9361) );
  NAND3_X1 U435 ( .A1(n7419), .A2(n429), .A3(n428), .ZN(n9300) );
  NOR2_X1 U908 ( .A1(n7545), .A2(n7546), .ZN(n8959) );
  BUF_X1 U12626 ( .A(n5556), .Z(n19716) );
  NAND2_X1 U1903 ( .A1(n7706), .A2(n20293), .ZN(n8974) );
  AND2_X1 U453 ( .A1(n7734), .A2(n7735), .ZN(n9249) );
  NAND2_X1 U5590 ( .A1(n1158), .A2(n1160), .ZN(n7866) );
  NAND2_X1 U5242 ( .A1(n1422), .A2(n1839), .ZN(n9528) );
  AND2_X1 U1700 ( .A1(n9137), .A2(n8445), .ZN(n9134) );
  OR2_X1 U449 ( .A1(n8698), .A2(n9163), .ZN(n8613) );
  MUX2_X1 U378 ( .A(n7842), .B(n7841), .S(n8623), .Z(n9420) );
  AND2_X1 U315 ( .A1(n19596), .A2(n19595), .ZN(n9862) );
  OAI211_X1 U413 ( .C1(n8947), .C2(n7613), .A(n7612), .B(n7611), .ZN(n10054)
         );
  NAND2_X1 U297 ( .A1(n8447), .A2(n8448), .ZN(n10303) );
  OR2_X1 U1109 ( .A1(n2746), .A2(n2747), .ZN(n8593) );
  OAI211_X1 U9119 ( .C1(n9451), .C2(n9094), .A(n9093), .B(n9092), .ZN(n10027)
         );
  OAI21_X1 U857 ( .B1(n1255), .B2(n1257), .A(n1254), .ZN(n9697) );
  OR2_X1 U1689 ( .A1(n1738), .A2(n1737), .ZN(n9600) );
  OAI21_X1 U756 ( .B1(n8523), .B2(n8522), .A(n8521), .ZN(n10551) );
  OAI211_X1 U3170 ( .C1(n8866), .C2(n8869), .A(n8123), .B(n8122), .ZN(n10271)
         );
  NAND3_X1 U467 ( .A1(n1766), .A2(n8038), .A3(n8039), .ZN(n10270) );
  MUX2_X1 U400 ( .A(n9223), .B(n9222), .S(n1428), .Z(n10473) );
  OAI21_X1 U928 ( .B1(n8587), .B2(n8588), .A(n2351), .ZN(n10367) );
  NAND2_X1 U320 ( .A1(n8465), .A2(n8464), .ZN(n10557) );
  NAND2_X1 U2099 ( .A1(n9044), .A2(n1932), .ZN(n10046) );
  INV_X1 U2674 ( .A(n10598), .ZN(n10514) );
  OR2_X1 U476 ( .A1(n8863), .A2(n8864), .ZN(n9391) );
  OR2_X1 U44 ( .A1(n9584), .A2(n9583), .ZN(n1032) );
  AOI21_X1 U1867 ( .B1(n8976), .B2(n8977), .A(n8975), .ZN(n9692) );
  OAI21_X1 U249 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n10558) );
  XNOR2_X1 U13694 ( .A(n9798), .B(n9797), .ZN(n11267) );
  XNOR2_X1 U1651 ( .A(n8821), .B(n8822), .ZN(n11170) );
  XNOR2_X1 U1079 ( .A(n10538), .B(n10539), .ZN(n11186) );
  XNOR2_X1 U983 ( .A(n8536), .B(n8535), .ZN(n11528) );
  XNOR2_X1 U157 ( .A(n550), .B(n9859), .ZN(n9883) );
  XNOR2_X1 U303 ( .A(n9708), .B(n9707), .ZN(n11330) );
  BUF_X1 U8787 ( .A(n11240), .Z(n10798) );
  XNOR2_X1 U829 ( .A(n9541), .B(n9540), .ZN(n11142) );
  XNOR2_X1 U13456 ( .A(n10520), .B(n10521), .ZN(n11035) );
  BUF_X1 U364 ( .A(n9545), .Z(n937) );
  XNOR2_X1 U52 ( .A(n10460), .B(n10459), .ZN(n10845) );
  BUF_X1 U505 ( .A(n10060), .Z(n11480) );
  BUF_X1 U19745 ( .A(n10742), .Z(n10936) );
  BUF_X1 U890 ( .A(n11104), .Z(n11041) );
  OR2_X1 U17 ( .A1(n10966), .A2(n3361), .ZN(n12220) );
  OAI211_X1 U398 ( .C1(n11282), .C2(n10695), .A(n1847), .B(n1848), .ZN(n180)
         );
  MUX2_X1 U14071 ( .A(n11537), .B(n11536), .S(n11535), .Z(n11543) );
  OAI21_X1 U331 ( .B1(n9747), .B2(n9746), .A(n9745), .ZN(n12009) );
  OR2_X1 U238 ( .A1(n12552), .A2(n12548), .ZN(n12542) );
  NAND2_X1 U639 ( .A1(n10759), .A2(n2522), .ZN(n2523) );
  NOR2_X1 U3573 ( .A1(n10857), .A2(n11378), .ZN(n2606) );
  AOI21_X1 U1559 ( .B1(n1498), .B2(n1497), .A(n606), .ZN(n11841) );
  AND2_X1 U845 ( .A1(n9973), .A2(n2704), .ZN(n12005) );
  AND2_X1 U1574 ( .A1(n1804), .A2(n11453), .ZN(n12460) );
  AND2_X1 U1567 ( .A1(n11252), .A2(n1599), .ZN(n12381) );
  INV_X1 U844 ( .A(n12005), .ZN(n201) );
  AND2_X1 U1533 ( .A1(n3613), .A2(n3616), .ZN(n11977) );
  NAND2_X1 U661 ( .A1(n10067), .A2(n1418), .ZN(n12499) );
  NAND2_X1 U8172 ( .A1(n11517), .A2(n11518), .ZN(n12533) );
  AND3_X1 U1540 ( .A1(n3630), .A2(n965), .A3(n3629), .ZN(n12338) );
  AOI21_X1 U1563 ( .B1(n11498), .B2(n11497), .A(n11496), .ZN(n12162) );
  NOR2_X1 U527 ( .A1(n12207), .A2(n12208), .ZN(n12065) );
  NAND2_X1 U1090 ( .A1(n10669), .A2(n1917), .ZN(n12443) );
  CLKBUF_X1 U564 ( .A(n12631), .Z(n20184) );
  AND2_X2 U2888 ( .A1(n724), .A2(n721), .ZN(n12500) );
  NAND2_X1 U2198 ( .A1(n371), .A2(n373), .ZN(n12502) );
  OR3_X1 U18272 ( .A1(n12595), .A2(n12589), .A3(n12202), .ZN(n12203) );
  OAI21_X1 U35 ( .B1(n10837), .B2(n10836), .A(n10835), .ZN(n12200) );
  NOR2_X1 U2771 ( .A1(n12374), .A2(n12269), .ZN(n12377) );
  NAND2_X1 U967 ( .A1(n313), .A2(n3480), .ZN(n12537) );
  OR3_X1 U8432 ( .A1(n12338), .A2(n12336), .A3(n12335), .ZN(n12343) );
  BUF_X1 U11582 ( .A(n13702), .Z(n20155) );
  OAI21_X1 U414 ( .B1(n12134), .B2(n11590), .A(n11589), .ZN(n13425) );
  AND3_X1 U25 ( .A1(n513), .A2(n512), .A3(n33), .ZN(n13018) );
  AOI21_X1 U853 ( .B1(n12052), .B2(n12051), .A(n12050), .ZN(n13260) );
  OAI211_X1 U14726 ( .C1(n11807), .C2(n12537), .A(n11806), .B(n11805), .ZN(
        n19892) );
  NOR2_X1 U1504 ( .A1(n9622), .A2(n9621), .ZN(n12696) );
  NOR2_X1 U1503 ( .A1(n11858), .A2(n11857), .ZN(n12471) );
  OR2_X1 U5499 ( .A1(n12432), .A2(n12431), .ZN(n12433) );
  MUX2_X1 U2769 ( .A(n12239), .B(n12238), .S(n12606), .Z(n13755) );
  NAND3_X1 U535 ( .A1(n3631), .A2(n3633), .A3(n11601), .ZN(n13368) );
  AND3_X1 U109 ( .A1(n588), .A2(n1116), .A3(n1117), .ZN(n13042) );
  AND2_X1 U1522 ( .A1(n1258), .A2(n1224), .ZN(n1260) );
  MUX2_X1 U426 ( .A(n11584), .B(n11583), .S(n12040), .Z(n12863) );
  AOI22_X1 U4524 ( .A1(n12502), .A2(n12503), .B1(n12501), .B2(n201), .ZN(
        n13468) );
  OAI211_X1 U14123 ( .C1(n11617), .C2(n11616), .A(n11615), .B(n11614), .ZN(
        n13774) );
  MUX2_X1 U1784 ( .A(n11678), .B(n11677), .S(n11820), .Z(n13687) );
  NAND2_X1 U2381 ( .A1(n458), .A2(n11723), .ZN(n13517) );
  OAI21_X1 U3612 ( .B1(n12610), .B2(n11630), .A(n3761), .ZN(n13580) );
  AND2_X1 U236 ( .A1(n19557), .A2(n19555), .ZN(n13643) );
  XNOR2_X1 U91 ( .A(n3364), .B(n3363), .ZN(n14663) );
  XNOR2_X1 U886 ( .A(n13487), .B(n13488), .ZN(n14747) );
  XNOR2_X1 U992 ( .A(n13084), .B(n13083), .ZN(n15120) );
  XNOR2_X1 U48 ( .A(n11715), .B(n11716), .ZN(n14593) );
  XNOR2_X1 U811 ( .A(n13220), .B(n13219), .ZN(n14547) );
  XNOR2_X1 U17534 ( .A(n13593), .B(n13594), .ZN(n14394) );
  BUF_X1 U1444 ( .A(n14388), .Z(n14723) );
  OAI21_X1 U3282 ( .B1(n14307), .B2(n14499), .A(n3034), .ZN(n13975) );
  MUX2_X1 U9597 ( .A(n14794), .B(n14793), .S(n2412), .Z(n15815) );
  OAI21_X1 U1781 ( .B1(n14174), .B2(n774), .A(n14173), .ZN(n15309) );
  AND4_X1 U2442 ( .A1(n3245), .A2(n3244), .A3(n2839), .A4(n13016), .ZN(n15684)
         );
  AND3_X1 U4983 ( .A1(n1292), .A2(n1294), .A3(n1024), .ZN(n15898) );
  NAND2_X1 U9571 ( .A1(n1625), .A2(n1624), .ZN(n15551) );
  AND3_X1 U596 ( .A1(n2775), .A2(n2774), .A3(n2773), .ZN(n15187) );
  BUF_X1 U3071 ( .A(n15341), .Z(n19888) );
  CLKBUF_X1 U119 ( .A(n14902), .Z(n20147) );
  NAND3_X1 U216 ( .A1(n3539), .A2(n3538), .A3(n14080), .ZN(n15521) );
  NAND3_X1 U247 ( .A1(n14008), .A2(n36), .A3(n35), .ZN(n15698) );
  BUF_X1 U591 ( .A(n14997), .Z(n15257) );
  NOR2_X1 U2573 ( .A1(n13683), .A2(n530), .ZN(n15228) );
  OAI21_X1 U3104 ( .B1(n14025), .B2(n2626), .A(n14024), .ZN(n15754) );
  NOR2_X2 U16201 ( .A1(n20182), .A2(n15803), .ZN(n15802) );
  NOR2_X1 U3125 ( .A1(n15819), .A2(n2114), .ZN(n17110) );
  NAND2_X1 U15730 ( .A1(n13917), .A2(n13916), .ZN(n16931) );
  AND2_X1 U1280 ( .A1(n3103), .A2(n14900), .ZN(n17377) );
  XNOR2_X1 U16292 ( .A(n14885), .B(n14884), .ZN(n17210) );
  XNOR2_X1 U11687 ( .A(n16986), .B(n16985), .ZN(n18025) );
  BUF_X1 U1331 ( .A(n19737), .Z(n18103) );
  OR2_X1 U990 ( .A1(n17654), .A2(n20004), .ZN(n19399) );
  AOI21_X1 U86 ( .B1(n17516), .B2(n17515), .A(n17514), .ZN(n18512) );
  OR2_X1 U1224 ( .A1(n1712), .A2(n3485), .ZN(n18376) );
  NOR2_X1 U1565 ( .A1(n17675), .A2(n17674), .ZN(n19278) );
  AOI22_X1 U19528 ( .A1(n19406), .A2(n19405), .B1(n19403), .B2(n19404), .ZN(
        n19432) );
  OAI211_X1 U1041 ( .C1(n19400), .C2(n19399), .A(n19398), .B(n19397), .ZN(
        n19441) );
  OR2_X1 U1294 ( .A1(n18117), .A2(n18116), .ZN(n18634) );
  AND2_X1 U204 ( .A1(n17659), .A2(n17658), .ZN(n19246) );
  NAND3_X1 U19739 ( .A1(n17722), .A2(n17721), .A3(n17720), .ZN(n19032) );
  AND3_X1 U18641 ( .A1(n17963), .A2(n17962), .A3(n17961), .ZN(n18671) );
  NAND2_X1 U256 ( .A1(n17560), .A2(n18211), .ZN(n18625) );
  NOR2_X1 U3061 ( .A1(n19283), .A2(n19282), .ZN(n19304) );
  NAND3_X4 U758 ( .A1(n5885), .A2(n2928), .A3(n4057), .ZN(n6046) );
  OR2_X1 U7690 ( .A1(n4550), .A2(n3094), .ZN(n5768) );
  INV_X1 U6884 ( .A(n7862), .ZN(n3775) );
  CLKBUF_X1 U2538 ( .A(n8060), .Z(n7893) );
  AND3_X1 U1759 ( .A1(n7876), .A2(n7599), .A3(n7598), .ZN(n8945) );
  INV_X2 U411 ( .A(n9151), .ZN(n9145) );
  INV_X1 U7986 ( .A(n9291), .ZN(n9579) );
  INV_X2 U12080 ( .A(n8596), .ZN(n8933) );
  BUF_X1 U1708 ( .A(n8419), .Z(n9137) );
  INV_X1 U973 ( .A(n11290), .ZN(n19506) );
  INV_X1 U13915 ( .A(n12280), .ZN(n12040) );
  NAND3_X1 U734 ( .A1(n1315), .A2(n1318), .A3(n1314), .ZN(n12642) );
  NAND2_X1 U6827 ( .A1(n12785), .A2(n12784), .ZN(n13312) );
  NOR2_X1 U1062 ( .A1(n2806), .A2(n13890), .ZN(n15857) );
  AND2_X2 U516 ( .A1(n6361), .A2(n6360), .ZN(n8884) );
  NOR2_X2 U308 ( .A1(n14317), .A2(n14318), .ZN(n14903) );
  OR2_X2 U5498 ( .A1(n12433), .A2(n1550), .ZN(n13747) );
  AND2_X2 U690 ( .A1(n3850), .A2(n3849), .ZN(n6064) );
  OR2_X2 U8110 ( .A1(n8909), .A2(n8908), .ZN(n8917) );
  MUX2_X2 U4285 ( .A(n7955), .B(n7954), .S(n7953), .Z(n9167) );
  AND3_X2 U1427 ( .A1(n18236), .A2(n18235), .A3(n18234), .ZN(n18762) );
  NAND3_X2 U513 ( .A1(n662), .A2(n4556), .A3(n661), .ZN(n5802) );
  AND2_X2 U99 ( .A1(n20027), .A2(n20026), .ZN(n12429) );
  AND2_X2 U191 ( .A1(n760), .A2(n761), .ZN(n5201) );
  XNOR2_X2 U831 ( .A(n6399), .B(n6400), .ZN(n8365) );
  NAND2_X2 U524 ( .A1(n3407), .A2(n5521), .ZN(n6736) );
  AND2_X2 U1654 ( .A1(n2617), .A2(n969), .ZN(n10105) );
  OAI211_X2 U624 ( .C1(n12388), .C2(n12470), .A(n1946), .B(n1945), .ZN(n12992)
         );
  OR2_X2 U637 ( .A1(n3332), .A2(n3331), .ZN(n15007) );
  NAND2_X2 U1923 ( .A1(n20292), .A2(n667), .ZN(n670) );
  OR2_X2 U495 ( .A1(n11740), .A2(n11744), .ZN(n12274) );
  XNOR2_X2 U11214 ( .A(n7192), .B(n7191), .ZN(n8315) );
  AND3_X2 U878 ( .A1(n2150), .A2(n8835), .A3(n8834), .ZN(n9934) );
  XNOR2_X2 U672 ( .A(Key[147]), .B(Plaintext[147]), .ZN(n4204) );
  BUF_X2 U617 ( .A(n17758), .Z(n18753) );
  AOI21_X2 U19616 ( .B1(n12276), .B2(n12300), .A(n1872), .ZN(n19883) );
  INV_X2 U10046 ( .A(n5556), .ZN(n8411) );
  AND3_X2 U869 ( .A1(n1719), .A2(n1720), .A3(n452), .ZN(n5320) );
  BUF_X2 U18489 ( .A(n16743), .Z(n20267) );
  AOI22_X2 U18497 ( .A1(n1682), .A2(n15588), .B1(n14040), .B2(n15755), .ZN(
        n16743) );
  OR2_X2 U175 ( .A1(n5121), .A2(n5120), .ZN(n5917) );
  NAND2_X2 U2954 ( .A1(n1825), .A2(n7977), .ZN(n8569) );
  OAI211_X2 U104 ( .C1(n14219), .C2(n3697), .A(n14217), .B(n14218), .ZN(n15405) );
  AND4_X2 U4733 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n12237) );
  AOI21_X2 U16465 ( .B1(n15063), .B2(n15064), .A(n15062), .ZN(n16690) );
  OAI21_X2 U193 ( .B1(n11040), .B2(n11039), .A(n3459), .ZN(n12261) );
  BUF_X2 U12047 ( .A(n10761), .Z(n11544) );
  NAND3_X2 U2636 ( .A1(n566), .A2(n2866), .A3(n2868), .ZN(n657) );
  AND2_X2 U2413 ( .A1(n3251), .A2(n475), .ZN(n9564) );
  NAND2_X2 U7561 ( .A1(n17077), .A2(n1109), .ZN(n19165) );
  INV_X2 U542 ( .A(n15495), .ZN(n3431) );
  BUF_X2 U1358 ( .A(n14722), .Z(n19843) );
  AND2_X2 U7845 ( .A1(n3289), .A2(n4109), .ZN(n5815) );
  XNOR2_X2 U5497 ( .A(n6424), .B(n6425), .ZN(n7748) );
  OAI211_X2 U860 ( .C1(n8260), .C2(n8259), .A(n8258), .B(n8257), .ZN(n8276) );
  OR2_X2 U965 ( .A1(n5414), .A2(n5413), .ZN(n7014) );
  BUF_X2 U882 ( .A(n8156), .Z(n9338) );
  OR2_X2 U2351 ( .A1(n12408), .A2(n12389), .ZN(n12412) );
  NOR2_X2 U180 ( .A1(n9382), .A2(n9381), .ZN(n10579) );
  MUX2_X2 U1735 ( .A(n8907), .B(n8911), .S(n8910), .Z(n8923) );
  NAND4_X2 U1871 ( .A1(n4212), .A2(n2718), .A3(n4211), .A4(n4210), .ZN(n6489)
         );
  BUF_X2 U855 ( .A(n4656), .Z(n164) );
  BUF_X2 U1042 ( .A(n18709), .Z(n18781) );
  NAND3_X2 U7624 ( .A1(n9561), .A2(n9562), .A3(n3023), .ZN(n11829) );
  AND3_X2 U350 ( .A1(n16268), .A2(n16267), .A3(n1248), .ZN(n19208) );
  XNOR2_X2 U113 ( .A(n16723), .B(n16722), .ZN(n18961) );
  OAI211_X2 U14379 ( .C1(n11959), .C2(n11958), .A(n11957), .B(n11956), .ZN(
        n13736) );
  NAND2_X2 U7643 ( .A1(n15591), .A2(n15590), .ZN(n16928) );
  OAI211_X2 U5813 ( .C1(n8299), .C2(n5963), .A(n19578), .B(n19577), .ZN(n9234)
         );
  OR2_X2 U1889 ( .A1(n4273), .A2(n4272), .ZN(n5622) );
  AND3_X2 U1484 ( .A1(n17844), .A2(n17843), .A3(n17842), .ZN(n19067) );
  XNOR2_X2 U986 ( .A(Key[67]), .B(Plaintext[67]), .ZN(n4840) );
  NAND2_X2 U421 ( .A1(n2481), .A2(n4884), .ZN(n7188) );
  OR2_X2 U1588 ( .A1(n11248), .A2(n11247), .ZN(n12269) );
  INV_X2 U450 ( .A(n13514), .ZN(n13397) );
  MUX2_X2 U4825 ( .A(n11676), .B(n11675), .S(n11674), .Z(n13514) );
  NOR2_X2 U16518 ( .A1(n6188), .A2(n6187), .ZN(n6967) );
  OAI21_X2 U1377 ( .B1(n15419), .B2(n15910), .A(n2577), .ZN(n16236) );
  XNOR2_X2 U684 ( .A(Key[12]), .B(Plaintext[12]), .ZN(n4982) );
  BUF_X2 U336 ( .A(n6344), .Z(n8359) );
  OAI21_X2 U1861 ( .B1(n5254), .B2(n5367), .A(n5253), .ZN(n6977) );
  BUF_X2 U980 ( .A(n5117), .Z(n19508) );
  XNOR2_X2 U1458 ( .A(n12847), .B(n12848), .ZN(n14453) );
  MUX2_X2 U2463 ( .A(n10820), .B(n10819), .S(n11365), .Z(n11811) );
  OR2_X2 U1440 ( .A1(n19442), .A2(n19441), .ZN(n19425) );
  NAND3_X2 U1857 ( .A1(n1563), .A2(n4025), .A3(n1561), .ZN(n6745) );
  BUF_X2 U2484 ( .A(n6702), .Z(n8114) );
  NAND2_X2 U1134 ( .A1(n434), .A2(n432), .ZN(n6044) );
  BUF_X2 U762 ( .A(n3897), .Z(n4988) );
  OAI211_X2 U1664 ( .C1(n8683), .C2(n9149), .A(n392), .B(n391), .ZN(n9777) );
  NAND2_X2 U343 ( .A1(n2111), .A2(n2110), .ZN(n17275) );
  NOR2_X2 U1994 ( .A1(n5679), .A2(n5678), .ZN(n19764) );
  XNOR2_X2 U8985 ( .A(Key[117]), .B(Plaintext[117]), .ZN(n4439) );
  NAND4_X2 U11737 ( .A1(n7941), .A2(n7940), .A3(n7939), .A4(n7938), .ZN(n8786)
         );
  NAND2_X2 U1734 ( .A1(n13804), .A2(n67), .ZN(n15442) );
  BUF_X2 U873 ( .A(n10048), .Z(n19990) );
  MUX2_X2 U865 ( .A(n7401), .B(n7400), .S(n8026), .Z(n8596) );
  BUF_X2 U335 ( .A(n9919), .Z(n11219) );
  AND2_X2 U276 ( .A1(n2859), .A2(n2856), .ZN(n12440) );
  NOR2_X2 U1361 ( .A1(n485), .A2(n11774), .ZN(n13539) );
  NAND3_X2 U1928 ( .A1(n523), .A2(n973), .A3(n4225), .ZN(n5825) );
  BUF_X1 U933 ( .A(n4686), .Z(n176) );
  XNOR2_X2 U1466 ( .A(n13208), .B(n13209), .ZN(n14656) );
  BUF_X2 U985 ( .A(n11325), .Z(n191) );
  BUF_X2 U15 ( .A(n15153), .Z(n16015) );
  AND2_X2 U1300 ( .A1(n15253), .A2(n15254), .ZN(n18427) );
  BUF_X2 U341 ( .A(n12973), .Z(n14637) );
  NOR2_X2 U1581 ( .A1(n10994), .A2(n10993), .ZN(n12576) );
  AND3_X2 U4814 ( .A1(n20030), .A2(n3178), .A3(n14054), .ZN(n15266) );
  XNOR2_X2 U2315 ( .A(n2036), .B(Key[29]), .ZN(n4887) );
  AOI21_X2 U1418 ( .B1(n14538), .B2(n13179), .A(n13178), .ZN(n14866) );
  OAI21_X2 U563 ( .B1(n11262), .B2(n11261), .A(n11260), .ZN(n12373) );
  XNOR2_X2 U17057 ( .A(n16028), .B(n16029), .ZN(n17896) );
  OR2_X2 U1858 ( .A1(n3936), .A2(n3935), .ZN(n6693) );
  BUF_X2 U18850 ( .A(n7115), .Z(n6478) );
  CLKBUF_X3 U430 ( .A(n14052), .Z(n14359) );
  OR2_X2 U366 ( .A1(n8422), .A2(n8421), .ZN(n1960) );
  NAND2_X2 U701 ( .A1(n1518), .A2(n1519), .ZN(n15577) );
  AND2_X2 U718 ( .A1(n2930), .A2(n2933), .ZN(n9210) );
  AOI21_X2 U676 ( .B1(n14399), .B2(n14398), .A(n14397), .ZN(n15627) );
  AOI21_X2 U599 ( .B1(n10656), .B2(n2231), .A(n3219), .ZN(n12417) );
  XNOR2_X2 U833 ( .A(n8607), .B(n8608), .ZN(n11550) );
  BUF_X2 U748 ( .A(n17261), .Z(n947) );
  NOR2_X2 U1897 ( .A1(n9002), .A2(n20037), .ZN(n10026) );
  NAND2_X2 U1299 ( .A1(n16451), .A2(n19695), .ZN(n18555) );
  OR2_X2 U3742 ( .A1(n5027), .A2(n5026), .ZN(n3309) );
  OR2_X2 U8495 ( .A1(n4744), .A2(n4745), .ZN(n4559) );
  XNOR2_X2 U8827 ( .A(Key[148]), .B(Plaintext[148]), .ZN(n4745) );
  AND3_X2 U590 ( .A1(n14832), .A2(n14831), .A3(n2779), .ZN(n15581) );
  OR2_X2 U4523 ( .A1(n5408), .A2(n3959), .ZN(n5572) );
  CLKBUF_X2 U5036 ( .A(n5005), .Z(n4248) );
  AND2_X1 U1922 ( .A1(n4009), .A2(n4008), .ZN(n5395) );
  MUX2_X1 U6914 ( .A(n8089), .B(n8088), .S(n20254), .Z(n9333) );
  BUF_X1 U801 ( .A(n10194), .Z(n11265) );
  BUF_X1 U1623 ( .A(n10450), .Z(n11202) );
  INV_X1 U1596 ( .A(n10785), .ZN(n1039) );
  OR2_X1 U1825 ( .A1(n11328), .A2(n11244), .ZN(n11375) );
  BUF_X2 U680 ( .A(n11563), .Z(n11782) );
  BUF_X2 U5 ( .A(n12290), .Z(n182) );
  OAI211_X1 U221 ( .C1(n12082), .C2(n11608), .A(n11607), .B(n11606), .ZN(
        n13277) );
  AND2_X1 U1491 ( .A1(n1509), .A2(n1513), .ZN(n13344) );
  AND3_X1 U1487 ( .A1(n19527), .A2(n852), .A3(n851), .ZN(n13126) );
  BUF_X2 U2456 ( .A(n12842), .Z(n15336) );
  AND3_X1 U895 ( .A1(n3644), .A2(n3643), .A3(n15757), .ZN(n15756) );
  AND3_X1 U2841 ( .A1(n1368), .A2(n14661), .A3(n681), .ZN(n15574) );
  BUF_X1 U530 ( .A(n15994), .Z(n17330) );
  OR2_X1 U4090 ( .A1(n17063), .A2(n17840), .ZN(n3287) );
  NAND3_X1 U6 ( .A1(n2144), .A2(n5779), .A3(n146), .ZN(n6839) );
  BUF_X2 U16 ( .A(n4882), .Z(n5741) );
  AND3_X2 U18 ( .A1(n7438), .A2(n20029), .A3(n7440), .ZN(n9602) );
  MUX2_X2 U23 ( .A(n3208), .B(n18237), .S(n18240), .Z(n3206) );
  NAND2_X2 U27 ( .A1(n20690), .A2(n1481), .ZN(n9922) );
  OR2_X2 U40 ( .A1(n3563), .A2(n3564), .ZN(n6155) );
  NOR2_X2 U42 ( .A1(n16441), .A2(n16440), .ZN(n18567) );
  AND2_X2 U58 ( .A1(n12037), .A2(n12036), .ZN(n11717) );
  NAND2_X2 U67 ( .A1(n4710), .A2(n20679), .ZN(n6184) );
  NOR2_X2 U77 ( .A1(n12524), .A2(n12167), .ZN(n12522) );
  AOI21_X2 U82 ( .B1(n9133), .B2(n9132), .A(n9131), .ZN(n19945) );
  XNOR2_X2 U87 ( .A(n13441), .B(n13442), .ZN(n14555) );
  BUF_X2 U98 ( .A(n4868), .Z(n20357) );
  NAND2_X2 U108 ( .A1(n515), .A2(n20649), .ZN(n7240) );
  XNOR2_X2 U114 ( .A(n10512), .B(n10511), .ZN(n11037) );
  AND2_X2 U126 ( .A1(n2578), .A2(n15906), .ZN(n15912) );
  BUF_X2 U145 ( .A(n17935), .Z(n18357) );
  OAI21_X1 U148 ( .B1(n3081), .B2(n17507), .A(n3080), .ZN(n18467) );
  XNOR2_X1 U159 ( .A(n15249), .B(n19893), .ZN(n15968) );
  OAI21_X1 U171 ( .B1(n11771), .B2(n12292), .A(n11770), .ZN(n13255) );
  BUF_X1 U181 ( .A(n7764), .Z(n20358) );
  BUF_X1 U183 ( .A(n7764), .Z(n20360) );
  OAI211_X1 U192 ( .C1(n4743), .C2(n5055), .A(n4742), .B(n4741), .ZN(n6104) );
  XNOR2_X1 U215 ( .A(n16877), .B(n16876), .ZN(n18977) );
  XOR2_X1 U223 ( .A(n7280), .B(n7281), .Z(n20347) );
  NOR2_X2 U246 ( .A1(n7429), .A2(n7428), .ZN(n9304) );
  XNOR2_X2 U260 ( .A(n10102), .B(n10101), .ZN(n19949) );
  OR2_X2 U262 ( .A1(n10983), .A2(n10984), .ZN(n11686) );
  AOI22_X2 U263 ( .A1(n11785), .A2(n11784), .B1(n920), .B2(n11783), .ZN(n13602) );
  XNOR2_X2 U268 ( .A(n2783), .B(n2784), .ZN(n14818) );
  OAI21_X2 U279 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(n868) );
  NOR2_X2 U285 ( .A1(n15144), .A2(n15143), .ZN(n19720) );
  BUF_X2 U296 ( .A(n17244), .Z(n20354) );
  OAI21_X2 U300 ( .B1(n19379), .B2(n19733), .A(n19378), .ZN(n19439) );
  MUX2_X2 U301 ( .A(n17709), .B(n17708), .S(n18941), .Z(n19047) );
  AND2_X2 U305 ( .A1(n3499), .A2(n10767), .ZN(n13617) );
  XNOR2_X2 U327 ( .A(Key[27]), .B(Plaintext[27]), .ZN(n4118) );
  XNOR2_X2 U332 ( .A(Key[109]), .B(Plaintext[109]), .ZN(n5086) );
  XNOR2_X2 U333 ( .A(n16833), .B(n16832), .ZN(n18270) );
  XNOR2_X2 U339 ( .A(n11818), .B(n11819), .ZN(n14627) );
  NAND2_X2 U342 ( .A1(n578), .A2(n6094), .ZN(n7026) );
  XNOR2_X2 U344 ( .A(n3994), .B(Key[58]), .ZN(n4684) );
  OAI21_X2 U346 ( .B1(n8391), .B2(n8392), .A(n8390), .ZN(n803) );
  NAND4_X2 U348 ( .A1(n9336), .A2(n9337), .A3(n9334), .A4(n9335), .ZN(n10248)
         );
  CLKBUF_X1 U372 ( .A(n18635), .Z(n20348) );
  BUF_X2 U374 ( .A(n18635), .Z(n20349) );
  XNOR2_X1 U376 ( .A(n16357), .B(n16356), .ZN(n18635) );
  OAI21_X2 U380 ( .B1(n15160), .B2(n13887), .A(n13886), .ZN(n16587) );
  OAI21_X2 U385 ( .B1(n3183), .B2(n972), .A(n3185), .ZN(n10280) );
  AOI22_X2 U392 ( .A1(n3943), .A2(n3942), .B1(n3941), .B2(n19581), .ZN(n5581)
         );
  AND2_X2 U399 ( .A1(n7875), .A2(n7874), .ZN(n8991) );
  XNOR2_X2 U402 ( .A(Key[44]), .B(Plaintext[44]), .ZN(n4482) );
  BUF_X2 U409 ( .A(n9250), .Z(n9252) );
  XNOR2_X2 U412 ( .A(Plaintext[38]), .B(Key[38]), .ZN(n4892) );
  XNOR2_X2 U429 ( .A(n6965), .B(n6964), .ZN(n7972) );
  NAND3_X2 U442 ( .A1(n2025), .A2(n7465), .A3(n2024), .ZN(n10482) );
  OAI211_X2 U455 ( .C1(n5660), .C2(n4776), .A(n4775), .B(n368), .ZN(n7384) );
  XNOR2_X2 U477 ( .A(n6683), .B(n6684), .ZN(n8261) );
  AOI21_X2 U480 ( .B1(n13880), .B2(n13879), .A(n13878), .ZN(n15195) );
  CLKBUF_X1 U482 ( .A(n12421), .Z(n20350) );
  BUF_X1 U485 ( .A(n12421), .Z(n20351) );
  BUF_X1 U486 ( .A(n12421), .Z(n20352) );
  NAND2_X2 U490 ( .A1(n787), .A2(n15404), .ZN(n16568) );
  XNOR2_X2 U492 ( .A(n6238), .B(n6239), .ZN(n7936) );
  AOI22_X2 U499 ( .A1(n1591), .A2(n12615), .B1(n874), .B2(n12242), .ZN(n11983)
         );
  NAND2_X2 U506 ( .A1(n8739), .A2(n3504), .ZN(n9902) );
  NOR2_X2 U523 ( .A1(n13055), .A2(n13056), .ZN(n15454) );
  NAND3_X2 U531 ( .A1(n697), .A2(n12132), .A3(n695), .ZN(n13250) );
  AND2_X2 U538 ( .A1(n8715), .A2(n8714), .ZN(n9646) );
  XNOR2_X2 U543 ( .A(n2990), .B(Key[142]), .ZN(n5018) );
  XNOR2_X2 U548 ( .A(Key[133]), .B(Plaintext[133]), .ZN(n5022) );
  XNOR2_X2 U556 ( .A(n12560), .B(n12561), .ZN(n14790) );
  NOR2_X2 U562 ( .A1(n10311), .A2(n10312), .ZN(n12332) );
  OAI21_X2 U600 ( .B1(n9517), .B2(n1670), .A(n1669), .ZN(n11670) );
  MUX2_X2 U601 ( .A(n8404), .B(n8403), .S(n9166), .Z(n10472) );
  OAI21_X2 U602 ( .B1(n14004), .B2(n14003), .A(n14002), .ZN(n15695) );
  OAI211_X2 U610 ( .C1(n31), .C2(n5470), .A(n5469), .B(n5468), .ZN(n7263) );
  XNOR2_X2 U629 ( .A(n13450), .B(n13449), .ZN(n14554) );
  OAI211_X2 U633 ( .C1(n20439), .C2(n4822), .A(n5948), .B(n4821), .ZN(n6918)
         );
  NAND2_X2 U640 ( .A1(n15913), .A2(n1152), .ZN(n16225) );
  XNOR2_X2 U645 ( .A(Key[92]), .B(Plaintext[92]), .ZN(n5092) );
  BUF_X1 U660 ( .A(n17244), .Z(n20353) );
  XNOR2_X1 U662 ( .A(n15998), .B(n15176), .ZN(n17244) );
  OAI21_X2 U681 ( .B1(n4051), .B2(n3259), .A(n4050), .ZN(n6042) );
  XNOR2_X2 U688 ( .A(Key[160]), .B(Plaintext[160]), .ZN(n4574) );
  OAI21_X2 U691 ( .B1(n10940), .B2(n10939), .A(n10938), .ZN(n12228) );
  XNOR2_X2 U693 ( .A(Key[36]), .B(Plaintext[36]), .ZN(n4136) );
  XNOR2_X2 U694 ( .A(n7195), .B(n6300), .ZN(n6824) );
  NAND2_X2 U699 ( .A1(n5206), .A2(n1474), .ZN(n7195) );
  MUX2_X2 U708 ( .A(n4813), .B(n4812), .S(n5080), .Z(n6097) );
  XNOR2_X2 U711 ( .A(n6543), .B(n6544), .ZN(n8232) );
  NOR2_X2 U722 ( .A1(n5679), .A2(n5678), .ZN(n19765) );
  XNOR2_X2 U728 ( .A(n9732), .B(n9731), .ZN(n11397) );
  XNOR2_X2 U730 ( .A(n10169), .B(n10170), .ZN(n11106) );
  XNOR2_X2 U738 ( .A(Key[59]), .B(Plaintext[59]), .ZN(n3996) );
  BUF_X2 U742 ( .A(n12831), .Z(n13544) );
  XNOR2_X2 U747 ( .A(n13814), .B(n13813), .ZN(n14601) );
  NAND2_X2 U749 ( .A1(n8746), .A2(n19604), .ZN(n10213) );
  CLKBUF_X1 U750 ( .A(n4868), .Z(n20355) );
  CLKBUF_X1 U761 ( .A(n4868), .Z(n20356) );
  XNOR2_X1 U765 ( .A(n3982), .B(Key[65]), .ZN(n4868) );
  NAND3_X2 U776 ( .A1(n1437), .A2(n14297), .A3(n14298), .ZN(n16755) );
  AND3_X2 U781 ( .A1(n709), .A2(n711), .A3(n710), .ZN(n9107) );
  NAND4_X2 U785 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n6917)
         );
  XNOR2_X2 U788 ( .A(n13245), .B(n13246), .ZN(n14570) );
  OAI21_X2 U802 ( .B1(n10754), .B2(n10753), .A(n10752), .ZN(n12407) );
  XNOR2_X2 U804 ( .A(Key[47]), .B(Plaintext[47]), .ZN(n4479) );
  OAI211_X2 U815 ( .C1(n12199), .C2(n13907), .A(n12198), .B(n12197), .ZN(
        n15769) );
  NOR2_X2 U816 ( .A1(n14322), .A2(n3149), .ZN(n15553) );
  NOR2_X2 U817 ( .A1(n18050), .A2(n18049), .ZN(n3030) );
  XNOR2_X2 U819 ( .A(Key[158]), .B(Plaintext[158]), .ZN(n4576) );
  AOI21_X2 U825 ( .B1(n12000), .B2(n11999), .A(n2658), .ZN(n13081) );
  OR2_X2 U832 ( .A1(n3323), .A2(n3322), .ZN(n5691) );
  OAI211_X2 U835 ( .C1(n4523), .C2(n4191), .A(n4190), .B(n4189), .ZN(n5425) );
  NAND2_X2 U836 ( .A1(n3334), .A2(n3336), .ZN(n8998) );
  XNOR2_X2 U838 ( .A(n10378), .B(n10377), .ZN(n11133) );
  OAI21_X2 U840 ( .B1(n8476), .B2(n8974), .A(n577), .ZN(n10281) );
  XNOR2_X2 U863 ( .A(n1088), .B(Key[64]), .ZN(n4652) );
  XNOR2_X2 U875 ( .A(Key[3]), .B(Plaintext[3]), .ZN(n4623) );
  OAI211_X2 U881 ( .C1(n5935), .C2(n5934), .A(n5932), .B(n19), .ZN(n6768) );
  OAI21_X2 U883 ( .B1(n9012), .B2(n9013), .A(n9011), .ZN(n10008) );
  XNOR2_X2 U884 ( .A(Key[50]), .B(Plaintext[50]), .ZN(n4907) );
  NOR2_X2 U896 ( .A1(n11892), .A2(n11891), .ZN(n12267) );
  OAI21_X2 U900 ( .B1(n13132), .B2(n14263), .A(n13133), .ZN(n15683) );
  XNOR2_X2 U903 ( .A(n10155), .B(n10156), .ZN(n11105) );
  AOI21_X2 U913 ( .B1(n2002), .B2(n14438), .A(n14437), .ZN(n15297) );
  AOI22_X2 U917 ( .A1(n7847), .A2(n8217), .B1(n7648), .B2(n7647), .ZN(n8742)
         );
  AOI22_X2 U918 ( .A1(n13935), .A2(n13934), .B1(n20453), .B2(n13936), .ZN(
        n15505) );
  OAI21_X2 U925 ( .B1(n20435), .B2(n14969), .A(n14967), .ZN(n17366) );
  XNOR2_X2 U930 ( .A(n17371), .B(n17372), .ZN(n18260) );
  OAI211_X2 U931 ( .C1(n7712), .C2(n8363), .A(n7710), .B(n7711), .ZN(n8879) );
  AND3_X2 U938 ( .A1(n2863), .A2(n3777), .A3(n10070), .ZN(n13588) );
  NOR2_X2 U943 ( .A1(n15118), .A2(n15117), .ZN(n17111) );
  OAI21_X2 U964 ( .B1(n14687), .B2(n859), .A(n14686), .ZN(n16853) );
  AND2_X2 U968 ( .A1(n370), .A2(n11531), .ZN(n9933) );
  XNOR2_X2 U970 ( .A(n8440), .B(n8441), .ZN(n11527) );
  BUF_X1 U979 ( .A(n7764), .Z(n20359) );
  XNOR2_X1 U982 ( .A(n6243), .B(n6242), .ZN(n7764) );
  BUF_X2 U996 ( .A(n18377), .Z(n20361) );
  INV_X1 U997 ( .A(n15454), .ZN(n20362) );
  INV_X1 U1000 ( .A(n14452), .ZN(n14448) );
  INV_X1 U1004 ( .A(n12533), .ZN(n20363) );
  INV_X1 U1018 ( .A(n180), .ZN(n1371) );
  XNOR2_X1 U1030 ( .A(n7131), .B(n7132), .ZN(n7953) );
  BUF_X1 U1040 ( .A(n5118), .Z(n169) );
  CLKBUF_X1 U1054 ( .A(Key[54]), .Z(n20593) );
  CLKBUF_X1 U1060 ( .A(Key[142]), .Z(n20672) );
  CLKBUF_X1 U1080 ( .A(Key[179]), .Z(n18278) );
  BUF_X1 U1081 ( .A(Key[100]), .Z(n20682) );
  BUF_X1 U1083 ( .A(Key[51]), .Z(n2445) );
  CLKBUF_X1 U1087 ( .A(Key[33]), .Z(n18084) );
  CLKBUF_X1 U1091 ( .A(Key[137]), .Z(n2317) );
  AND2_X1 U1106 ( .A1(n16075), .A2(n16076), .ZN(n20460) );
  INV_X1 U1124 ( .A(n19284), .ZN(n20364) );
  OAI21_X1 U1130 ( .B1(n17555), .B2(n18106), .A(n17554), .ZN(n18622) );
  AND3_X1 U1140 ( .A1(n17971), .A2(n17970), .A3(n17969), .ZN(n18672) );
  NAND3_X1 U1149 ( .A1(n17702), .A2(n17703), .A3(n1921), .ZN(n19046) );
  AND3_X1 U1189 ( .A1(n2662), .A2(n2664), .A3(n2660), .ZN(n19682) );
  OR2_X1 U1196 ( .A1(n16815), .A2(n16814), .ZN(n19668) );
  AOI21_X1 U1215 ( .B1(n17159), .B2(n17158), .A(n17157), .ZN(n19656) );
  INV_X1 U1260 ( .A(n18585), .ZN(n20365) );
  BUF_X2 U1273 ( .A(n17497), .Z(n19815) );
  BUF_X1 U1276 ( .A(n17695), .Z(n18962) );
  BUF_X2 U1286 ( .A(n19371), .Z(n19666) );
  XNOR2_X1 U1290 ( .A(n16299), .B(n16298), .ZN(n19403) );
  OR2_X1 U1291 ( .A1(n3710), .A2(n15421), .ZN(n15917) );
  AND2_X1 U1305 ( .A1(n15676), .A2(n15443), .ZN(n20647) );
  NAND3_X1 U1323 ( .A1(n700), .A2(n12927), .A3(n12928), .ZN(n15379) );
  AND2_X1 U1326 ( .A1(n2920), .A2(n20624), .ZN(n15459) );
  NAND2_X1 U1329 ( .A1(n13910), .A2(n2654), .ZN(n2655) );
  NOR2_X1 U1372 ( .A1(n13998), .A2(n13999), .ZN(n20449) );
  OR2_X1 U1373 ( .A1(n14666), .A2(n14667), .ZN(n14315) );
  XNOR2_X1 U1394 ( .A(n2095), .B(n13854), .ZN(n20513) );
  XNOR2_X1 U1404 ( .A(n11318), .B(n11317), .ZN(n14778) );
  XNOR2_X1 U1419 ( .A(n13107), .B(n13106), .ZN(n13981) );
  OAI21_X1 U1425 ( .B1(n12684), .B2(n11613), .A(n11612), .ZN(n13707) );
  OR2_X1 U1428 ( .A1(n11692), .A2(n11646), .ZN(n1951) );
  OR2_X1 U1430 ( .A1(n11464), .A2(n12524), .ZN(n11793) );
  CLKBUF_X1 U1434 ( .A(n12639), .Z(n922) );
  AND2_X1 U1456 ( .A1(n10933), .A2(n3105), .ZN(n20583) );
  MUX2_X1 U1489 ( .A(n10832), .B(n10831), .S(n11420), .Z(n20430) );
  NAND3_X1 U1512 ( .A1(n10707), .A2(n20522), .A3(n20521), .ZN(n12630) );
  OR2_X1 U1530 ( .A1(n10705), .A2(n10951), .ZN(n20522) );
  OR2_X1 U1541 ( .A1(n10708), .A2(n11011), .ZN(n20521) );
  BUF_X2 U1542 ( .A(n11144), .Z(n20366) );
  XNOR2_X1 U1548 ( .A(n9460), .B(n9461), .ZN(n10953) );
  AND2_X1 U1555 ( .A1(n20646), .A2(n506), .ZN(n8746) );
  INV_X1 U1573 ( .A(n9794), .ZN(n20608) );
  OR2_X1 U1578 ( .A1(n363), .A2(n362), .ZN(n10237) );
  OR2_X1 U1584 ( .A1(n8484), .A2(n8602), .ZN(n20659) );
  OR2_X1 U1591 ( .A1(n1507), .A2(n9453), .ZN(n401) );
  AND3_X2 U1600 ( .A1(n1679), .A2(n1678), .A3(n1677), .ZN(n1507) );
  NAND4_X1 U1668 ( .A1(n3581), .A2(n7483), .A3(n7484), .A4(n7482), .ZN(n8812)
         );
  INV_X1 U1669 ( .A(n8208), .ZN(n20585) );
  XNOR2_X1 U1687 ( .A(n6335), .B(n6336), .ZN(n8354) );
  CLKBUF_X1 U1690 ( .A(n6887), .Z(n20455) );
  XNOR2_X1 U1701 ( .A(n6317), .B(n6316), .ZN(n7981) );
  INV_X1 U1705 ( .A(n7479), .ZN(n20367) );
  NAND3_X1 U1731 ( .A1(n2555), .A2(n5459), .A3(n2556), .ZN(n7070) );
  NAND3_X1 U1749 ( .A1(n20411), .A2(n20410), .A3(n4097), .ZN(n5989) );
  NAND2_X1 U1752 ( .A1(n4375), .A2(n4369), .ZN(n5720) );
  INV_X1 U1791 ( .A(n5914), .ZN(n20368) );
  OR2_X1 U1793 ( .A1(n4424), .A2(n4423), .ZN(n20655) );
  OR2_X1 U1797 ( .A1(n4098), .A2(n5024), .ZN(n20411) );
  OR2_X1 U1816 ( .A1(n4711), .A2(n4769), .ZN(n20679) );
  OR2_X1 U1818 ( .A1(n4481), .A2(n3967), .ZN(n20606) );
  XNOR2_X1 U1837 ( .A(n20635), .B(Key[56]), .ZN(n3995) );
  XNOR2_X1 U1845 ( .A(n3970), .B(Key[37]), .ZN(n4960) );
  XNOR2_X1 U1850 ( .A(n3869), .B(Key[31]), .ZN(n4474) );
  OR2_X1 U1866 ( .A1(n2490), .A2(n4987), .ZN(n2489) );
  BUF_X1 U1876 ( .A(n4060), .Z(n4588) );
  AND2_X1 U1904 ( .A1(n3527), .A2(n5685), .ZN(n20553) );
  INV_X1 U1913 ( .A(n6156), .ZN(n20403) );
  AND2_X1 U1952 ( .A1(n5971), .A2(n5699), .ZN(n20674) );
  OAI211_X1 U1960 ( .C1(n5056), .C2(n4739), .A(n4590), .B(n4588), .ZN(n5885)
         );
  INV_X1 U1965 ( .A(n2454), .ZN(n20551) );
  OR2_X1 U1997 ( .A1(n3948), .A2(n4350), .ZN(n4256) );
  BUF_X1 U1999 ( .A(n6404), .Z(n19855) );
  AND2_X1 U2027 ( .A1(n7633), .A2(n20511), .ZN(n20586) );
  AND2_X1 U2028 ( .A1(n19922), .A2(n8205), .ZN(n20584) );
  OR2_X1 U2037 ( .A1(n20177), .A2(n8387), .ZN(n7685) );
  BUF_X1 U2056 ( .A(n8380), .Z(n163) );
  INV_X1 U2058 ( .A(n7953), .ZN(n20013) );
  OR2_X1 U2059 ( .A1(n8744), .A2(n8602), .ZN(n20646) );
  INV_X1 U2110 ( .A(n7590), .ZN(n20651) );
  BUF_X1 U2117 ( .A(n8004), .Z(n8312) );
  AND2_X1 U2119 ( .A1(n19565), .A2(n20554), .ZN(n2888) );
  CLKBUF_X1 U2123 ( .A(n8993), .Z(n19732) );
  INV_X1 U2133 ( .A(n20010), .ZN(n9090) );
  OR2_X1 U2136 ( .A1(n9250), .A2(n9249), .ZN(n9260) );
  OR2_X1 U2139 ( .A1(n9313), .A2(n9228), .ZN(n9227) );
  NOR2_X1 U2140 ( .A1(n20659), .A2(n8485), .ZN(n8486) );
  NAND2_X1 U2158 ( .A1(n10329), .A2(n10328), .ZN(n10052) );
  INV_X1 U2162 ( .A(n8593), .ZN(n10620) );
  AND2_X1 U2170 ( .A1(n8734), .A2(n8499), .ZN(n8334) );
  OAI211_X1 U2190 ( .C1(n8278), .C2(n8279), .A(n8433), .B(n8277), .ZN(n10431)
         );
  AOI21_X1 U2191 ( .B1(n11281), .B2(n11284), .A(n19817), .ZN(n20641) );
  OAI21_X1 U2192 ( .B1(n10719), .B2(n1988), .A(n11192), .ZN(n20561) );
  XNOR2_X1 U2223 ( .A(n8481), .B(n8480), .ZN(n11521) );
  OR2_X1 U2226 ( .A1(n19983), .A2(n11186), .ZN(n20591) );
  AND2_X1 U2240 ( .A1(n19864), .A2(n11513), .ZN(n20560) );
  BUF_X1 U2245 ( .A(n10259), .Z(n11886) );
  INV_X1 U2261 ( .A(n20496), .ZN(n20660) );
  INV_X1 U2266 ( .A(n3401), .ZN(n11722) );
  NOR2_X1 U2286 ( .A1(n10750), .A2(n10749), .ZN(n12408) );
  NOR2_X1 U2322 ( .A1(n12149), .A2(n20618), .ZN(n19558) );
  BUF_X1 U2354 ( .A(n12021), .Z(n20191) );
  AND2_X1 U2361 ( .A1(n11695), .A2(n953), .ZN(n20644) );
  AND3_X2 U2364 ( .A1(n10714), .A2(n10715), .A3(n10713), .ZN(n11618) );
  XNOR2_X1 U2380 ( .A(n13398), .B(n13422), .ZN(n13649) );
  OR2_X1 U2384 ( .A1(n14482), .A2(n14171), .ZN(n14485) );
  XNOR2_X1 U2392 ( .A(n12968), .B(n12967), .ZN(n14512) );
  AND2_X1 U2411 ( .A1(n13556), .A2(n2921), .ZN(n20624) );
  INV_X1 U2418 ( .A(n13931), .ZN(n14339) );
  BUF_X1 U2433 ( .A(n14820), .Z(n912) );
  CLKBUF_X1 U2434 ( .A(n14087), .Z(n19821) );
  NOR2_X1 U2437 ( .A1(n13317), .A2(n14705), .ZN(n13318) );
  NAND2_X1 U2482 ( .A1(n20609), .A2(n19613), .ZN(n15583) );
  OAI211_X1 U2485 ( .C1(n20513), .C2(n2682), .A(n2666), .B(n13855), .ZN(n15443) );
  OR2_X1 U2489 ( .A1(n15677), .A2(n15228), .ZN(n15445) );
  OR2_X1 U2495 ( .A1(n14667), .A2(n14663), .ZN(n13166) );
  MUX2_X1 U2502 ( .A(n14618), .B(n14617), .S(n20112), .Z(n14631) );
  NOR2_X1 U2510 ( .A1(n14670), .A2(n14671), .ZN(n860) );
  INV_X1 U2517 ( .A(n20101), .ZN(n20391) );
  XNOR2_X1 U2521 ( .A(n14956), .B(n16711), .ZN(n17026) );
  OR2_X1 U2541 ( .A1(n17530), .A2(n19110), .ZN(n20661) );
  CLKBUF_X1 U2546 ( .A(n17836), .Z(n20423) );
  XNOR2_X1 U2556 ( .A(n16040), .B(n16041), .ZN(n19707) );
  CLKBUF_X1 U2557 ( .A(n16166), .Z(n16480) );
  AND2_X1 U2563 ( .A1(n811), .A2(n814), .ZN(n20654) );
  NOR2_X1 U2571 ( .A1(n18036), .A2(n18035), .ZN(n18857) );
  CLKBUF_X1 U2617 ( .A(Key[119]), .Z(n17999) );
  INV_X1 U2624 ( .A(n2067), .ZN(n16788) );
  XOR2_X1 U2632 ( .A(Key[176]), .B(Plaintext[176]), .Z(n20369) );
  NAND3_X1 U2634 ( .A1(n2120), .A2(n18932), .A3(n18029), .ZN(n20370) );
  OR2_X1 U2652 ( .A1(n14214), .A2(n15071), .ZN(n20371) );
  XOR2_X1 U2656 ( .A(n17035), .B(n17270), .Z(n20372) );
  INV_X1 U2657 ( .A(n5741), .ZN(n20568) );
  AND2_X1 U2679 ( .A1(n19856), .A2(n8001), .ZN(n20373) );
  INV_X1 U2690 ( .A(n6155), .ZN(n20405) );
  AND2_X1 U2708 ( .A1(n8095), .A2(n7632), .ZN(n20374) );
  OR2_X1 U2727 ( .A1(n10654), .A2(n19872), .ZN(n20375) );
  XOR2_X1 U2734 ( .A(n13373), .B(n13372), .Z(n20376) );
  XOR2_X1 U2777 ( .A(n2095), .B(n13854), .Z(n20377) );
  XOR2_X1 U2779 ( .A(n13622), .B(n18988), .Z(n20378) );
  OR2_X1 U2789 ( .A1(n15535), .A2(n15895), .ZN(n20379) );
  XOR2_X1 U2791 ( .A(n12983), .B(n12982), .Z(n20380) );
  INV_X1 U2821 ( .A(n14778), .ZN(n20408) );
  AND2_X1 U2835 ( .A1(n19940), .A2(n14499), .ZN(n20381) );
  AND2_X1 U2837 ( .A1(n19439), .A2(n19440), .ZN(n20382) );
  AND2_X1 U2838 ( .A1(n19170), .A2(n20394), .ZN(n20383) );
  AND2_X1 U2879 ( .A1(n20396), .A2(n20393), .ZN(n20384) );
  OAI21_X2 U2880 ( .B1(n2671), .B2(n2670), .A(n20385), .ZN(n6101) );
  NAND2_X1 U2889 ( .A1(n4800), .A2(n5043), .ZN(n20385) );
  XNOR2_X1 U2891 ( .A(n20386), .B(n311), .ZN(Ciphertext[14]) );
  NAND2_X1 U2905 ( .A1(n20549), .A2(n15930), .ZN(n20386) );
  NAND3_X2 U2915 ( .A1(n20387), .A2(n7055), .A3(n92), .ZN(n9038) );
  NAND2_X1 U2923 ( .A1(n91), .A2(n90), .ZN(n20387) );
  NAND2_X1 U2941 ( .A1(n6041), .A2(n1214), .ZN(n6043) );
  NAND2_X2 U2973 ( .A1(n1320), .A2(n4043), .ZN(n6041) );
  OR2_X2 U2974 ( .A1(n7630), .A2(n7629), .ZN(n8482) );
  NAND2_X1 U2980 ( .A1(n7626), .A2(n1335), .ZN(n7630) );
  NAND3_X1 U2981 ( .A1(n241), .A2(n20390), .A3(n20388), .ZN(n1700) );
  NAND2_X1 U2995 ( .A1(n20389), .A2(n14547), .ZN(n20388) );
  INV_X1 U3002 ( .A(n20471), .ZN(n20389) );
  OR2_X1 U3012 ( .A1(n14548), .A2(n14547), .ZN(n20390) );
  AND3_X2 U3051 ( .A1(n14068), .A2(n14067), .A3(n2528), .ZN(n864) );
  NAND2_X1 U3052 ( .A1(n3479), .A2(n3478), .ZN(n12531) );
  NAND2_X1 U3063 ( .A1(n20392), .A2(n20391), .ZN(n17950) );
  NAND2_X1 U3066 ( .A1(n18131), .A2(n19744), .ZN(n20392) );
  OAI21_X1 U3067 ( .B1(n9365), .B2(n9366), .A(n9364), .ZN(n598) );
  NAND2_X1 U3091 ( .A1(n8958), .A2(n8960), .ZN(n9366) );
  NAND3_X1 U3094 ( .A1(n20412), .A2(n3346), .A3(n3217), .ZN(n18009) );
  NAND3_X1 U3173 ( .A1(n17951), .A2(n17953), .A3(n17952), .ZN(n18667) );
  AND3_X2 U3175 ( .A1(n2106), .A2(n11135), .A3(n11134), .ZN(n12386) );
  NAND2_X1 U3177 ( .A1(n20395), .A2(n20394), .ZN(n20393) );
  INV_X1 U3178 ( .A(n2368), .ZN(n20394) );
  INV_X1 U3194 ( .A(n18156), .ZN(n20395) );
  NAND2_X1 U3240 ( .A1(n16159), .A2(n20383), .ZN(n20396) );
  XNOR2_X1 U3283 ( .A(n20397), .B(n18066), .ZN(Ciphertext[115]) );
  NAND2_X1 U3301 ( .A1(n2399), .A2(n18063), .ZN(n20397) );
  NAND2_X1 U3334 ( .A1(n19993), .A2(n18061), .ZN(n19035) );
  INV_X1 U3358 ( .A(n792), .ZN(n5613) );
  NAND2_X1 U3395 ( .A1(n6153), .A2(n5611), .ZN(n792) );
  NAND2_X1 U3420 ( .A1(n10989), .A2(n10988), .ZN(n11683) );
  NAND2_X1 U3443 ( .A1(n5956), .A2(n20398), .ZN(n941) );
  NOR2_X1 U3507 ( .A1(n367), .A2(n145), .ZN(n20398) );
  XNOR2_X1 U3514 ( .A(n20399), .B(n15579), .ZN(n15586) );
  XNOR2_X1 U3587 ( .A(n15571), .B(n17407), .ZN(n20399) );
  NAND2_X1 U3588 ( .A1(n20401), .A2(n20400), .ZN(n3401) );
  NAND2_X1 U3589 ( .A1(n10702), .A2(n20366), .ZN(n20400) );
  NAND2_X1 U3594 ( .A1(n10703), .A2(n11140), .ZN(n20401) );
  NAND2_X1 U3597 ( .A1(n5247), .A2(n20402), .ZN(n7254) );
  NAND3_X1 U3604 ( .A1(n20406), .A2(n20404), .A3(n20403), .ZN(n20402) );
  NAND2_X1 U3672 ( .A1(n20405), .A2(n6150), .ZN(n20404) );
  NAND2_X1 U3690 ( .A1(n6151), .A2(n6155), .ZN(n20406) );
  NAND2_X1 U3691 ( .A1(n20409), .A2(n20407), .ZN(n14856) );
  NAND2_X1 U3708 ( .A1(n11320), .A2(n20408), .ZN(n20407) );
  NAND2_X1 U3711 ( .A1(n11319), .A2(n14778), .ZN(n20409) );
  NAND3_X1 U3723 ( .A1(n20043), .A2(n4098), .A3(n5029), .ZN(n20410) );
  NAND2_X1 U3764 ( .A1(n20013), .A2(n7952), .ZN(n7813) );
  BUF_X1 U3783 ( .A(n14781), .Z(n20518) );
  NAND2_X1 U3805 ( .A1(n17490), .A2(n3347), .ZN(n20412) );
  NAND2_X1 U3837 ( .A1(n12095), .A2(n12430), .ZN(n3514) );
  NAND3_X1 U3846 ( .A1(n8727), .A2(n1023), .A3(n20413), .ZN(n1268) );
  NAND2_X1 U3956 ( .A1(n8726), .A2(n9361), .ZN(n20413) );
  NOR2_X2 U3957 ( .A1(n14047), .A2(n20414), .ZN(n15845) );
  NAND2_X1 U3993 ( .A1(n340), .A2(n341), .ZN(n20414) );
  NAND2_X1 U4028 ( .A1(n14405), .A2(n14148), .ZN(n14010) );
  AOI22_X2 U4029 ( .A1(n14183), .A2(n14182), .B1(n14450), .B2(n14181), .ZN(
        n15310) );
  NAND3_X1 U4057 ( .A1(n1213), .A2(n12335), .A3(n11992), .ZN(n11993) );
  OAI211_X2 U4066 ( .C1(n8754), .C2(n8933), .A(n20416), .B(n20415), .ZN(n9952)
         );
  NAND2_X1 U4072 ( .A1(n8750), .A2(n8933), .ZN(n20415) );
  NAND2_X1 U4076 ( .A1(n8751), .A2(n8752), .ZN(n20416) );
  OR2_X1 U4117 ( .A1(n8065), .A2(n1431), .ZN(n20505) );
  AND3_X1 U4120 ( .A1(n13958), .A2(n13956), .A3(n402), .ZN(n19739) );
  XNOR2_X1 U4141 ( .A(n15347), .B(n15346), .ZN(n17501) );
  INV_X1 U4144 ( .A(n19668), .ZN(n20417) );
  AND2_X1 U4162 ( .A1(n14516), .A2(n20206), .ZN(n20636) );
  NAND3_X1 U4180 ( .A1(n20370), .A2(n20613), .A3(n20612), .ZN(n20418) );
  AOI21_X2 U4214 ( .B1(n15605), .B2(n15274), .A(n15011), .ZN(n15935) );
  NAND3_X1 U4262 ( .A1(n20370), .A2(n20613), .A3(n20612), .ZN(n18868) );
  NOR2_X2 U4270 ( .A1(n20419), .A2(n20420), .ZN(n16844) );
  AND2_X1 U4272 ( .A1(n15203), .A2(n16126), .ZN(n20419) );
  NAND2_X1 U4340 ( .A1(n57), .A2(n55), .ZN(n20420) );
  XOR2_X1 U4356 ( .A(n16884), .B(n16883), .Z(n20421) );
  NAND2_X1 U4360 ( .A1(n17313), .A2(n17312), .ZN(n20422) );
  OR2_X1 U4408 ( .A1(n9274), .A2(n885), .ZN(n20554) );
  XNOR2_X1 U4469 ( .A(n16143), .B(n16144), .ZN(n17836) );
  OR2_X1 U4477 ( .A1(n20286), .A2(n19094), .ZN(n2196) );
  OR2_X1 U4498 ( .A1(n20142), .A2(n19031), .ZN(n20528) );
  XNOR2_X1 U4587 ( .A(n13117), .B(n13116), .ZN(n20424) );
  XNOR2_X1 U4635 ( .A(n5297), .B(n6835), .ZN(n8303) );
  XNOR2_X1 U4636 ( .A(n16392), .B(n20426), .ZN(n20425) );
  XOR2_X1 U4638 ( .A(n16840), .B(n16651), .Z(n20426) );
  XNOR2_X1 U4643 ( .A(n11756), .B(n11755), .ZN(n14807) );
  XNOR2_X1 U4644 ( .A(n20425), .B(n16395), .ZN(n19658) );
  XNOR2_X1 U4646 ( .A(n16150), .B(n16149), .ZN(n17715) );
  NOR2_X2 U4658 ( .A1(n16728), .A2(n16729), .ZN(n16780) );
  OAI21_X1 U4672 ( .B1(n15429), .B2(n15428), .A(n15427), .ZN(n15534) );
  AND2_X1 U4677 ( .A1(n9444), .A2(n9443), .ZN(n20427) );
  AND2_X1 U4709 ( .A1(n9444), .A2(n9443), .ZN(n11650) );
  OR2_X1 U4710 ( .A1(n20182), .A2(n15371), .ZN(n20428) );
  BUF_X1 U4717 ( .A(n17572), .Z(n20429) );
  MUX2_X1 U4736 ( .A(n10832), .B(n10831), .S(n11420), .Z(n12594) );
  INV_X1 U4749 ( .A(n5081), .ZN(n20431) );
  AND2_X1 U4760 ( .A1(n12129), .A2(n12126), .ZN(n696) );
  BUF_X1 U4765 ( .A(n14714), .Z(n19862) );
  MUX2_X1 U4770 ( .A(n14860), .B(n14861), .S(n15237), .Z(n14862) );
  INV_X1 U4782 ( .A(n15237), .ZN(n1458) );
  INV_X1 U4792 ( .A(n18382), .ZN(n20611) );
  NOR2_X1 U4809 ( .A1(n19599), .A2(n15180), .ZN(n15186) );
  AND2_X1 U4810 ( .A1(n15656), .A2(n15659), .ZN(n20565) );
  OR2_X1 U4816 ( .A1(n11981), .A2(n20430), .ZN(n20543) );
  NOR2_X1 U4830 ( .A1(n12644), .A2(n12643), .ZN(n13154) );
  XNOR2_X1 U4831 ( .A(n16204), .B(n16203), .ZN(n20432) );
  INV_X1 U4834 ( .A(n214), .ZN(n20433) );
  OAI21_X1 U4860 ( .B1(n17474), .B2(n18539), .A(n17473), .ZN(n18511) );
  AOI22_X1 U4879 ( .A1(n17614), .A2(n17613), .B1(n17612), .B2(n17611), .ZN(
        n20434) );
  NAND2_X1 U4883 ( .A1(n19573), .A2(n14960), .ZN(n16927) );
  NOR2_X1 U4898 ( .A1(n15672), .A2(n20151), .ZN(n15438) );
  NOR2_X1 U4946 ( .A1(n17551), .A2(n17550), .ZN(n18630) );
  AOI22_X1 U4948 ( .A1(n15562), .A2(n15558), .B1(n15510), .B2(n15509), .ZN(
        n20435) );
  MUX2_X1 U4949 ( .A(n9252), .B(n8971), .S(n670), .Z(n7736) );
  XNOR2_X1 U4991 ( .A(n16548), .B(n16547), .ZN(n20436) );
  INV_X1 U5027 ( .A(n18376), .ZN(n20437) );
  CLKBUF_X1 U5029 ( .A(Key[36]), .Z(n620) );
  CLKBUF_X1 U5035 ( .A(n18257), .Z(n20438) );
  INV_X1 U5038 ( .A(n19658), .ZN(n17956) );
  OR2_X1 U5082 ( .A1(n5663), .A2(n5952), .ZN(n20439) );
  OR2_X1 U5095 ( .A1(n5663), .A2(n5952), .ZN(n5661) );
  OAI21_X1 U5099 ( .B1(n12358), .B2(n12357), .A(n12356), .ZN(n20440) );
  OAI21_X1 U5100 ( .B1(n12358), .B2(n12357), .A(n12356), .ZN(n13826) );
  INV_X1 U5110 ( .A(n15228), .ZN(n15679) );
  OR2_X1 U5121 ( .A1(n17208), .A2(n17210), .ZN(n20633) );
  NAND3_X1 U5135 ( .A1(n14933), .A2(n14932), .A3(n460), .ZN(n16602) );
  AND2_X1 U5147 ( .A1(n17565), .A2(n17471), .ZN(n18538) );
  OR2_X1 U5153 ( .A1(n14836), .A2(n15813), .ZN(n579) );
  AOI22_X1 U5184 ( .A1(n5038), .A2(n5039), .B1(n5036), .B2(n5037), .ZN(n6025)
         );
  XNOR2_X1 U5210 ( .A(n6452), .B(n6451), .ZN(n20441) );
  XNOR2_X1 U5215 ( .A(n12906), .B(n13848), .ZN(n20442) );
  XNOR2_X1 U5222 ( .A(n12983), .B(n12982), .ZN(n20443) );
  OAI211_X1 U5228 ( .C1(n18658), .C2(n18659), .A(n20581), .B(n20580), .ZN(
        n18661) );
  CLKBUF_X1 U5231 ( .A(n19276), .Z(n20444) );
  INV_X1 U5258 ( .A(n8831), .ZN(n8829) );
  NAND2_X2 U5285 ( .A1(n1725), .A2(n7535), .ZN(n8736) );
  NAND3_X1 U5292 ( .A1(n17148), .A2(n3065), .A3(n3064), .ZN(n20445) );
  NAND3_X1 U5293 ( .A1(n17148), .A2(n3065), .A3(n3064), .ZN(n18585) );
  OAI21_X1 U5295 ( .B1(n14343), .B2(n14106), .A(n14105), .ZN(n15746) );
  OR2_X1 U5302 ( .A1(n4898), .A2(n20446), .ZN(n2573) );
  NOR2_X1 U5318 ( .A1(n4899), .A2(n4962), .ZN(n20446) );
  OR2_X1 U5329 ( .A1(n16795), .A2(n20648), .ZN(n1337) );
  CLKBUF_X1 U5356 ( .A(n1205), .Z(n20447) );
  BUF_X1 U5364 ( .A(n19274), .Z(n20448) );
  MUX2_X1 U5365 ( .A(n19675), .B(n3347), .S(n17154), .Z(n16247) );
  NOR2_X1 U5401 ( .A1(n11062), .A2(n11726), .ZN(n20623) );
  OR3_X1 U5429 ( .A1(n15857), .A2(n15329), .A3(n15327), .ZN(n15331) );
  OR2_X1 U5438 ( .A1(n15863), .A2(n15857), .ZN(n15332) );
  OAI21_X1 U5439 ( .B1(n2581), .B2(n15870), .A(n15305), .ZN(n20450) );
  OAI21_X1 U5526 ( .B1(n2581), .B2(n15870), .A(n15305), .ZN(n16555) );
  XNOR2_X1 U5537 ( .A(n13373), .B(n13372), .ZN(n20451) );
  NOR2_X1 U5538 ( .A1(n15906), .A2(n2723), .ZN(n15417) );
  XNOR2_X1 U5551 ( .A(n17050), .B(n17049), .ZN(n20452) );
  XNOR2_X1 U5582 ( .A(n17050), .B(n17049), .ZN(n18937) );
  NAND2_X1 U5585 ( .A1(n7850), .A2(n7849), .ZN(n9265) );
  XNOR2_X1 U5646 ( .A(n13467), .B(n20285), .ZN(n20453) );
  XNOR2_X1 U5656 ( .A(n13467), .B(n20285), .ZN(n14426) );
  XNOR2_X1 U5662 ( .A(n11103), .B(n11102), .ZN(n20454) );
  XOR2_X1 U5699 ( .A(n9977), .B(n9937), .Z(n20456) );
  OR2_X1 U5748 ( .A1(n12876), .A2(n19485), .ZN(n14341) );
  OR2_X1 U5759 ( .A1(n14335), .A2(n19485), .ZN(n20665) );
  AND2_X1 U5789 ( .A1(n20340), .A2(n382), .ZN(n20457) );
  AND2_X1 U5818 ( .A1(n20340), .A2(n382), .ZN(n20458) );
  AND2_X1 U5844 ( .A1(n20340), .A2(n382), .ZN(n12455) );
  CLKBUF_X1 U5850 ( .A(n4864), .Z(n20459) );
  XNOR2_X1 U5863 ( .A(n3984), .B(Key[62]), .ZN(n4864) );
  AND2_X1 U5868 ( .A1(n16075), .A2(n16076), .ZN(n18327) );
  XNOR2_X1 U5873 ( .A(n4059), .B(Key[127]), .ZN(n20461) );
  INV_X1 U5892 ( .A(n11686), .ZN(n20462) );
  XNOR2_X1 U5900 ( .A(n4059), .B(Key[127]), .ZN(n5052) );
  AOI22_X2 U5901 ( .A1(n15550), .A2(n15410), .B1(n15409), .B2(n15551), .ZN(
        n2973) );
  OR2_X1 U5929 ( .A1(n19174), .A2(n19170), .ZN(n18161) );
  OAI211_X1 U5942 ( .C1(n19880), .C2(n19710), .A(n8655), .B(n8654), .ZN(n10589) );
  AOI22_X1 U5961 ( .A1(n9269), .A2(n19880), .B1(n9267), .B2(n9268), .ZN(n9270)
         );
  XNOR2_X1 U5965 ( .A(n15613), .B(n15612), .ZN(n20463) );
  XNOR2_X1 U5976 ( .A(n15613), .B(n15612), .ZN(n19383) );
  OAI211_X1 U5977 ( .C1(n7779), .C2(n8312), .A(n7778), .B(n7777), .ZN(n9176)
         );
  NAND2_X2 U5993 ( .A1(n17598), .A2(n17597), .ZN(n19292) );
  XNOR2_X1 U5997 ( .A(Key[119]), .B(Plaintext[119]), .ZN(n20464) );
  XNOR2_X1 U6001 ( .A(n4465), .B(n4466), .ZN(n20465) );
  XNOR2_X1 U6027 ( .A(n4465), .B(n4466), .ZN(n8062) );
  CLKBUF_X1 U6033 ( .A(n14127), .Z(n20466) );
  AND3_X1 U6047 ( .A1(n19151), .A2(n19144), .A3(n19134), .ZN(n3141) );
  INV_X1 U6057 ( .A(n15380), .ZN(n20467) );
  BUF_X1 U6075 ( .A(n10683), .Z(n20468) );
  BUF_X1 U6076 ( .A(n13396), .Z(n20469) );
  OAI22_X1 U6091 ( .A1(n12492), .A2(n12491), .B1(n12489), .B2(n12490), .ZN(
        n13396) );
  XOR2_X1 U6117 ( .A(n9474), .B(n9473), .Z(n20470) );
  XNOR2_X1 U6146 ( .A(n13214), .B(n13213), .ZN(n20471) );
  INV_X1 U6162 ( .A(n888), .ZN(n20539) );
  INV_X1 U6167 ( .A(n8846), .ZN(n20472) );
  XNOR2_X1 U6169 ( .A(n12943), .B(n12942), .ZN(n20473) );
  BUF_X1 U6197 ( .A(n15130), .Z(n20474) );
  OAI21_X1 U6202 ( .B1(n14513), .B2(n14512), .A(n14511), .ZN(n15130) );
  AND3_X1 U6241 ( .A1(n17722), .A2(n17721), .A3(n17720), .ZN(n20475) );
  OAI211_X1 U6264 ( .C1(n11545), .C2(n10889), .A(n258), .B(n20681), .ZN(n509)
         );
  OR2_X1 U6291 ( .A1(n6904), .A2(n7903), .ZN(n19582) );
  OAI21_X1 U6299 ( .B1(n12572), .B2(n12573), .A(n12571), .ZN(n13479) );
  OR2_X1 U6309 ( .A1(n15588), .A2(n15760), .ZN(n20667) );
  BUF_X1 U6321 ( .A(n16992), .Z(n17102) );
  BUF_X1 U6354 ( .A(n9834), .Z(n20476) );
  OAI211_X1 U6365 ( .C1(n8073), .C2(n8202), .A(n20020), .B(n8072), .ZN(n9834)
         );
  NOR2_X1 U6370 ( .A1(n15215), .A2(n15214), .ZN(n20477) );
  NOR2_X1 U6371 ( .A1(n15215), .A2(n15214), .ZN(n20478) );
  NOR2_X1 U6384 ( .A1(n15215), .A2(n15214), .ZN(n17123) );
  NAND2_X1 U6403 ( .A1(n14072), .A2(n20525), .ZN(n16593) );
  XNOR2_X1 U6421 ( .A(n9097), .B(n9096), .ZN(n20479) );
  XNOR2_X1 U6425 ( .A(n9097), .B(n9096), .ZN(n10968) );
  AND2_X1 U6450 ( .A1(n20671), .A2(n1376), .ZN(n12465) );
  INV_X1 U6478 ( .A(n14228), .ZN(n20480) );
  NAND2_X1 U6503 ( .A1(n20032), .A2(n15448), .ZN(n20481) );
  NAND2_X1 U6510 ( .A1(n20032), .A2(n15448), .ZN(n16965) );
  OAI211_X1 U6521 ( .C1(n2911), .C2(n3305), .A(n3754), .B(n2910), .ZN(n20482)
         );
  OAI211_X1 U6541 ( .C1(n2911), .C2(n3305), .A(n3754), .B(n2910), .ZN(n13534)
         );
  MUX2_X1 U6566 ( .A(n7495), .B(n7494), .S(n8165), .Z(n9047) );
  AND2_X2 U6568 ( .A1(n3354), .A2(n3355), .ZN(n10030) );
  NOR2_X1 U6576 ( .A1(n8856), .A2(n8855), .ZN(n20483) );
  NOR2_X1 U6590 ( .A1(n8856), .A2(n8855), .ZN(n20484) );
  MUX2_X1 U6603 ( .A(n8854), .B(n8853), .S(n9038), .Z(n8855) );
  BUF_X1 U6622 ( .A(n8041), .Z(n20485) );
  AOI22_X1 U6623 ( .A1(n11334), .A2(n11333), .B1(n11332), .B2(n11331), .ZN(
        n20486) );
  AOI22_X1 U6629 ( .A1(n11334), .A2(n11333), .B1(n11332), .B2(n11331), .ZN(
        n12152) );
  XNOR2_X1 U6701 ( .A(Key[176]), .B(Plaintext[176]), .ZN(n20487) );
  XNOR2_X1 U6704 ( .A(n16332), .B(n16333), .ZN(n20488) );
  XNOR2_X1 U6740 ( .A(n16332), .B(n16333), .ZN(n17558) );
  NOR2_X1 U6762 ( .A1(n19418), .A2(n19439), .ZN(n20571) );
  CLKBUF_X1 U6823 ( .A(n10808), .Z(n10788) );
  NAND3_X2 U6841 ( .A1(n11700), .A2(n3783), .A3(n3780), .ZN(n13222) );
  OR2_X1 U6879 ( .A1(n12644), .A2(n12643), .ZN(n20489) );
  AND2_X2 U6925 ( .A1(n16473), .A2(n16472), .ZN(n20139) );
  XNOR2_X1 U6936 ( .A(n7245), .B(n7244), .ZN(n20490) );
  XNOR2_X1 U6944 ( .A(n7245), .B(n7244), .ZN(n7797) );
  XNOR2_X1 U6945 ( .A(n9824), .B(n10126), .ZN(n19829) );
  NAND3_X2 U7011 ( .A1(n14865), .A2(n1443), .A3(n1444), .ZN(n17339) );
  BUF_X1 U7031 ( .A(n10210), .Z(n20491) );
  INV_X1 U7038 ( .A(n12313), .ZN(n20618) );
  INV_X1 U7070 ( .A(n3305), .ZN(n20524) );
  OAI211_X1 U7156 ( .C1(n20230), .C2(n18541), .A(n17486), .B(n17485), .ZN(
        n20492) );
  OAI211_X1 U7161 ( .C1(n20230), .C2(n18541), .A(n17486), .B(n17485), .ZN(
        n18519) );
  INV_X1 U7222 ( .A(n8100), .ZN(n20493) );
  XNOR2_X1 U7226 ( .A(n17035), .B(n17270), .ZN(n20494) );
  NAND3_X2 U7227 ( .A1(n14870), .A2(n14869), .A3(n14868), .ZN(n17270) );
  OR2_X1 U7252 ( .A1(n15030), .A2(n15029), .ZN(n15033) );
  XOR2_X1 U7274 ( .A(n6533), .B(n6532), .Z(n20495) );
  XOR2_X1 U7276 ( .A(n9631), .B(n9630), .Z(n20496) );
  BUF_X1 U7309 ( .A(n12372), .Z(n20497) );
  XNOR2_X1 U7313 ( .A(n20664), .B(n13300), .ZN(n20498) );
  XNOR2_X1 U7356 ( .A(n16897), .B(n16896), .ZN(n20499) );
  XNOR2_X1 U7360 ( .A(n16897), .B(n16896), .ZN(n18978) );
  XNOR2_X1 U7361 ( .A(n2833), .B(n2832), .ZN(n20500) );
  XNOR2_X1 U7366 ( .A(n2833), .B(n2832), .ZN(n14801) );
  XNOR2_X1 U7387 ( .A(n17018), .B(n17017), .ZN(n20501) );
  INV_X1 U7404 ( .A(n15469), .ZN(n20502) );
  INV_X1 U7407 ( .A(n20502), .ZN(n20503) );
  XOR2_X1 U7408 ( .A(n4728), .B(n4729), .Z(n20504) );
  XNOR2_X1 U7410 ( .A(n15974), .B(n15973), .ZN(n20506) );
  XNOR2_X1 U7414 ( .A(n15974), .B(n15973), .ZN(n20507) );
  OR2_X1 U7430 ( .A1(n16728), .A2(n16729), .ZN(n20508) );
  MUX2_X1 U7491 ( .A(n12887), .B(n12886), .S(n14468), .Z(n15028) );
  OAI211_X1 U7498 ( .C1(n4631), .C2(n4630), .A(n4629), .B(n4628), .ZN(n20509)
         );
  INV_X1 U7517 ( .A(n19284), .ZN(n20510) );
  BUF_X1 U7538 ( .A(n19092), .Z(n19911) );
  XOR2_X1 U7580 ( .A(n6597), .B(n6596), .Z(n20511) );
  BUF_X1 U7582 ( .A(n17872), .Z(n20512) );
  XNOR2_X1 U7660 ( .A(n15983), .B(n15982), .ZN(n17872) );
  NOR2_X2 U7740 ( .A1(n129), .A2(n14291), .ZN(n15896) );
  OR2_X1 U7741 ( .A1(n19388), .A2(n19389), .ZN(n651) );
  XNOR2_X1 U7794 ( .A(n15978), .B(n15977), .ZN(n20514) );
  OAI21_X1 U7818 ( .B1(n17609), .B2(n19404), .A(n17608), .ZN(n20515) );
  OAI21_X1 U7822 ( .B1(n17609), .B2(n19404), .A(n17608), .ZN(n19302) );
  XNOR2_X1 U7823 ( .A(n8172), .B(n8173), .ZN(n20516) );
  XNOR2_X1 U7841 ( .A(n8172), .B(n8173), .ZN(n1654) );
  XNOR2_X1 U7903 ( .A(n9789), .B(n9790), .ZN(n20517) );
  XNOR2_X1 U7985 ( .A(n10795), .B(n10794), .ZN(n14781) );
  BUF_X1 U8013 ( .A(n16577), .Z(n20519) );
  MUX2_X1 U8082 ( .A(n9065), .B(n8542), .S(n9834), .Z(n8074) );
  NAND2_X1 U8111 ( .A1(n3785), .A2(n20520), .ZN(n8128) );
  NAND3_X1 U8144 ( .A1(n1452), .A2(n1453), .A3(n3784), .ZN(n20520) );
  NAND2_X1 U8170 ( .A1(n19737), .A2(n19658), .ZN(n17553) );
  AND3_X2 U8184 ( .A1(n2315), .A2(n7604), .A3(n7605), .ZN(n8941) );
  NAND2_X1 U8265 ( .A1(n11465), .A2(n1514), .ZN(n1513) );
  NAND3_X1 U8272 ( .A1(n12393), .A2(n12394), .A3(n12396), .ZN(n2539) );
  NOR2_X1 U8282 ( .A1(n12237), .A2(n20523), .ZN(n3762) );
  NAND2_X1 U8291 ( .A1(n12606), .A2(n20524), .ZN(n20523) );
  OAI21_X1 U8326 ( .B1(n14070), .B2(n15505), .A(n1758), .ZN(n20525) );
  NAND2_X1 U8337 ( .A1(n20526), .A2(n8189), .ZN(n9221) );
  OR2_X1 U8339 ( .A1(n8191), .A2(n8190), .ZN(n20526) );
  NAND3_X1 U8344 ( .A1(n5776), .A2(n5777), .A3(n1214), .ZN(n5779) );
  NAND2_X1 U8379 ( .A1(n1089), .A2(n13868), .ZN(n3034) );
  XNOR2_X1 U8391 ( .A(n20527), .B(n18209), .ZN(Ciphertext[114]) );
  NAND3_X1 U8411 ( .A1(n18207), .A2(n18206), .A3(n20528), .ZN(n20527) );
  INV_X1 U8418 ( .A(n2548), .ZN(n3074) );
  AND2_X1 U8446 ( .A1(n20529), .A2(n2548), .ZN(n7441) );
  XNOR2_X2 U8488 ( .A(n7342), .B(n7341), .ZN(n2548) );
  INV_X1 U8515 ( .A(n7585), .ZN(n20529) );
  NAND2_X1 U8524 ( .A1(n20530), .A2(n9327), .ZN(n9078) );
  OAI21_X1 U8583 ( .B1(n20008), .B2(n9333), .A(n9076), .ZN(n20530) );
  OAI211_X2 U8590 ( .C1(n3925), .C2(n4527), .A(n4525), .B(n20531), .ZN(n5765)
         );
  NAND2_X1 U8593 ( .A1(n4521), .A2(n3925), .ZN(n20531) );
  NAND2_X1 U8637 ( .A1(n2829), .A2(n19673), .ZN(n2828) );
  NAND2_X1 U8648 ( .A1(n3693), .A2(n18622), .ZN(n2829) );
  NAND3_X1 U8662 ( .A1(n1412), .A2(n15079), .A3(n20532), .ZN(n16600) );
  NAND2_X1 U8717 ( .A1(n15417), .A2(n20533), .ZN(n20532) );
  INV_X1 U8734 ( .A(n15007), .ZN(n20533) );
  XNOR2_X1 U8803 ( .A(n13817), .B(n20378), .ZN(n12286) );
  NAND2_X1 U8846 ( .A1(n18131), .A2(n18130), .ZN(n17556) );
  XNOR2_X2 U8927 ( .A(n17437), .B(n17436), .ZN(n18131) );
  NAND2_X1 U8936 ( .A1(n1567), .A2(n8676), .ZN(n8671) );
  NAND2_X1 U8969 ( .A1(n4366), .A2(n4010), .ZN(n4012) );
  XNOR2_X2 U8993 ( .A(n16703), .B(n16704), .ZN(n18966) );
  OAI21_X1 U9113 ( .B1(n19488), .B2(n14011), .A(n14611), .ZN(n14013) );
  XNOR2_X2 U9123 ( .A(n12160), .B(n12161), .ZN(n19488) );
  AND3_X2 U9130 ( .A1(n20021), .A2(n3392), .A3(n15663), .ZN(n16295) );
  OAI21_X1 U9132 ( .B1(n18051), .B2(n20535), .A(n20534), .ZN(n20052) );
  OR2_X1 U9219 ( .A1(n18052), .A2(n19989), .ZN(n20534) );
  INV_X1 U9352 ( .A(n19989), .ZN(n20535) );
  NAND3_X1 U9376 ( .A1(n20536), .A2(n7808), .A3(n8031), .ZN(n1657) );
  NAND2_X1 U9403 ( .A1(n463), .A2(n461), .ZN(n20536) );
  NAND2_X1 U9407 ( .A1(n20537), .A2(n18430), .ZN(n18435) );
  NAND2_X1 U9530 ( .A1(n3512), .A2(n18429), .ZN(n20537) );
  OAI21_X1 U9677 ( .B1(n18467), .B2(n20139), .A(n17726), .ZN(n18429) );
  OAI211_X1 U9700 ( .C1(n19505), .C2(n19719), .A(n20539), .B(n20538), .ZN(
        n2492) );
  NAND2_X1 U9701 ( .A1(n19505), .A2(n3051), .ZN(n20538) );
  AND2_X2 U9754 ( .A1(n20541), .A2(n20540), .ZN(n16963) );
  NAND2_X1 U9757 ( .A1(n2279), .A2(n15687), .ZN(n20540) );
  NAND2_X1 U9765 ( .A1(n20542), .A2(n15454), .ZN(n20541) );
  NAND2_X1 U9789 ( .A1(n15450), .A2(n15451), .ZN(n20542) );
  NAND3_X1 U9812 ( .A1(n8703), .A2(n8155), .A3(n9567), .ZN(n8170) );
  NAND2_X1 U10002 ( .A1(n14260), .A2(n19652), .ZN(n14265) );
  NAND2_X1 U10005 ( .A1(n9053), .A2(n1752), .ZN(n1750) );
  NAND2_X1 U10058 ( .A1(n20544), .A2(n20543), .ZN(n13103) );
  NAND2_X1 U10095 ( .A1(n20626), .A2(n12593), .ZN(n20544) );
  NAND2_X1 U10102 ( .A1(n18341), .A2(n18344), .ZN(n18290) );
  NAND2_X1 U10218 ( .A1(n12060), .A2(n563), .ZN(n12064) );
  NAND2_X1 U10291 ( .A1(n20371), .A2(n20545), .ZN(n14221) );
  NOR2_X1 U10402 ( .A1(n15408), .A2(n15546), .ZN(n20545) );
  NAND2_X1 U10473 ( .A1(n8540), .A2(n2173), .ZN(n10604) );
  NAND2_X1 U10488 ( .A1(n14280), .A2(n14281), .ZN(n14282) );
  NAND2_X1 U10767 ( .A1(n14555), .A2(n14556), .ZN(n14281) );
  INV_X1 U10835 ( .A(n5648), .ZN(n5650) );
  NAND2_X1 U10848 ( .A1(n5443), .A2(n5643), .ZN(n5648) );
  INV_X1 U10888 ( .A(n8537), .ZN(n8539) );
  NAND2_X1 U10912 ( .A1(n8866), .A2(n9326), .ZN(n8537) );
  NAND2_X1 U11051 ( .A1(n13273), .A2(n20546), .ZN(n13276) );
  INV_X1 U11166 ( .A(n20547), .ZN(n20546) );
  OAI21_X1 U11200 ( .B1(n13274), .B2(n13275), .A(n13272), .ZN(n20547) );
  NAND2_X1 U11269 ( .A1(n900), .A2(n20548), .ZN(n1584) );
  NAND2_X1 U11270 ( .A1(n8245), .A2(n8251), .ZN(n20548) );
  NAND2_X1 U11356 ( .A1(n2018), .A2(n2019), .ZN(n20549) );
  NAND2_X1 U11363 ( .A1(n20072), .A2(n17507), .ZN(n1899) );
  NAND3_X1 U11425 ( .A1(n15042), .A2(n942), .A3(n15567), .ZN(n1177) );
  AND2_X1 U11434 ( .A1(n888), .A2(n11491), .ZN(n11070) );
  NAND2_X1 U11447 ( .A1(n16211), .A2(n20550), .ZN(n17729) );
  NAND2_X1 U11448 ( .A1(n17163), .A2(n17565), .ZN(n20550) );
  OAI22_X1 U11487 ( .A1(n18502), .A2(n18501), .B1(n18499), .B2(n18500), .ZN(
        n1843) );
  NOR2_X1 U11508 ( .A1(n15400), .A2(n15898), .ZN(n15891) );
  NAND3_X1 U11520 ( .A1(n4251), .A2(n19539), .A3(n4250), .ZN(n99) );
  XNOR2_X1 U11522 ( .A(n20552), .B(n20551), .ZN(n7210) );
  NAND2_X1 U11524 ( .A1(n3528), .A2(n20553), .ZN(n20552) );
  NAND3_X1 U11538 ( .A1(n8947), .A2(n8730), .A3(n8940), .ZN(n20614) );
  AND2_X2 U11595 ( .A1(n2319), .A2(n2360), .ZN(n12095) );
  OR2_X1 U11617 ( .A1(n8129), .A2(n1507), .ZN(n8563) );
  OR2_X1 U11663 ( .A1(n11035), .A2(n10783), .ZN(n11437) );
  OAI21_X1 U11693 ( .B1(n14598), .B2(n14395), .A(n14596), .ZN(n3757) );
  NAND2_X1 U11694 ( .A1(n14154), .A2(n14393), .ZN(n14596) );
  NAND2_X1 U11755 ( .A1(n19652), .A2(n14261), .ZN(n14543) );
  NAND2_X1 U11788 ( .A1(n19404), .A2(n16306), .ZN(n17607) );
  NAND3_X1 U11790 ( .A1(n20306), .A2(n20307), .A3(n17688), .ZN(n19034) );
  XNOR2_X1 U11792 ( .A(n20556), .B(n20555), .ZN(Ciphertext[70]) );
  INV_X1 U11873 ( .A(n17989), .ZN(n20555) );
  NAND3_X1 U11923 ( .A1(n17988), .A2(n3829), .A3(n17987), .ZN(n20556) );
  NAND2_X1 U11924 ( .A1(n15110), .A2(n14461), .ZN(n15292) );
  NOR2_X2 U11980 ( .A1(n14471), .A2(n14470), .ZN(n15110) );
  NAND2_X1 U11993 ( .A1(n6950), .A2(n2961), .ZN(n9164) );
  NAND2_X1 U12032 ( .A1(n8609), .A2(n8696), .ZN(n8610) );
  AND2_X2 U12052 ( .A1(n2390), .A2(n2391), .ZN(n14461) );
  NAND2_X1 U12084 ( .A1(n8372), .A2(n8370), .ZN(n7705) );
  NAND3_X1 U12099 ( .A1(n8883), .A2(n8881), .A3(n8882), .ZN(n20690) );
  XNOR2_X2 U12104 ( .A(n20558), .B(n20557), .ZN(n11231) );
  XNOR2_X1 U12109 ( .A(n9880), .B(n10580), .ZN(n20557) );
  XNOR2_X1 U12115 ( .A(n10004), .B(n9877), .ZN(n20558) );
  NAND3_X1 U12116 ( .A1(n20559), .A2(n8557), .A3(n8558), .ZN(n1186) );
  NAND2_X1 U12128 ( .A1(n8556), .A2(n9107), .ZN(n20559) );
  NAND2_X1 U12146 ( .A1(n6133), .A2(n5691), .ZN(n5692) );
  OAI21_X1 U12191 ( .B1(n259), .B2(n20560), .A(n20640), .ZN(n11517) );
  NAND2_X1 U12195 ( .A1(n10722), .A2(n20561), .ZN(n12648) );
  NAND2_X1 U12198 ( .A1(n9319), .A2(n1855), .ZN(n9323) );
  OAI21_X1 U12254 ( .B1(n15649), .B2(n15257), .A(n20562), .ZN(n14583) );
  NAND3_X1 U12261 ( .A1(n15257), .A2(n15831), .A3(n20563), .ZN(n20562) );
  INV_X1 U12307 ( .A(n15643), .ZN(n20563) );
  AOI22_X1 U12308 ( .A1(n20594), .A2(n7608), .B1(n8730), .B2(n8729), .ZN(n7612) );
  INV_X1 U12312 ( .A(n5666), .ZN(n20616) );
  NAND2_X1 U12375 ( .A1(n17699), .A2(n18928), .ZN(n1921) );
  NAND2_X1 U12376 ( .A1(n20564), .A2(n19534), .ZN(n19627) );
  NAND2_X1 U12388 ( .A1(n19288), .A2(n19304), .ZN(n20564) );
  NAND2_X1 U12409 ( .A1(n15246), .A2(n20565), .ZN(n15247) );
  NAND3_X2 U12419 ( .A1(n5499), .A2(n20567), .A3(n20566), .ZN(n7230) );
  NAND2_X1 U12465 ( .A1(n1353), .A2(n5498), .ZN(n20566) );
  NAND2_X1 U12528 ( .A1(n5496), .A2(n20568), .ZN(n20567) );
  NAND3_X1 U12609 ( .A1(n15568), .A2(n20569), .A3(n20428), .ZN(n15570) );
  NAND2_X1 U12721 ( .A1(n15565), .A2(n15804), .ZN(n20569) );
  NAND2_X1 U12737 ( .A1(n3712), .A2(n3713), .ZN(n11222) );
  AND2_X2 U12878 ( .A1(n20570), .A2(n3646), .ZN(n13624) );
  NAND2_X1 U12880 ( .A1(n2804), .A2(n3649), .ZN(n20570) );
  OAI21_X1 U12885 ( .B1(n20382), .B2(n20571), .A(n19434), .ZN(n20316) );
  NAND2_X1 U12989 ( .A1(n20574), .A2(n20572), .ZN(n19378) );
  NAND2_X1 U12993 ( .A1(n20573), .A2(n19375), .ZN(n20572) );
  NAND2_X1 U13100 ( .A1(n19374), .A2(n19733), .ZN(n20573) );
  NAND2_X1 U13172 ( .A1(n19377), .A2(n19666), .ZN(n20574) );
  OR2_X1 U13410 ( .A1(n15453), .A2(n19978), .ZN(n15786) );
  NAND3_X1 U13512 ( .A1(n1329), .A2(n1327), .A3(n20575), .ZN(n12543) );
  NAND3_X1 U13541 ( .A1(n20660), .A2(n764), .A3(n11383), .ZN(n20575) );
  XNOR2_X1 U13585 ( .A(n20576), .B(n2395), .ZN(Ciphertext[170]) );
  NAND3_X1 U13588 ( .A1(n18166), .A2(n2226), .A3(n2227), .ZN(n20576) );
  NAND2_X1 U13698 ( .A1(n19881), .A2(n8375), .ZN(n6733) );
  NAND2_X1 U13723 ( .A1(n20577), .A2(n12098), .ZN(n13065) );
  NOR2_X1 U13754 ( .A1(n20579), .A2(n20578), .ZN(n20577) );
  NOR2_X1 U13758 ( .A1(n12428), .A2(n3649), .ZN(n20578) );
  INV_X1 U13777 ( .A(n12097), .ZN(n20579) );
  NOR2_X1 U13810 ( .A1(n13742), .A2(n13743), .ZN(n15677) );
  NAND2_X1 U13863 ( .A1(n18653), .A2(n18654), .ZN(n20580) );
  NAND2_X1 U13868 ( .A1(n18655), .A2(n18656), .ZN(n20581) );
  XNOR2_X1 U13885 ( .A(n20582), .B(n18148), .ZN(Ciphertext[59]) );
  NAND4_X1 U13934 ( .A1(n20629), .A2(n2830), .A3(n2828), .A4(n18147), .ZN(
        n20582) );
  NAND2_X1 U13936 ( .A1(n9529), .A2(n9528), .ZN(n9527) );
  NAND2_X1 U14000 ( .A1(n8721), .A2(n9357), .ZN(n9529) );
  NAND2_X1 U14001 ( .A1(n19511), .A2(n19395), .ZN(n19631) );
  NAND3_X1 U14021 ( .A1(n1459), .A2(n3104), .A3(n20583), .ZN(n12047) );
  OAI21_X1 U14064 ( .B1(n20585), .B2(n20584), .A(n585), .ZN(n20035) );
  OAI21_X1 U14073 ( .B1(n11282), .B2(n11281), .A(n20641), .ZN(n1498) );
  NAND3_X1 U14075 ( .A1(n18319), .A2(n19174), .A3(n1035), .ZN(n18322) );
  NAND2_X1 U14246 ( .A1(n88), .A2(n8075), .ZN(n10552) );
  OR2_X1 U14262 ( .A1(n19185), .A2(n20642), .ZN(n19186) );
  NAND2_X1 U14342 ( .A1(n20586), .A2(n8209), .ZN(n7434) );
  NAND2_X1 U14346 ( .A1(n9006), .A2(n8890), .ZN(n1672) );
  NAND2_X1 U14391 ( .A1(n20589), .A2(n20587), .ZN(n7997) );
  NAND2_X1 U14415 ( .A1(n7989), .A2(n20588), .ZN(n20587) );
  INV_X1 U14446 ( .A(n8705), .ZN(n20588) );
  NAND2_X1 U14482 ( .A1(n7988), .A2(n8705), .ZN(n20589) );
  NAND3_X2 U14497 ( .A1(n15542), .A2(n15541), .A3(n20379), .ZN(n16181) );
  OAI21_X1 U14530 ( .B1(n11187), .B2(n20591), .A(n20590), .ZN(n11196) );
  NAND2_X1 U14562 ( .A1(n11189), .A2(n19983), .ZN(n20590) );
  NAND2_X1 U14563 ( .A1(n20592), .A2(n2981), .ZN(n2980) );
  NAND2_X1 U14589 ( .A1(n18145), .A2(n18641), .ZN(n20592) );
  NAND3_X1 U14716 ( .A1(n6051), .A2(n6052), .A3(n6050), .ZN(n6053) );
  NAND2_X1 U14717 ( .A1(n11637), .A2(n20430), .ZN(n11979) );
  NAND2_X1 U14724 ( .A1(n19879), .A2(n15666), .ZN(n15771) );
  NAND2_X1 U14728 ( .A1(n722), .A2(n723), .ZN(n721) );
  NOR2_X1 U14823 ( .A1(n317), .A2(n8945), .ZN(n20594) );
  OR2_X1 U14826 ( .A1(n11528), .A2(n11526), .ZN(n20279) );
  NAND2_X1 U14878 ( .A1(n10863), .A2(n11387), .ZN(n10867) );
  OAI211_X1 U14890 ( .C1(n11544), .C2(n11549), .A(n20595), .B(n11550), .ZN(
        n10762) );
  NAND2_X1 U15069 ( .A1(n11544), .A2(n10926), .ZN(n20595) );
  NAND2_X1 U15088 ( .A1(n20596), .A2(n8057), .ZN(n2750) );
  OAI211_X1 U15131 ( .C1(n8054), .C2(n19802), .A(n3472), .B(n8052), .ZN(n20596) );
  XNOR2_X2 U15133 ( .A(n20598), .B(n20597), .ZN(n11546) );
  XNOR2_X1 U15134 ( .A(n9261), .B(n8635), .ZN(n20597) );
  XNOR2_X1 U15174 ( .A(n8627), .B(n9508), .ZN(n20598) );
  NAND3_X1 U15203 ( .A1(n1232), .A2(n4814), .A3(n5069), .ZN(n19612) );
  NAND2_X1 U15294 ( .A1(n20600), .A2(n20599), .ZN(n10991) );
  NAND2_X1 U15314 ( .A1(n11870), .A2(n11390), .ZN(n20599) );
  NAND2_X1 U15325 ( .A1(n20160), .A2(n20601), .ZN(n20600) );
  INV_X1 U15369 ( .A(n11389), .ZN(n20601) );
  NAND2_X1 U15370 ( .A1(n16659), .A2(n1115), .ZN(n16661) );
  NAND2_X1 U15399 ( .A1(n10653), .A2(n20375), .ZN(n11602) );
  NAND2_X1 U15546 ( .A1(n19679), .A2(n19757), .ZN(n18216) );
  OAI21_X1 U15576 ( .B1(n16780), .B2(n19143), .A(n20602), .ZN(n17810) );
  NAND2_X1 U15621 ( .A1(n16780), .A2(n19135), .ZN(n20602) );
  NAND2_X1 U15669 ( .A1(n5141), .A2(n20603), .ZN(n5143) );
  NAND3_X1 U15717 ( .A1(n6054), .A2(n5139), .A3(n5559), .ZN(n20603) );
  OAI21_X1 U15726 ( .B1(n12184), .B2(n12185), .A(n20604), .ZN(n12745) );
  NAND2_X1 U15731 ( .A1(n20201), .A2(n12181), .ZN(n20604) );
  NAND3_X1 U15776 ( .A1(n9169), .A2(n9170), .A3(n1211), .ZN(n10329) );
  XNOR2_X1 U15778 ( .A(n20605), .B(n2193), .ZN(Ciphertext[126]) );
  NAND3_X1 U15795 ( .A1(n2196), .A2(n2197), .A3(n2195), .ZN(n20605) );
  AOI22_X1 U15802 ( .A1(n12066), .A2(n12213), .B1(n12210), .B2(n12189), .ZN(
        n12068) );
  NAND2_X1 U15807 ( .A1(n236), .A2(n20451), .ZN(n14412) );
  NAND3_X1 U15812 ( .A1(n20645), .A2(n4384), .A3(n20606), .ZN(n3684) );
  NAND2_X1 U15857 ( .A1(n905), .A2(n8741), .ZN(n8951) );
  OR2_X1 U15947 ( .A1(n7629), .A2(n7630), .ZN(n905) );
  NAND2_X1 U15982 ( .A1(n14285), .A2(n20607), .ZN(n1437) );
  NOR2_X1 U16003 ( .A1(n14296), .A2(n15898), .ZN(n20607) );
  NAND3_X1 U16004 ( .A1(n8929), .A2(n8931), .A3(n8933), .ZN(n8935) );
  XNOR2_X1 U16082 ( .A(n9792), .B(n20608), .ZN(n9796) );
  NAND2_X1 U16095 ( .A1(n11632), .A2(n11633), .ZN(n12616) );
  NOR2_X1 U16096 ( .A1(n20040), .A2(n14817), .ZN(n20609) );
  OAI211_X1 U16101 ( .C1(n20437), .C2(n20361), .A(n18384), .B(n20610), .ZN(
        n595) );
  NAND2_X1 U16102 ( .A1(n20361), .A2(n20611), .ZN(n20610) );
  NAND3_X1 U16110 ( .A1(n4641), .A2(n4646), .A3(n4647), .ZN(n4148) );
  NAND2_X1 U16122 ( .A1(n18028), .A2(n18931), .ZN(n20612) );
  NAND2_X1 U16123 ( .A1(n18027), .A2(n20207), .ZN(n20613) );
  NAND2_X1 U16134 ( .A1(n20614), .A2(n318), .ZN(n8948) );
  OR2_X1 U16137 ( .A1(n5116), .A2(n5115), .ZN(n1914) );
  NAND2_X1 U16155 ( .A1(n1575), .A2(n9452), .ZN(n8885) );
  NAND2_X1 U16185 ( .A1(n5665), .A2(n20615), .ZN(n6735) );
  NAND2_X1 U16203 ( .A1(n20616), .A2(n5661), .ZN(n20615) );
  NAND2_X2 U16269 ( .A1(n20617), .A2(n3758), .ZN(n15275) );
  NAND2_X1 U16277 ( .A1(n3757), .A2(n14394), .ZN(n20617) );
  NAND2_X1 U16278 ( .A1(n12153), .A2(n20486), .ZN(n12149) );
  NAND3_X1 U16313 ( .A1(n2437), .A2(n15444), .A3(n2438), .ZN(n20032) );
  OAI211_X2 U16318 ( .C1(n20235), .C2(n9612), .A(n20620), .B(n20619), .ZN(
        n11951) );
  NAND2_X1 U16348 ( .A1(n9609), .A2(n11292), .ZN(n20619) );
  NAND2_X1 U16350 ( .A1(n9610), .A2(n11404), .ZN(n20620) );
  NAND3_X1 U16351 ( .A1(n20621), .A2(n15226), .A3(n15779), .ZN(n14870) );
  NAND2_X1 U16365 ( .A1(n15685), .A2(n15783), .ZN(n20621) );
  OR2_X1 U16366 ( .A1(n7952), .A2(n7481), .ZN(n7814) );
  AOI22_X2 U16381 ( .A1(n19387), .A2(n19386), .B1(n19385), .B2(n19384), .ZN(
        n19442) );
  NOR2_X1 U16408 ( .A1(n11903), .A2(n12148), .ZN(n11904) );
  NOR2_X2 U16409 ( .A1(n11345), .A2(n11344), .ZN(n12148) );
  NAND2_X1 U16410 ( .A1(n3451), .A2(n5074), .ZN(n4459) );
  NAND2_X1 U16423 ( .A1(n3270), .A2(n3272), .ZN(n447) );
  AND2_X2 U16476 ( .A1(n20623), .A2(n20622), .ZN(n13321) );
  NAND2_X1 U16560 ( .A1(n11063), .A2(n12267), .ZN(n20622) );
  NAND2_X1 U16566 ( .A1(n9059), .A2(n9031), .ZN(n8573) );
  NAND3_X1 U16580 ( .A1(n18749), .A2(n18711), .A3(n18773), .ZN(n18712) );
  NAND2_X1 U16596 ( .A1(n8712), .A2(n9233), .ZN(n8412) );
  NOR2_X1 U16601 ( .A1(n19716), .A2(n9234), .ZN(n8712) );
  NAND2_X1 U16640 ( .A1(n20625), .A2(n1929), .ZN(n10567) );
  OAI22_X1 U16645 ( .A1(n8673), .A2(n8674), .B1(n9021), .B2(n8676), .ZN(n20625) );
  NOR2_X2 U16681 ( .A1(n9184), .A2(n9185), .ZN(n10571) );
  NAND2_X1 U16687 ( .A1(n11979), .A2(n11978), .ZN(n20626) );
  AOI22_X2 U16707 ( .A1(n8759), .A2(n9273), .B1(n20627), .B2(n8991), .ZN(n9894) );
  OAI21_X1 U16708 ( .B1(n9277), .B2(n9275), .A(n19732), .ZN(n20627) );
  NAND2_X1 U16709 ( .A1(n20628), .A2(n2294), .ZN(n6942) );
  NAND2_X1 U16725 ( .A1(n3700), .A2(n5751), .ZN(n20628) );
  NAND2_X1 U16726 ( .A1(n20039), .A2(n2829), .ZN(n20629) );
  NAND2_X1 U16764 ( .A1(n12065), .A2(n12211), .ZN(n11814) );
  OAI211_X2 U16766 ( .C1(n5980), .C2(n5155), .A(n5153), .B(n20630), .ZN(n7232)
         );
  NAND2_X1 U16771 ( .A1(n3767), .A2(n6075), .ZN(n20630) );
  XNOR2_X1 U16778 ( .A(n20631), .B(n18316), .ZN(Ciphertext[177]) );
  NAND2_X1 U17000 ( .A1(n18315), .A2(n20632), .ZN(n20631) );
  AND2_X1 U17016 ( .A1(n18314), .A2(n18313), .ZN(n20632) );
  NAND2_X1 U17017 ( .A1(n20634), .A2(n20633), .ZN(n15026) );
  XNOR2_X2 U17111 ( .A(n14971), .B(n14970), .ZN(n17208) );
  NAND2_X1 U17192 ( .A1(n16465), .A2(n17210), .ZN(n20634) );
  AND3_X2 U17193 ( .A1(n10762), .A2(n10763), .A3(n10764), .ZN(n12389) );
  INV_X1 U17194 ( .A(Plaintext[56]), .ZN(n20635) );
  NAND2_X1 U17198 ( .A1(n14515), .A2(n20636), .ZN(n15125) );
  OAI22_X1 U17239 ( .A1(n7861), .A2(n8083), .B1(n20638), .B2(n20637), .ZN(
        n1159) );
  INV_X1 U17265 ( .A(n20495), .ZN(n20637) );
  NAND2_X1 U17341 ( .A1(n6539), .A2(n20108), .ZN(n20638) );
  NAND3_X1 U17392 ( .A1(n20640), .A2(n10936), .A3(n20639), .ZN(n725) );
  INV_X1 U17396 ( .A(n11573), .ZN(n20639) );
  INV_X1 U17431 ( .A(n20106), .ZN(n20640) );
  NAND2_X1 U17432 ( .A1(n14624), .A2(n14627), .ZN(n13856) );
  NAND2_X1 U17498 ( .A1(n15474), .A2(n12659), .ZN(n12662) );
  NOR2_X1 U17514 ( .A1(n19183), .A2(n19212), .ZN(n20642) );
  XNOR2_X1 U17568 ( .A(n20643), .B(n18717), .ZN(Ciphertext[78]) );
  NAND4_X1 U17659 ( .A1(n18714), .A2(n18713), .A3(n18715), .A4(n18712), .ZN(
        n20643) );
  XNOR2_X1 U17662 ( .A(n13138), .B(n13339), .ZN(n13139) );
  AOI21_X2 U17686 ( .B1(n11696), .B2(n12399), .A(n20644), .ZN(n13339) );
  OAI211_X2 U17749 ( .C1(n14753), .C2(n14430), .A(n14428), .B(n14429), .ZN(
        n15296) );
  NAND2_X1 U17750 ( .A1(n4480), .A2(n3967), .ZN(n20645) );
  NAND2_X1 U17751 ( .A1(n12473), .A2(n19833), .ZN(n12484) );
  NAND2_X1 U17793 ( .A1(n20058), .A2(n20060), .ZN(n19492) );
  XNOR2_X1 U17800 ( .A(n20664), .B(n13300), .ZN(n14707) );
  NOR2_X1 U17833 ( .A1(n15679), .A2(n20647), .ZN(n15231) );
  INV_X1 U18067 ( .A(n16165), .ZN(n20648) );
  NAND2_X1 U18128 ( .A1(n17498), .A2(n15485), .ZN(n16795) );
  XNOR2_X2 U18308 ( .A(n10440), .B(n10439), .ZN(n11445) );
  NAND2_X1 U18337 ( .A1(n343), .A2(n6097), .ZN(n20649) );
  NAND2_X1 U18353 ( .A1(n20689), .A2(n789), .ZN(n787) );
  NAND3_X1 U18386 ( .A1(n138), .A2(n1775), .A3(n1772), .ZN(n137) );
  NAND3_X1 U18392 ( .A1(n267), .A2(n266), .A3(n9242), .ZN(n3288) );
  OAI211_X2 U18394 ( .C1(n8431), .C2(n9218), .A(n8429), .B(n8430), .ZN(n10072)
         );
  NAND3_X1 U18401 ( .A1(n7587), .A2(n7588), .A3(n20650), .ZN(n8644) );
  NAND2_X1 U18459 ( .A1(n20373), .A2(n20651), .ZN(n20650) );
  NAND2_X1 U18476 ( .A1(n7603), .A2(n7795), .ZN(n7605) );
  NAND2_X1 U18482 ( .A1(n19403), .A2(n19402), .ZN(n17649) );
  OAI211_X2 U18490 ( .C1(n15890), .C2(n14913), .A(n14911), .B(n20652), .ZN(
        n17378) );
  NAND2_X1 U18555 ( .A1(n15890), .A2(n20006), .ZN(n20652) );
  NAND3_X1 U18633 ( .A1(n14666), .A2(n14535), .A3(n14662), .ZN(n14313) );
  XNOR2_X2 U18634 ( .A(n13177), .B(n13176), .ZN(n14662) );
  NAND2_X1 U18636 ( .A1(n20367), .A2(n7953), .ZN(n7818) );
  NAND2_X1 U18655 ( .A1(n14623), .A2(n14626), .ZN(n14625) );
  NAND3_X1 U18683 ( .A1(n20653), .A2(n12919), .A3(n14443), .ZN(n2775) );
  NAND2_X1 U18684 ( .A1(n14439), .A2(n14168), .ZN(n20653) );
  INV_X1 U18698 ( .A(n18500), .ZN(n17737) );
  NAND2_X2 U18706 ( .A1(n816), .A2(n20654), .ZN(n18500) );
  NAND2_X1 U18751 ( .A1(n4422), .A2(n20655), .ZN(n6119) );
  NAND2_X1 U18766 ( .A1(n12129), .A2(n11586), .ZN(n699) );
  NAND2_X1 U18778 ( .A1(n3487), .A2(n3488), .ZN(n12129) );
  OR2_X1 U18827 ( .A1(n6138), .A2(n5859), .ZN(n20333) );
  OAI21_X1 U18829 ( .B1(n7836), .B2(n7958), .A(n20656), .ZN(n8911) );
  NAND2_X1 U18830 ( .A1(n20165), .A2(n7836), .ZN(n20656) );
  AOI21_X1 U18853 ( .B1(n5900), .B2(n6087), .A(n5908), .ZN(n1466) );
  OAI22_X2 U18899 ( .A1(n1164), .A2(n7283), .B1(n7812), .B2(n7811), .ZN(n8890)
         );
  NAND2_X1 U18932 ( .A1(n6155), .A2(n5612), .ZN(n5610) );
  OAI211_X2 U18935 ( .C1(n7992), .C2(n8015), .A(n20657), .B(n7472), .ZN(n8813)
         );
  NAND2_X1 U18944 ( .A1(n3243), .A2(n7994), .ZN(n20657) );
  NAND2_X1 U18959 ( .A1(n1902), .A2(n2970), .ZN(n12036) );
  NAND2_X1 U18962 ( .A1(n14572), .A2(n14573), .ZN(n14741) );
  AND2_X2 U19077 ( .A1(n20658), .A2(n3672), .ZN(n6410) );
  NAND2_X1 U19087 ( .A1(n4502), .A2(n3674), .ZN(n20658) );
  NAND2_X1 U19088 ( .A1(n8734), .A2(n8923), .ZN(n8498) );
  NAND2_X1 U19109 ( .A1(n45), .A2(n44), .ZN(n8) );
  AND3_X2 U19125 ( .A1(n15833), .A2(n15834), .A3(n15835), .ZN(n16975) );
  NAND3_X1 U19126 ( .A1(n19911), .A2(n17529), .A3(n20661), .ZN(n17532) );
  NAND2_X1 U19128 ( .A1(n4147), .A2(n4148), .ZN(n4149) );
  NAND3_X1 U19209 ( .A1(n2492), .A2(n20663), .A3(n20662), .ZN(n12513) );
  NAND2_X1 U19398 ( .A1(n10623), .A2(n888), .ZN(n20662) );
  NAND2_X1 U19406 ( .A1(n3814), .A2(n913), .ZN(n20663) );
  OAI22_X1 U19407 ( .A1(n11911), .A2(n12812), .B1(n11912), .B2(n12490), .ZN(
        n11913) );
  NAND2_X1 U19474 ( .A1(n3586), .A2(n12807), .ZN(n11911) );
  XNOR2_X1 U19487 ( .A(n6563), .B(n7117), .ZN(n3570) );
  INV_X1 U19518 ( .A(n16465), .ZN(n16660) );
  XNOR2_X2 U19519 ( .A(n14995), .B(n14994), .ZN(n16465) );
  NOR2_X2 U19520 ( .A1(n14445), .A2(n1722), .ZN(n15294) );
  INV_X1 U19542 ( .A(n14998), .ZN(n15832) );
  NAND2_X1 U19543 ( .A1(n15828), .A2(n19891), .ZN(n14998) );
  XNOR2_X1 U19544 ( .A(n13463), .B(n13298), .ZN(n20664) );
  NAND3_X1 U19589 ( .A1(n14339), .A2(n14049), .A3(n20665), .ZN(n12802) );
  NAND2_X1 U19601 ( .A1(n14335), .A2(n13930), .ZN(n14049) );
  NAND2_X1 U19605 ( .A1(n15469), .A2(n15465), .ZN(n15340) );
  NAND2_X1 U19625 ( .A1(n20666), .A2(n8869), .ZN(n8465) );
  NAND2_X1 U19626 ( .A1(n9326), .A2(n9076), .ZN(n20666) );
  AOI22_X2 U19655 ( .A1(n2109), .A2(n15343), .B1(n15342), .B2(n19888), .ZN(
        n19889) );
  NAND2_X1 U19675 ( .A1(n1507), .A2(n20010), .ZN(n1652) );
  NOR2_X2 U19684 ( .A1(n6320), .A2(n6319), .ZN(n20010) );
  NAND2_X1 U19703 ( .A1(n15990), .A2(n20667), .ZN(n15591) );
  NAND3_X1 U19704 ( .A1(n1469), .A2(n13959), .A3(n13960), .ZN(n20119) );
  NAND2_X1 U19713 ( .A1(n14666), .A2(n14663), .ZN(n14314) );
  NAND3_X1 U19744 ( .A1(n6055), .A2(n20669), .A3(n20668), .ZN(n385) );
  NAND2_X1 U19750 ( .A1(n6057), .A2(n5891), .ZN(n20668) );
  NAND2_X1 U19767 ( .A1(n906), .A2(n20670), .ZN(n20669) );
  INV_X1 U19777 ( .A(n5304), .ZN(n20670) );
  NAND2_X1 U19790 ( .A1(n20358), .A2(n7932), .ZN(n7760) );
  NAND2_X1 U19794 ( .A1(n12507), .A2(n12506), .ZN(n1609) );
  NAND3_X1 U19806 ( .A1(n11019), .A2(n11020), .A3(n12500), .ZN(n11021) );
  NAND3_X1 U19807 ( .A1(n20299), .A2(n1378), .A3(n20300), .ZN(n20671) );
  AND2_X2 U19819 ( .A1(n20683), .A2(n20684), .ZN(n9039) );
  NAND2_X1 U19823 ( .A1(n5623), .A2(n6129), .ZN(n1770) );
  AOI21_X2 U19825 ( .B1(n4279), .B2(n3682), .A(n19559), .ZN(n5623) );
  OAI21_X1 U19828 ( .B1(n20674), .B2(n5525), .A(n20673), .ZN(n1170) );
  INV_X1 U19835 ( .A(n5294), .ZN(n20673) );
  NAND2_X1 U19840 ( .A1(n19201), .A2(n19842), .ZN(n19193) );
  NAND2_X1 U19845 ( .A1(n20675), .A2(n11326), .ZN(n11709) );
  OAI21_X1 U19856 ( .B1(n1124), .B2(n191), .A(n1122), .ZN(n20675) );
  NAND2_X1 U19858 ( .A1(n2246), .A2(n66), .ZN(n2814) );
  INV_X1 U19859 ( .A(n20676), .ZN(n19974) );
  XNOR2_X1 U19860 ( .A(n17415), .B(n17414), .ZN(n20676) );
  AND3_X2 U19861 ( .A1(n15528), .A2(n1337), .A3(n16443), .ZN(n15529) );
  NAND3_X1 U19862 ( .A1(n4736), .A2(n3903), .A3(n4737), .ZN(n3905) );
  NAND2_X1 U19863 ( .A1(n679), .A2(n2049), .ZN(n678) );
  NAND2_X1 U19864 ( .A1(n3031), .A2(n18869), .ZN(n679) );
  XNOR2_X2 U19865 ( .A(n7387), .B(n7388), .ZN(n8289) );
  NOR2_X2 U19866 ( .A1(n11084), .A2(n11085), .ZN(n13147) );
  INV_X1 U19867 ( .A(n20677), .ZN(n1894) );
  OAI21_X1 U19868 ( .B1(n6037), .B2(n6036), .A(n6035), .ZN(n20677) );
  NAND3_X1 U19869 ( .A1(n2166), .A2(n1416), .A3(n2165), .ZN(n8833) );
  NAND2_X1 U19870 ( .A1(n1642), .A2(n420), .ZN(n14735) );
  NAND2_X1 U19871 ( .A1(n4460), .A2(n20431), .ZN(n3189) );
  NAND2_X1 U19872 ( .A1(n14742), .A2(n14743), .ZN(n14745) );
  AOI21_X1 U19873 ( .B1(n20678), .B2(n7920), .A(n7768), .ZN(n6320) );
  NAND2_X1 U19874 ( .A1(n6299), .A2(n505), .ZN(n20678) );
  NAND2_X1 U19875 ( .A1(n19301), .A2(n20515), .ZN(n19303) );
  OAI21_X1 U19876 ( .B1(n20381), .B2(n14501), .A(n20680), .ZN(n14504) );
  NAND2_X1 U19877 ( .A1(n14502), .A2(n14501), .ZN(n20680) );
  OR2_X1 U19878 ( .A1(n11546), .A2(n10761), .ZN(n20681) );
  INV_X1 U19879 ( .A(n4043), .ZN(n1442) );
  NAND3_X1 U19880 ( .A1(n4042), .A2(n713), .A3(n5034), .ZN(n4043) );
  NAND2_X1 U19881 ( .A1(n9039), .A2(n8851), .ZN(n9045) );
  NAND2_X1 U19882 ( .A1(n7402), .A2(n7171), .ZN(n20683) );
  NAND2_X1 U19883 ( .A1(n7170), .A2(n7814), .ZN(n20684) );
  NAND3_X1 U19884 ( .A1(n20685), .A2(n2116), .A3(n8984), .ZN(n1157) );
  NAND2_X1 U19885 ( .A1(n9267), .A2(n2118), .ZN(n20685) );
  OAI211_X2 U19886 ( .C1(n9051), .C2(n9289), .A(n20686), .B(n839), .ZN(n9824)
         );
  NAND2_X1 U19887 ( .A1(n736), .A2(n19896), .ZN(n20686) );
  NAND2_X1 U19888 ( .A1(n2102), .A2(n2103), .ZN(n2101) );
  XNOR2_X1 U19889 ( .A(n20687), .B(n19273), .ZN(Ciphertext[166]) );
  NAND3_X1 U19890 ( .A1(n2262), .A2(n2261), .A3(n19272), .ZN(n20687) );
  NAND2_X1 U19891 ( .A1(n6049), .A2(n6048), .ZN(n2641) );
  OAI211_X2 U19892 ( .C1(n4509), .C2(n4574), .A(n3909), .B(n3910), .ZN(n6048)
         );
  NAND2_X2 U19893 ( .A1(n12459), .A2(n12460), .ZN(n12137) );
  NAND2_X1 U19894 ( .A1(n1943), .A2(n1944), .ZN(n12459) );
  NAND2_X1 U19895 ( .A1(n17968), .A2(n19943), .ZN(n2951) );
  NAND2_X1 U19896 ( .A1(n17558), .A2(n18114), .ZN(n17968) );
  NAND2_X1 U19897 ( .A1(n20338), .A2(n12104), .ZN(n1854) );
  XNOR2_X2 U19898 ( .A(n6758), .B(n6757), .ZN(n8387) );
  NAND2_X1 U19899 ( .A1(n20688), .A2(n14149), .ZN(n14152) );
  NAND2_X1 U19900 ( .A1(n14400), .A2(n14401), .ZN(n20688) );
  NAND2_X1 U19901 ( .A1(n2840), .A2(n7551), .ZN(n7552) );
  OR2_X1 U19902 ( .A1(n11376), .A2(n11330), .ZN(n1853) );
  INV_X1 U19903 ( .A(n15891), .ZN(n20689) );
  NAND3_X1 U19904 ( .A1(n360), .A2(n197), .A3(n15059), .ZN(n14988) );
  AND3_X2 U19905 ( .A1(n1700), .A2(n1697), .A3(n1696), .ZN(n15256) );
  OAI21_X1 U19906 ( .B1(n20374), .B2(n20691), .A(n8209), .ZN(n1910) );
  NOR2_X1 U19907 ( .A1(n8095), .A2(n7631), .ZN(n20691) );
  XNOR2_X1 U19908 ( .A(n20692), .B(n18379), .ZN(Ciphertext[7]) );
  NAND2_X1 U19909 ( .A1(n18378), .A2(n20693), .ZN(n20692) );
  OR2_X1 U19910 ( .A1(n18393), .A2(n1296), .ZN(n20693) );
  XNOR2_X1 U19911 ( .A(n13632), .B(n13633), .ZN(n13639) );
  NAND2_X1 U19912 ( .A1(n20362), .A2(n15686), .ZN(n15453) );
  NAND2_X1 U19913 ( .A1(n5520), .A2(n5927), .ZN(n5193) );
  NAND2_X1 U19914 ( .A1(n4809), .A2(n4810), .ZN(n4813) );
  NAND2_X1 U19915 ( .A1(n5074), .A2(n20431), .ZN(n4810) );
  NAND2_X1 U19916 ( .A1(n1831), .A2(n8660), .ZN(n1830) );
  NAND2_X1 U19917 ( .A1(n13053), .A2(n20694), .ZN(n13055) );
  NAND3_X1 U19918 ( .A1(n14307), .A2(n19940), .A3(n13040), .ZN(n20694) );
  OAI211_X1 U19919 ( .C1(n12275), .C2(n12028), .A(n11782), .B(n20695), .ZN(
        n2366) );
  NAND2_X1 U19920 ( .A1(n12275), .A2(n12029), .ZN(n20695) );
  AND3_X2 U19921 ( .A1(n20696), .A2(n1424), .A3(n449), .ZN(n9172) );
  NAND2_X1 U19922 ( .A1(n836), .A2(n837), .ZN(n20696) );
  OAI21_X1 U19923 ( .B1(n8616), .B2(n8763), .A(n20697), .ZN(n20054) );
  INV_X1 U19924 ( .A(n8693), .ZN(n20697) );
  XNOR2_X2 U19925 ( .A(n13197), .B(n13196), .ZN(n20266) );
  BUF_X2 U19926 ( .A(n17349), .Z(n19836) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;
  wire   n3;
  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFF_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CK(clk), .Q(reg_in[191]) );
  DFF_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CK(clk), .Q(reg_in[190]) );
  DFF_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CK(clk), .Q(reg_in[189]) );
  DFF_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CK(clk), .Q(reg_in[188]) );
  DFF_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CK(clk), .Q(reg_in[187]) );
  DFF_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CK(clk), .Q(reg_in[186]) );
  DFF_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CK(clk), .Q(reg_in[185]) );
  DFF_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CK(clk), .Q(reg_in[184]) );
  DFF_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CK(clk), .Q(reg_in[183]) );
  DFF_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CK(clk), .Q(reg_in[182]) );
  DFF_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CK(clk), .Q(reg_in[181]) );
  DFF_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CK(clk), .Q(reg_in[180]) );
  DFF_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CK(clk), .Q(reg_in[179]) );
  DFF_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CK(clk), .Q(reg_in[178]) );
  DFF_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CK(clk), .Q(reg_in[177]) );
  DFF_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CK(clk), .Q(reg_in[176]) );
  DFF_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CK(clk), .Q(reg_in[175]) );
  DFF_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CK(clk), .Q(reg_in[174]) );
  DFF_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CK(clk), .Q(reg_in[173]) );
  DFF_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CK(clk), .Q(reg_in[172]) );
  DFF_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CK(clk), .Q(reg_in[171]) );
  DFF_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CK(clk), .Q(reg_in[170]) );
  DFF_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CK(clk), .Q(reg_in[169]) );
  DFF_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CK(clk), .Q(reg_in[168]) );
  DFF_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CK(clk), .Q(reg_in[167]) );
  DFF_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CK(clk), .Q(reg_in[166]) );
  DFF_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CK(clk), .Q(reg_in[165]) );
  DFF_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CK(clk), .Q(reg_in[164]) );
  DFF_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CK(clk), .Q(reg_in[163]) );
  DFF_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CK(clk), .Q(reg_in[162]) );
  DFF_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CK(clk), .Q(reg_in[161]) );
  DFF_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CK(clk), .Q(reg_in[160]) );
  DFF_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CK(clk), .Q(reg_in[159]) );
  DFF_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CK(clk), .Q(reg_in[158]) );
  DFF_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CK(clk), .Q(reg_in[157]) );
  DFF_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CK(clk), .Q(reg_in[156]) );
  DFF_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CK(clk), .Q(reg_in[155]) );
  DFF_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CK(clk), .Q(reg_in[154]) );
  DFF_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CK(clk), .Q(reg_in[153]) );
  DFF_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CK(clk), .Q(reg_in[152]) );
  DFF_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CK(clk), .Q(reg_in[151]) );
  DFF_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CK(clk), .Q(reg_in[150]) );
  DFF_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CK(clk), .Q(reg_in[149]) );
  DFF_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CK(clk), .Q(reg_in[148]) );
  DFF_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CK(clk), .Q(reg_in[147]) );
  DFF_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CK(clk), .Q(reg_in[146]) );
  DFF_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CK(clk), .Q(reg_in[145]) );
  DFF_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CK(clk), .Q(reg_in[144]) );
  DFF_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CK(clk), .Q(reg_in[143]) );
  DFF_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CK(clk), .Q(reg_in[142]) );
  DFF_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CK(clk), .Q(reg_in[141]) );
  DFF_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CK(clk), .Q(reg_in[140]) );
  DFF_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CK(clk), .Q(reg_in[139]) );
  DFF_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CK(clk), .Q(reg_in[138]) );
  DFF_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CK(clk), .Q(reg_in[137]) );
  DFF_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CK(clk), .Q(reg_in[136]) );
  DFF_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CK(clk), .Q(reg_in[135]) );
  DFF_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CK(clk), .Q(reg_in[134]) );
  DFF_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CK(clk), .Q(reg_in[133]) );
  DFF_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CK(clk), .Q(reg_in[132]) );
  DFF_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CK(clk), .Q(reg_in[131]) );
  DFF_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CK(clk), .Q(reg_in[130]) );
  DFF_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CK(clk), .Q(reg_in[129]) );
  DFF_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CK(clk), .Q(reg_in[128]) );
  DFF_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CK(clk), .Q(reg_in[127]) );
  DFF_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CK(clk), .Q(reg_in[126]) );
  DFF_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CK(clk), .Q(reg_in[125]) );
  DFF_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CK(clk), .Q(reg_in[124]) );
  DFF_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CK(clk), .Q(reg_in[123]) );
  DFF_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CK(clk), .Q(reg_in[122]) );
  DFF_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CK(clk), .Q(reg_in[121]) );
  DFF_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CK(clk), .Q(reg_in[120]) );
  DFF_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CK(clk), .Q(reg_in[119]) );
  DFF_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CK(clk), .Q(reg_in[118]) );
  DFF_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CK(clk), .Q(reg_in[117]) );
  DFF_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CK(clk), .Q(reg_in[116]) );
  DFF_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CK(clk), .Q(reg_in[115]) );
  DFF_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CK(clk), .Q(reg_in[114]) );
  DFF_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CK(clk), .Q(reg_in[113]) );
  DFF_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CK(clk), .Q(reg_in[112]) );
  DFF_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CK(clk), .Q(reg_in[111]) );
  DFF_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CK(clk), .Q(reg_in[110]) );
  DFF_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CK(clk), .Q(reg_in[109]) );
  DFF_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CK(clk), .Q(reg_in[108]) );
  DFF_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CK(clk), .Q(reg_in[107]) );
  DFF_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CK(clk), .Q(reg_in[106]) );
  DFF_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CK(clk), .Q(reg_in[105]) );
  DFF_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CK(clk), .Q(reg_in[104]) );
  DFF_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CK(clk), .Q(reg_in[103]) );
  DFF_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CK(clk), .Q(reg_in[102]) );
  DFF_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CK(clk), .Q(reg_in[101]) );
  DFF_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CK(clk), .Q(reg_in[100]) );
  DFF_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CK(clk), .Q(reg_in[99]) );
  DFF_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CK(clk), .Q(reg_in[98]) );
  DFF_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CK(clk), .Q(reg_in[97]) );
  DFF_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CK(clk), .Q(reg_in[96]) );
  DFF_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CK(clk), .Q(reg_in[95]) );
  DFF_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CK(clk), .Q(reg_in[94]) );
  DFF_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CK(clk), .Q(reg_in[93]) );
  DFF_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CK(clk), .Q(reg_in[92]) );
  DFF_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CK(clk), .Q(reg_in[91]) );
  DFF_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CK(clk), .Q(reg_in[90]) );
  DFF_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CK(clk), .Q(reg_in[89]) );
  DFF_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CK(clk), .Q(reg_in[88]) );
  DFF_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CK(clk), .Q(reg_in[87]) );
  DFF_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CK(clk), .Q(reg_in[86]) );
  DFF_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CK(clk), .Q(reg_in[85]) );
  DFF_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CK(clk), .Q(reg_in[84]) );
  DFF_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CK(clk), .Q(reg_in[83]) );
  DFF_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CK(clk), .Q(reg_in[82]) );
  DFF_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CK(clk), .Q(reg_in[81]) );
  DFF_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CK(clk), .Q(reg_in[80]) );
  DFF_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CK(clk), .Q(reg_in[79]) );
  DFF_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CK(clk), .Q(reg_in[78]) );
  DFF_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CK(clk), .Q(reg_in[77]) );
  DFF_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CK(clk), .Q(reg_in[76]) );
  DFF_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CK(clk), .Q(reg_in[75]) );
  DFF_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CK(clk), .Q(reg_in[74]) );
  DFF_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CK(clk), .Q(reg_in[73]) );
  DFF_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CK(clk), .Q(reg_in[72]) );
  DFF_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CK(clk), .Q(reg_in[71]) );
  DFF_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CK(clk), .Q(reg_in[70]) );
  DFF_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CK(clk), .Q(reg_in[69]) );
  DFF_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CK(clk), .Q(reg_in[68]) );
  DFF_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CK(clk), .Q(reg_in[67]) );
  DFF_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CK(clk), .Q(reg_in[66]) );
  DFF_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CK(clk), .Q(reg_in[65]) );
  DFF_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CK(clk), .Q(reg_in[64]) );
  DFF_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CK(clk), .Q(reg_in[63]) );
  DFF_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CK(clk), .Q(reg_in[62]) );
  DFF_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CK(clk), .Q(reg_in[61]) );
  DFF_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CK(clk), .Q(reg_in[60]) );
  DFF_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CK(clk), .Q(reg_in[59]) );
  DFF_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CK(clk), .Q(reg_in[58]) );
  DFF_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CK(clk), .Q(reg_in[57]) );
  DFF_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CK(clk), .Q(reg_in[56]) );
  DFF_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CK(clk), .Q(reg_in[55]) );
  DFF_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CK(clk), .Q(reg_in[54]) );
  DFF_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CK(clk), .Q(reg_in[53]) );
  DFF_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CK(clk), .Q(reg_in[52]) );
  DFF_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CK(clk), .Q(reg_in[51]) );
  DFF_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CK(clk), .Q(reg_in[50]) );
  DFF_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CK(clk), .Q(reg_in[49]) );
  DFF_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CK(clk), .Q(reg_in[48]) );
  DFF_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CK(clk), .Q(reg_in[47]) );
  DFF_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CK(clk), .Q(reg_in[46]) );
  DFF_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CK(clk), .Q(reg_in[45]) );
  DFF_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CK(clk), .Q(reg_in[44]) );
  DFF_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CK(clk), .Q(reg_in[43]) );
  DFF_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CK(clk), .Q(reg_in[42]) );
  DFF_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CK(clk), .Q(reg_in[41]) );
  DFF_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CK(clk), .Q(reg_in[40]) );
  DFF_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CK(clk), .Q(reg_in[39]) );
  DFF_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CK(clk), .Q(reg_in[38]) );
  DFF_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CK(clk), .Q(reg_in[37]) );
  DFF_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CK(clk), .Q(reg_in[36]) );
  DFF_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CK(clk), .Q(reg_in[35]) );
  DFF_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CK(clk), .Q(reg_in[34]) );
  DFF_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CK(clk), .Q(reg_in[33]) );
  DFF_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CK(clk), .Q(reg_in[32]) );
  DFF_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CK(clk), .Q(reg_in[31]) );
  DFF_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CK(clk), .Q(reg_in[30]) );
  DFF_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CK(clk), .Q(reg_in[29]) );
  DFF_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CK(clk), .Q(reg_in[28]) );
  DFF_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CK(clk), .Q(reg_in[27]) );
  DFF_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CK(clk), .Q(reg_in[26]) );
  DFF_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CK(clk), .Q(reg_in[25]) );
  DFF_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CK(clk), .Q(reg_in[24]) );
  DFF_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CK(clk), .Q(reg_in[23]) );
  DFF_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CK(clk), .Q(reg_in[22]) );
  DFF_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CK(clk), .Q(reg_in[21]) );
  DFF_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CK(clk), .Q(reg_in[20]) );
  DFF_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CK(clk), .Q(reg_in[19]) );
  DFF_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CK(clk), .Q(reg_in[18]) );
  DFF_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CK(clk), .Q(reg_in[17]) );
  DFF_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CK(clk), .Q(reg_in[16]) );
  DFF_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CK(clk), .Q(reg_in[15]) );
  DFF_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CK(clk), .Q(reg_in[14]) );
  DFF_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CK(clk), .Q(reg_in[13]) );
  DFF_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CK(clk), .Q(reg_in[12]) );
  DFF_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CK(clk), .Q(reg_in[11]) );
  DFF_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CK(clk), .Q(reg_in[10]) );
  DFF_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CK(clk), .Q(reg_in[9]) );
  DFF_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CK(clk), .Q(reg_in[8]) );
  DFF_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CK(clk), .Q(reg_in[7]) );
  DFF_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CK(clk), .Q(reg_in[6]) );
  DFF_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CK(clk), .Q(reg_in[5]) );
  DFF_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CK(clk), .Q(reg_in[4]) );
  DFF_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CK(clk), .Q(reg_in[3]) );
  DFF_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CK(clk), .Q(reg_in[2]) );
  DFF_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CK(clk), .Q(reg_in[1]) );
  DFF_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CK(clk), .Q(reg_in[0]) );
  DFF_X1 \reg_key_reg[191]  ( .D(Key[191]), .CK(clk), .Q(reg_key[191]) );
  DFF_X1 \reg_key_reg[190]  ( .D(Key[190]), .CK(clk), .Q(reg_key[190]) );
  DFF_X1 \reg_key_reg[189]  ( .D(Key[189]), .CK(clk), .Q(reg_key[189]) );
  DFF_X1 \reg_key_reg[188]  ( .D(Key[188]), .CK(clk), .Q(reg_key[188]) );
  DFF_X1 \reg_key_reg[186]  ( .D(Key[186]), .CK(clk), .Q(n3) );
  DFF_X1 \reg_key_reg[184]  ( .D(Key[184]), .CK(clk), .Q(reg_key[184]) );
  DFF_X1 \reg_key_reg[181]  ( .D(Key[181]), .CK(clk), .Q(reg_key[181]) );
  DFF_X1 \reg_key_reg[180]  ( .D(Key[180]), .CK(clk), .Q(reg_key[180]) );
  DFF_X1 \reg_key_reg[178]  ( .D(Key[178]), .CK(clk), .Q(reg_key[178]) );
  DFF_X1 \reg_key_reg[177]  ( .D(Key[177]), .CK(clk), .Q(reg_key[177]) );
  DFF_X1 \reg_key_reg[176]  ( .D(Key[176]), .CK(clk), .Q(reg_key[176]) );
  DFF_X1 \reg_key_reg[175]  ( .D(Key[175]), .CK(clk), .Q(reg_key[175]) );
  DFF_X1 \reg_key_reg[174]  ( .D(Key[174]), .CK(clk), .Q(reg_key[174]) );
  DFF_X1 \reg_key_reg[173]  ( .D(Key[173]), .CK(clk), .Q(reg_key[173]) );
  DFF_X1 \reg_key_reg[172]  ( .D(Key[172]), .CK(clk), .Q(reg_key[172]) );
  DFF_X1 \reg_key_reg[170]  ( .D(Key[170]), .CK(clk), .Q(reg_key[170]) );
  DFF_X1 \reg_key_reg[169]  ( .D(Key[169]), .CK(clk), .Q(reg_key[169]) );
  DFF_X1 \reg_key_reg[168]  ( .D(Key[168]), .CK(clk), .Q(reg_key[168]) );
  DFF_X1 \reg_key_reg[167]  ( .D(Key[167]), .CK(clk), .Q(reg_key[167]) );
  DFF_X1 \reg_key_reg[164]  ( .D(Key[164]), .CK(clk), .Q(reg_key[164]) );
  DFF_X1 \reg_key_reg[163]  ( .D(Key[163]), .CK(clk), .Q(reg_key[163]) );
  DFF_X1 \reg_key_reg[162]  ( .D(Key[162]), .CK(clk), .Q(reg_key[162]) );
  DFF_X1 \reg_key_reg[161]  ( .D(Key[161]), .CK(clk), .Q(reg_key[161]) );
  DFF_X1 \reg_key_reg[160]  ( .D(Key[160]), .CK(clk), .Q(reg_key[160]) );
  DFF_X1 \reg_key_reg[159]  ( .D(Key[159]), .CK(clk), .Q(reg_key[159]) );
  DFF_X1 \reg_key_reg[158]  ( .D(Key[158]), .CK(clk), .Q(reg_key[158]) );
  DFF_X1 \reg_key_reg[157]  ( .D(Key[157]), .CK(clk), .Q(reg_key[157]) );
  DFF_X1 \reg_key_reg[156]  ( .D(Key[156]), .CK(clk), .Q(reg_key[156]) );
  DFF_X1 \reg_key_reg[155]  ( .D(Key[155]), .CK(clk), .Q(reg_key[155]) );
  DFF_X1 \reg_key_reg[154]  ( .D(Key[154]), .CK(clk), .Q(reg_key[154]) );
  DFF_X1 \reg_key_reg[153]  ( .D(Key[153]), .CK(clk), .Q(reg_key[153]) );
  DFF_X1 \reg_key_reg[152]  ( .D(Key[152]), .CK(clk), .Q(reg_key[152]) );
  DFF_X1 \reg_key_reg[151]  ( .D(Key[151]), .CK(clk), .Q(reg_key[151]) );
  DFF_X1 \reg_key_reg[149]  ( .D(Key[149]), .CK(clk), .Q(reg_key[149]) );
  DFF_X1 \reg_key_reg[148]  ( .D(Key[148]), .CK(clk), .Q(reg_key[148]) );
  DFF_X1 \reg_key_reg[147]  ( .D(Key[147]), .CK(clk), .Q(reg_key[147]) );
  DFF_X1 \reg_key_reg[146]  ( .D(Key[146]), .CK(clk), .Q(reg_key[146]) );
  DFF_X1 \reg_key_reg[145]  ( .D(Key[145]), .CK(clk), .Q(reg_key[145]) );
  DFF_X1 \reg_key_reg[144]  ( .D(Key[144]), .CK(clk), .Q(reg_key[144]) );
  DFF_X1 \reg_key_reg[143]  ( .D(Key[143]), .CK(clk), .Q(reg_key[143]) );
  DFF_X1 \reg_key_reg[142]  ( .D(Key[142]), .CK(clk), .Q(reg_key[142]) );
  DFF_X1 \reg_key_reg[141]  ( .D(Key[141]), .CK(clk), .Q(reg_key[141]) );
  DFF_X1 \reg_key_reg[140]  ( .D(Key[140]), .CK(clk), .Q(reg_key[140]) );
  DFF_X1 \reg_key_reg[139]  ( .D(Key[139]), .CK(clk), .Q(reg_key[139]) );
  DFF_X1 \reg_key_reg[138]  ( .D(Key[138]), .CK(clk), .Q(reg_key[138]) );
  DFF_X1 \reg_key_reg[137]  ( .D(Key[137]), .CK(clk), .Q(reg_key[137]) );
  DFF_X1 \reg_key_reg[136]  ( .D(Key[136]), .CK(clk), .Q(reg_key[136]) );
  DFF_X1 \reg_key_reg[135]  ( .D(Key[135]), .CK(clk), .Q(reg_key[135]) );
  DFF_X1 \reg_key_reg[133]  ( .D(Key[133]), .CK(clk), .Q(reg_key[133]) );
  DFF_X1 \reg_key_reg[132]  ( .D(Key[132]), .CK(clk), .Q(reg_key[132]) );
  DFF_X1 \reg_key_reg[131]  ( .D(Key[131]), .CK(clk), .Q(reg_key[131]) );
  DFF_X1 \reg_key_reg[130]  ( .D(Key[130]), .CK(clk), .Q(reg_key[130]) );
  DFF_X1 \reg_key_reg[129]  ( .D(Key[129]), .CK(clk), .Q(reg_key[129]) );
  DFF_X1 \reg_key_reg[128]  ( .D(Key[128]), .CK(clk), .Q(reg_key[128]) );
  DFF_X1 \reg_key_reg[127]  ( .D(Key[127]), .CK(clk), .Q(reg_key[127]) );
  DFF_X1 \reg_key_reg[125]  ( .D(Key[125]), .CK(clk), .Q(reg_key[125]) );
  DFF_X1 \reg_key_reg[124]  ( .D(Key[124]), .CK(clk), .Q(reg_key[124]) );
  DFF_X1 \reg_key_reg[123]  ( .D(Key[123]), .CK(clk), .Q(reg_key[123]) );
  DFF_X1 \reg_key_reg[122]  ( .D(Key[122]), .CK(clk), .Q(reg_key[122]) );
  DFF_X1 \reg_key_reg[121]  ( .D(Key[121]), .CK(clk), .Q(reg_key[121]) );
  DFF_X1 \reg_key_reg[120]  ( .D(Key[120]), .CK(clk), .Q(reg_key[120]) );
  DFF_X1 \reg_key_reg[119]  ( .D(Key[119]), .CK(clk), .Q(reg_key[119]) );
  DFF_X1 \reg_key_reg[118]  ( .D(Key[118]), .CK(clk), .Q(reg_key[118]) );
  DFF_X1 \reg_key_reg[117]  ( .D(Key[117]), .CK(clk), .Q(reg_key[117]) );
  DFF_X1 \reg_key_reg[116]  ( .D(Key[116]), .CK(clk), .Q(reg_key[116]) );
  DFF_X1 \reg_key_reg[115]  ( .D(Key[115]), .CK(clk), .Q(reg_key[115]) );
  DFF_X1 \reg_key_reg[114]  ( .D(Key[114]), .CK(clk), .Q(reg_key[114]) );
  DFF_X1 \reg_key_reg[112]  ( .D(Key[112]), .CK(clk), .Q(reg_key[112]) );
  DFF_X1 \reg_key_reg[111]  ( .D(Key[111]), .CK(clk), .Q(reg_key[111]) );
  DFF_X1 \reg_key_reg[109]  ( .D(Key[109]), .CK(clk), .Q(reg_key[109]) );
  DFF_X1 \reg_key_reg[108]  ( .D(Key[108]), .CK(clk), .Q(reg_key[108]) );
  DFF_X1 \reg_key_reg[106]  ( .D(Key[106]), .CK(clk), .Q(reg_key[106]) );
  DFF_X1 \reg_key_reg[104]  ( .D(Key[104]), .CK(clk), .Q(reg_key[104]) );
  DFF_X1 \reg_key_reg[103]  ( .D(Key[103]), .CK(clk), .Q(reg_key[103]) );
  DFF_X1 \reg_key_reg[102]  ( .D(Key[102]), .CK(clk), .Q(reg_key[102]) );
  DFF_X1 \reg_key_reg[101]  ( .D(Key[101]), .CK(clk), .Q(reg_key[101]) );
  DFF_X1 \reg_key_reg[100]  ( .D(Key[100]), .CK(clk), .Q(reg_key[100]) );
  DFF_X1 \reg_key_reg[99]  ( .D(Key[99]), .CK(clk), .Q(reg_key[99]) );
  DFF_X1 \reg_key_reg[98]  ( .D(Key[98]), .CK(clk), .Q(reg_key[98]) );
  DFF_X1 \reg_key_reg[97]  ( .D(Key[97]), .CK(clk), .Q(reg_key[97]) );
  DFF_X1 \reg_key_reg[96]  ( .D(Key[96]), .CK(clk), .Q(reg_key[96]) );
  DFF_X1 \reg_key_reg[95]  ( .D(Key[95]), .CK(clk), .Q(reg_key[95]) );
  DFF_X1 \reg_key_reg[94]  ( .D(Key[94]), .CK(clk), .Q(reg_key[94]) );
  DFF_X1 \reg_key_reg[93]  ( .D(Key[93]), .CK(clk), .Q(reg_key[93]) );
  DFF_X1 \reg_key_reg[92]  ( .D(Key[92]), .CK(clk), .Q(reg_key[92]) );
  DFF_X1 \reg_key_reg[91]  ( .D(Key[91]), .CK(clk), .Q(reg_key[91]) );
  DFF_X1 \reg_key_reg[90]  ( .D(Key[90]), .CK(clk), .Q(reg_key[90]) );
  DFF_X1 \reg_key_reg[88]  ( .D(Key[88]), .CK(clk), .Q(reg_key[88]) );
  DFF_X1 \reg_key_reg[85]  ( .D(Key[85]), .CK(clk), .Q(reg_key[85]) );
  DFF_X1 \reg_key_reg[84]  ( .D(Key[84]), .CK(clk), .Q(reg_key[84]) );
  DFF_X1 \reg_key_reg[82]  ( .D(Key[82]), .CK(clk), .Q(reg_key[82]) );
  DFF_X1 \reg_key_reg[81]  ( .D(Key[81]), .CK(clk), .Q(reg_key[81]) );
  DFF_X1 \reg_key_reg[80]  ( .D(Key[80]), .CK(clk), .Q(reg_key[80]) );
  DFF_X1 \reg_key_reg[78]  ( .D(Key[78]), .CK(clk), .Q(reg_key[78]) );
  DFF_X1 \reg_key_reg[76]  ( .D(Key[76]), .CK(clk), .Q(reg_key[76]) );
  DFF_X1 \reg_key_reg[75]  ( .D(Key[75]), .CK(clk), .Q(reg_key[75]) );
  DFF_X1 \reg_key_reg[74]  ( .D(Key[74]), .CK(clk), .Q(reg_key[74]) );
  DFF_X1 \reg_key_reg[73]  ( .D(Key[73]), .CK(clk), .Q(reg_key[73]) );
  DFF_X1 \reg_key_reg[72]  ( .D(Key[72]), .CK(clk), .Q(reg_key[72]) );
  DFF_X1 \reg_key_reg[70]  ( .D(Key[70]), .CK(clk), .Q(reg_key[70]) );
  DFF_X1 \reg_key_reg[69]  ( .D(Key[69]), .CK(clk), .Q(reg_key[69]) );
  DFF_X1 \reg_key_reg[67]  ( .D(Key[67]), .CK(clk), .Q(reg_key[67]) );
  DFF_X1 \reg_key_reg[66]  ( .D(Key[66]), .CK(clk), .Q(reg_key[66]) );
  DFF_X1 \reg_key_reg[61]  ( .D(Key[61]), .CK(clk), .Q(reg_key[61]) );
  DFF_X1 \reg_key_reg[59]  ( .D(Key[59]), .CK(clk), .Q(reg_key[59]) );
  DFF_X1 \reg_key_reg[58]  ( .D(Key[58]), .CK(clk), .Q(reg_key[58]) );
  DFF_X1 \reg_key_reg[57]  ( .D(Key[57]), .CK(clk), .Q(reg_key[57]) );
  DFF_X1 \reg_key_reg[55]  ( .D(Key[55]), .CK(clk), .Q(reg_key[55]) );
  DFF_X1 \reg_key_reg[54]  ( .D(Key[54]), .CK(clk), .Q(reg_key[54]) );
  DFF_X1 \reg_key_reg[53]  ( .D(Key[53]), .CK(clk), .Q(reg_key[53]) );
  DFF_X1 \reg_key_reg[51]  ( .D(Key[51]), .CK(clk), .Q(reg_key[51]) );
  DFF_X1 \reg_key_reg[50]  ( .D(Key[50]), .CK(clk), .Q(reg_key[50]) );
  DFF_X1 \reg_key_reg[49]  ( .D(Key[49]), .CK(clk), .Q(reg_key[49]) );
  DFF_X1 \reg_key_reg[48]  ( .D(Key[48]), .CK(clk), .Q(reg_key[48]) );
  DFF_X1 \reg_key_reg[47]  ( .D(Key[47]), .CK(clk), .Q(reg_key[47]) );
  DFF_X1 \reg_key_reg[45]  ( .D(Key[45]), .CK(clk), .Q(reg_key[45]) );
  DFF_X1 \reg_key_reg[44]  ( .D(Key[44]), .CK(clk), .Q(reg_key[44]) );
  DFF_X1 \reg_key_reg[43]  ( .D(Key[43]), .CK(clk), .Q(reg_key[43]) );
  DFF_X1 \reg_key_reg[42]  ( .D(Key[42]), .CK(clk), .Q(reg_key[42]) );
  DFF_X1 \reg_key_reg[40]  ( .D(Key[40]), .CK(clk), .Q(reg_key[40]) );
  DFF_X1 \reg_key_reg[39]  ( .D(Key[39]), .CK(clk), .Q(reg_key[39]) );
  DFF_X1 \reg_key_reg[38]  ( .D(Key[38]), .CK(clk), .Q(reg_key[38]) );
  DFF_X1 \reg_key_reg[36]  ( .D(Key[36]), .CK(clk), .Q(reg_key[36]) );
  DFF_X1 \reg_key_reg[35]  ( .D(Key[35]), .CK(clk), .Q(reg_key[35]) );
  DFF_X1 \reg_key_reg[34]  ( .D(Key[34]), .CK(clk), .Q(reg_key[34]) );
  DFF_X1 \reg_key_reg[33]  ( .D(Key[33]), .CK(clk), .Q(reg_key[33]) );
  DFF_X1 \reg_key_reg[32]  ( .D(Key[32]), .CK(clk), .Q(reg_key[32]) );
  DFF_X1 \reg_key_reg[31]  ( .D(Key[31]), .CK(clk), .Q(reg_key[31]) );
  DFF_X1 \reg_key_reg[30]  ( .D(Key[30]), .CK(clk), .Q(reg_key[30]) );
  DFF_X1 \reg_key_reg[29]  ( .D(Key[29]), .CK(clk), .Q(reg_key[29]) );
  DFF_X1 \reg_key_reg[27]  ( .D(Key[27]), .CK(clk), .Q(reg_key[27]) );
  DFF_X1 \reg_key_reg[26]  ( .D(Key[26]), .CK(clk), .Q(reg_key[26]) );
  DFF_X1 \reg_key_reg[25]  ( .D(Key[25]), .CK(clk), .Q(reg_key[25]) );
  DFF_X1 \reg_key_reg[24]  ( .D(Key[24]), .CK(clk), .Q(reg_key[24]) );
  DFF_X1 \reg_key_reg[22]  ( .D(Key[22]), .CK(clk), .Q(reg_key[22]) );
  DFF_X1 \reg_key_reg[21]  ( .D(Key[21]), .CK(clk), .Q(reg_key[21]) );
  DFF_X1 \reg_key_reg[20]  ( .D(Key[20]), .CK(clk), .Q(reg_key[20]) );
  DFF_X1 \reg_key_reg[19]  ( .D(Key[19]), .CK(clk), .Q(reg_key[19]) );
  DFF_X1 \reg_key_reg[18]  ( .D(Key[18]), .CK(clk), .Q(reg_key[18]) );
  DFF_X1 \reg_key_reg[17]  ( .D(Key[17]), .CK(clk), .Q(reg_key[17]) );
  DFF_X1 \reg_key_reg[16]  ( .D(Key[16]), .CK(clk), .Q(reg_key[16]) );
  DFF_X1 \reg_key_reg[15]  ( .D(Key[15]), .CK(clk), .Q(reg_key[15]) );
  DFF_X1 \reg_key_reg[14]  ( .D(Key[14]), .CK(clk), .Q(reg_key[14]) );
  DFF_X1 \reg_key_reg[12]  ( .D(Key[12]), .CK(clk), .Q(reg_key[12]) );
  DFF_X1 \reg_key_reg[11]  ( .D(Key[11]), .CK(clk), .Q(reg_key[11]) );
  DFF_X1 \reg_key_reg[10]  ( .D(Key[10]), .CK(clk), .Q(reg_key[10]) );
  DFF_X1 \reg_key_reg[9]  ( .D(Key[9]), .CK(clk), .Q(reg_key[9]) );
  DFF_X1 \reg_key_reg[8]  ( .D(Key[8]), .CK(clk), .Q(reg_key[8]) );
  DFF_X1 \reg_key_reg[7]  ( .D(Key[7]), .CK(clk), .Q(reg_key[7]) );
  DFF_X1 \reg_key_reg[6]  ( .D(Key[6]), .CK(clk), .Q(reg_key[6]) );
  DFF_X1 \reg_key_reg[5]  ( .D(Key[5]), .CK(clk), .Q(reg_key[5]) );
  DFF_X1 \reg_key_reg[4]  ( .D(Key[4]), .CK(clk), .Q(reg_key[4]) );
  DFF_X1 \reg_key_reg[3]  ( .D(Key[3]), .CK(clk), .Q(reg_key[3]) );
  DFF_X1 \reg_key_reg[2]  ( .D(Key[2]), .CK(clk), .Q(reg_key[2]) );
  DFF_X1 \reg_key_reg[1]  ( .D(Key[1]), .CK(clk), .Q(reg_key[1]) );
  DFF_X1 \reg_key_reg[0]  ( .D(Key[0]), .CK(clk), .Q(reg_key[0]) );
  DFF_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CK(clk), .Q(
        Ciphertext[191]) );
  DFF_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CK(clk), .Q(
        Ciphertext[190]) );
  DFF_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CK(clk), .Q(
        Ciphertext[189]) );
  DFF_X1 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CK(clk), .Q(
        Ciphertext[188]) );
  DFF_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CK(clk), .Q(
        Ciphertext[187]) );
  DFF_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CK(clk), .Q(
        Ciphertext[186]) );
  DFF_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CK(clk), .Q(
        Ciphertext[185]) );
  DFF_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CK(clk), .Q(
        Ciphertext[184]) );
  DFF_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CK(clk), .Q(
        Ciphertext[183]) );
  DFF_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CK(clk), .Q(
        Ciphertext[182]) );
  DFF_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CK(clk), .Q(
        Ciphertext[181]) );
  DFF_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CK(clk), .Q(
        Ciphertext[180]) );
  DFF_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CK(clk), .Q(
        Ciphertext[179]) );
  DFF_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CK(clk), .Q(
        Ciphertext[178]) );
  DFF_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CK(clk), .Q(
        Ciphertext[177]) );
  DFF_X1 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CK(clk), .Q(
        Ciphertext[176]) );
  DFF_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CK(clk), .Q(
        Ciphertext[175]) );
  DFF_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CK(clk), .Q(
        Ciphertext[174]) );
  DFF_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CK(clk), .Q(
        Ciphertext[173]) );
  DFF_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CK(clk), .Q(
        Ciphertext[172]) );
  DFF_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CK(clk), .Q(
        Ciphertext[171]) );
  DFF_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CK(clk), .Q(
        Ciphertext[170]) );
  DFF_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CK(clk), .Q(
        Ciphertext[169]) );
  DFF_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CK(clk), .Q(
        Ciphertext[168]) );
  DFF_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CK(clk), .Q(
        Ciphertext[167]) );
  DFF_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CK(clk), .Q(
        Ciphertext[166]) );
  DFF_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CK(clk), .Q(
        Ciphertext[165]) );
  DFF_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CK(clk), .Q(
        Ciphertext[164]) );
  DFF_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CK(clk), .Q(
        Ciphertext[162]) );
  DFF_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CK(clk), .Q(
        Ciphertext[161]) );
  DFF_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CK(clk), .Q(
        Ciphertext[159]) );
  DFF_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CK(clk), .Q(
        Ciphertext[158]) );
  DFF_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CK(clk), .Q(
        Ciphertext[157]) );
  DFF_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CK(clk), .Q(
        Ciphertext[155]) );
  DFF_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CK(clk), .Q(
        Ciphertext[154]) );
  DFF_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CK(clk), .Q(
        Ciphertext[153]) );
  DFF_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CK(clk), .Q(
        Ciphertext[152]) );
  DFF_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CK(clk), .Q(
        Ciphertext[151]) );
  DFF_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CK(clk), .Q(
        Ciphertext[150]) );
  DFF_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CK(clk), .Q(
        Ciphertext[149]) );
  DFF_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CK(clk), .Q(
        Ciphertext[148]) );
  DFF_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CK(clk), .Q(
        Ciphertext[147]) );
  DFF_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CK(clk), .Q(
        Ciphertext[146]) );
  DFF_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CK(clk), .Q(
        Ciphertext[145]) );
  DFF_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CK(clk), .Q(
        Ciphertext[144]) );
  DFF_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CK(clk), .Q(
        Ciphertext[143]) );
  DFF_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CK(clk), .Q(
        Ciphertext[142]) );
  DFF_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CK(clk), .Q(
        Ciphertext[141]) );
  DFF_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CK(clk), .Q(
        Ciphertext[140]) );
  DFF_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CK(clk), .Q(
        Ciphertext[139]) );
  DFF_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CK(clk), .Q(
        Ciphertext[138]) );
  DFF_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CK(clk), .Q(
        Ciphertext[137]) );
  DFF_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CK(clk), .Q(
        Ciphertext[136]) );
  DFF_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CK(clk), .Q(
        Ciphertext[135]) );
  DFF_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CK(clk), .Q(
        Ciphertext[134]) );
  DFF_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CK(clk), .Q(
        Ciphertext[133]) );
  DFF_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CK(clk), .Q(
        Ciphertext[132]) );
  DFF_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CK(clk), .Q(
        Ciphertext[131]) );
  DFF_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CK(clk), .Q(
        Ciphertext[130]) );
  DFF_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CK(clk), .Q(
        Ciphertext[129]) );
  DFF_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CK(clk), .Q(
        Ciphertext[128]) );
  DFF_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CK(clk), .Q(
        Ciphertext[127]) );
  DFF_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CK(clk), .Q(
        Ciphertext[126]) );
  DFF_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CK(clk), .Q(
        Ciphertext[125]) );
  DFF_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CK(clk), .Q(
        Ciphertext[124]) );
  DFF_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CK(clk), .Q(
        Ciphertext[123]) );
  DFF_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CK(clk), .Q(
        Ciphertext[122]) );
  DFF_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CK(clk), .Q(
        Ciphertext[121]) );
  DFF_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CK(clk), .Q(
        Ciphertext[120]) );
  DFF_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CK(clk), .Q(
        Ciphertext[119]) );
  DFF_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CK(clk), .Q(
        Ciphertext[118]) );
  DFF_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CK(clk), .Q(
        Ciphertext[117]) );
  DFF_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CK(clk), .Q(
        Ciphertext[116]) );
  DFF_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CK(clk), .Q(
        Ciphertext[114]) );
  DFF_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CK(clk), .Q(
        Ciphertext[113]) );
  DFF_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CK(clk), .Q(
        Ciphertext[112]) );
  DFF_X1 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CK(clk), .Q(
        Ciphertext[111]) );
  DFF_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CK(clk), .Q(
        Ciphertext[110]) );
  DFF_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CK(clk), .Q(
        Ciphertext[109]) );
  DFF_X1 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CK(clk), .Q(
        Ciphertext[108]) );
  DFF_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CK(clk), .Q(
        Ciphertext[107]) );
  DFF_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CK(clk), .Q(
        Ciphertext[106]) );
  DFF_X1 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CK(clk), .Q(
        Ciphertext[105]) );
  DFF_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CK(clk), .Q(
        Ciphertext[104]) );
  DFF_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CK(clk), .Q(
        Ciphertext[103]) );
  DFF_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CK(clk), .Q(
        Ciphertext[102]) );
  DFF_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CK(clk), .Q(
        Ciphertext[101]) );
  DFF_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CK(clk), .Q(
        Ciphertext[100]) );
  DFF_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CK(clk), .Q(Ciphertext[98])
         );
  DFF_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CK(clk), .Q(Ciphertext[97])
         );
  DFF_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CK(clk), .Q(Ciphertext[96])
         );
  DFF_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CK(clk), .Q(Ciphertext[95])
         );
  DFF_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CK(clk), .Q(Ciphertext[94])
         );
  DFF_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CK(clk), .Q(Ciphertext[93])
         );
  DFF_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CK(clk), .Q(Ciphertext[91])
         );
  DFF_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CK(clk), .Q(Ciphertext[90])
         );
  DFF_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CK(clk), .Q(Ciphertext[89])
         );
  DFF_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CK(clk), .Q(Ciphertext[88])
         );
  DFF_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CK(clk), .Q(Ciphertext[86])
         );
  DFF_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CK(clk), .Q(Ciphertext[85])
         );
  DFF_X1 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CK(clk), .Q(Ciphertext[84])
         );
  DFF_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CK(clk), .Q(Ciphertext[83])
         );
  DFF_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CK(clk), .Q(Ciphertext[82])
         );
  DFF_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CK(clk), .Q(Ciphertext[81])
         );
  DFF_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CK(clk), .Q(Ciphertext[80])
         );
  DFF_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CK(clk), .Q(Ciphertext[78])
         );
  DFF_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CK(clk), .Q(Ciphertext[77])
         );
  DFF_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CK(clk), .Q(Ciphertext[76])
         );
  DFF_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CK(clk), .Q(Ciphertext[75])
         );
  DFF_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CK(clk), .Q(Ciphertext[74])
         );
  DFF_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CK(clk), .Q(Ciphertext[73])
         );
  DFF_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CK(clk), .Q(Ciphertext[72])
         );
  DFF_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CK(clk), .Q(Ciphertext[71])
         );
  DFF_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CK(clk), .Q(Ciphertext[70])
         );
  DFF_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CK(clk), .Q(Ciphertext[69])
         );
  DFF_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CK(clk), .Q(Ciphertext[68])
         );
  DFF_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CK(clk), .Q(Ciphertext[67])
         );
  DFF_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CK(clk), .Q(Ciphertext[66])
         );
  DFF_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CK(clk), .Q(Ciphertext[65])
         );
  DFF_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CK(clk), .Q(Ciphertext[64])
         );
  DFF_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CK(clk), .Q(Ciphertext[63])
         );
  DFF_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CK(clk), .Q(Ciphertext[62])
         );
  DFF_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CK(clk), .Q(Ciphertext[61])
         );
  DFF_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CK(clk), .Q(Ciphertext[60])
         );
  DFF_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CK(clk), .Q(Ciphertext[59])
         );
  DFF_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CK(clk), .Q(Ciphertext[57])
         );
  DFF_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CK(clk), .Q(Ciphertext[56])
         );
  DFF_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CK(clk), .Q(Ciphertext[55])
         );
  DFF_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CK(clk), .Q(Ciphertext[54])
         );
  DFF_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CK(clk), .Q(Ciphertext[53])
         );
  DFF_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CK(clk), .Q(Ciphertext[52])
         );
  DFF_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CK(clk), .Q(Ciphertext[51])
         );
  DFF_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CK(clk), .Q(Ciphertext[50])
         );
  DFF_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CK(clk), .Q(Ciphertext[49])
         );
  DFF_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CK(clk), .Q(Ciphertext[48])
         );
  DFF_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CK(clk), .Q(Ciphertext[47])
         );
  DFF_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CK(clk), .Q(Ciphertext[46])
         );
  DFF_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CK(clk), .Q(Ciphertext[45])
         );
  DFF_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CK(clk), .Q(Ciphertext[44])
         );
  DFF_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CK(clk), .Q(Ciphertext[43])
         );
  DFF_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CK(clk), .Q(Ciphertext[42])
         );
  DFF_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CK(clk), .Q(Ciphertext[41])
         );
  DFF_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CK(clk), .Q(Ciphertext[39])
         );
  DFF_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CK(clk), .Q(Ciphertext[38])
         );
  DFF_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CK(clk), .Q(Ciphertext[37])
         );
  DFF_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CK(clk), .Q(Ciphertext[36])
         );
  DFF_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CK(clk), .Q(Ciphertext[35])
         );
  DFF_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CK(clk), .Q(Ciphertext[34])
         );
  DFF_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CK(clk), .Q(Ciphertext[32])
         );
  DFF_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CK(clk), .Q(Ciphertext[31])
         );
  DFF_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CK(clk), .Q(Ciphertext[30])
         );
  DFF_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CK(clk), .Q(Ciphertext[29])
         );
  DFF_X1 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CK(clk), .Q(Ciphertext[28])
         );
  DFF_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CK(clk), .Q(Ciphertext[27])
         );
  DFF_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CK(clk), .Q(Ciphertext[26])
         );
  DFF_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CK(clk), .Q(Ciphertext[25])
         );
  DFF_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CK(clk), .Q(Ciphertext[24])
         );
  DFF_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CK(clk), .Q(Ciphertext[23])
         );
  DFF_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CK(clk), .Q(Ciphertext[22])
         );
  DFF_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CK(clk), .Q(Ciphertext[21])
         );
  DFF_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CK(clk), .Q(Ciphertext[20])
         );
  DFF_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CK(clk), .Q(Ciphertext[19])
         );
  DFF_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CK(clk), .Q(Ciphertext[18])
         );
  DFF_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CK(clk), .Q(Ciphertext[17])
         );
  DFF_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CK(clk), .Q(Ciphertext[16])
         );
  DFF_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CK(clk), .Q(Ciphertext[15])
         );
  DFF_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CK(clk), .Q(Ciphertext[14])
         );
  DFF_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CK(clk), .Q(Ciphertext[13])
         );
  DFF_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CK(clk), .Q(Ciphertext[11])
         );
  DFF_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CK(clk), .Q(Ciphertext[10])
         );
  DFF_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CK(clk), .Q(Ciphertext[9]) );
  DFF_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CK(clk), .Q(Ciphertext[7]) );
  DFF_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CK(clk), .Q(Ciphertext[6]) );
  DFF_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CK(clk), .Q(Ciphertext[5]) );
  DFF_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CK(clk), .Q(Ciphertext[4]) );
  DFF_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CK(clk), .Q(Ciphertext[2]) );
  DFF_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CK(clk), .Q(Ciphertext[1]) );
  DFF_X1 \reg_key_reg[179]  ( .D(Key[179]), .CK(clk), .Q(reg_key[179]) );
  DFF_X1 \reg_key_reg[62]  ( .D(Key[62]), .CK(clk), .Q(reg_key[62]) );
  DFF_X1 \reg_key_reg[113]  ( .D(Key[113]), .CK(clk), .Q(reg_key[113]) );
  DFF_X1 \reg_key_reg[79]  ( .D(Key[79]), .CK(clk), .Q(reg_key[79]) );
  DFF_X1 \reg_key_reg[183]  ( .D(Key[183]), .CK(clk), .Q(reg_key[183]) );
  DFF_X1 \reg_key_reg[166]  ( .D(Key[166]), .CK(clk), .Q(reg_key[166]) );
  DFF_X1 \reg_key_reg[107]  ( .D(Key[107]), .CK(clk), .Q(reg_key[107]) );
  DFF_X1 \reg_key_reg[56]  ( .D(Key[56]), .CK(clk), .Q(reg_key[56]) );
  DFF_X1 \reg_key_reg[187]  ( .D(Key[187]), .CK(clk), .Q(reg_key[187]) );
  DFF_X1 \reg_key_reg[77]  ( .D(Key[77]), .CK(clk), .Q(reg_key[77]) );
  DFF_X1 \reg_key_reg[23]  ( .D(Key[23]), .CK(clk), .Q(reg_key[23]) );
  DFFRS_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CK(clk), .RN(1'b1), .SN(1'b1), .Q(Ciphertext[3]) );
  DFF_X1 \reg_key_reg[83]  ( .D(Key[83]), .CK(clk), .Q(reg_key[83]) );
  DFF_X1 \reg_key_reg[71]  ( .D(Key[71]), .CK(clk), .Q(reg_key[71]) );
  DFF_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CK(clk), .Q(
        Ciphertext[156]) );
  DFF_X1 \reg_key_reg[68]  ( .D(Key[68]), .CK(clk), .Q(reg_key[68]) );
  DFF_X1 \reg_key_reg[171]  ( .D(Key[171]), .CK(clk), .Q(reg_key[171]) );
  DFF_X1 \reg_key_reg[13]  ( .D(Key[13]), .CK(clk), .Q(reg_key[13]) );
  DFF_X1 \reg_key_reg[165]  ( .D(Key[165]), .CK(clk), .Q(reg_key[165]) );
  DFF_X1 \reg_key_reg[64]  ( .D(Key[64]), .CK(clk), .Q(reg_key[64]) );
  DFF_X1 \reg_key_reg[63]  ( .D(Key[63]), .CK(clk), .Q(reg_key[63]) );
  DFF_X1 \reg_key_reg[126]  ( .D(Key[126]), .CK(clk), .Q(reg_key[126]) );
  DFF_X1 \reg_key_reg[185]  ( .D(Key[185]), .CK(clk), .Q(reg_key[185]) );
  DFF_X1 \reg_key_reg[134]  ( .D(Key[134]), .CK(clk), .Q(reg_key[134]) );
  DFF_X1 \reg_key_reg[182]  ( .D(Key[182]), .CK(clk), .Q(reg_key[182]) );
  DFF_X1 \reg_key_reg[65]  ( .D(Key[65]), .CK(clk), .Q(reg_key[65]) );
  DFF_X1 \reg_key_reg[37]  ( .D(Key[37]), .CK(clk), .Q(reg_key[37]) );
  DFF_X1 \reg_key_reg[89]  ( .D(Key[89]), .CK(clk), .Q(reg_key[89]) );
  DFF_X1 \reg_key_reg[105]  ( .D(Key[105]), .CK(clk), .Q(reg_key[105]) );
  DFF_X1 \reg_key_reg[110]  ( .D(Key[110]), .CK(clk), .Q(reg_key[110]) );
  DFF_X1 \reg_key_reg[52]  ( .D(Key[52]), .CK(clk), .Q(reg_key[52]) );
  DFF_X1 \reg_key_reg[86]  ( .D(Key[86]), .CK(clk), .Q(reg_key[86]) );
  DFF_X1 \reg_key_reg[28]  ( .D(Key[28]), .CK(clk), .Q(reg_key[28]) );
  DFF_X1 \reg_key_reg[150]  ( .D(Key[150]), .CK(clk), .Q(reg_key[150]) );
  DFF_X1 \reg_key_reg[87]  ( .D(Key[87]), .CK(clk), .Q(reg_key[87]) );
  DFF_X1 \reg_key_reg[46]  ( .D(Key[46]), .CK(clk), .Q(reg_key[46]) );
  DFF_X1 \reg_key_reg[41]  ( .D(Key[41]), .CK(clk), .Q(reg_key[41]) );
  DFF_X2 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CK(clk), .Q(
        Ciphertext[115]) );
  DFF_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CK(clk), .Q(Ciphertext[33])
         );
  DFF_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CK(clk), .Q(Ciphertext[79])
         );
  DFF_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CK(clk), .Q(Ciphertext[87])
         );
  DFFRS_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Ciphertext[58]) );
  DFF_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CK(clk), .Q(Ciphertext[0]) );
  DFF_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CK(clk), .Q(Ciphertext[92])
         );
  DFF_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CK(clk), .Q(
        Ciphertext[160]) );
  SPEEDY_Rounds5_0 SPEEDY_instance ( .Plaintext(reg_in), .Key({
        reg_key[191:187], n3, reg_key[185:0]}), .Ciphertext(reg_out) );
  DFFRS_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Ciphertext[99]) );
  DFFS_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CK(clk), .SN(1'b1), .Q(
        Ciphertext[163]) );
  DFFRS_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CK(clk), .RN(1'b1), .SN(
        1'b1), .Q(Ciphertext[12]) );
  DFF_X2 \reg_key_reg[60]  ( .D(Key[60]), .CK(clk), .Q(reg_key[60]) );
  DFF_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CK(clk), .Q(Ciphertext[8]) );
  DFF_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CK(clk), .Q(Ciphertext[40])
         );
endmodule

